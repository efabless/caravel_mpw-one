magic
tech sky130A
magscale 1 2
timestamp 1606716760
<< checkpaint >>
rect -1260 -1260 170854 14285
<< locali >>
rect 23397 12087 23431 12937
rect 55229 12835 55263 12937
rect 24317 12087 24351 12665
rect 30849 12087 30883 12801
rect 32413 12801 32631 12835
rect 32413 12767 32447 12801
rect 32321 12087 32355 12325
rect 32413 12291 32447 12461
rect 32505 12155 32539 12733
rect 32597 12427 32631 12801
rect 41429 12801 41521 12835
rect 41429 12767 41463 12801
rect 56425 12767 56459 12937
rect 57931 12733 58081 12767
rect 67683 12733 67741 12767
rect 35633 12529 36587 12563
rect 35633 12427 35667 12529
rect 36553 12495 36587 12529
rect 32597 12393 32689 12427
rect 32597 12087 32631 12325
rect 35725 12223 35759 12393
rect 36461 12291 36495 12461
rect 32321 12053 32631 12087
rect 39865 12087 39899 12733
rect 41613 12563 41647 12665
rect 41463 12529 41647 12563
rect 46305 12155 46339 12733
rect 55815 12665 56091 12699
rect 50905 12495 50939 12597
rect 55781 12087 55815 12529
rect 55965 12291 55999 12597
rect 56057 12291 56091 12665
rect 58357 12291 58391 12461
rect 65717 12223 65751 12461
rect 77953 12087 77987 12733
rect 125183 12189 125517 12223
rect 122665 12121 122849 12155
rect 122665 12087 122699 12121
rect 56701 11679 56735 11849
rect 70777 11679 70811 11849
rect 148609 11747 148643 11849
rect 11161 11135 11195 11305
rect 28917 11135 28951 11305
rect 33793 11135 33827 11305
rect 43453 11135 43487 11305
rect 38669 10999 38703 11101
rect 40233 10999 40267 11101
rect 55781 11067 55815 11237
rect 55873 11135 55907 11237
rect 57345 11135 57379 11237
rect 60289 11135 60323 11237
rect 69489 11135 69523 11237
rect 69857 11067 69891 11305
rect 74181 11135 74215 11305
rect 101137 11067 101171 11305
rect 104633 11135 104667 11305
rect 112913 11135 112947 11305
rect 121469 11135 121503 11305
rect 123033 11067 123067 11237
rect 123585 11135 123619 11237
rect 126345 11067 126379 11169
rect 27721 10455 27755 10625
rect 55781 10591 55815 10693
rect 71881 10523 71915 10625
rect 24133 10047 24167 10217
rect 19901 9911 19935 10013
rect 30665 9979 30699 10149
rect 35633 10047 35667 10217
rect 36001 9979 36035 10081
rect 40969 10047 41003 10217
rect 41245 10115 41279 10217
rect 39313 9911 39347 10013
rect 42349 9979 42383 10149
rect 49065 10047 49099 10217
rect 52193 10047 52227 10217
rect 56183 10081 56241 10115
rect 57713 9911 57747 10081
rect 58725 9911 58759 10013
rect 59001 9911 59035 10081
rect 60381 9979 60415 10217
rect 73169 10047 73203 10149
rect 70133 9911 70167 10013
rect 73445 9911 73479 10149
rect 80069 9911 80103 10081
rect 98469 9911 98503 10217
rect 112821 9979 112855 10217
rect 119445 10047 119479 10217
rect 124689 10047 124723 10149
rect 125793 10047 125827 10217
rect 151921 9979 151955 10217
rect 54125 9367 54159 9537
rect 112545 9367 112579 9537
rect 18521 8959 18555 9061
rect 23581 9027 23615 9129
rect 28273 8959 28307 9129
rect 51917 8959 51951 9129
rect 58633 9027 58667 9129
rect 108221 9027 108255 9129
rect 21005 8823 21039 8925
rect 50813 8823 50847 8925
rect 109325 8823 109359 9061
rect 122941 8959 122975 9061
rect 37473 8347 37507 8449
rect 98101 8347 98135 8517
rect 113281 8347 113315 8585
rect 26617 7871 26651 8041
rect 39497 7871 39531 8041
rect 49341 7803 49375 7973
rect 59277 7871 59311 7973
rect 63141 7939 63175 8041
rect 64061 7803 64095 7905
rect 49341 7769 49433 7803
rect 99757 7599 99791 7769
rect 9689 7259 9723 7361
rect 20545 7191 20579 7361
rect 37381 7191 37415 7429
rect 42717 7191 42751 7361
rect 57069 6851 57103 6953
rect 33609 6715 33643 6817
rect 37841 6647 37875 6817
rect 45661 6715 45695 6817
rect 48329 6647 48363 6749
rect 51825 6715 51859 6817
rect 79977 6715 80011 6885
rect 80989 6715 81023 6953
rect 56609 6171 56643 6409
rect 81265 6103 81299 6205
rect 22753 5559 22787 5661
rect 31125 5627 31159 5865
rect 33425 5763 33459 5865
rect 46213 5695 46247 5865
rect 50445 5695 50479 5865
rect 55321 5627 55355 5729
rect 56885 5559 56919 5865
rect 58449 5763 58483 5865
rect 95065 5831 95099 6409
rect 94881 5729 94973 5763
rect 93133 5287 93167 5457
rect 26617 4607 26651 4777
rect 33149 4539 33183 4709
rect 33241 4607 33275 4709
rect 47869 4539 47903 4641
rect 49065 4471 49099 4573
rect 49525 4539 49559 4777
rect 54677 4607 54711 4777
rect 94881 4743 94915 5729
rect 94973 5083 95007 5525
rect 99021 5491 99055 5525
rect 99021 5457 99297 5491
rect 99389 5287 99423 5457
rect 99389 5253 100067 5287
rect 100033 4539 100067 5253
rect 100217 5151 100251 7837
rect 101781 7803 101815 7973
rect 101873 7735 101907 7973
rect 102977 7735 103011 7905
rect 110429 7803 110463 7905
rect 113925 7735 113959 7837
rect 101413 7259 101447 7633
rect 101505 5627 101539 6817
rect 120457 6783 120491 6953
rect 123493 6647 123527 6749
rect 102609 5559 102643 5661
rect 111165 5559 111199 5661
rect 105737 4471 105771 4777
rect 7389 3519 7423 3621
rect 26157 3383 26191 3689
rect 29377 3519 29411 3689
rect 45661 3383 45695 3485
rect 49065 3451 49099 3621
rect 49525 3519 49559 3689
rect 51733 3519 51767 3689
rect 58449 3519 58483 3689
rect 61853 3383 61887 3689
rect 64061 3383 64095 3621
rect 71973 3383 72007 3485
rect 23305 2975 23339 3077
rect 61301 2907 61335 2941
rect 61243 2873 61335 2907
rect 73261 2839 73295 3009
rect 22569 2431 22603 2601
rect 24685 2431 24719 2601
rect 39589 2499 39623 2601
rect 43361 2431 43395 2601
rect 44925 2431 44959 2601
rect 21465 2295 21499 2397
rect 26617 2295 26651 2397
rect 60381 2295 60415 2601
rect 66729 2295 66763 2397
rect 69489 2295 69523 2397
rect 74825 2363 74859 2601
rect 83657 2295 83691 2397
rect 21005 1751 21039 1921
rect 42993 1751 43027 1989
rect 73721 1751 73755 1921
rect 73813 1819 73847 1921
rect 80437 1819 80471 1921
rect 83657 1751 83691 1921
rect 86693 1751 86727 1853
rect 100033 1819 100067 2533
rect 99389 1785 100067 1819
rect 98653 1547 98687 1649
rect 99389 1615 99423 1785
rect 46305 1343 46339 1513
rect 61117 1411 61151 1513
rect 72709 1411 72743 1513
rect 84761 1343 84795 1445
rect 19809 1207 19843 1309
rect 30573 1207 30607 1309
rect 33057 1207 33091 1309
rect 59093 1207 59127 1309
rect 100861 1071 100895 3417
rect 122113 3383 122147 3485
rect 107577 2839 107611 3077
rect 130025 2839 130059 3077
rect 139041 2839 139075 3009
rect 104023 2601 104115 2635
rect 104081 2295 104115 2601
rect 109693 2295 109727 2397
rect 111349 2295 111383 2601
rect 111901 2295 111935 2397
rect 112913 2295 112947 2397
rect 117605 2295 117639 2397
rect 126253 2295 126287 2397
rect 127725 2363 127759 2533
rect 127817 2295 127851 2465
rect 118341 1819 118375 1989
rect 124873 1751 124907 1921
rect 132233 1207 132267 1309
rect 133555 969 133647 1003
rect 3433 867 3467 969
rect 16773 731 16807 833
rect 38485 731 38519 969
rect 48789 799 48823 969
rect 52653 731 52687 833
rect 103989 799 104023 969
rect 120917 663 120951 833
rect 128645 663 128679 833
rect 131405 663 131439 833
rect 133613 663 133647 969
rect 136373 799 136407 969
rect 166641 867 166675 969
rect 138857 663 138891 833
rect 42441 391 42475 425
rect 42165 357 42475 391
rect 42165 119 42199 357
rect 36679 85 41061 119
rect 36461 51 36495 85
rect 42257 51 42291 85
rect 50997 51 51031 425
rect 111349 119 111383 289
rect 36461 17 42291 51
rect 49927 17 51031 51
rect 111257 51 111291 85
rect 111441 51 111475 289
rect 134165 119 134199 289
rect 111257 17 111475 51
<< viali >>
rect 23397 12937 23431 12971
rect 55229 12937 55263 12971
rect 30849 12801 30883 12835
rect 23397 12053 23431 12087
rect 24317 12665 24351 12699
rect 24317 12053 24351 12087
rect 32413 12733 32447 12767
rect 32505 12733 32539 12767
rect 32413 12461 32447 12495
rect 30849 12053 30883 12087
rect 32321 12325 32355 12359
rect 32413 12257 32447 12291
rect 41521 12801 41555 12835
rect 55229 12801 55263 12835
rect 56425 12937 56459 12971
rect 39865 12733 39899 12767
rect 41429 12733 41463 12767
rect 46305 12733 46339 12767
rect 56425 12733 56459 12767
rect 57897 12733 57931 12767
rect 58081 12733 58115 12767
rect 67649 12733 67683 12767
rect 67741 12733 67775 12767
rect 77953 12733 77987 12767
rect 36461 12461 36495 12495
rect 36553 12461 36587 12495
rect 32689 12393 32723 12427
rect 35633 12393 35667 12427
rect 35725 12393 35759 12427
rect 32505 12121 32539 12155
rect 32597 12325 32631 12359
rect 36461 12257 36495 12291
rect 35725 12189 35759 12223
rect 41613 12665 41647 12699
rect 41429 12529 41463 12563
rect 55781 12665 55815 12699
rect 50905 12597 50939 12631
rect 55965 12597 55999 12631
rect 50905 12461 50939 12495
rect 55781 12529 55815 12563
rect 46305 12121 46339 12155
rect 39865 12053 39899 12087
rect 55965 12257 55999 12291
rect 56057 12257 56091 12291
rect 58357 12461 58391 12495
rect 58357 12257 58391 12291
rect 65717 12461 65751 12495
rect 65717 12189 65751 12223
rect 55781 12053 55815 12087
rect 125149 12189 125183 12223
rect 125517 12189 125551 12223
rect 77953 12053 77987 12087
rect 122849 12121 122883 12155
rect 122665 12053 122699 12087
rect 32137 11849 32171 11883
rect 56701 11849 56735 11883
rect 63233 11849 63267 11883
rect 70777 11849 70811 11883
rect 73905 11849 73939 11883
rect 79057 11849 79091 11883
rect 83289 11849 83323 11883
rect 108313 11849 108347 11883
rect 118801 11849 118835 11883
rect 148609 11849 148643 11883
rect 5089 11781 5123 11815
rect 26893 11781 26927 11815
rect 29745 11781 29779 11815
rect 34713 11781 34747 11815
rect 35817 11781 35851 11815
rect 37565 11781 37599 11815
rect 4813 11713 4847 11747
rect 7757 11713 7791 11747
rect 22385 11713 22419 11747
rect 24041 11713 24075 11747
rect 26801 11713 26835 11747
rect 29101 11713 29135 11747
rect 32505 11713 32539 11747
rect 35357 11713 35391 11747
rect 38209 11713 38243 11747
rect 38577 11713 38611 11747
rect 41061 11713 41095 11747
rect 46121 11713 46155 11747
rect 46765 11713 46799 11747
rect 47685 11713 47719 11747
rect 48973 11713 49007 11747
rect 49617 11713 49651 11747
rect 53297 11713 53331 11747
rect 53757 11713 53791 11747
rect 56149 11713 56183 11747
rect 56517 11713 56551 11747
rect 57805 11713 57839 11747
rect 58081 11713 58115 11747
rect 61485 11713 61519 11747
rect 61945 11713 61979 11747
rect 64705 11713 64739 11747
rect 65165 11713 65199 11747
rect 69213 11713 69247 11747
rect 69673 11713 69707 11747
rect 73445 11781 73479 11815
rect 96905 11781 96939 11815
rect 134993 11781 135027 11815
rect 71789 11713 71823 11747
rect 72341 11713 72375 11747
rect 73353 11713 73387 11747
rect 74825 11713 74859 11747
rect 75193 11713 75227 11747
rect 76205 11713 76239 11747
rect 76665 11713 76699 11747
rect 77493 11713 77527 11747
rect 78965 11713 78999 11747
rect 82093 11713 82127 11747
rect 83197 11713 83231 11747
rect 84209 11713 84243 11747
rect 87153 11713 87187 11747
rect 90649 11713 90683 11747
rect 93317 11713 93351 11747
rect 96353 11713 96387 11747
rect 98193 11713 98227 11747
rect 101045 11713 101079 11747
rect 103161 11713 103195 11747
rect 104725 11713 104759 11747
rect 106657 11713 106691 11747
rect 107761 11713 107795 11747
rect 110061 11713 110095 11747
rect 113005 11713 113039 11747
rect 116133 11713 116167 11747
rect 118249 11713 118283 11747
rect 118341 11713 118375 11747
rect 121837 11713 121871 11747
rect 123125 11713 123159 11747
rect 123217 11713 123251 11747
rect 124137 11713 124171 11747
rect 127909 11713 127943 11747
rect 128829 11713 128863 11747
rect 129289 11713 129323 11747
rect 129841 11713 129875 11747
rect 133245 11713 133279 11747
rect 134533 11713 134567 11747
rect 135545 11713 135579 11747
rect 137385 11713 137419 11747
rect 138397 11713 138431 11747
rect 138489 11713 138523 11747
rect 141341 11713 141375 11747
rect 142077 11713 142111 11747
rect 143549 11713 143583 11747
rect 146861 11713 146895 11747
rect 147321 11713 147355 11747
rect 148609 11713 148643 11747
rect 150541 11713 150575 11747
rect 151645 11713 151679 11747
rect 154497 11713 154531 11747
rect 156237 11713 156271 11747
rect 157349 11713 157383 11747
rect 157809 11713 157843 11747
rect 160201 11713 160235 11747
rect 161949 11713 161983 11747
rect 163053 11713 163087 11747
rect 163513 11713 163547 11747
rect 165905 11713 165939 11747
rect 165997 11713 166031 11747
rect 3341 11645 3375 11679
rect 6193 11645 6227 11679
rect 19257 11645 19291 11679
rect 20821 11645 20855 11679
rect 21833 11645 21867 11679
rect 24133 11645 24167 11679
rect 27721 11645 27755 11679
rect 36277 11645 36311 11679
rect 37013 11645 37047 11679
rect 41981 11645 42015 11679
rect 45937 11645 45971 11679
rect 49341 11645 49375 11679
rect 50077 11645 50111 11679
rect 50537 11645 50571 11679
rect 51825 11645 51859 11679
rect 54861 11645 54895 11679
rect 55413 11645 55447 11679
rect 56701 11645 56735 11679
rect 56977 11645 57011 11679
rect 59093 11645 59127 11679
rect 67833 11645 67867 11679
rect 69949 11645 69983 11679
rect 70501 11645 70535 11679
rect 70777 11645 70811 11679
rect 72157 11645 72191 11679
rect 77585 11645 77619 11679
rect 79517 11645 79551 11679
rect 80529 11645 80563 11679
rect 81541 11645 81575 11679
rect 84301 11645 84335 11679
rect 86049 11645 86083 11679
rect 91753 11645 91787 11679
rect 93133 11645 93167 11679
rect 93685 11645 93719 11679
rect 94605 11645 94639 11679
rect 99205 11645 99239 11679
rect 99665 11645 99699 11679
rect 101965 11645 101999 11679
rect 102057 11645 102091 11679
rect 104633 11645 104667 11679
rect 108957 11645 108991 11679
rect 111717 11645 111751 11679
rect 113097 11645 113131 11679
rect 114569 11645 114603 11679
rect 115857 11645 115891 11679
rect 120273 11645 120307 11679
rect 121285 11645 121319 11679
rect 124229 11645 124263 11679
rect 126345 11645 126379 11679
rect 127357 11645 127391 11679
rect 131681 11645 131715 11679
rect 132693 11645 132727 11679
rect 138857 11645 138891 11679
rect 140237 11645 140271 11679
rect 141249 11645 141283 11679
rect 144561 11645 144595 11679
rect 146585 11645 146619 11679
rect 148793 11645 148827 11679
rect 156981 11645 157015 11679
rect 158361 11645 158395 11679
rect 164801 11645 164835 11679
rect 166365 11645 166399 11679
rect 7665 11577 7699 11611
rect 110245 11577 110279 11611
rect 129933 11577 129967 11611
rect 134625 11577 134659 11611
rect 143641 11577 143675 11611
rect 150633 11577 150667 11611
rect 152105 11577 152139 11611
rect 156337 11577 156371 11611
rect 160293 11577 160327 11611
rect 4169 11509 4203 11543
rect 5825 11509 5859 11543
rect 9597 11509 9631 11543
rect 20177 11509 20211 11543
rect 27261 11509 27295 11543
rect 40693 11509 40727 11543
rect 52469 11509 52503 11543
rect 53113 11509 53147 11543
rect 55965 11509 55999 11543
rect 57621 11509 57655 11543
rect 59737 11509 59771 11543
rect 61301 11509 61335 11543
rect 64521 11509 64555 11543
rect 69029 11509 69063 11543
rect 70961 11509 70995 11543
rect 72801 11509 72835 11543
rect 74733 11509 74767 11543
rect 76297 11509 76331 11543
rect 77033 11509 77067 11543
rect 80161 11509 80195 11543
rect 87245 11509 87279 11543
rect 95525 11509 95559 11543
rect 96445 11509 96479 11543
rect 98285 11509 98319 11543
rect 106749 11509 106783 11543
rect 107117 11509 107151 11543
rect 107853 11509 107887 11543
rect 111257 11509 111291 11543
rect 116501 11509 116535 11543
rect 117973 11509 118007 11543
rect 124689 11509 124723 11543
rect 128921 11509 128955 11543
rect 130393 11509 130427 11543
rect 134349 11509 134383 11543
rect 135637 11509 135671 11543
rect 136005 11509 136039 11543
rect 137477 11509 137511 11543
rect 138121 11509 138155 11543
rect 144009 11509 144043 11543
rect 146953 11509 146987 11543
rect 151001 11509 151035 11543
rect 151737 11509 151771 11543
rect 154589 11509 154623 11543
rect 157441 11509 157475 11543
rect 162041 11509 162075 11543
rect 163145 11509 163179 11543
rect 4813 11305 4847 11339
rect 11161 11305 11195 11339
rect 11437 11305 11471 11339
rect 16497 11305 16531 11339
rect 22385 11305 22419 11339
rect 23581 11305 23615 11339
rect 28917 11305 28951 11339
rect 29193 11305 29227 11339
rect 29469 11305 29503 11339
rect 30113 11305 30147 11339
rect 33241 11305 33275 11339
rect 33793 11305 33827 11339
rect 34069 11305 34103 11339
rect 39681 11305 39715 11339
rect 42901 11305 42935 11339
rect 43453 11305 43487 11339
rect 43729 11305 43763 11339
rect 69857 11305 69891 11339
rect 70777 11305 70811 11339
rect 72341 11305 72375 11339
rect 74181 11305 74215 11339
rect 74457 11305 74491 11339
rect 75009 11305 75043 11339
rect 75377 11305 75411 11339
rect 77677 11305 77711 11339
rect 77953 11305 77987 11339
rect 78965 11305 78999 11339
rect 82001 11305 82035 11339
rect 83013 11305 83047 11339
rect 83381 11305 83415 11339
rect 84761 11305 84795 11339
rect 87153 11305 87187 11339
rect 98193 11305 98227 11339
rect 101137 11305 101171 11339
rect 101413 11305 101447 11339
rect 104081 11305 104115 11339
rect 104633 11305 104667 11339
rect 104909 11305 104943 11339
rect 105277 11305 105311 11339
rect 106565 11305 106599 11339
rect 112913 11305 112947 11339
rect 113189 11305 113223 11339
rect 121285 11305 121319 11339
rect 121469 11305 121503 11339
rect 121745 11305 121779 11339
rect 122021 11305 122055 11339
rect 123125 11305 123159 11339
rect 124229 11305 124263 11339
rect 127725 11305 127759 11339
rect 130485 11305 130519 11339
rect 132509 11305 132543 11339
rect 133245 11305 133279 11339
rect 136097 11305 136131 11339
rect 137477 11305 137511 11339
rect 141065 11305 141099 11339
rect 156245 11305 156279 11339
rect 160201 11305 160235 11339
rect 162317 11305 162351 11339
rect 165905 11305 165939 11339
rect 7205 11237 7239 11271
rect 2237 11169 2271 11203
rect 4537 11169 4571 11203
rect 7665 11169 7699 11203
rect 9505 11169 9539 11203
rect 10977 11169 11011 11203
rect 16037 11237 16071 11271
rect 24225 11237 24259 11271
rect 24593 11237 24627 11271
rect 26617 11237 26651 11271
rect 21189 11169 21223 11203
rect 27261 11169 27295 11203
rect 28273 11169 28307 11203
rect 30757 11237 30791 11271
rect 32137 11169 32171 11203
rect 35541 11169 35575 11203
rect 37013 11169 37047 11203
rect 38025 11169 38059 11203
rect 49157 11237 49191 11271
rect 50997 11237 51031 11271
rect 51641 11237 51675 11271
rect 55781 11237 55815 11271
rect 4169 11101 4203 11135
rect 5733 11101 5767 11135
rect 7297 11101 7331 11135
rect 8033 11101 8067 11135
rect 11069 11101 11103 11135
rect 11161 11101 11195 11135
rect 14565 11101 14599 11135
rect 16129 11101 16163 11135
rect 20177 11101 20211 11135
rect 21741 11101 21775 11135
rect 22109 11101 22143 11135
rect 23765 11101 23799 11135
rect 28825 11101 28859 11135
rect 28917 11101 28951 11135
rect 30297 11101 30331 11135
rect 31217 11101 31251 11135
rect 32045 11101 32079 11135
rect 33609 11101 33643 11135
rect 33793 11101 33827 11135
rect 34529 11101 34563 11135
rect 36093 11101 36127 11135
rect 38485 11101 38519 11135
rect 38669 11101 38703 11135
rect 40049 11101 40083 11135
rect 40233 11101 40267 11135
rect 40969 11101 41003 11135
rect 41613 11101 41647 11135
rect 42073 11101 42107 11135
rect 43269 11101 43303 11135
rect 43453 11101 43487 11135
rect 45845 11101 45879 11135
rect 46029 11101 46063 11135
rect 46305 11101 46339 11135
rect 47133 11101 47167 11135
rect 49709 11101 49743 11135
rect 50997 11101 51031 11135
rect 52469 11101 52503 11135
rect 52561 11101 52595 11135
rect 52929 11101 52963 11135
rect 53297 11101 53331 11135
rect 55137 11101 55171 11135
rect 55321 11101 55355 11135
rect 55505 11101 55539 11135
rect 11989 11033 12023 11067
rect 13461 11033 13495 11067
rect 14289 11033 14323 11067
rect 18889 11033 18923 11067
rect 19993 11033 20027 11067
rect 25789 11033 25823 11067
rect 32413 11033 32447 11067
rect 34437 11033 34471 11067
rect 36461 11033 36495 11067
rect 38945 11033 38979 11067
rect 24685 10965 24719 10999
rect 38669 10965 38703 10999
rect 55873 11237 55907 11271
rect 57345 11237 57379 11271
rect 57621 11237 57655 11271
rect 59553 11237 59587 11271
rect 60289 11237 60323 11271
rect 60565 11237 60599 11271
rect 61117 11237 61151 11271
rect 68753 11237 68787 11271
rect 69489 11237 69523 11271
rect 69765 11237 69799 11271
rect 55873 11101 55907 11135
rect 56057 11101 56091 11135
rect 56425 11101 56459 11135
rect 56793 11101 56827 11135
rect 56885 11101 56919 11135
rect 57253 11101 57287 11135
rect 57345 11101 57379 11135
rect 59737 11101 59771 11135
rect 60197 11101 60231 11135
rect 60289 11101 60323 11135
rect 60933 11101 60967 11135
rect 61301 11101 61335 11135
rect 61761 11101 61795 11135
rect 62129 11101 62163 11135
rect 63601 11101 63635 11135
rect 64705 11101 64739 11135
rect 66085 11101 66119 11135
rect 67649 11101 67683 11135
rect 68569 11101 68603 11135
rect 68937 11101 68971 11135
rect 69397 11101 69431 11135
rect 69489 11101 69523 11135
rect 72525 11169 72559 11203
rect 73537 11169 73571 11203
rect 76389 11237 76423 11271
rect 85405 11237 85439 11271
rect 92949 11237 92983 11271
rect 96997 11237 97031 11271
rect 100953 11237 100987 11271
rect 78321 11169 78355 11203
rect 80437 11169 80471 11203
rect 81725 11169 81759 11203
rect 84393 11169 84427 11203
rect 93133 11169 93167 11203
rect 94145 11169 94179 11203
rect 95525 11169 95559 11203
rect 99481 11169 99515 11203
rect 70133 11101 70167 11135
rect 70685 11101 70719 11135
rect 71237 11101 71271 11135
rect 71697 11101 71731 11135
rect 74089 11101 74123 11135
rect 74181 11101 74215 11135
rect 74917 11101 74951 11135
rect 75745 11101 75779 11135
rect 76297 11101 76331 11135
rect 76849 11101 76883 11135
rect 77309 11101 77343 11135
rect 77861 11101 77895 11135
rect 79425 11101 79459 11135
rect 80989 11101 81023 11135
rect 81909 11101 81943 11135
rect 82369 11101 82403 11135
rect 82921 11101 82955 11135
rect 83749 11101 83783 11135
rect 83933 11101 83967 11135
rect 84945 11101 84979 11135
rect 94697 11101 94731 11135
rect 96629 11101 96663 11135
rect 97365 11101 97399 11135
rect 100769 11101 100803 11135
rect 101873 11169 101907 11203
rect 103161 11169 103195 11203
rect 108129 11237 108163 11271
rect 112729 11237 112763 11271
rect 105645 11169 105679 11203
rect 106657 11169 106691 11203
rect 110889 11169 110923 11203
rect 111257 11169 111291 11203
rect 113557 11169 113591 11203
rect 115029 11169 115063 11203
rect 116593 11169 116627 11203
rect 117973 11169 118007 11203
rect 118985 11169 119019 11203
rect 103437 11101 103471 11135
rect 104357 11101 104391 11135
rect 104633 11101 104667 11135
rect 108221 11101 108255 11135
rect 108589 11101 108623 11135
rect 109969 11101 110003 11135
rect 110521 11101 110555 11135
rect 112821 11101 112855 11135
rect 112913 11101 112947 11135
rect 114477 11101 114511 11135
rect 115397 11101 115431 11135
rect 115581 11101 115615 11135
rect 117145 11101 117179 11135
rect 119537 11101 119571 11135
rect 119905 11101 119939 11135
rect 121193 11101 121227 11135
rect 121469 11101 121503 11135
rect 123033 11237 123067 11271
rect 123401 11237 123435 11271
rect 123585 11237 123619 11271
rect 123861 11237 123895 11271
rect 126161 11237 126195 11271
rect 128553 11237 128587 11271
rect 139317 11237 139351 11271
rect 150449 11237 150483 11271
rect 125333 11169 125367 11203
rect 126345 11169 126379 11203
rect 126897 11169 126931 11203
rect 129657 11169 129691 11203
rect 132877 11169 132911 11203
rect 135269 11169 135303 11203
rect 141157 11169 141191 11203
rect 142353 11169 142387 11203
rect 144653 11169 144687 11203
rect 146493 11169 146527 11203
rect 147505 11169 147539 11203
rect 149529 11169 149563 11203
rect 150541 11169 150575 11203
rect 151553 11169 151587 11203
rect 157901 11169 157935 11203
rect 163881 11169 163915 11203
rect 166089 11169 166123 11203
rect 167101 11169 167135 11203
rect 123309 11101 123343 11135
rect 123585 11101 123619 11135
rect 124321 11101 124355 11135
rect 125885 11101 125919 11135
rect 40509 11033 40543 11067
rect 44649 11033 44683 11067
rect 49617 11033 49651 11067
rect 53573 11033 53607 11067
rect 53941 11033 53975 11067
rect 55781 11033 55815 11067
rect 57989 11033 58023 11067
rect 62589 11033 62623 11067
rect 65625 11033 65659 11067
rect 69857 11033 69891 11067
rect 74825 11033 74859 11067
rect 81357 11033 81391 11067
rect 84025 11033 84059 11067
rect 85037 11033 85071 11067
rect 87521 11033 87555 11067
rect 91753 11033 91787 11067
rect 92029 11033 92063 11067
rect 95065 11033 95099 11067
rect 101137 11033 101171 11067
rect 103805 11033 103839 11067
rect 104449 11033 104483 11067
rect 110061 11033 110095 11067
rect 114385 11033 114419 11067
rect 117513 11033 117547 11067
rect 120273 11033 120307 11067
rect 122205 11033 122239 11067
rect 123033 11033 123067 11067
rect 126805 11101 126839 11135
rect 127265 11101 127299 11135
rect 128645 11101 128679 11135
rect 130209 11101 130243 11135
rect 131037 11101 131071 11135
rect 131497 11101 131531 11135
rect 132417 11101 132451 11135
rect 134257 11101 134291 11135
rect 135821 11101 135855 11135
rect 136649 11101 136683 11135
rect 137109 11101 137143 11135
rect 138029 11101 138063 11135
rect 139133 11101 139167 11135
rect 139869 11101 139903 11135
rect 142261 11101 142295 11135
rect 142997 11101 143031 11135
rect 143365 11101 143399 11135
rect 143641 11101 143675 11135
rect 145021 11101 145055 11135
rect 145481 11101 145515 11135
rect 147597 11101 147631 11135
rect 148333 11101 148367 11135
rect 151645 11101 151679 11135
rect 152381 11101 152415 11135
rect 156889 11101 156923 11135
rect 157993 11101 158027 11135
rect 158729 11101 158763 11135
rect 162869 11101 162903 11135
rect 163973 11101 164007 11135
rect 164709 11101 164743 11135
rect 167193 11101 167227 11135
rect 167929 11101 167963 11135
rect 126345 11033 126379 11067
rect 126621 11033 126655 11067
rect 131129 11033 131163 11067
rect 131957 11033 131991 11067
rect 136741 11033 136775 11067
rect 140237 11033 140271 11067
rect 152933 11033 152967 11067
rect 154497 11033 154531 11067
rect 161857 11033 161891 11067
rect 162685 11033 162719 11067
rect 40233 10965 40267 10999
rect 40785 10965 40819 10999
rect 46765 10965 46799 10999
rect 48237 10965 48271 10999
rect 54493 10965 54527 10999
rect 58081 10965 58115 10999
rect 58541 10965 58575 10999
rect 62497 10965 62531 10999
rect 65073 10965 65107 10999
rect 85957 10965 85991 10999
rect 90373 10965 90407 10999
rect 109049 10965 109083 10999
rect 114569 10965 114603 10999
rect 155141 10965 155175 10999
rect 159281 10965 159315 10999
rect 6285 10761 6319 10795
rect 10149 10761 10183 10795
rect 23581 10761 23615 10795
rect 60657 10761 60691 10795
rect 72065 10761 72099 10795
rect 75101 10761 75135 10795
rect 78321 10761 78355 10795
rect 83105 10761 83139 10795
rect 86969 10761 87003 10795
rect 90465 10761 90499 10795
rect 91017 10761 91051 10795
rect 94605 10761 94639 10795
rect 118525 10761 118559 10795
rect 124781 10761 124815 10795
rect 128185 10761 128219 10795
rect 131957 10761 131991 10795
rect 24501 10693 24535 10727
rect 30849 10693 30883 10727
rect 32413 10693 32447 10727
rect 34529 10693 34563 10727
rect 45385 10693 45419 10727
rect 47409 10693 47443 10727
rect 55781 10693 55815 10727
rect 56057 10693 56091 10727
rect 82645 10693 82679 10727
rect 135269 10693 135303 10727
rect 139501 10693 139535 10727
rect 4353 10625 4387 10659
rect 4721 10625 4755 10659
rect 5089 10625 5123 10659
rect 9321 10625 9355 10659
rect 12633 10625 12667 10659
rect 14197 10625 14231 10659
rect 18705 10625 18739 10659
rect 19717 10625 19751 10659
rect 21281 10625 21315 10659
rect 21649 10625 21683 10659
rect 24409 10625 24443 10659
rect 25881 10625 25915 10659
rect 26065 10625 26099 10659
rect 27445 10625 27479 10659
rect 27721 10625 27755 10659
rect 29009 10625 29043 10659
rect 29285 10625 29319 10659
rect 30757 10625 30791 10659
rect 32229 10625 32263 10659
rect 35173 10625 35207 10659
rect 37473 10625 37507 10659
rect 41153 10625 41187 10659
rect 42717 10625 42751 10659
rect 46397 10625 46431 10659
rect 47133 10625 47167 10659
rect 47961 10625 47995 10659
rect 49525 10625 49559 10659
rect 51089 10625 51123 10659
rect 51733 10625 51767 10659
rect 52561 10625 52595 10659
rect 53297 10625 53331 10659
rect 54953 10625 54987 10659
rect 55505 10625 55539 10659
rect 3341 10557 3375 10591
rect 6745 10557 6779 10591
rect 7757 10557 7791 10591
rect 16221 10557 16255 10591
rect 17325 10557 17359 10591
rect 20729 10557 20763 10591
rect 9229 10489 9263 10523
rect 14105 10489 14139 10523
rect 18613 10489 18647 10523
rect 57161 10625 57195 10659
rect 58725 10625 58759 10659
rect 59829 10625 59863 10659
rect 60289 10625 60323 10659
rect 62221 10625 62255 10659
rect 66269 10625 66303 10659
rect 68661 10625 68695 10659
rect 69397 10625 69431 10659
rect 70225 10625 70259 10659
rect 71789 10625 71823 10659
rect 71881 10625 71915 10659
rect 73629 10625 73663 10659
rect 73997 10625 74031 10659
rect 75009 10625 75043 10659
rect 77677 10625 77711 10659
rect 79057 10625 79091 10659
rect 81725 10625 81759 10659
rect 82553 10625 82587 10659
rect 83565 10625 83599 10659
rect 85773 10625 85807 10659
rect 86509 10625 86543 10659
rect 87061 10625 87095 10659
rect 88349 10625 88383 10659
rect 88901 10625 88935 10659
rect 93777 10625 93811 10659
rect 98929 10625 98963 10659
rect 103805 10625 103839 10659
rect 106197 10625 106231 10659
rect 108773 10625 108807 10659
rect 111349 10625 111383 10659
rect 114661 10625 114695 10659
rect 117237 10625 117271 10659
rect 121101 10625 121135 10659
rect 122849 10625 122883 10659
rect 124689 10625 124723 10659
rect 127265 10625 127299 10659
rect 128093 10625 128127 10659
rect 130669 10625 130703 10659
rect 134073 10625 134107 10659
rect 135177 10625 135211 10659
rect 137293 10625 137327 10659
rect 139041 10625 139075 10659
rect 142169 10625 142203 10659
rect 144929 10625 144963 10659
rect 145665 10625 145699 10659
rect 147873 10625 147907 10659
rect 150909 10625 150943 10659
rect 153209 10625 153243 10659
rect 155969 10625 156003 10659
rect 158453 10625 158487 10659
rect 159557 10625 159591 10659
rect 161121 10625 161155 10659
rect 162869 10625 162903 10659
rect 164341 10625 164375 10659
rect 166733 10625 166767 10659
rect 36093 10557 36127 10591
rect 37105 10557 37139 10591
rect 38025 10557 38059 10591
rect 38485 10557 38519 10591
rect 42441 10557 42475 10591
rect 44281 10557 44315 10591
rect 46029 10557 46063 10591
rect 48973 10557 49007 10591
rect 51365 10557 51399 10591
rect 55781 10557 55815 10591
rect 59921 10557 59955 10591
rect 61117 10557 61151 10591
rect 63233 10557 63267 10591
rect 64889 10557 64923 10591
rect 76205 10557 76239 10591
rect 77401 10557 77435 10591
rect 80161 10557 80195 10591
rect 81173 10557 81207 10591
rect 84669 10557 84703 10591
rect 85681 10557 85715 10591
rect 88073 10557 88107 10591
rect 92213 10557 92247 10591
rect 93225 10557 93259 10591
rect 95893 10557 95927 10591
rect 97365 10557 97399 10591
rect 98469 10557 98503 10591
rect 99757 10557 99791 10591
rect 102241 10557 102275 10591
rect 103253 10557 103287 10591
rect 104633 10557 104667 10591
rect 106105 10557 106139 10591
rect 107669 10557 107703 10591
rect 110061 10557 110095 10591
rect 113281 10557 113315 10591
rect 114753 10557 114787 10591
rect 115673 10557 115707 10591
rect 116685 10557 116719 10591
rect 119537 10557 119571 10591
rect 120549 10557 120583 10591
rect 125701 10557 125735 10591
rect 126713 10557 126747 10591
rect 129565 10557 129599 10591
rect 130577 10557 130611 10591
rect 132969 10557 133003 10591
rect 134165 10557 134199 10591
rect 136189 10557 136223 10591
rect 137201 10557 137235 10591
rect 139133 10557 139167 10591
rect 140973 10557 141007 10591
rect 143825 10557 143859 10591
rect 146401 10557 146435 10591
rect 149345 10557 149379 10591
rect 152013 10557 152047 10591
rect 154773 10557 154807 10591
rect 156153 10557 156187 10591
rect 159465 10557 159499 10591
rect 162133 10557 162167 10591
rect 163237 10557 163271 10591
rect 164249 10557 164283 10591
rect 165629 10557 165663 10591
rect 166641 10557 166675 10591
rect 46489 10489 46523 10523
rect 58449 10489 58483 10523
rect 66177 10489 66211 10523
rect 68753 10489 68787 10523
rect 71513 10489 71547 10523
rect 71881 10489 71915 10523
rect 73537 10489 73571 10523
rect 83657 10489 83691 10523
rect 108957 10489 108991 10523
rect 111533 10489 111567 10523
rect 142261 10489 142295 10523
rect 145113 10489 145147 10523
rect 147873 10489 147907 10523
rect 150817 10489 150851 10523
rect 153301 10489 153335 10523
rect 3985 10421 4019 10455
rect 27353 10421 27387 10455
rect 27721 10421 27755 10455
rect 27905 10421 27939 10455
rect 32689 10421 32723 10455
rect 35541 10421 35575 10455
rect 49985 10421 50019 10455
rect 52009 10421 52043 10455
rect 52653 10421 52687 10455
rect 55045 10421 55079 10455
rect 56333 10421 56367 10455
rect 61669 10421 61703 10455
rect 72433 10421 72467 10455
rect 74457 10421 74491 10455
rect 79149 10421 79183 10455
rect 94145 10421 94179 10455
rect 111901 10421 111935 10455
rect 112913 10421 112947 10455
rect 121377 10421 121411 10455
rect 122573 10421 122607 10455
rect 122941 10421 122975 10455
rect 127633 10421 127667 10455
rect 128553 10421 128587 10455
rect 132417 10421 132451 10455
rect 133705 10421 133739 10455
rect 138029 10421 138063 10455
rect 140421 10421 140455 10455
rect 157993 10421 158027 10455
rect 160477 10421 160511 10455
rect 5365 10217 5399 10251
rect 8309 10217 8343 10251
rect 9229 10217 9263 10251
rect 12633 10217 12667 10251
rect 14013 10217 14047 10251
rect 17325 10217 17359 10251
rect 18705 10217 18739 10251
rect 19717 10217 19751 10251
rect 24133 10217 24167 10251
rect 24409 10217 24443 10251
rect 30849 10217 30883 10251
rect 34713 10217 34747 10251
rect 35633 10217 35667 10251
rect 35909 10217 35943 10251
rect 40325 10217 40359 10251
rect 40969 10217 41003 10251
rect 41061 10217 41095 10251
rect 41245 10217 41279 10251
rect 41521 10217 41555 10251
rect 48053 10217 48087 10251
rect 48329 10217 48363 10251
rect 49065 10217 49099 10251
rect 49341 10217 49375 10251
rect 50905 10217 50939 10251
rect 52193 10217 52227 10251
rect 53573 10217 53607 10251
rect 55137 10217 55171 10251
rect 55413 10217 55447 10251
rect 60381 10217 60415 10251
rect 60841 10217 60875 10251
rect 65257 10217 65291 10251
rect 68753 10217 68787 10251
rect 69397 10217 69431 10251
rect 70317 10217 70351 10251
rect 70777 10217 70811 10251
rect 74825 10217 74859 10251
rect 75561 10217 75595 10251
rect 76389 10217 76423 10251
rect 76757 10217 76791 10251
rect 78229 10217 78263 10251
rect 78413 10217 78447 10251
rect 79057 10217 79091 10251
rect 80253 10217 80287 10251
rect 80437 10217 80471 10251
rect 81541 10217 81575 10251
rect 82737 10217 82771 10251
rect 83565 10217 83599 10251
rect 84669 10217 84703 10251
rect 89453 10217 89487 10251
rect 95893 10217 95927 10251
rect 98009 10217 98043 10251
rect 98377 10217 98411 10251
rect 98469 10217 98503 10251
rect 99573 10217 99607 10251
rect 107669 10217 107703 10251
rect 108957 10217 108991 10251
rect 111441 10217 111475 10251
rect 112821 10217 112855 10251
rect 117145 10217 117179 10251
rect 119445 10217 119479 10251
rect 119537 10217 119571 10251
rect 123125 10217 123159 10251
rect 124965 10217 124999 10251
rect 125793 10217 125827 10251
rect 125977 10217 126011 10251
rect 127357 10217 127391 10251
rect 127909 10217 127943 10251
rect 130301 10217 130335 10251
rect 134257 10217 134291 10251
rect 135269 10217 135303 10251
rect 137477 10217 137511 10251
rect 149069 10217 149103 10251
rect 151921 10217 151955 10251
rect 152105 10217 152139 10251
rect 153301 10217 153335 10251
rect 155325 10217 155359 10251
rect 156337 10217 156371 10251
rect 157901 10217 157935 10251
rect 159833 10217 159867 10251
rect 162685 10217 162719 10251
rect 165077 10217 165111 10251
rect 165629 10217 165663 10251
rect 166917 10217 166951 10251
rect 4169 10081 4203 10115
rect 7113 10081 7147 10115
rect 19073 10081 19107 10115
rect 20177 10081 20211 10115
rect 21189 10081 21223 10115
rect 25605 10149 25639 10183
rect 27077 10149 27111 10183
rect 28917 10149 28951 10183
rect 30665 10149 30699 10183
rect 34897 10149 34931 10183
rect 24777 10081 24811 10115
rect 27445 10081 27479 10115
rect 3985 10013 4019 10047
rect 4537 10013 4571 10047
rect 6101 10013 6135 10047
rect 7665 10013 7699 10047
rect 19901 10013 19935 10047
rect 21741 10013 21775 10047
rect 22109 10013 22143 10047
rect 23581 10013 23615 10047
rect 23673 10013 23707 10047
rect 24041 10013 24075 10047
rect 24133 10013 24167 10047
rect 26617 10013 26651 10047
rect 26709 10013 26743 10047
rect 27813 10013 27847 10047
rect 27905 10013 27939 10047
rect 28273 10013 28307 10047
rect 28641 10013 28675 10047
rect 32597 10013 32631 10047
rect 32689 10013 32723 10047
rect 33057 10013 33091 10047
rect 35081 10013 35115 10047
rect 35541 10013 35575 10047
rect 35633 10013 35667 10047
rect 36001 10081 36035 10115
rect 37473 10081 37507 10115
rect 37657 10081 37691 10115
rect 38669 10081 38703 10115
rect 30665 9945 30699 9979
rect 41245 10081 41279 10115
rect 42349 10149 42383 10183
rect 39221 10013 39255 10047
rect 39313 10013 39347 10047
rect 40693 10013 40727 10047
rect 40969 10013 41003 10047
rect 36001 9945 36035 9979
rect 49709 10149 49743 10183
rect 49893 10149 49927 10183
rect 56149 10081 56183 10115
rect 56241 10081 56275 10115
rect 57713 10081 57747 10115
rect 45845 10013 45879 10047
rect 46213 10013 46247 10047
rect 46581 10013 46615 10047
rect 46949 10013 46983 10047
rect 48421 10013 48455 10047
rect 48973 10013 49007 10047
rect 49065 10013 49099 10047
rect 49985 10013 50019 10047
rect 50537 10013 50571 10047
rect 51641 10013 51675 10047
rect 51733 10013 51767 10047
rect 52101 10013 52135 10047
rect 52193 10013 52227 10047
rect 52469 10013 52503 10047
rect 55597 10013 55631 10047
rect 56057 10013 56091 10047
rect 56425 10013 56459 10047
rect 57161 10013 57195 10047
rect 57253 10013 57287 10047
rect 57529 10013 57563 10047
rect 42349 9945 42383 9979
rect 47317 9945 47351 9979
rect 53297 9945 53331 9979
rect 59001 10081 59035 10115
rect 58725 10013 58759 10047
rect 57989 9945 58023 9979
rect 59277 10013 59311 10047
rect 59645 10013 59679 10047
rect 59829 10013 59863 10047
rect 60197 10013 60231 10047
rect 73169 10149 73203 10183
rect 68937 10081 68971 10115
rect 72065 10081 72099 10115
rect 73445 10149 73479 10183
rect 79425 10149 79459 10183
rect 91937 10149 91971 10183
rect 97549 10149 97583 10183
rect 73261 10081 73295 10115
rect 60473 10013 60507 10047
rect 61025 10013 61059 10047
rect 62037 10013 62071 10047
rect 70133 10013 70167 10047
rect 70869 10013 70903 10047
rect 71421 10013 71455 10047
rect 71697 10013 71731 10047
rect 72433 10013 72467 10047
rect 72617 10013 72651 10047
rect 72801 10013 72835 10047
rect 73169 10013 73203 10047
rect 60381 9945 60415 9979
rect 5089 9877 5123 9911
rect 6009 9877 6043 9911
rect 8033 9877 8067 9911
rect 16405 9877 16439 9911
rect 19901 9877 19935 9911
rect 29101 9877 29135 9911
rect 30297 9877 30331 9911
rect 32137 9877 32171 9911
rect 33425 9877 33459 9911
rect 36277 9877 36311 9911
rect 39313 9877 39347 9911
rect 39589 9877 39623 9911
rect 42625 9877 42659 9911
rect 43177 9877 43211 9911
rect 51181 9877 51215 9911
rect 52837 9877 52871 9911
rect 54309 9877 54343 9911
rect 56793 9877 56827 9911
rect 57713 9877 57747 9911
rect 58541 9877 58575 9911
rect 58725 9877 58759 9911
rect 58909 9877 58943 9911
rect 59001 9877 59035 9911
rect 63049 9877 63083 9911
rect 66269 9877 66303 9911
rect 70133 9877 70167 9911
rect 79793 10081 79827 10115
rect 80069 10081 80103 10115
rect 83013 10081 83047 10115
rect 83933 10081 83967 10115
rect 85037 10081 85071 10115
rect 86049 10081 86083 10115
rect 88533 10081 88567 10115
rect 90465 10081 90499 10115
rect 94145 10081 94179 10115
rect 96077 10081 96111 10115
rect 74089 10013 74123 10047
rect 74181 10013 74215 10047
rect 74365 10013 74399 10047
rect 75193 10013 75227 10047
rect 76297 10013 76331 10047
rect 77309 10013 77343 10047
rect 77769 10013 77803 10047
rect 78321 10013 78355 10047
rect 79333 10013 79367 10047
rect 77401 9945 77435 9979
rect 80345 10013 80379 10047
rect 80805 10013 80839 10047
rect 81909 10013 81943 10047
rect 82369 10013 82403 10047
rect 82921 10013 82955 10047
rect 86601 10013 86635 10047
rect 87521 10013 87555 10047
rect 88993 10013 89027 10047
rect 91937 10013 91971 10047
rect 92305 10013 92339 10047
rect 93133 10013 93167 10047
rect 94237 10013 94271 10047
rect 94973 10013 95007 10047
rect 97641 10013 97675 10047
rect 82001 9945 82035 9979
rect 98929 10081 98963 10115
rect 99665 10081 99699 10115
rect 100861 10081 100895 10115
rect 102241 10081 102275 10115
rect 102701 10081 102735 10115
rect 107025 10081 107059 10115
rect 108129 10081 108163 10115
rect 110429 10081 110463 10115
rect 110981 10081 111015 10115
rect 101229 10013 101263 10047
rect 101597 10013 101631 10047
rect 114293 10081 114327 10115
rect 115581 10081 115615 10115
rect 116593 10081 116627 10115
rect 117605 10081 117639 10115
rect 124689 10149 124723 10183
rect 125333 10149 125367 10183
rect 122205 10081 122239 10115
rect 146217 10149 146251 10183
rect 150725 10149 150759 10183
rect 126897 10081 126931 10115
rect 129013 10081 129047 10115
rect 130485 10081 130519 10115
rect 131221 10081 131255 10115
rect 132417 10081 132451 10115
rect 133429 10081 133463 10115
rect 136281 10081 136315 10115
rect 136741 10081 136775 10115
rect 139041 10081 139075 10115
rect 141433 10081 141467 10115
rect 142261 10081 142295 10115
rect 151645 10081 151679 10115
rect 112913 10013 112947 10047
rect 114385 10013 114419 10047
rect 114753 10013 114787 10047
rect 119077 10013 119111 10047
rect 119445 10013 119479 10047
rect 120089 10013 120123 10047
rect 121193 10013 121227 10047
rect 122757 10013 122791 10047
rect 124413 10013 124447 10047
rect 124689 10013 124723 10047
rect 125425 10013 125459 10047
rect 125793 10013 125827 10047
rect 126805 10013 126839 10047
rect 128001 10013 128035 10047
rect 129565 10013 129599 10047
rect 130393 10013 130427 10047
rect 130853 10013 130887 10047
rect 133521 10013 133555 10047
rect 134809 10013 134843 10047
rect 135637 10013 135671 10047
rect 138029 10013 138063 10047
rect 139133 10013 139167 10047
rect 140421 10013 140455 10047
rect 141525 10013 141559 10047
rect 142629 10013 142663 10047
rect 144745 10013 144779 10047
rect 146309 10013 146343 10047
rect 149253 10013 149287 10047
rect 150357 10013 150391 10047
rect 156981 10081 157015 10115
rect 157993 10081 158027 10115
rect 159373 10081 159407 10115
rect 160477 10081 160511 10115
rect 161489 10081 161523 10115
rect 162869 10081 162903 10115
rect 163881 10081 163915 10115
rect 166089 10081 166123 10115
rect 159557 10013 159591 10047
rect 161581 10013 161615 10047
rect 162317 10013 162351 10047
rect 163973 10013 164007 10047
rect 164709 10013 164743 10047
rect 109969 9945 110003 9979
rect 112821 9945 112855 9979
rect 115213 9945 115247 9979
rect 125517 9945 125551 9979
rect 134901 9945 134935 9979
rect 139869 9945 139903 9979
rect 143641 9945 143675 9979
rect 147781 9945 147815 9979
rect 148701 9945 148735 9979
rect 151921 9945 151955 9979
rect 152657 9945 152691 9979
rect 73445 9877 73479 9911
rect 73629 9877 73663 9911
rect 76113 9877 76147 9911
rect 80069 9877 80103 9911
rect 86969 9877 87003 9911
rect 87245 9877 87279 9911
rect 92765 9877 92799 9911
rect 98469 9877 98503 9911
rect 103253 9877 103287 9911
rect 103805 9877 103839 9911
rect 104633 9877 104667 9911
rect 106013 9877 106047 9911
rect 116041 9877 116075 9911
rect 120825 9877 120859 9911
rect 124505 9877 124539 9911
rect 126253 9877 126287 9911
rect 129933 9877 129967 9911
rect 144193 9877 144227 9911
rect 144561 9877 144595 9911
rect 146677 9877 146711 9911
rect 146953 9877 146987 9911
rect 147137 9877 147171 9911
rect 148149 9877 148183 9911
rect 151093 9877 151127 9911
rect 151553 9877 151587 9911
rect 153669 9877 153703 9911
rect 154865 9877 154899 9911
rect 155877 9877 155911 9911
rect 7113 9673 7147 9707
rect 27629 9673 27663 9707
rect 28549 9673 28583 9707
rect 32321 9673 32355 9707
rect 49801 9673 49835 9707
rect 64245 9673 64279 9707
rect 85129 9673 85163 9707
rect 93317 9673 93351 9707
rect 132141 9673 132175 9707
rect 141065 9673 141099 9707
rect 144009 9673 144043 9707
rect 148241 9673 148275 9707
rect 153025 9673 153059 9707
rect 6101 9605 6135 9639
rect 15301 9605 15335 9639
rect 21373 9605 21407 9639
rect 34713 9605 34747 9639
rect 37933 9605 37967 9639
rect 41245 9605 41279 9639
rect 48053 9605 48087 9639
rect 48513 9605 48547 9639
rect 54677 9605 54711 9639
rect 57253 9605 57287 9639
rect 60657 9605 60691 9639
rect 63233 9605 63267 9639
rect 70225 9605 70259 9639
rect 70869 9605 70903 9639
rect 71237 9605 71271 9639
rect 72341 9605 72375 9639
rect 79701 9605 79735 9639
rect 101597 9605 101631 9639
rect 111165 9605 111199 9639
rect 112821 9605 112855 9639
rect 113373 9605 113407 9639
rect 126897 9605 126931 9639
rect 127817 9605 127851 9639
rect 133153 9605 133187 9639
rect 135177 9605 135211 9639
rect 137753 9605 137787 9639
rect 139225 9605 139259 9639
rect 151829 9605 151863 9639
rect 160017 9605 160051 9639
rect 162133 9605 162167 9639
rect 18797 9537 18831 9571
rect 19809 9537 19843 9571
rect 20545 9537 20579 9571
rect 24869 9537 24903 9571
rect 24961 9537 24995 9571
rect 25329 9537 25363 9571
rect 26433 9537 26467 9571
rect 26893 9537 26927 9571
rect 27261 9537 27295 9571
rect 30757 9537 30791 9571
rect 31493 9537 31527 9571
rect 36369 9537 36403 9571
rect 36829 9537 36863 9571
rect 38577 9537 38611 9571
rect 40417 9537 40451 9571
rect 40877 9537 40911 9571
rect 41889 9537 41923 9571
rect 42073 9537 42107 9571
rect 42441 9537 42475 9571
rect 46581 9537 46615 9571
rect 47133 9537 47167 9571
rect 51089 9537 51123 9571
rect 51733 9537 51767 9571
rect 53297 9537 53331 9571
rect 54033 9537 54067 9571
rect 54125 9537 54159 9571
rect 55137 9537 55171 9571
rect 55505 9537 55539 9571
rect 57805 9537 57839 9571
rect 58265 9537 58299 9571
rect 58633 9537 58667 9571
rect 59369 9537 59403 9571
rect 59829 9537 59863 9571
rect 62221 9537 62255 9571
rect 69213 9537 69247 9571
rect 74365 9537 74399 9571
rect 74733 9537 74767 9571
rect 76389 9537 76423 9571
rect 80713 9537 80747 9571
rect 81909 9537 81943 9571
rect 82921 9537 82955 9571
rect 86601 9537 86635 9571
rect 88165 9537 88199 9571
rect 91477 9537 91511 9571
rect 92765 9537 92799 9571
rect 97917 9537 97951 9571
rect 100401 9537 100435 9571
rect 104725 9537 104759 9571
rect 109601 9537 109635 9571
rect 112545 9537 112579 9571
rect 115213 9537 115247 9571
rect 120457 9537 120491 9571
rect 121469 9537 121503 9571
rect 123033 9537 123067 9571
rect 125977 9537 126011 9571
rect 126805 9537 126839 9571
rect 131129 9537 131163 9571
rect 131589 9537 131623 9571
rect 143181 9537 143215 9571
rect 147965 9537 147999 9571
rect 148793 9537 148827 9571
rect 150173 9537 150207 9571
rect 150633 9537 150667 9571
rect 154313 9537 154347 9571
rect 155877 9537 155911 9571
rect 159189 9537 159223 9571
rect 164341 9537 164375 9571
rect 165077 9537 165111 9571
rect 165629 9537 165663 9571
rect 166917 9537 166951 9571
rect 3985 9469 4019 9503
rect 15577 9469 15611 9503
rect 17785 9469 17819 9503
rect 20821 9469 20855 9503
rect 22937 9469 22971 9503
rect 51089 9401 51123 9435
rect 74549 9469 74583 9503
rect 80805 9469 80839 9503
rect 87613 9469 87647 9503
rect 88993 9469 89027 9503
rect 89913 9469 89947 9503
rect 90281 9469 90315 9503
rect 92489 9469 92523 9503
rect 93869 9469 93903 9503
rect 96445 9469 96479 9503
rect 97457 9469 97491 9503
rect 98837 9469 98871 9503
rect 99849 9469 99883 9503
rect 103161 9469 103195 9503
rect 104173 9469 104207 9503
rect 108129 9469 108163 9503
rect 109141 9469 109175 9503
rect 54953 9401 54987 9435
rect 83013 9401 83047 9435
rect 114017 9469 114051 9503
rect 115949 9469 115983 9503
rect 116409 9469 116443 9503
rect 118893 9469 118927 9503
rect 119905 9469 119939 9503
rect 122481 9469 122515 9503
rect 124413 9469 124447 9503
rect 125425 9469 125459 9503
rect 129381 9469 129415 9503
rect 129749 9469 129783 9503
rect 130761 9469 130795 9503
rect 141617 9469 141651 9503
rect 143089 9469 143123 9503
rect 145021 9469 145055 9503
rect 146401 9469 146435 9503
rect 147873 9469 147907 9503
rect 148701 9469 148735 9503
rect 152013 9469 152047 9503
rect 155693 9469 155727 9503
rect 157625 9469 157659 9503
rect 158729 9469 158763 9503
rect 160569 9469 160603 9503
rect 161029 9469 161063 9503
rect 163237 9469 163271 9503
rect 164249 9469 164283 9503
rect 166641 9469 166675 9503
rect 115305 9401 115339 9435
rect 150265 9401 150299 9435
rect 4537 9333 4571 9367
rect 6561 9333 6595 9367
rect 19901 9333 19935 9367
rect 21833 9333 21867 9367
rect 26065 9333 26099 9367
rect 26249 9333 26283 9367
rect 30849 9333 30883 9367
rect 39037 9333 39071 9367
rect 40233 9333 40267 9367
rect 42809 9333 42843 9367
rect 46581 9333 46615 9367
rect 53389 9333 53423 9367
rect 54125 9333 54159 9367
rect 54401 9333 54435 9367
rect 56793 9333 56827 9367
rect 57621 9333 57655 9367
rect 59185 9333 59219 9367
rect 76481 9333 76515 9367
rect 82001 9333 82035 9367
rect 88533 9333 88567 9367
rect 94329 9333 94363 9367
rect 112545 9333 112579 9367
rect 121285 9333 121319 9367
rect 127541 9333 127575 9367
rect 156245 9333 156279 9367
rect 157257 9333 157291 9367
rect 159557 9333 159591 9367
rect 3893 9129 3927 9163
rect 17509 9129 17543 9163
rect 19901 9129 19935 9163
rect 20269 9129 20303 9163
rect 21281 9129 21315 9163
rect 23581 9129 23615 9163
rect 24869 9129 24903 9163
rect 25329 9129 25363 9163
rect 25881 9129 25915 9163
rect 28273 9129 28307 9163
rect 28549 9129 28583 9163
rect 30941 9129 30975 9163
rect 39221 9129 39255 9163
rect 42441 9129 42475 9163
rect 43729 9129 43763 9163
rect 51917 9129 51951 9163
rect 52193 9129 52227 9163
rect 55873 9129 55907 9163
rect 57897 9129 57931 9163
rect 58633 9129 58667 9163
rect 59277 9129 59311 9163
rect 59921 9129 59955 9163
rect 74365 9129 74399 9163
rect 75377 9129 75411 9163
rect 76849 9129 76883 9163
rect 80713 9129 80747 9163
rect 83197 9129 83231 9163
rect 86969 9129 87003 9163
rect 92121 9129 92155 9163
rect 96813 9129 96847 9163
rect 98193 9129 98227 9163
rect 108221 9129 108255 9163
rect 108313 9129 108347 9163
rect 121009 9129 121043 9163
rect 124597 9129 124631 9163
rect 127081 9129 127115 9163
rect 145941 9129 145975 9163
rect 154405 9129 154439 9163
rect 157165 9129 157199 9163
rect 165813 9129 165847 9163
rect 18521 9061 18555 9095
rect 18797 9061 18831 9095
rect 3985 8993 4019 9027
rect 4997 8993 5031 9027
rect 6377 8993 6411 9027
rect 7389 8993 7423 9027
rect 16313 8993 16347 9027
rect 22845 8993 22879 9027
rect 23581 8993 23615 9027
rect 24225 8993 24259 9027
rect 31677 9061 31711 9095
rect 47133 9061 47167 9095
rect 29009 8993 29043 9027
rect 34989 8993 35023 9027
rect 36829 8993 36863 9027
rect 37013 8993 37047 9027
rect 40417 8993 40451 9027
rect 41889 8993 41923 9027
rect 46397 8993 46431 9027
rect 47501 8993 47535 9027
rect 50077 8993 50111 9027
rect 54125 9061 54159 9095
rect 55045 9061 55079 9095
rect 63233 9061 63267 9095
rect 82461 9061 82495 9095
rect 52653 8993 52687 9027
rect 53573 8993 53607 9027
rect 55597 8993 55631 9027
rect 57345 8993 57379 9027
rect 58633 8993 58667 9027
rect 58909 8993 58943 9027
rect 64153 8993 64187 9027
rect 71881 8993 71915 9027
rect 72893 8993 72927 9027
rect 73905 8993 73939 9027
rect 74917 8993 74951 9027
rect 76297 8993 76331 9027
rect 80069 8993 80103 9027
rect 82829 8993 82863 9027
rect 85405 8993 85439 9027
rect 88533 8993 88567 9027
rect 90925 8993 90959 9027
rect 93133 8993 93167 9027
rect 95341 8993 95375 9027
rect 97825 8993 97859 9027
rect 99757 8993 99791 9027
rect 104357 8993 104391 9027
rect 107853 8993 107887 9027
rect 108221 8993 108255 9027
rect 109325 9061 109359 9095
rect 5089 8925 5123 8959
rect 7941 8925 7975 8959
rect 15301 8925 15335 8959
rect 16865 8925 16899 8959
rect 17693 8925 17727 8959
rect 18061 8925 18095 8959
rect 18429 8925 18463 8959
rect 18521 8925 18555 8959
rect 20177 8925 20211 8959
rect 20913 8925 20947 8959
rect 21005 8925 21039 8959
rect 21833 8925 21867 8959
rect 23397 8925 23431 8959
rect 26065 8925 26099 8959
rect 26525 8925 26559 8959
rect 27721 8925 27755 8959
rect 27813 8925 27847 8959
rect 28181 8925 28215 8959
rect 28273 8925 28307 8959
rect 38117 8925 38151 8959
rect 38761 8925 38795 8959
rect 39957 8925 39991 8959
rect 40325 8925 40359 8959
rect 40785 8925 40819 8959
rect 41153 8925 41187 8959
rect 42809 8925 42843 8959
rect 42993 8925 43027 8959
rect 43361 8925 43395 8959
rect 50813 8925 50847 8959
rect 50997 8925 51031 8959
rect 51365 8925 51399 8959
rect 51457 8925 51491 8959
rect 51825 8925 51859 8959
rect 51917 8925 51951 8959
rect 52561 8925 52595 8959
rect 54309 8925 54343 8959
rect 54769 8925 54803 8959
rect 56241 8925 56275 8959
rect 56609 8925 56643 8959
rect 56977 8925 57011 8959
rect 58081 8925 58115 8959
rect 58357 8925 58391 8959
rect 63049 8925 63083 8959
rect 63417 8925 63451 8959
rect 63693 8925 63727 8959
rect 81909 8925 81943 8959
rect 87521 8925 87555 8959
rect 89085 8925 89119 8959
rect 89913 8925 89947 8959
rect 91477 8925 91511 8959
rect 94329 8925 94363 8959
rect 95893 8925 95927 8959
rect 96721 8925 96755 8959
rect 98561 8925 98595 8959
rect 98745 8925 98779 8959
rect 100309 8925 100343 8959
rect 8309 8857 8343 8891
rect 26893 8857 26927 8891
rect 57713 8857 57747 8891
rect 61485 8857 61519 8891
rect 82001 8857 82035 8891
rect 86417 8857 86451 8891
rect 87245 8857 87279 8891
rect 101137 8857 101171 8891
rect 103345 8857 103379 8891
rect 122941 9061 122975 9095
rect 123217 9061 123251 9095
rect 147965 9061 147999 9095
rect 150817 9061 150851 9095
rect 163513 9061 163547 9095
rect 112269 8993 112303 9027
rect 113925 8993 113959 9027
rect 114385 8993 114419 9027
rect 115581 8993 115615 9027
rect 116593 8993 116627 9027
rect 122297 8993 122331 9027
rect 124137 8993 124171 9027
rect 127541 8993 127575 9027
rect 128553 8993 128587 9027
rect 129473 8993 129507 9027
rect 131129 8993 131163 9027
rect 138029 8993 138063 9027
rect 139041 8993 139075 9027
rect 142537 8993 142571 9027
rect 144653 8993 144687 9027
rect 148793 8993 148827 9027
rect 149345 8993 149379 9027
rect 151737 8993 151771 9027
rect 153117 8993 153151 9027
rect 156061 8993 156095 9027
rect 158637 8993 158671 9027
rect 160477 8993 160511 9027
rect 161489 8993 161523 9027
rect 163605 8993 163639 9027
rect 164617 8993 164651 9027
rect 117145 8925 117179 8959
rect 118801 8925 118835 8959
rect 119261 8925 119295 8959
rect 121285 8925 121319 8959
rect 122573 8925 122607 8959
rect 122941 8925 122975 8959
rect 129105 8925 129139 8959
rect 129933 8925 129967 8959
rect 131405 8925 131439 8959
rect 131773 8925 131807 8959
rect 140053 8925 140087 8959
rect 141065 8925 141099 8959
rect 142353 8925 142387 8959
rect 143365 8925 143399 8959
rect 146493 8925 146527 8959
rect 148057 8925 148091 8959
rect 150909 8925 150943 8959
rect 153301 8925 153335 8959
rect 154865 8925 154899 8959
rect 155969 8925 156003 8959
rect 156705 8925 156739 8959
rect 157257 8925 157291 8959
rect 158545 8925 158579 8959
rect 162041 8925 162075 8959
rect 164709 8925 164743 8959
rect 165445 8925 165479 8959
rect 142997 8857 143031 8891
rect 163145 8857 163179 8891
rect 166089 8857 166123 8891
rect 5825 8789 5859 8823
rect 17233 8789 17267 8823
rect 19533 8789 19567 8823
rect 21005 8789 21039 8823
rect 21649 8789 21683 8823
rect 23765 8789 23799 8823
rect 27261 8789 27295 8823
rect 33977 8789 34011 8823
rect 41521 8789 41555 8823
rect 48421 8789 48455 8823
rect 50537 8789 50571 8823
rect 50813 8789 50847 8823
rect 59461 8789 59495 8823
rect 60473 8789 60507 8823
rect 89453 8789 89487 8823
rect 91845 8789 91879 8823
rect 92765 8789 92799 8823
rect 96261 8789 96295 8823
rect 96629 8789 96663 8823
rect 97273 8789 97307 8823
rect 100585 8789 100619 8823
rect 101045 8789 101079 8823
rect 102885 8789 102919 8823
rect 104909 8789 104943 8823
rect 106473 8789 106507 8823
rect 109325 8789 109359 8823
rect 109509 8789 109543 8823
rect 115305 8789 115339 8823
rect 117513 8789 117547 8823
rect 120273 8789 120307 8823
rect 123585 8789 123619 8823
rect 125425 8789 125459 8823
rect 125977 8789 126011 8823
rect 129749 8789 129783 8823
rect 140881 8789 140915 8823
rect 143641 8789 143675 8823
rect 146309 8789 146343 8823
rect 148425 8789 148459 8823
rect 151277 8789 151311 8823
rect 153669 8789 153703 8823
rect 153945 8789 153979 8823
rect 159189 8789 159223 8823
rect 162317 8789 162351 8823
rect 166917 8789 166951 8823
rect 5549 8585 5583 8619
rect 6377 8585 6411 8619
rect 27445 8585 27479 8619
rect 41521 8585 41555 8619
rect 50997 8585 51031 8619
rect 51641 8585 51675 8619
rect 57989 8585 58023 8619
rect 59461 8585 59495 8619
rect 65257 8585 65291 8619
rect 73445 8585 73479 8619
rect 74457 8585 74491 8619
rect 80161 8585 80195 8619
rect 90005 8585 90039 8619
rect 94789 8585 94823 8619
rect 98377 8585 98411 8619
rect 113281 8585 113315 8619
rect 122297 8585 122331 8619
rect 124689 8585 124723 8619
rect 128093 8585 128127 8619
rect 139685 8585 139719 8619
rect 142169 8585 142203 8619
rect 145297 8585 145331 8619
rect 157625 8585 157659 8619
rect 18705 8517 18739 8551
rect 37749 8517 37783 8551
rect 42533 8517 42567 8551
rect 49617 8517 49651 8551
rect 57713 8517 57747 8551
rect 85681 8517 85715 8551
rect 98101 8517 98135 8551
rect 101505 8517 101539 8551
rect 5181 8449 5215 8483
rect 14841 8449 14875 8483
rect 15853 8449 15887 8483
rect 16405 8449 16439 8483
rect 17325 8449 17359 8483
rect 17877 8449 17911 8483
rect 19809 8449 19843 8483
rect 20269 8449 20303 8483
rect 21097 8449 21131 8483
rect 21833 8449 21867 8483
rect 23121 8449 23155 8483
rect 23673 8449 23707 8483
rect 25053 8449 25087 8483
rect 25237 8449 25271 8483
rect 25605 8449 25639 8483
rect 34805 8449 34839 8483
rect 35173 8449 35207 8483
rect 35541 8449 35575 8483
rect 36737 8449 36771 8483
rect 37381 8449 37415 8483
rect 37473 8449 37507 8483
rect 38669 8449 38703 8483
rect 39773 8449 39807 8483
rect 40141 8449 40175 8483
rect 40509 8449 40543 8483
rect 48881 8449 48915 8483
rect 49341 8449 49375 8483
rect 52285 8449 52319 8483
rect 52745 8449 52779 8483
rect 55137 8449 55171 8483
rect 55597 8449 55631 8483
rect 56609 8449 56643 8483
rect 57345 8449 57379 8483
rect 58633 8449 58667 8483
rect 59001 8449 59035 8483
rect 60197 8449 60231 8483
rect 60289 8449 60323 8483
rect 60473 8449 60507 8483
rect 64429 8449 64463 8483
rect 83473 8449 83507 8483
rect 89269 8449 89303 8483
rect 91661 8449 91695 8483
rect 92857 8449 92891 8483
rect 94421 8449 94455 8483
rect 97641 8449 97675 8483
rect 3617 8381 3651 8415
rect 4629 8381 4663 8415
rect 13277 8381 13311 8415
rect 14289 8381 14323 8415
rect 16037 8381 16071 8415
rect 20913 8381 20947 8415
rect 21465 8381 21499 8415
rect 26433 8381 26467 8415
rect 37013 8381 37047 8415
rect 46673 8381 46707 8415
rect 53573 8381 53607 8415
rect 55873 8381 55907 8415
rect 58725 8381 58759 8415
rect 62865 8381 62899 8415
rect 63877 8381 63911 8415
rect 71789 8381 71823 8415
rect 79057 8381 79091 8415
rect 82001 8381 82035 8415
rect 83013 8381 83047 8415
rect 86693 8381 86727 8415
rect 87705 8381 87739 8415
rect 90281 8381 90315 8415
rect 91293 8381 91327 8415
rect 93869 8381 93903 8415
rect 96077 8381 96111 8415
rect 98469 8449 98503 8483
rect 100033 8449 100067 8483
rect 103069 8449 103103 8483
rect 104633 8449 104667 8483
rect 107117 8449 107151 8483
rect 108497 8449 108531 8483
rect 99481 8381 99515 8415
rect 104081 8381 104115 8415
rect 108129 8381 108163 8415
rect 114385 8449 114419 8483
rect 121377 8449 121411 8483
rect 125701 8449 125735 8483
rect 126805 8449 126839 8483
rect 131037 8449 131071 8483
rect 142353 8449 142387 8483
rect 143917 8449 143951 8483
rect 146396 8449 146430 8483
rect 147781 8449 147815 8483
rect 148241 8449 148275 8483
rect 150817 8449 150851 8483
rect 152381 8449 152415 8483
rect 153945 8449 153979 8483
rect 154773 8449 154807 8483
rect 156061 8449 156095 8483
rect 156613 8449 156647 8483
rect 160753 8449 160787 8483
rect 165629 8449 165663 8483
rect 113373 8381 113407 8415
rect 115949 8381 115983 8415
rect 116409 8381 116443 8415
rect 119905 8381 119939 8415
rect 120917 8381 120951 8415
rect 126713 8381 126747 8415
rect 129565 8381 129599 8415
rect 130577 8381 130611 8415
rect 132693 8381 132727 8415
rect 141341 8381 141375 8415
rect 141801 8381 141835 8415
rect 143549 8381 143583 8415
rect 147413 8381 147447 8415
rect 149253 8381 149287 8415
rect 150541 8381 150575 8415
rect 153393 8381 153427 8415
rect 155969 8381 156003 8415
rect 159465 8381 159499 8415
rect 160477 8381 160511 8415
rect 161397 8381 161431 8415
rect 161857 8381 161891 8415
rect 163513 8381 163547 8415
rect 164525 8381 164559 8415
rect 17417 8313 17451 8347
rect 19625 8313 19659 8347
rect 20637 8313 20671 8347
rect 22109 8313 22143 8347
rect 23029 8313 23063 8347
rect 23949 8313 23983 8347
rect 37473 8313 37507 8347
rect 48697 8313 48731 8347
rect 52101 8313 52135 8347
rect 54953 8313 54987 8347
rect 56701 8313 56735 8347
rect 88993 8313 89027 8347
rect 95617 8313 95651 8347
rect 97365 8313 97399 8347
rect 98101 8313 98135 8347
rect 100309 8313 100343 8347
rect 113281 8313 113315 8347
rect 154313 8313 154347 8347
rect 158545 8313 158579 8347
rect 165813 8313 165847 8347
rect 25973 8245 26007 8279
rect 45753 8245 45787 8279
rect 54401 8245 54435 8279
rect 61025 8245 61059 8279
rect 79517 8245 79551 8279
rect 83841 8245 83875 8279
rect 87521 8245 87555 8279
rect 98009 8245 98043 8279
rect 112269 8245 112303 8279
rect 133153 8245 133187 8279
rect 145021 8245 145055 8279
rect 151185 8245 151219 8279
rect 15853 8041 15887 8075
rect 16681 8041 16715 8075
rect 18061 8041 18095 8075
rect 18337 8041 18371 8075
rect 20545 8041 20579 8075
rect 21833 8041 21867 8075
rect 23949 8041 23983 8075
rect 25145 8041 25179 8075
rect 25605 8041 25639 8075
rect 26617 8041 26651 8075
rect 26893 8041 26927 8075
rect 34805 8041 34839 8075
rect 35541 8041 35575 8075
rect 39405 8041 39439 8075
rect 39497 8041 39531 8075
rect 39957 8041 39991 8075
rect 49985 8041 50019 8075
rect 52745 8041 52779 8075
rect 53021 8041 53055 8075
rect 55689 8041 55723 8075
rect 59001 8041 59035 8075
rect 60197 8041 60231 8075
rect 60565 8041 60599 8075
rect 63141 8041 63175 8075
rect 63233 8041 63267 8075
rect 71697 8041 71731 8075
rect 87245 8041 87279 8075
rect 92673 8041 92707 8075
rect 103069 8041 103103 8075
rect 107117 8041 107151 8075
rect 108497 8041 108531 8075
rect 125977 8041 126011 8075
rect 129565 8041 129599 8075
rect 147229 8041 147263 8075
rect 152473 8041 152507 8075
rect 155233 8041 155267 8075
rect 166181 8041 166215 8075
rect 2789 7973 2823 8007
rect 25881 7973 25915 8007
rect 4629 7905 4663 7939
rect 6009 7905 6043 7939
rect 15117 7905 15151 7939
rect 16129 7905 16163 7939
rect 19625 7905 19659 7939
rect 23121 7905 23155 7939
rect 27353 7905 27387 7939
rect 38117 7905 38151 7939
rect 39037 7905 39071 7939
rect 41245 7973 41279 8007
rect 49341 7973 49375 8007
rect 49617 7973 49651 8007
rect 59277 7973 59311 8007
rect 42625 7905 42659 7939
rect 45753 7905 45787 7939
rect 46765 7905 46799 7939
rect 3617 7837 3651 7871
rect 5181 7837 5215 7871
rect 14841 7837 14875 7871
rect 18613 7837 18647 7871
rect 18889 7837 18923 7871
rect 19257 7837 19291 7871
rect 20453 7837 20487 7871
rect 21189 7837 21223 7871
rect 22109 7837 22143 7871
rect 23673 7837 23707 7871
rect 25789 7837 25823 7871
rect 26525 7837 26559 7871
rect 26617 7837 26651 7871
rect 35909 7837 35943 7871
rect 36737 7837 36771 7871
rect 37105 7837 37139 7871
rect 38669 7837 38703 7871
rect 39497 7837 39531 7871
rect 40141 7837 40175 7871
rect 40601 7837 40635 7871
rect 40969 7837 41003 7871
rect 47317 7837 47351 7871
rect 48789 7837 48823 7871
rect 48881 7837 48915 7871
rect 49249 7837 49283 7871
rect 57989 7905 58023 7939
rect 89821 7973 89855 8007
rect 101781 7973 101815 8007
rect 61025 7905 61059 7939
rect 62129 7905 62163 7939
rect 63141 7905 63175 7939
rect 63417 7905 63451 7939
rect 64061 7905 64095 7939
rect 71789 7905 71823 7939
rect 72801 7905 72835 7939
rect 79425 7905 79459 7939
rect 80437 7905 80471 7939
rect 81909 7905 81943 7939
rect 82369 7905 82403 7939
rect 83473 7905 83507 7939
rect 84485 7905 84519 7939
rect 86417 7905 86451 7939
rect 87521 7905 87555 7939
rect 88533 7905 88567 7939
rect 89913 7905 89947 7939
rect 91109 7905 91143 7939
rect 50077 7837 50111 7871
rect 51549 7837 51583 7871
rect 51733 7837 51767 7871
rect 52101 7837 52135 7871
rect 54401 7837 54435 7871
rect 54585 7837 54619 7871
rect 54953 7837 54987 7871
rect 55321 7837 55355 7871
rect 56793 7837 56827 7871
rect 56977 7837 57011 7871
rect 58357 7837 58391 7871
rect 59277 7837 59311 7871
rect 62589 7837 62623 7871
rect 62957 7837 62991 7871
rect 73353 7837 73387 7871
rect 80897 7837 80931 7871
rect 81265 7837 81299 7871
rect 84761 7837 84795 7871
rect 85313 7837 85347 7871
rect 89085 7837 89119 7871
rect 91477 7837 91511 7871
rect 100217 7837 100251 7871
rect 17509 7769 17543 7803
rect 24501 7769 24535 7803
rect 34897 7769 34931 7803
rect 36369 7769 36403 7803
rect 39773 7769 39807 7803
rect 49433 7769 49467 7803
rect 55965 7769 55999 7803
rect 64061 7769 64095 7803
rect 64245 7769 64279 7803
rect 91845 7769 91879 7803
rect 99757 7769 99791 7803
rect 2237 7701 2271 7735
rect 3065 7701 3099 7735
rect 5549 7701 5583 7735
rect 8953 7701 8987 7735
rect 13369 7701 13403 7735
rect 13461 7701 13495 7735
rect 19901 7701 19935 7735
rect 41429 7701 41463 7735
rect 47593 7701 47627 7735
rect 56425 7701 56459 7735
rect 59461 7701 59495 7735
rect 68845 7701 68879 7735
rect 73721 7701 73755 7735
rect 83381 7701 83415 7735
rect 89453 7701 89487 7735
rect 99757 7565 99791 7599
rect 45845 7497 45879 7531
rect 83381 7497 83415 7531
rect 18705 7429 18739 7463
rect 20821 7429 20855 7463
rect 34161 7429 34195 7463
rect 37381 7429 37415 7463
rect 42441 7429 42475 7463
rect 48789 7429 48823 7463
rect 49249 7429 49283 7463
rect 50997 7429 51031 7463
rect 51549 7429 51583 7463
rect 52837 7429 52871 7463
rect 53849 7429 53883 7463
rect 54861 7429 54895 7463
rect 60933 7429 60967 7463
rect 90465 7429 90499 7463
rect 91293 7429 91327 7463
rect 91753 7429 91787 7463
rect 5089 7361 5123 7395
rect 9505 7361 9539 7395
rect 9689 7361 9723 7395
rect 14105 7361 14139 7395
rect 15669 7361 15703 7395
rect 17693 7361 17727 7395
rect 19717 7361 19751 7395
rect 20453 7361 20487 7395
rect 20545 7361 20579 7395
rect 21557 7361 21591 7395
rect 22017 7361 22051 7395
rect 22385 7361 22419 7395
rect 25053 7361 25087 7395
rect 36277 7361 36311 7395
rect 36645 7361 36679 7395
rect 3617 7293 3651 7327
rect 4629 7293 4663 7327
rect 5549 7293 5583 7327
rect 7941 7293 7975 7327
rect 8953 7293 8987 7327
rect 13093 7293 13127 7327
rect 15209 7293 15243 7327
rect 16037 7293 16071 7327
rect 20085 7293 20119 7327
rect 9689 7225 9723 7259
rect 23673 7293 23707 7327
rect 24685 7293 24719 7327
rect 26525 7293 26559 7327
rect 37289 7293 37323 7327
rect 21189 7225 21223 7259
rect 36093 7225 36127 7259
rect 37841 7361 37875 7395
rect 38301 7361 38335 7395
rect 41337 7361 41371 7395
rect 42717 7361 42751 7395
rect 46857 7361 46891 7395
rect 47961 7361 47995 7395
rect 56609 7361 56643 7395
rect 57345 7361 57379 7395
rect 59829 7361 59863 7395
rect 68845 7361 68879 7395
rect 70133 7361 70167 7395
rect 81357 7361 81391 7395
rect 89361 7361 89395 7395
rect 38577 7293 38611 7327
rect 39773 7293 39807 7327
rect 40785 7293 40819 7327
rect 41613 7293 41647 7327
rect 42901 7293 42935 7327
rect 44281 7293 44315 7327
rect 48145 7293 48179 7327
rect 58449 7293 58483 7327
rect 59461 7293 59495 7327
rect 69857 7293 69891 7327
rect 79793 7293 79827 7327
rect 80805 7293 80839 7327
rect 86785 7293 86819 7327
rect 87797 7293 87831 7327
rect 89085 7293 89119 7327
rect 89729 7293 89763 7327
rect 56701 7225 56735 7259
rect 9781 7157 9815 7191
rect 20545 7157 20579 7191
rect 21373 7157 21407 7191
rect 23121 7157 23155 7191
rect 33977 7157 34011 7191
rect 37381 7157 37415 7191
rect 37657 7157 37691 7191
rect 42717 7157 42751 7191
rect 44925 7157 44959 7191
rect 52101 7157 52135 7191
rect 57621 7157 57655 7191
rect 58357 7157 58391 7191
rect 60289 7157 60323 7191
rect 81909 7157 81943 7191
rect 14013 6953 14047 6987
rect 23673 6953 23707 6987
rect 26433 6953 26467 6987
rect 38485 6953 38519 6987
rect 39405 6953 39439 6987
rect 46857 6953 46891 6987
rect 51089 6953 51123 6987
rect 57069 6953 57103 6987
rect 57345 6953 57379 6987
rect 58909 6953 58943 6987
rect 68845 6953 68879 6987
rect 70133 6953 70167 6987
rect 80989 6953 81023 6987
rect 5733 6885 5767 6919
rect 10241 6885 10275 6919
rect 22753 6885 22787 6919
rect 37105 6885 37139 6919
rect 41153 6885 41187 6919
rect 42717 6885 42751 6919
rect 79977 6885 80011 6919
rect 3433 6817 3467 6851
rect 3893 6817 3927 6851
rect 6377 6817 6411 6851
rect 7849 6817 7883 6851
rect 8309 6817 8343 6851
rect 8769 6817 8803 6851
rect 8953 6817 8987 6851
rect 13461 6817 13495 6851
rect 14289 6817 14323 6851
rect 14565 6817 14599 6851
rect 15577 6817 15611 6851
rect 19073 6817 19107 6851
rect 19901 6817 19935 6851
rect 20453 6817 20487 6851
rect 21005 6817 21039 6851
rect 23857 6817 23891 6851
rect 26525 6817 26559 6851
rect 27537 6817 27571 6851
rect 33609 6817 33643 6851
rect 34069 6817 34103 6851
rect 34805 6817 34839 6851
rect 37841 6817 37875 6851
rect 4353 6749 4387 6783
rect 4445 6749 4479 6783
rect 6009 6749 6043 6783
rect 10517 6749 10551 6783
rect 16129 6749 16163 6783
rect 18061 6749 18095 6783
rect 21465 6749 21499 6783
rect 22569 6749 22603 6783
rect 23305 6749 23339 6783
rect 27997 6749 28031 6783
rect 33977 6749 34011 6783
rect 34437 6749 34471 6783
rect 36277 6749 36311 6783
rect 37289 6749 37323 6783
rect 37749 6749 37783 6783
rect 16497 6681 16531 6715
rect 33609 6681 33643 6715
rect 35265 6681 35299 6715
rect 36737 6681 36771 6715
rect 45661 6817 45695 6851
rect 39773 6749 39807 6783
rect 39865 6749 39899 6783
rect 41337 6749 41371 6783
rect 42717 6749 42751 6783
rect 43361 6749 43395 6783
rect 43729 6749 43763 6783
rect 44925 6749 44959 6783
rect 45109 6749 45143 6783
rect 45477 6749 45511 6783
rect 51825 6817 51859 6851
rect 52101 6817 52135 6851
rect 54401 6817 54435 6851
rect 56885 6817 56919 6851
rect 57069 6817 57103 6851
rect 59921 6817 59955 6851
rect 60933 6817 60967 6851
rect 79609 6817 79643 6851
rect 45845 6749 45879 6783
rect 48329 6749 48363 6783
rect 49985 6749 50019 6783
rect 51273 6749 51307 6783
rect 51549 6749 51583 6783
rect 45661 6681 45695 6715
rect 55413 6749 55447 6783
rect 57621 6749 57655 6783
rect 57805 6749 57839 6783
rect 58173 6749 58207 6783
rect 58449 6749 58483 6783
rect 61485 6749 61519 6783
rect 61853 6749 61887 6783
rect 51825 6681 51859 6715
rect 80069 6817 80103 6851
rect 79977 6681 80011 6715
rect 83197 6885 83231 6919
rect 87797 6885 87831 6919
rect 81909 6817 81943 6851
rect 88165 6817 88199 6851
rect 88349 6817 88383 6851
rect 89361 6817 89395 6851
rect 91753 6817 91787 6851
rect 83013 6749 83047 6783
rect 83749 6749 83783 6783
rect 89913 6749 89947 6783
rect 80989 6681 81023 6715
rect 90281 6681 90315 6715
rect 10885 6613 10919 6647
rect 21281 6613 21315 6647
rect 25053 6613 25087 6647
rect 28457 6613 28491 6647
rect 37841 6613 37875 6647
rect 38025 6613 38059 6647
rect 38853 6613 38887 6647
rect 41705 6613 41739 6647
rect 46305 6613 46339 6647
rect 48329 6613 48363 6647
rect 48513 6613 48547 6647
rect 56425 6613 56459 6647
rect 59829 6613 59863 6647
rect 65073 6613 65107 6647
rect 69581 6613 69615 6647
rect 81173 6613 81207 6647
rect 4261 6409 4295 6443
rect 21833 6409 21867 6443
rect 36553 6409 36587 6443
rect 39773 6409 39807 6443
rect 53941 6409 53975 6443
rect 56609 6409 56643 6443
rect 56701 6409 56735 6443
rect 60105 6409 60139 6443
rect 81357 6409 81391 6443
rect 87981 6409 88015 6443
rect 95065 6409 95099 6443
rect 37565 6341 37599 6375
rect 55505 6341 55539 6375
rect 9045 6273 9079 6307
rect 21097 6273 21131 6307
rect 24041 6273 24075 6307
rect 26065 6273 26099 6307
rect 26157 6273 26191 6307
rect 26525 6273 26559 6307
rect 29837 6273 29871 6307
rect 30297 6273 30331 6307
rect 35725 6273 35759 6307
rect 41705 6273 41739 6307
rect 43269 6273 43303 6307
rect 47225 6273 47259 6307
rect 51273 6273 51307 6307
rect 52653 6273 52687 6307
rect 3249 6205 3283 6239
rect 5917 6205 5951 6239
rect 6101 6205 6135 6239
rect 7481 6205 7515 6239
rect 8585 6205 8619 6239
rect 9873 6205 9907 6239
rect 10425 6205 10459 6239
rect 16037 6205 16071 6239
rect 19533 6205 19567 6239
rect 20545 6205 20579 6239
rect 23397 6205 23431 6239
rect 27353 6205 27387 6239
rect 34161 6205 34195 6239
rect 35173 6205 35207 6239
rect 42717 6205 42751 6239
rect 45661 6205 45695 6239
rect 46673 6205 46707 6239
rect 52285 6205 52319 6239
rect 57713 6273 57747 6307
rect 59277 6273 59311 6307
rect 64521 6273 64555 6307
rect 66085 6273 66119 6307
rect 69949 6273 69983 6307
rect 71513 6273 71547 6307
rect 91845 6273 91879 6307
rect 65533 6205 65567 6239
rect 70961 6205 70995 6239
rect 81265 6205 81299 6239
rect 86509 6205 86543 6239
rect 87521 6205 87555 6239
rect 88993 6205 89027 6239
rect 90281 6205 90315 6239
rect 91293 6205 91327 6239
rect 56609 6137 56643 6171
rect 59001 6137 59035 6171
rect 3709 6069 3743 6103
rect 21373 6069 21407 6103
rect 36093 6069 36127 6103
rect 81265 6069 81299 6103
rect 9229 5865 9263 5899
rect 12357 5865 12391 5899
rect 15945 5865 15979 5899
rect 19533 5865 19567 5899
rect 20913 5865 20947 5899
rect 23397 5865 23431 5899
rect 25605 5865 25639 5899
rect 30297 5865 30331 5899
rect 31125 5865 31159 5899
rect 11897 5797 11931 5831
rect 26893 5797 26927 5831
rect 2237 5729 2271 5763
rect 3433 5729 3467 5763
rect 4445 5729 4479 5763
rect 5825 5729 5859 5763
rect 6929 5729 6963 5763
rect 7757 5729 7791 5763
rect 10425 5729 10459 5763
rect 16037 5729 16071 5763
rect 17049 5729 17083 5763
rect 19073 5729 19107 5763
rect 21097 5729 21131 5763
rect 22109 5729 22143 5763
rect 4997 5661 5031 5695
rect 7389 5661 7423 5695
rect 11989 5661 12023 5695
rect 17601 5661 17635 5695
rect 17969 5661 18003 5695
rect 22661 5661 22695 5695
rect 22753 5661 22787 5695
rect 24041 5661 24075 5695
rect 24501 5661 24535 5695
rect 26433 5661 26467 5695
rect 5365 5593 5399 5627
rect 33425 5865 33459 5899
rect 33701 5865 33735 5899
rect 46213 5865 46247 5899
rect 46397 5865 46431 5899
rect 50445 5865 50479 5899
rect 50721 5865 50755 5899
rect 56885 5865 56919 5899
rect 57437 5865 57471 5899
rect 57897 5865 57931 5899
rect 58449 5865 58483 5899
rect 58725 5865 58759 5899
rect 64521 5865 64555 5899
rect 69949 5865 69983 5899
rect 90281 5865 90315 5899
rect 42993 5797 43027 5831
rect 33149 5729 33183 5763
rect 33425 5729 33459 5763
rect 35173 5729 35207 5763
rect 37013 5729 37047 5763
rect 41521 5729 41555 5763
rect 41981 5729 42015 5763
rect 49893 5797 49927 5831
rect 51181 5729 51215 5763
rect 51641 5729 51675 5763
rect 52653 5729 52687 5763
rect 54493 5729 54527 5763
rect 55321 5729 55355 5763
rect 56057 5729 56091 5763
rect 34069 5661 34103 5695
rect 34161 5661 34195 5695
rect 35633 5661 35667 5695
rect 45937 5661 45971 5695
rect 46213 5661 46247 5695
rect 50261 5661 50295 5695
rect 50445 5661 50479 5695
rect 55137 5661 55171 5695
rect 56701 5661 56735 5695
rect 23489 5593 23523 5627
rect 25789 5593 25823 5627
rect 31125 5593 31159 5627
rect 36093 5593 36127 5627
rect 45293 5593 45327 5627
rect 55321 5593 55355 5627
rect 89453 5797 89487 5831
rect 95065 5797 95099 5831
rect 58449 5729 58483 5763
rect 87521 5729 87555 5763
rect 88717 5729 88751 5763
rect 94973 5729 95007 5763
rect 57161 5661 57195 5695
rect 57713 5661 57747 5695
rect 89085 5661 89119 5695
rect 91753 5593 91787 5627
rect 8033 5525 8067 5559
rect 22753 5525 22787 5559
rect 23029 5525 23063 5559
rect 47041 5525 47075 5559
rect 55597 5525 55631 5559
rect 56885 5525 56919 5559
rect 59093 5525 59127 5559
rect 65901 5525 65935 5559
rect 71329 5525 71363 5559
rect 90741 5525 90775 5559
rect 91661 5525 91695 5559
rect 93133 5457 93167 5491
rect 7297 5321 7331 5355
rect 45753 5321 45787 5355
rect 18889 5253 18923 5287
rect 20269 5253 20303 5287
rect 26249 5253 26283 5287
rect 89729 5253 89763 5287
rect 93133 5253 93167 5287
rect 3433 5185 3467 5219
rect 4997 5185 5031 5219
rect 5365 5185 5399 5219
rect 16221 5185 16255 5219
rect 18429 5185 18463 5219
rect 21465 5185 21499 5219
rect 24501 5185 24535 5219
rect 34805 5185 34839 5219
rect 46397 5185 46431 5219
rect 47685 5185 47719 5219
rect 48329 5185 48363 5219
rect 49893 5185 49927 5219
rect 54125 5185 54159 5219
rect 57253 5185 57287 5219
rect 89361 5185 89395 5219
rect 90741 5185 90775 5219
rect 91753 5185 91787 5219
rect 4445 5117 4479 5151
rect 15577 5117 15611 5151
rect 21281 5117 21315 5151
rect 22937 5117 22971 5151
rect 23949 5117 23983 5151
rect 25329 5117 25363 5151
rect 46121 5117 46155 5151
rect 49249 5117 49283 5151
rect 53481 5117 53515 5151
rect 86785 5117 86819 5151
rect 87797 5117 87831 5151
rect 89269 5117 89303 5151
rect 90833 5117 90867 5151
rect 24869 5049 24903 5083
rect 90557 5049 90591 5083
rect 18061 4981 18095 5015
rect 34437 4981 34471 5015
rect 56885 4981 56919 5015
rect 91845 4981 91879 5015
rect 3525 4777 3559 4811
rect 16037 4777 16071 4811
rect 17325 4777 17359 4811
rect 21649 4777 21683 4811
rect 22569 4777 22603 4811
rect 22937 4777 22971 4811
rect 26617 4777 26651 4811
rect 26893 4777 26927 4811
rect 49525 4777 49559 4811
rect 49709 4777 49743 4811
rect 53665 4777 53699 4811
rect 54677 4777 54711 4811
rect 54953 4777 54987 4811
rect 88625 4777 88659 4811
rect 91845 4777 91879 4811
rect 4997 4641 5031 4675
rect 21005 4641 21039 4675
rect 22017 4641 22051 4675
rect 23029 4641 23063 4675
rect 24041 4641 24075 4675
rect 25789 4641 25823 4675
rect 30573 4709 30607 4743
rect 33149 4709 33183 4743
rect 3985 4573 4019 4607
rect 5549 4573 5583 4607
rect 16865 4573 16899 4607
rect 17969 4573 18003 4607
rect 18797 4573 18831 4607
rect 24593 4573 24627 4607
rect 26341 4573 26375 4607
rect 26617 4573 26651 4607
rect 30113 4573 30147 4607
rect 32965 4573 32999 4607
rect 33241 4709 33275 4743
rect 33425 4709 33459 4743
rect 34621 4709 34655 4743
rect 39773 4641 39807 4675
rect 46581 4641 46615 4675
rect 47869 4641 47903 4675
rect 33241 4573 33275 4607
rect 40233 4573 40267 4607
rect 40785 4573 40819 4607
rect 5917 4505 5951 4539
rect 29469 4505 29503 4539
rect 32321 4505 32355 4539
rect 33149 4505 33183 4539
rect 48881 4573 48915 4607
rect 49065 4573 49099 4607
rect 47869 4505 47903 4539
rect 48053 4505 48087 4539
rect 48237 4505 48271 4539
rect 94973 5525 95007 5559
rect 99021 5525 99055 5559
rect 99297 5457 99331 5491
rect 99389 5457 99423 5491
rect 94973 5049 95007 5083
rect 55965 4709 55999 4743
rect 56793 4709 56827 4743
rect 57161 4709 57195 4743
rect 90281 4709 90315 4743
rect 92673 4709 92707 4743
rect 94881 4709 94915 4743
rect 87797 4641 87831 4675
rect 88257 4641 88291 4675
rect 88809 4641 88843 4675
rect 53849 4573 53883 4607
rect 54493 4573 54527 4607
rect 54677 4573 54711 4607
rect 55781 4573 55815 4607
rect 90373 4573 90407 4607
rect 91753 4573 91787 4607
rect 101781 7769 101815 7803
rect 101873 7973 101907 8007
rect 148885 7973 148919 8007
rect 156797 7973 156831 8007
rect 164801 7973 164835 8007
rect 102977 7905 103011 7939
rect 103345 7905 103379 7939
rect 110429 7905 110463 7939
rect 112269 7905 112303 7939
rect 113281 7905 113315 7939
rect 117329 7905 117363 7939
rect 119997 7905 120031 7939
rect 120457 7905 120491 7939
rect 125517 7905 125551 7939
rect 127449 7905 127483 7939
rect 128737 7905 128771 7939
rect 129749 7905 129783 7939
rect 130761 7905 130795 7939
rect 133061 7905 133095 7939
rect 134073 7905 134107 7939
rect 140697 7905 140731 7939
rect 141801 7905 141835 7939
rect 142813 7905 142847 7939
rect 145021 7905 145055 7939
rect 146033 7905 146067 7939
rect 147413 7905 147447 7939
rect 150909 7905 150943 7939
rect 154037 7905 154071 7939
rect 159373 7905 159407 7939
rect 161121 7905 161155 7939
rect 162133 7905 162167 7939
rect 166733 7905 166767 7939
rect 113833 7837 113867 7871
rect 113925 7837 113959 7871
rect 116317 7837 116351 7871
rect 117881 7837 117915 7871
rect 118157 7837 118191 7871
rect 134257 7837 134291 7871
rect 134901 7837 134935 7871
rect 143365 7837 143399 7871
rect 146401 7837 146435 7871
rect 146861 7837 146895 7871
rect 148977 7837 149011 7871
rect 149713 7837 149747 7871
rect 149897 7837 149931 7871
rect 151001 7837 151035 7871
rect 151737 7837 151771 7871
rect 153025 7837 153059 7871
rect 154589 7837 154623 7871
rect 155509 7837 155543 7871
rect 156981 7837 157015 7871
rect 158269 7837 158303 7871
rect 158361 7837 158395 7871
rect 159741 7837 159775 7871
rect 160201 7837 160235 7871
rect 162225 7837 162259 7871
rect 162961 7837 162995 7871
rect 163513 7837 163547 7871
rect 164617 7837 164651 7871
rect 165353 7837 165387 7871
rect 110429 7769 110463 7803
rect 121285 7769 121319 7803
rect 143733 7769 143767 7803
rect 157441 7769 157475 7803
rect 101873 7701 101907 7735
rect 102333 7701 102367 7735
rect 102977 7701 103011 7735
rect 104449 7701 104483 7735
rect 113925 7701 113959 7735
rect 114201 7701 114235 7735
rect 118985 7701 119019 7735
rect 121837 7701 121871 7735
rect 127081 7701 127115 7735
rect 131221 7701 131255 7735
rect 144101 7701 144135 7735
rect 149345 7701 149379 7735
rect 152933 7701 152967 7735
rect 154957 7701 154991 7735
rect 160753 7701 160787 7735
rect 163421 7701 163455 7735
rect 165813 7701 165847 7735
rect 101413 7633 101447 7667
rect 142445 7497 142479 7531
rect 145205 7497 145239 7531
rect 147045 7497 147079 7531
rect 147505 7497 147539 7531
rect 149897 7497 149931 7531
rect 150449 7497 150483 7531
rect 156153 7497 156187 7531
rect 158729 7497 158763 7531
rect 159465 7497 159499 7531
rect 166273 7497 166307 7531
rect 151461 7429 151495 7463
rect 156705 7429 156739 7463
rect 102609 7361 102643 7395
rect 103989 7361 104023 7395
rect 114937 7361 114971 7395
rect 115305 7361 115339 7395
rect 117145 7361 117179 7395
rect 118985 7361 119019 7395
rect 120549 7361 120583 7395
rect 122941 7361 122975 7395
rect 123217 7361 123251 7395
rect 126897 7361 126931 7395
rect 133337 7361 133371 7395
rect 144377 7361 144411 7395
rect 149345 7361 149379 7395
rect 155877 7361 155911 7395
rect 161029 7361 161063 7395
rect 161765 7361 161799 7395
rect 164985 7361 165019 7395
rect 113373 7293 113407 7327
rect 114385 7293 114419 7327
rect 115765 7293 115799 7327
rect 116777 7293 116811 7327
rect 119997 7293 120031 7327
rect 121377 7293 121411 7327
rect 122389 7293 122423 7327
rect 125425 7293 125459 7327
rect 126437 7293 126471 7327
rect 127541 7293 127575 7327
rect 127817 7293 127851 7327
rect 129933 7293 129967 7327
rect 130209 7293 130243 7327
rect 132233 7293 132267 7327
rect 133429 7293 133463 7327
rect 142813 7293 142847 7327
rect 143825 7293 143859 7327
rect 148057 7293 148091 7327
rect 149529 7293 149563 7327
rect 153301 7293 153335 7327
rect 154313 7293 154347 7327
rect 155325 7293 155359 7327
rect 159925 7293 159959 7327
rect 161121 7293 161155 7327
rect 162777 7293 162811 7327
rect 163881 7293 163915 7327
rect 164893 7293 164927 7327
rect 101413 7225 101447 7259
rect 103897 7225 103931 7259
rect 134901 7157 134935 7191
rect 141801 7157 141835 7191
rect 153025 7157 153059 7191
rect 163513 7157 163547 7191
rect 113373 6953 113407 6987
rect 118985 6953 119019 6987
rect 120457 6953 120491 6987
rect 121377 6953 121411 6987
rect 132233 6953 132267 6987
rect 155233 6953 155267 6987
rect 163329 6953 163363 6987
rect 102793 6885 102827 6919
rect 103989 6885 104023 6919
rect 114753 6885 114787 6919
rect 101505 6817 101539 6851
rect 112177 6817 112211 6851
rect 115397 6817 115431 6851
rect 128737 6885 128771 6919
rect 136189 6885 136223 6919
rect 143089 6885 143123 6919
rect 154313 6885 154347 6919
rect 162409 6885 162443 6919
rect 164801 6885 164835 6919
rect 122849 6817 122883 6851
rect 125425 6817 125459 6851
rect 125885 6817 125919 6851
rect 127449 6817 127483 6851
rect 129841 6817 129875 6851
rect 130853 6817 130887 6851
rect 133061 6817 133095 6851
rect 141801 6817 141835 6851
rect 146033 6817 146067 6851
rect 148149 6817 148183 6851
rect 148609 6817 148643 6851
rect 151829 6817 151863 6851
rect 156521 6817 156555 6851
rect 160017 6817 160051 6851
rect 160477 6817 160511 6851
rect 163513 6817 163547 6851
rect 102333 6749 102367 6783
rect 113465 6749 113499 6783
rect 114661 6749 114695 6783
rect 120089 6749 120123 6783
rect 120457 6749 120491 6783
rect 121101 6749 121135 6783
rect 121837 6749 121871 6783
rect 123401 6749 123435 6783
rect 123493 6749 123527 6783
rect 128553 6749 128587 6783
rect 129289 6749 129323 6783
rect 131129 6749 131163 6783
rect 131681 6749 131715 6783
rect 134901 6749 134935 6783
rect 136005 6749 136039 6783
rect 136741 6749 136775 6783
rect 142905 6749 142939 6783
rect 143641 6749 143675 6783
rect 150541 6749 150575 6783
rect 150633 6749 150667 6783
rect 152105 6749 152139 6783
rect 152473 6749 152507 6783
rect 153025 6749 153059 6783
rect 154129 6749 154163 6783
rect 154865 6749 154899 6783
rect 160937 6749 160971 6783
rect 161121 6749 161155 6783
rect 162501 6749 162535 6783
rect 164617 6749 164651 6783
rect 165721 6749 165755 6783
rect 162961 6681 162995 6715
rect 113005 6613 113039 6647
rect 115765 6613 115799 6647
rect 117145 6613 117179 6647
rect 120641 6613 120675 6647
rect 123493 6613 123527 6647
rect 123769 6613 123803 6647
rect 126805 6613 126839 6647
rect 133521 6613 133555 6647
rect 144561 6613 144595 6647
rect 149345 6613 149379 6647
rect 155509 6613 155543 6647
rect 155969 6613 156003 6647
rect 165353 6613 165387 6647
rect 159741 6409 159775 6443
rect 161489 6409 161523 6443
rect 162501 6409 162535 6443
rect 135821 6341 135855 6375
rect 142169 6341 142203 6375
rect 142813 6341 142847 6375
rect 143181 6341 143215 6375
rect 150817 6341 150851 6375
rect 155785 6341 155819 6375
rect 156797 6341 156831 6375
rect 122481 6273 122515 6307
rect 149989 6273 150023 6307
rect 153117 6273 153151 6307
rect 154865 6273 154899 6307
rect 164985 6273 165019 6307
rect 113373 6205 113407 6239
rect 115213 6205 115247 6239
rect 120917 6205 120951 6239
rect 121929 6205 121963 6239
rect 122941 6205 122975 6239
rect 123309 6205 123343 6239
rect 129105 6205 129139 6239
rect 148425 6205 148459 6239
rect 149437 6205 149471 6239
rect 153393 6205 153427 6239
rect 158269 6205 158303 6239
rect 163881 6205 163915 6239
rect 166273 6205 166307 6239
rect 154681 6137 154715 6171
rect 165169 6137 165203 6171
rect 156337 6069 156371 6103
rect 163605 6069 163639 6103
rect 116317 5865 116351 5899
rect 128921 5865 128955 5899
rect 148425 5865 148459 5899
rect 152933 5865 152967 5899
rect 158269 5865 158303 5899
rect 159281 5865 159315 5899
rect 163513 5865 163547 5899
rect 154497 5797 154531 5831
rect 115213 5729 115247 5763
rect 123861 5729 123895 5763
rect 129013 5729 129047 5763
rect 130025 5729 130059 5763
rect 148793 5729 148827 5763
rect 151001 5729 151035 5763
rect 156797 5729 156831 5763
rect 162593 5729 162627 5763
rect 163605 5729 163639 5763
rect 164709 5729 164743 5763
rect 102333 5661 102367 5695
rect 102609 5661 102643 5695
rect 110889 5661 110923 5695
rect 111165 5661 111199 5695
rect 114661 5661 114695 5695
rect 116225 5661 116259 5695
rect 121009 5661 121043 5695
rect 121837 5661 121871 5695
rect 122849 5661 122883 5695
rect 124413 5661 124447 5695
rect 130577 5661 130611 5695
rect 153025 5661 153059 5695
rect 154589 5661 154623 5695
rect 155785 5661 155819 5695
rect 157349 5661 157383 5695
rect 157625 5661 157659 5695
rect 158177 5661 158211 5695
rect 158637 5661 158671 5695
rect 159189 5661 159223 5695
rect 159649 5661 159683 5695
rect 165077 5661 165111 5695
rect 165445 5661 165479 5695
rect 101505 5593 101539 5627
rect 114753 5593 114787 5627
rect 116777 5593 116811 5627
rect 102425 5525 102459 5559
rect 102609 5525 102643 5559
rect 102885 5525 102919 5559
rect 110981 5525 111015 5559
rect 111165 5525 111199 5559
rect 111441 5525 111475 5559
rect 122389 5525 122423 5559
rect 124781 5525 124815 5559
rect 130945 5525 130979 5559
rect 150081 5525 150115 5559
rect 152013 5525 152047 5559
rect 154865 5525 154899 5559
rect 155325 5525 155359 5559
rect 165813 5525 165847 5559
rect 105921 5321 105955 5355
rect 127817 5321 127851 5355
rect 145849 5321 145883 5355
rect 164709 5321 164743 5355
rect 104633 5185 104667 5219
rect 105829 5185 105863 5219
rect 110245 5185 110279 5219
rect 115305 5185 115339 5219
rect 127725 5185 127759 5219
rect 145757 5185 145791 5219
rect 152933 5185 152967 5219
rect 154497 5185 154531 5219
rect 156613 5185 156647 5219
rect 158269 5185 158303 5219
rect 159557 5185 159591 5219
rect 164617 5185 164651 5219
rect 100217 5117 100251 5151
rect 103069 5117 103103 5151
rect 104081 5117 104115 5151
rect 110337 5117 110371 5151
rect 153945 5117 153979 5151
rect 155325 5117 155359 5151
rect 156521 5117 156555 5151
rect 159281 5117 159315 5151
rect 115397 5049 115431 5083
rect 104449 4777 104483 4811
rect 105737 4777 105771 4811
rect 121929 4777 121963 4811
rect 129197 4777 129231 4811
rect 130209 4777 130243 4811
rect 131221 4777 131255 4811
rect 147321 4777 147355 4811
rect 150173 4777 150207 4811
rect 151737 4777 151771 4811
rect 153393 4777 153427 4811
rect 154037 4777 154071 4811
rect 155877 4777 155911 4811
rect 156613 4777 156647 4811
rect 158269 4777 158303 4811
rect 163237 4777 163271 4811
rect 102885 4641 102919 4675
rect 103345 4641 103379 4675
rect 49525 4505 49559 4539
rect 90833 4505 90867 4539
rect 100033 4505 100067 4539
rect 150633 4641 150667 4675
rect 152933 4641 152967 4675
rect 155233 4641 155267 4675
rect 156797 4641 156831 4675
rect 121837 4573 121871 4607
rect 129105 4573 129139 4607
rect 130117 4573 130151 4607
rect 131129 4573 131163 4607
rect 147221 4573 147255 4607
rect 150081 4573 150115 4607
rect 151645 4573 151679 4607
rect 153945 4573 153979 4607
rect 155785 4573 155819 4607
rect 163145 4573 163179 4607
rect 129657 4505 129691 4539
rect 145849 4505 145883 4539
rect 147781 4505 147815 4539
rect 154497 4505 154531 4539
rect 7205 4437 7239 4471
rect 16681 4437 16715 4471
rect 18061 4437 18095 4471
rect 24961 4437 24995 4471
rect 49065 4437 49099 4471
rect 49249 4437 49283 4471
rect 92305 4437 92339 4471
rect 105737 4437 105771 4471
rect 105921 4437 105955 4471
rect 110245 4437 110279 4471
rect 115397 4437 115431 4471
rect 122389 4437 122423 4471
rect 127817 4437 127851 4471
rect 130669 4437 130703 4471
rect 131681 4437 131715 4471
rect 152197 4437 152231 4471
rect 154865 4437 154899 4471
rect 156337 4437 156371 4471
rect 159557 4437 159591 4471
rect 163605 4437 163639 4471
rect 164709 4437 164743 4471
rect 3525 4233 3559 4267
rect 3985 4233 4019 4267
rect 61209 4233 61243 4267
rect 62313 4233 62347 4267
rect 68477 4233 68511 4267
rect 114845 4233 114879 4267
rect 153485 4233 153519 4267
rect 9597 4165 9631 4199
rect 53665 4165 53699 4199
rect 88165 4165 88199 4199
rect 115949 4165 115983 4199
rect 124689 4165 124723 4199
rect 137937 4165 137971 4199
rect 7665 4097 7699 4131
rect 18889 4097 18923 4131
rect 24041 4097 24075 4131
rect 24685 4097 24719 4131
rect 25145 4097 25179 4131
rect 26249 4097 26283 4131
rect 32689 4097 32723 4131
rect 41705 4097 41739 4131
rect 47961 4097 47995 4131
rect 49617 4097 49651 4131
rect 52653 4097 52687 4131
rect 55321 4097 55355 4131
rect 61117 4097 61151 4131
rect 62221 4097 62255 4131
rect 62773 4097 62807 4131
rect 63233 4097 63267 4131
rect 63325 4097 63359 4131
rect 68385 4097 68419 4131
rect 69949 4097 69983 4131
rect 70041 4097 70075 4131
rect 70961 4097 70995 4131
rect 71053 4097 71087 4131
rect 71973 4097 72007 4131
rect 72065 4097 72099 4131
rect 89177 4097 89211 4131
rect 90281 4097 90315 4131
rect 91753 4097 91787 4131
rect 102333 4097 102367 4131
rect 106565 4097 106599 4131
rect 106657 4097 106691 4131
rect 107761 4097 107795 4131
rect 107853 4097 107887 4131
rect 113749 4097 113783 4131
rect 114753 4097 114787 4131
rect 115857 4097 115891 4131
rect 119537 4097 119571 4131
rect 121561 4097 121595 4131
rect 124597 4097 124631 4131
rect 125609 4097 125643 4131
rect 125701 4097 125735 4131
rect 126897 4097 126931 4131
rect 126989 4097 127023 4131
rect 130209 4097 130243 4131
rect 130301 4097 130335 4131
rect 131313 4097 131347 4131
rect 131405 4097 131439 4131
rect 148149 4097 148183 4131
rect 148241 4097 148275 4131
rect 150081 4097 150115 4131
rect 155049 4097 155083 4131
rect 156061 4097 156095 4131
rect 156153 4097 156187 4131
rect 158453 4097 158487 4131
rect 158545 4097 158579 4131
rect 160201 4097 160235 4131
rect 161213 4097 161247 4131
rect 162225 4097 162259 4131
rect 165537 4097 165571 4131
rect 165629 4097 165663 4131
rect 4537 4029 4571 4063
rect 6101 4029 6135 4063
rect 7113 4029 7147 4063
rect 18245 4029 18279 4063
rect 21097 4029 21131 4063
rect 21189 4029 21223 4063
rect 25605 4029 25639 4063
rect 32321 4029 32355 4063
rect 41061 4029 41095 4063
rect 49249 4029 49283 4063
rect 52009 4029 52043 4063
rect 54677 4029 54711 4063
rect 90373 4029 90407 4063
rect 91845 4029 91879 4063
rect 155141 4029 155175 4063
rect 160293 4029 160327 4063
rect 161305 4029 161339 4063
rect 162317 4029 162351 4063
rect 119629 3961 119663 3995
rect 121653 3961 121687 3995
rect 46029 3893 46063 3927
rect 47961 3893 47995 3927
rect 89269 3893 89303 3927
rect 102425 3893 102459 3927
rect 113833 3893 113867 3927
rect 126437 3893 126471 3927
rect 150173 3893 150207 3927
rect 6653 3689 6687 3723
rect 7205 3689 7239 3723
rect 8033 3689 8067 3723
rect 9413 3689 9447 3723
rect 18705 3689 18739 3723
rect 24225 3689 24259 3723
rect 25053 3689 25087 3723
rect 26157 3689 26191 3723
rect 26341 3689 26375 3723
rect 27997 3689 28031 3723
rect 29377 3689 29411 3723
rect 29653 3689 29687 3723
rect 48053 3689 48087 3723
rect 49525 3689 49559 3723
rect 49617 3689 49651 3723
rect 51089 3689 51123 3723
rect 51733 3689 51767 3723
rect 51825 3689 51859 3723
rect 55413 3689 55447 3723
rect 58265 3689 58299 3723
rect 58449 3689 58483 3723
rect 58725 3689 58759 3723
rect 61301 3689 61335 3723
rect 61853 3689 61887 3723
rect 89177 3689 89211 3723
rect 92673 3689 92707 3723
rect 113833 3689 113867 3723
rect 121929 3689 121963 3723
rect 124965 3689 124999 3723
rect 126437 3689 126471 3723
rect 130853 3689 130887 3723
rect 133521 3689 133555 3723
rect 164249 3689 164283 3723
rect 165537 3689 165571 3723
rect 7389 3621 7423 3655
rect 5733 3553 5767 3587
rect 7573 3553 7607 3587
rect 9597 3553 9631 3587
rect 10609 3553 10643 3587
rect 18245 3553 18279 3587
rect 21925 3553 21959 3587
rect 4721 3485 4755 3519
rect 6285 3485 6319 3519
rect 7113 3485 7147 3519
rect 7389 3485 7423 3519
rect 11161 3485 11195 3519
rect 17785 3485 17819 3519
rect 21097 3485 21131 3519
rect 21189 3485 21223 3519
rect 21557 3485 21591 3519
rect 23029 3485 23063 3519
rect 24593 3485 24627 3519
rect 3709 3417 3743 3451
rect 4537 3417 4571 3451
rect 7021 3417 7055 3451
rect 11529 3417 11563 3451
rect 17141 3417 17175 3451
rect 22385 3417 22419 3451
rect 32689 3621 32723 3655
rect 49065 3621 49099 3655
rect 41521 3553 41555 3587
rect 43361 3553 43395 3587
rect 44465 3553 44499 3587
rect 46857 3553 46891 3587
rect 27537 3485 27571 3519
rect 29193 3485 29227 3519
rect 29377 3485 29411 3519
rect 37013 3485 37047 3519
rect 37473 3485 37507 3519
rect 38025 3485 38059 3519
rect 43913 3485 43947 3519
rect 45661 3485 45695 3519
rect 45845 3485 45879 3519
rect 46121 3485 46155 3519
rect 46489 3485 46523 3519
rect 48881 3485 48915 3519
rect 26893 3417 26927 3451
rect 28549 3417 28583 3451
rect 11989 3349 12023 3383
rect 23489 3349 23523 3383
rect 25881 3349 25915 3383
rect 26157 3349 26191 3383
rect 56057 3621 56091 3655
rect 52377 3553 52411 3587
rect 61761 3621 61795 3655
rect 49249 3485 49283 3519
rect 49525 3485 49559 3519
rect 51457 3485 51491 3519
rect 51733 3485 51767 3519
rect 54309 3485 54343 3519
rect 55045 3485 55079 3519
rect 55965 3485 55999 3519
rect 56425 3485 56459 3519
rect 58173 3485 58207 3519
rect 58449 3485 58483 3519
rect 61117 3485 61151 3519
rect 61209 3485 61243 3519
rect 48237 3417 48271 3451
rect 49065 3417 49099 3451
rect 54401 3417 54435 3451
rect 63877 3621 63911 3655
rect 64061 3621 64095 3655
rect 69489 3621 69523 3655
rect 71789 3621 71823 3655
rect 72249 3621 72283 3655
rect 89453 3621 89487 3655
rect 90281 3621 90315 3655
rect 146033 3621 146067 3655
rect 149989 3621 150023 3655
rect 150817 3621 150851 3655
rect 63325 3553 63359 3587
rect 62865 3485 62899 3519
rect 63785 3485 63819 3519
rect 62129 3417 62163 3451
rect 68109 3553 68143 3587
rect 72801 3553 72835 3587
rect 130301 3553 130335 3587
rect 67557 3485 67591 3519
rect 67649 3485 67683 3519
rect 68937 3485 68971 3519
rect 70685 3485 70719 3519
rect 71697 3485 71731 3519
rect 71973 3485 72007 3519
rect 72709 3485 72743 3519
rect 73169 3485 73203 3519
rect 88257 3485 88291 3519
rect 89361 3485 89395 3519
rect 90373 3485 90407 3519
rect 91753 3485 91787 3519
rect 102333 3485 102367 3519
rect 102793 3485 102827 3519
rect 121837 3485 121871 3519
rect 122113 3485 122147 3519
rect 124873 3485 124907 3519
rect 125333 3485 125367 3519
rect 126345 3485 126379 3519
rect 130761 3485 130795 3519
rect 131313 3485 131347 3519
rect 133429 3485 133463 3519
rect 133889 3485 133923 3519
rect 138673 3485 138707 3519
rect 139133 3485 139167 3519
rect 145941 3485 145975 3519
rect 146493 3485 146527 3519
rect 149897 3485 149931 3519
rect 151553 3485 151587 3519
rect 164157 3485 164191 3519
rect 164617 3485 164651 3519
rect 70777 3417 70811 3451
rect 71237 3417 71271 3451
rect 91845 3417 91879 3451
rect 100861 3417 100895 3451
rect 103161 3417 103195 3451
rect 106657 3417 106691 3451
rect 45661 3349 45695 3383
rect 56977 3349 57011 3383
rect 59461 3349 59495 3383
rect 61853 3349 61887 3383
rect 62497 3349 62531 3383
rect 64061 3349 64095 3383
rect 64337 3349 64371 3383
rect 66545 3349 66579 3383
rect 68477 3349 68511 3383
rect 69029 3349 69063 3383
rect 70041 3349 70075 3383
rect 71513 3349 71547 3383
rect 71973 3349 72007 3383
rect 72617 3349 72651 3383
rect 73721 3349 73755 3383
rect 88349 3349 88383 3383
rect 88809 3349 88843 3383
rect 89913 3349 89947 3383
rect 90465 3349 90499 3383
rect 90925 3349 90959 3383
rect 92305 3349 92339 3383
rect 21925 3145 21959 3179
rect 44833 3145 44867 3179
rect 46489 3145 46523 3179
rect 47593 3145 47627 3179
rect 56701 3145 56735 3179
rect 57345 3145 57379 3179
rect 61393 3145 61427 3179
rect 62313 3145 62347 3179
rect 63417 3145 63451 3179
rect 64429 3145 64463 3179
rect 73537 3145 73571 3179
rect 88441 3145 88475 3179
rect 19901 3077 19935 3111
rect 23305 3077 23339 3111
rect 24961 3077 24995 3111
rect 28549 3077 28583 3111
rect 45385 3077 45419 3111
rect 53573 3077 53607 3111
rect 58725 3077 58759 3111
rect 3617 3009 3651 3043
rect 4721 3009 4755 3043
rect 7665 3009 7699 3043
rect 8493 3009 8527 3043
rect 9781 3009 9815 3043
rect 11713 3009 11747 3043
rect 13277 3009 13311 3043
rect 18429 3009 18463 3043
rect 20545 3009 20579 3043
rect 21833 3009 21867 3043
rect 24041 3009 24075 3043
rect 25605 3009 25639 3043
rect 27445 3009 27479 3043
rect 29193 3009 29227 3043
rect 30941 3009 30975 3043
rect 36737 3009 36771 3043
rect 40325 3009 40359 3043
rect 41337 3009 41371 3043
rect 43729 3009 43763 3043
rect 44097 3009 44131 3043
rect 44465 3009 44499 3043
rect 45569 3009 45603 3043
rect 47501 3009 47535 3043
rect 48789 3009 48823 3043
rect 54217 3009 54251 3043
rect 55137 3009 55171 3043
rect 56609 3009 56643 3043
rect 58633 3009 58667 3043
rect 60289 3009 60323 3043
rect 60381 3009 60415 3043
rect 60749 3009 60783 3043
rect 61117 3009 61151 3043
rect 62221 3009 62255 3043
rect 63325 3009 63359 3043
rect 64337 3009 64371 3043
rect 68477 3009 68511 3043
rect 69489 3009 69523 3043
rect 70501 3009 70535 3043
rect 71513 3009 71547 3043
rect 71605 3009 71639 3043
rect 73261 3009 73295 3043
rect 73445 3009 73479 3043
rect 87337 3009 87371 3043
rect 88349 3009 88383 3043
rect 90373 3009 90407 3043
rect 91845 3009 91879 3043
rect 92213 3009 92247 3043
rect 2605 2941 2639 2975
rect 6101 2941 6135 2975
rect 12725 2941 12759 2975
rect 18061 2941 18095 2975
rect 23305 2941 23339 2975
rect 23397 2941 23431 2975
rect 30573 2941 30607 2975
rect 36185 2941 36219 2975
rect 38945 2941 38979 2975
rect 39773 2941 39807 2975
rect 42717 2941 42751 2975
rect 57621 2941 57655 2975
rect 61301 2941 61335 2975
rect 65349 2941 65383 2975
rect 66729 2941 66763 2975
rect 4905 2873 4939 2907
rect 7389 2873 7423 2907
rect 9965 2873 9999 2907
rect 27905 2873 27939 2907
rect 56057 2873 56091 2907
rect 61209 2873 61243 2907
rect 70593 2873 70627 2907
rect 74457 2941 74491 2975
rect 76205 2941 76239 2975
rect 76757 2941 76791 2975
rect 77217 2941 77251 2975
rect 80897 2941 80931 2975
rect 83105 2941 83139 2975
rect 86325 2941 86359 2975
rect 91385 2941 91419 2975
rect 5549 2805 5583 2839
rect 19073 2805 19107 2839
rect 25973 2805 26007 2839
rect 27537 2805 27571 2839
rect 41429 2805 41463 2839
rect 48881 2805 48915 2839
rect 54585 2805 54619 2839
rect 55229 2805 55263 2839
rect 68569 2805 68603 2839
rect 69581 2805 69615 2839
rect 73261 2805 73295 2839
rect 87429 2805 87463 2839
rect 3709 2601 3743 2635
rect 3893 2601 3927 2635
rect 4721 2601 4755 2635
rect 8493 2601 8527 2635
rect 11989 2601 12023 2635
rect 22569 2601 22603 2635
rect 22845 2601 22879 2635
rect 23765 2601 23799 2635
rect 24685 2601 24719 2635
rect 24961 2601 24995 2635
rect 25421 2601 25455 2635
rect 27261 2601 27295 2635
rect 29653 2601 29687 2635
rect 30941 2601 30975 2635
rect 39589 2601 39623 2635
rect 40233 2601 40267 2635
rect 41429 2601 41463 2635
rect 43177 2601 43211 2635
rect 43361 2601 43395 2635
rect 43637 2601 43671 2635
rect 44925 2601 44959 2635
rect 45569 2601 45603 2635
rect 47501 2601 47535 2635
rect 49065 2601 49099 2635
rect 52837 2601 52871 2635
rect 53297 2601 53331 2635
rect 53665 2601 53699 2635
rect 55229 2601 55263 2635
rect 56701 2601 56735 2635
rect 57253 2601 57287 2635
rect 58725 2601 58759 2635
rect 60381 2601 60415 2635
rect 60933 2601 60967 2635
rect 61301 2601 61335 2635
rect 62681 2601 62715 2635
rect 63509 2601 63543 2635
rect 63693 2601 63727 2635
rect 64521 2601 64555 2635
rect 66545 2601 66579 2635
rect 67557 2601 67591 2635
rect 68569 2601 68603 2635
rect 70133 2601 70167 2635
rect 70501 2601 70535 2635
rect 71605 2601 71639 2635
rect 71881 2601 71915 2635
rect 73537 2601 73571 2635
rect 74273 2601 74307 2635
rect 74641 2601 74675 2635
rect 74825 2601 74859 2635
rect 75101 2601 75135 2635
rect 80805 2601 80839 2635
rect 82001 2601 82035 2635
rect 83473 2601 83507 2635
rect 86969 2601 87003 2635
rect 87337 2601 87371 2635
rect 87613 2601 87647 2635
rect 88441 2601 88475 2635
rect 90281 2601 90315 2635
rect 18337 2533 18371 2567
rect 19993 2533 20027 2567
rect 21649 2533 21683 2567
rect 2237 2465 2271 2499
rect 4813 2465 4847 2499
rect 5825 2465 5859 2499
rect 9597 2465 9631 2499
rect 10701 2465 10735 2499
rect 11621 2465 11655 2499
rect 23857 2465 23891 2499
rect 28365 2465 28399 2499
rect 29285 2465 29319 2499
rect 39589 2465 39623 2499
rect 45201 2465 45235 2499
rect 46029 2465 46063 2499
rect 46765 2465 46799 2499
rect 54033 2465 54067 2499
rect 3801 2397 3835 2431
rect 4261 2397 4295 2431
rect 6377 2397 6411 2431
rect 9689 2397 9723 2431
rect 11253 2397 11287 2431
rect 18521 2397 18555 2431
rect 18889 2397 18923 2431
rect 19257 2397 19291 2431
rect 20269 2397 20303 2431
rect 21189 2397 21223 2431
rect 21465 2397 21499 2431
rect 22385 2397 22419 2431
rect 22569 2397 22603 2431
rect 24501 2397 24535 2431
rect 24685 2397 24719 2431
rect 25789 2397 25823 2431
rect 26157 2397 26191 2431
rect 26525 2397 26559 2431
rect 26617 2397 26651 2431
rect 27353 2397 27387 2431
rect 28917 2397 28951 2431
rect 36553 2397 36587 2431
rect 38945 2397 38979 2431
rect 39129 2397 39163 2431
rect 39497 2397 39531 2431
rect 39865 2397 39899 2431
rect 43085 2397 43119 2431
rect 43361 2397 43395 2431
rect 44097 2397 44131 2431
rect 44465 2397 44499 2431
rect 44741 2397 44775 2431
rect 44925 2397 44959 2431
rect 45937 2397 45971 2431
rect 46397 2397 46431 2431
rect 49893 2397 49927 2431
rect 50261 2397 50295 2431
rect 50905 2397 50939 2431
rect 52745 2397 52779 2431
rect 54585 2397 54619 2431
rect 56241 2397 56275 2431
rect 57161 2397 57195 2431
rect 57713 2397 57747 2431
rect 58173 2397 58207 2431
rect 60105 2397 60139 2431
rect 6745 2329 6779 2363
rect 9229 2329 9263 2363
rect 12081 2329 12115 2363
rect 13093 2329 13127 2363
rect 44005 2329 44039 2363
rect 59461 2329 59495 2363
rect 65073 2465 65107 2499
rect 68017 2465 68051 2499
rect 60473 2397 60507 2431
rect 61117 2397 61151 2431
rect 62589 2397 62623 2431
rect 63049 2397 63083 2431
rect 63601 2397 63635 2431
rect 66453 2397 66487 2431
rect 66729 2397 66763 2431
rect 67465 2397 67499 2431
rect 69213 2397 69247 2431
rect 69489 2397 69523 2431
rect 70685 2397 70719 2431
rect 71789 2397 71823 2431
rect 73445 2397 73479 2431
rect 74549 2397 74583 2431
rect 100033 2533 100067 2567
rect 85405 2465 85439 2499
rect 89821 2465 89855 2499
rect 90373 2465 90407 2499
rect 91385 2465 91419 2499
rect 76573 2397 76607 2431
rect 76665 2397 76699 2431
rect 76849 2397 76883 2431
rect 77309 2397 77343 2431
rect 79333 2397 79367 2431
rect 80713 2397 80747 2431
rect 81173 2397 81207 2431
rect 81909 2397 81943 2431
rect 82369 2397 82403 2431
rect 83381 2397 83415 2431
rect 83657 2397 83691 2431
rect 86417 2397 86451 2431
rect 87521 2397 87555 2431
rect 88533 2397 88567 2431
rect 91937 2397 91971 2431
rect 92213 2397 92247 2431
rect 71237 2329 71271 2363
rect 74825 2329 74859 2363
rect 86509 2329 86543 2363
rect 88073 2329 88107 2363
rect 7205 2261 7239 2295
rect 7757 2261 7791 2295
rect 19625 2261 19659 2295
rect 20453 2261 20487 2295
rect 21465 2261 21499 2295
rect 22201 2261 22235 2295
rect 26617 2261 26651 2295
rect 26893 2261 26927 2295
rect 30297 2261 30331 2295
rect 55873 2261 55907 2295
rect 60381 2261 60415 2295
rect 62313 2261 62347 2295
rect 64153 2261 64187 2295
rect 66729 2261 66763 2295
rect 67005 2261 67039 2295
rect 69305 2261 69339 2295
rect 69489 2261 69523 2295
rect 69765 2261 69799 2295
rect 70777 2261 70811 2295
rect 72341 2261 72375 2295
rect 73997 2261 74031 2295
rect 83657 2261 83691 2295
rect 83933 2261 83967 2295
rect 88625 2261 88659 2295
rect 89085 2261 89119 2295
rect 6285 2057 6319 2091
rect 17325 2057 17359 2091
rect 42809 2057 42843 2091
rect 44189 2057 44223 2091
rect 48973 2057 49007 2091
rect 60381 2057 60415 2091
rect 63877 2057 63911 2091
rect 65165 2057 65199 2091
rect 66821 2057 66855 2091
rect 70041 2057 70075 2091
rect 71053 2057 71087 2091
rect 73537 2057 73571 2091
rect 77585 2057 77619 2091
rect 78045 2057 78079 2091
rect 79149 2057 79183 2091
rect 79517 2057 79551 2091
rect 82277 2057 82311 2091
rect 83105 2057 83139 2091
rect 84761 2057 84795 2091
rect 85773 2057 85807 2091
rect 88901 2057 88935 2091
rect 42073 1989 42107 2023
rect 42993 1989 43027 2023
rect 51181 1989 51215 2023
rect 54033 1989 54067 2023
rect 61669 1989 61703 2023
rect 63693 1989 63727 2023
rect 73077 1989 73111 2023
rect 4813 1921 4847 1955
rect 8217 1921 8251 1955
rect 10793 1921 10827 1955
rect 20913 1921 20947 1955
rect 21005 1921 21039 1955
rect 25237 1921 25271 1955
rect 26709 1921 26743 1955
rect 30021 1921 30055 1955
rect 30113 1921 30147 1955
rect 30481 1921 30515 1955
rect 2237 1853 2271 1887
rect 3249 1853 3283 1887
rect 4261 1853 4295 1887
rect 6653 1853 6687 1887
rect 7665 1853 7699 1887
rect 9229 1853 9263 1887
rect 10241 1853 10275 1887
rect 11161 1853 11195 1887
rect 11713 1853 11747 1887
rect 15117 1853 15151 1887
rect 18337 1853 18371 1887
rect 19349 1853 19383 1887
rect 20361 1853 20395 1887
rect 21741 1853 21775 1887
rect 23673 1853 23707 1887
rect 24685 1853 24719 1887
rect 26065 1853 26099 1887
rect 28549 1853 28583 1887
rect 30757 1853 30791 1887
rect 31309 1853 31343 1887
rect 32321 1853 32355 1887
rect 34529 1853 34563 1887
rect 35541 1853 35575 1887
rect 35909 1853 35943 1887
rect 37197 1853 37231 1887
rect 43729 1921 43763 1955
rect 45569 1921 45603 1955
rect 46121 1921 46155 1955
rect 47777 1921 47811 1955
rect 48789 1921 48823 1955
rect 53665 1921 53699 1955
rect 55229 1921 55263 1955
rect 57897 1921 57931 1955
rect 59001 1921 59035 1955
rect 59553 1921 59587 1955
rect 60013 1921 60047 1955
rect 60565 1921 60599 1955
rect 61301 1921 61335 1955
rect 62497 1921 62531 1955
rect 62865 1921 62899 1955
rect 63785 1921 63819 1955
rect 64245 1921 64279 1955
rect 65073 1921 65107 1955
rect 66729 1921 66763 1955
rect 68109 1921 68143 1955
rect 68569 1921 68603 1955
rect 68845 1921 68879 1955
rect 69949 1921 69983 1955
rect 70961 1921 70995 1955
rect 72341 1921 72375 1955
rect 73445 1921 73479 1955
rect 73721 1921 73755 1955
rect 52193 1853 52227 1887
rect 53205 1853 53239 1887
rect 54585 1853 54619 1887
rect 57437 1853 57471 1887
rect 60933 1853 60967 1887
rect 62589 1853 62623 1887
rect 68201 1853 68235 1887
rect 72433 1853 72467 1887
rect 73813 1921 73847 1955
rect 76665 1921 76699 1955
rect 77493 1921 77527 1955
rect 79057 1921 79091 1955
rect 80437 1921 80471 1955
rect 80897 1921 80931 1955
rect 81357 1921 81391 1955
rect 82185 1921 82219 1955
rect 83381 1921 83415 1955
rect 83657 1921 83691 1955
rect 84669 1921 84703 1955
rect 85681 1921 85715 1955
rect 86877 1921 86911 1955
rect 88257 1921 88291 1955
rect 91937 1921 91971 1955
rect 75101 1853 75135 1887
rect 76113 1853 76147 1887
rect 77033 1853 77067 1887
rect 73813 1785 73847 1819
rect 80989 1853 81023 1887
rect 83473 1853 83507 1887
rect 80437 1785 80471 1819
rect 84393 1853 84427 1887
rect 86693 1853 86727 1887
rect 90373 1853 90407 1887
rect 91385 1853 91419 1887
rect 88165 1785 88199 1819
rect 5181 1717 5215 1751
rect 21005 1717 21039 1751
rect 21281 1717 21315 1751
rect 22569 1717 22603 1751
rect 42993 1717 43027 1751
rect 43545 1717 43579 1751
rect 44465 1717 44499 1751
rect 47409 1717 47443 1751
rect 55597 1717 55631 1751
rect 57161 1717 57195 1751
rect 59093 1717 59127 1751
rect 67649 1717 67683 1751
rect 71697 1717 71731 1751
rect 73721 1717 73755 1751
rect 73997 1717 74031 1751
rect 83657 1717 83691 1751
rect 83933 1717 83967 1751
rect 86693 1717 86727 1751
rect 98653 1649 98687 1683
rect 99389 1581 99423 1615
rect 3801 1513 3835 1547
rect 7205 1513 7239 1547
rect 9229 1513 9263 1547
rect 10517 1513 10551 1547
rect 15117 1513 15151 1547
rect 25053 1513 25087 1547
rect 26801 1513 26835 1547
rect 28273 1513 28307 1547
rect 30481 1513 30515 1547
rect 46305 1513 46339 1547
rect 46489 1513 46523 1547
rect 49617 1513 49651 1547
rect 57069 1513 57103 1547
rect 58817 1513 58851 1547
rect 61117 1513 61151 1547
rect 61393 1513 61427 1547
rect 62129 1513 62163 1547
rect 63325 1513 63359 1547
rect 70041 1513 70075 1547
rect 72709 1513 72743 1547
rect 75193 1513 75227 1547
rect 81633 1513 81667 1547
rect 84853 1513 84887 1547
rect 91201 1513 91235 1547
rect 98653 1513 98687 1547
rect 23857 1445 23891 1479
rect 33885 1445 33919 1479
rect 5365 1377 5399 1411
rect 9505 1377 9539 1411
rect 11621 1377 11655 1411
rect 16221 1377 16255 1411
rect 21189 1377 21223 1411
rect 22569 1377 22603 1411
rect 29377 1377 29411 1411
rect 32413 1377 32447 1411
rect 41521 1377 41555 1411
rect 43729 1377 43763 1411
rect 55229 1445 55263 1479
rect 84761 1445 84795 1479
rect 46673 1377 46707 1411
rect 60841 1377 60875 1411
rect 61117 1377 61151 1411
rect 62865 1377 62899 1411
rect 65625 1377 65659 1411
rect 67373 1377 67407 1411
rect 68569 1377 68603 1411
rect 72709 1377 72743 1411
rect 72985 1377 73019 1411
rect 74365 1377 74399 1411
rect 77309 1377 77343 1411
rect 83013 1377 83047 1411
rect 84209 1377 84243 1411
rect 86325 1377 86359 1411
rect 88901 1377 88935 1411
rect 89913 1377 89947 1411
rect 92213 1377 92247 1411
rect 4353 1309 4387 1343
rect 5917 1309 5951 1343
rect 7757 1309 7791 1343
rect 10609 1309 10643 1343
rect 12173 1309 12207 1343
rect 15209 1309 15243 1343
rect 16773 1309 16807 1343
rect 18889 1309 18923 1343
rect 19533 1309 19567 1343
rect 19809 1309 19843 1343
rect 20177 1309 20211 1343
rect 21741 1309 21775 1343
rect 22109 1309 22143 1343
rect 23673 1309 23707 1343
rect 26157 1309 26191 1343
rect 26525 1309 26559 1343
rect 27353 1309 27387 1343
rect 28365 1309 28399 1343
rect 29929 1309 29963 1343
rect 30573 1309 30607 1343
rect 31125 1309 31159 1343
rect 31401 1309 31435 1343
rect 32965 1309 32999 1343
rect 33057 1309 33091 1343
rect 33609 1309 33643 1343
rect 33793 1309 33827 1343
rect 34529 1309 34563 1343
rect 35357 1309 35391 1343
rect 35725 1309 35759 1343
rect 36093 1309 36127 1343
rect 37013 1309 37047 1343
rect 37381 1309 37415 1343
rect 37749 1309 37783 1343
rect 38117 1309 38151 1343
rect 39221 1309 39255 1343
rect 40141 1309 40175 1343
rect 42717 1309 42751 1343
rect 44281 1309 44315 1343
rect 45109 1309 45143 1343
rect 45293 1309 45327 1343
rect 46121 1309 46155 1343
rect 46305 1309 46339 1343
rect 48881 1309 48915 1343
rect 49801 1309 49835 1343
rect 50445 1309 50479 1343
rect 50905 1309 50939 1343
rect 52009 1309 52043 1343
rect 52469 1309 52503 1343
rect 53573 1309 53607 1343
rect 53849 1309 53883 1343
rect 54217 1309 54251 1343
rect 54585 1309 54619 1343
rect 54953 1309 54987 1343
rect 55597 1309 55631 1343
rect 55781 1309 55815 1343
rect 56149 1309 56183 1343
rect 56977 1309 57011 1343
rect 57529 1309 57563 1343
rect 58357 1309 58391 1343
rect 59093 1309 59127 1343
rect 59461 1309 59495 1343
rect 60565 1309 60599 1343
rect 61761 1309 61795 1343
rect 62313 1309 62347 1343
rect 63601 1309 63635 1343
rect 63785 1309 63819 1343
rect 63969 1309 64003 1343
rect 64429 1309 64463 1343
rect 65073 1309 65107 1343
rect 65993 1309 66027 1343
rect 66545 1309 66579 1343
rect 66637 1309 66671 1343
rect 67557 1309 67591 1343
rect 69029 1309 69063 1343
rect 70961 1309 70995 1343
rect 71513 1309 71547 1343
rect 71789 1309 71823 1343
rect 72065 1309 72099 1343
rect 72433 1309 72467 1343
rect 72893 1309 72927 1343
rect 74549 1309 74583 1343
rect 76113 1309 76147 1343
rect 76297 1309 76331 1343
rect 77861 1309 77895 1343
rect 79333 1309 79367 1343
rect 79425 1309 79459 1343
rect 79609 1309 79643 1343
rect 80069 1309 80103 1343
rect 80621 1309 80655 1343
rect 81909 1309 81943 1343
rect 84577 1309 84611 1343
rect 84761 1309 84795 1343
rect 85405 1309 85439 1343
rect 86417 1309 86451 1343
rect 87245 1309 87279 1343
rect 87521 1309 87555 1343
rect 88441 1309 88475 1343
rect 90465 1309 90499 1343
rect 90741 1309 90775 1343
rect 91293 1309 91327 1343
rect 91753 1309 91787 1343
rect 3341 1241 3375 1275
rect 4169 1241 4203 1275
rect 19257 1241 19291 1275
rect 25329 1241 25363 1275
rect 34897 1241 34931 1275
rect 36461 1241 36495 1275
rect 39865 1241 39899 1275
rect 48237 1241 48271 1275
rect 49341 1241 49375 1275
rect 57989 1241 58023 1275
rect 69489 1241 69523 1275
rect 80713 1241 80747 1275
rect 81357 1241 81391 1275
rect 82369 1241 82403 1275
rect 85957 1241 85991 1275
rect 86969 1241 87003 1275
rect 2237 1173 2271 1207
rect 6285 1173 6319 1207
rect 6745 1173 6779 1207
rect 8309 1173 8343 1207
rect 12541 1173 12575 1207
rect 13001 1173 13035 1207
rect 17141 1173 17175 1207
rect 19809 1173 19843 1207
rect 19901 1173 19935 1207
rect 24501 1173 24535 1207
rect 30573 1173 30607 1207
rect 30849 1173 30883 1207
rect 33057 1173 33091 1207
rect 33333 1173 33367 1207
rect 44649 1173 44683 1207
rect 47593 1173 47627 1207
rect 56517 1173 56551 1207
rect 59093 1173 59127 1207
rect 59185 1173 59219 1207
rect 65165 1173 65199 1207
rect 67097 1173 67131 1207
rect 74917 1173 74951 1207
rect 78229 1173 78263 1207
rect 78965 1173 78999 1207
rect 80529 1173 80563 1207
rect 82001 1173 82035 1207
rect 82737 1173 82771 1207
rect 85497 1173 85531 1207
rect 86509 1173 86543 1207
rect 87613 1173 87647 1207
rect 88073 1173 88107 1207
rect 91385 1173 91419 1207
rect 150449 3417 150483 3451
rect 151645 3417 151679 3451
rect 155141 3417 155175 3451
rect 158545 3417 158579 3451
rect 102425 3349 102459 3383
rect 103345 3349 103379 3383
rect 107853 3349 107887 3383
rect 114845 3349 114879 3383
rect 115949 3349 115983 3383
rect 119629 3349 119663 3383
rect 121653 3349 121687 3383
rect 122113 3349 122147 3383
rect 122389 3349 122423 3383
rect 124597 3349 124631 3383
rect 125793 3349 125827 3383
rect 126989 3349 127023 3383
rect 131681 3349 131715 3383
rect 137293 3349 137327 3383
rect 138765 3349 138799 3383
rect 148241 3349 148275 3383
rect 152105 3349 152139 3383
rect 156153 3349 156187 3383
rect 159649 3349 159683 3383
rect 160293 3349 160327 3383
rect 161397 3349 161431 3383
rect 162317 3349 162351 3383
rect 133245 3145 133279 3179
rect 134257 3145 134291 3179
rect 145389 3145 145423 3179
rect 154313 3145 154347 3179
rect 155325 3145 155359 3179
rect 156337 3145 156371 3179
rect 159557 3145 159591 3179
rect 160753 3145 160787 3179
rect 164065 3145 164099 3179
rect 165077 3145 165111 3179
rect 107577 3077 107611 3111
rect 107853 3077 107887 3111
rect 130025 3077 130059 3111
rect 102333 3009 102367 3043
rect 102793 3009 102827 3043
rect 103337 3009 103371 3043
rect 104357 2941 104391 2975
rect 103437 2873 103471 2907
rect 107761 3009 107795 3043
rect 109601 3009 109635 3043
rect 109693 3009 109727 3043
rect 110889 3009 110923 3043
rect 113649 3009 113683 3043
rect 117145 3009 117179 3043
rect 122389 3009 122423 3043
rect 122481 3009 122515 3043
rect 126345 3009 126379 3043
rect 127909 3009 127943 3043
rect 126437 2941 126471 2975
rect 128001 2941 128035 2975
rect 113741 2873 113775 2907
rect 133153 3009 133187 3043
rect 134165 3009 134199 3043
rect 136649 3009 136683 3043
rect 137753 3009 137787 3043
rect 138765 3009 138799 3043
rect 139041 3009 139075 3043
rect 145297 3009 145331 3043
rect 149069 3009 149103 3043
rect 154221 3009 154255 3043
rect 155233 3009 155267 3043
rect 156245 3009 156279 3043
rect 159465 3009 159499 3043
rect 160661 3009 160695 3043
rect 163973 3009 164007 3043
rect 164985 3009 165019 3043
rect 165445 3009 165479 3043
rect 137845 2873 137879 2907
rect 139777 2941 139811 2975
rect 141433 2941 141467 2975
rect 143181 2941 143215 2975
rect 158269 2941 158303 2975
rect 162041 2941 162075 2975
rect 102425 2805 102459 2839
rect 103253 2805 103287 2839
rect 103897 2805 103931 2839
rect 107577 2805 107611 2839
rect 110981 2805 111015 2839
rect 117237 2805 117271 2839
rect 130025 2805 130059 2839
rect 136741 2805 136775 2839
rect 138857 2805 138891 2839
rect 139041 2805 139075 2839
rect 139317 2805 139351 2839
rect 149161 2805 149195 2839
rect 164709 2805 164743 2839
rect 103989 2601 104023 2635
rect 104173 2601 104207 2635
rect 108497 2601 108531 2635
rect 109509 2601 109543 2635
rect 109877 2601 109911 2635
rect 110705 2601 110739 2635
rect 111349 2601 111383 2635
rect 111533 2601 111567 2635
rect 112729 2601 112763 2635
rect 113741 2601 113775 2635
rect 114569 2601 114603 2635
rect 117237 2601 117271 2635
rect 118433 2601 118467 2635
rect 120825 2601 120859 2635
rect 122389 2601 122423 2635
rect 123769 2601 123803 2635
rect 124965 2601 124999 2635
rect 126069 2601 126103 2635
rect 126897 2601 126931 2635
rect 127541 2601 127575 2635
rect 161765 2601 161799 2635
rect 162777 2601 162811 2635
rect 103345 2465 103379 2499
rect 102333 2397 102367 2431
rect 103805 2397 103839 2431
rect 108405 2397 108439 2431
rect 109417 2397 109451 2431
rect 109693 2397 109727 2431
rect 110613 2397 110647 2431
rect 111165 2397 111199 2431
rect 127725 2533 127759 2567
rect 155877 2533 155911 2567
rect 157349 2533 157383 2567
rect 158453 2533 158487 2567
rect 160201 2533 160235 2567
rect 111625 2397 111659 2431
rect 111901 2397 111935 2431
rect 112637 2397 112671 2431
rect 112913 2397 112947 2431
rect 113649 2397 113683 2431
rect 116225 2397 116259 2431
rect 117329 2397 117363 2431
rect 117605 2397 117639 2431
rect 118341 2397 118375 2431
rect 118893 2397 118927 2431
rect 120733 2397 120767 2431
rect 123677 2397 123711 2431
rect 124873 2397 124907 2431
rect 125977 2397 126011 2431
rect 126253 2397 126287 2431
rect 127449 2397 127483 2431
rect 127725 2329 127759 2363
rect 127817 2465 127851 2499
rect 139685 2465 139719 2499
rect 142905 2465 142939 2499
rect 145389 2465 145423 2499
rect 146401 2465 146435 2499
rect 147781 2465 147815 2499
rect 148793 2465 148827 2499
rect 149989 2465 150023 2499
rect 151001 2465 151035 2499
rect 159465 2465 159499 2499
rect 127909 2397 127943 2431
rect 130209 2397 130243 2431
rect 130301 2397 130335 2431
rect 134993 2397 135027 2431
rect 135085 2397 135119 2431
rect 136373 2397 136407 2431
rect 137569 2397 137603 2431
rect 138397 2397 138431 2431
rect 138673 2397 138707 2431
rect 140237 2397 140271 2431
rect 140513 2397 140547 2431
rect 142813 2397 142847 2431
rect 145297 2397 145331 2431
rect 146309 2397 146343 2431
rect 146769 2397 146803 2431
rect 147689 2397 147723 2431
rect 148149 2397 148183 2431
rect 148701 2397 148735 2431
rect 149897 2397 149931 2431
rect 150909 2397 150943 2431
rect 151369 2397 151403 2431
rect 151921 2397 151955 2431
rect 152381 2397 152415 2431
rect 155785 2397 155819 2431
rect 156613 2397 156647 2431
rect 157257 2397 157291 2431
rect 158361 2397 158395 2431
rect 158821 2397 158855 2431
rect 159373 2397 159407 2431
rect 159833 2397 159867 2431
rect 161673 2397 161707 2431
rect 162133 2397 162167 2431
rect 162685 2397 162719 2431
rect 163145 2397 163179 2431
rect 164617 2397 164651 2431
rect 130669 2329 130703 2363
rect 135453 2329 135487 2363
rect 137293 2329 137327 2363
rect 138029 2329 138063 2363
rect 149161 2329 149195 2363
rect 152013 2329 152047 2363
rect 156337 2329 156371 2363
rect 165445 2329 165479 2363
rect 104081 2261 104115 2295
rect 105001 2261 105035 2295
rect 107761 2261 107795 2295
rect 108957 2261 108991 2295
rect 109693 2261 109727 2295
rect 110337 2261 110371 2295
rect 111349 2261 111383 2295
rect 111717 2261 111751 2295
rect 111901 2261 111935 2295
rect 112177 2261 112211 2295
rect 112913 2261 112947 2295
rect 113189 2261 113223 2295
rect 114201 2261 114235 2295
rect 116317 2261 116351 2295
rect 116777 2261 116811 2295
rect 117421 2261 117455 2295
rect 117605 2261 117639 2295
rect 117881 2261 117915 2295
rect 119353 2261 119387 2295
rect 121193 2261 121227 2295
rect 124229 2261 124263 2295
rect 125425 2261 125459 2295
rect 126253 2261 126287 2295
rect 126529 2261 126563 2295
rect 127817 2261 127851 2295
rect 128369 2261 128403 2295
rect 133245 2261 133279 2295
rect 134165 2261 134199 2295
rect 136465 2261 136499 2295
rect 136833 2261 136867 2295
rect 137661 2261 137695 2295
rect 141065 2261 141099 2295
rect 143365 2261 143399 2295
rect 145757 2261 145791 2295
rect 146125 2261 146159 2295
rect 149621 2261 149655 2295
rect 150449 2261 150483 2295
rect 154313 2261 154347 2295
rect 155233 2261 155267 2295
rect 157717 2261 157751 2295
rect 160661 2261 160695 2295
rect 164065 2261 164099 2295
rect 103253 2057 103287 2091
rect 106565 2057 106599 2091
rect 107853 2057 107887 2091
rect 130853 2057 130887 2091
rect 139041 2057 139075 2091
rect 139593 2057 139627 2091
rect 141157 2057 141191 2091
rect 146033 2057 146067 2091
rect 150357 2057 150391 2091
rect 153761 2057 153795 2091
rect 154773 2057 154807 2091
rect 155785 2057 155819 2091
rect 160937 2057 160971 2091
rect 162041 2057 162075 2091
rect 163973 2057 164007 2091
rect 117789 1989 117823 2023
rect 118341 1989 118375 2023
rect 119077 1989 119111 2023
rect 121101 1989 121135 2023
rect 122941 1989 122975 2023
rect 124689 1989 124723 2023
rect 136373 1989 136407 2023
rect 139317 1989 139351 2023
rect 152749 1989 152783 2023
rect 102333 1921 102367 1955
rect 103713 1921 103747 1955
rect 105277 1921 105311 1955
rect 106473 1921 106507 1955
rect 107761 1921 107795 1955
rect 108773 1921 108807 1955
rect 111349 1921 111383 1955
rect 112177 1921 112211 1955
rect 112637 1921 112671 1955
rect 115397 1921 115431 1955
rect 116225 1921 116259 1955
rect 117697 1921 117731 1955
rect 104725 1853 104759 1887
rect 108865 1853 108899 1887
rect 109785 1853 109819 1887
rect 110797 1853 110831 1887
rect 113833 1853 113867 1887
rect 114845 1853 114879 1887
rect 116317 1853 116351 1887
rect 118985 1921 119019 1955
rect 119997 1921 120031 1955
rect 121009 1921 121043 1955
rect 122849 1921 122883 1955
rect 124597 1921 124631 1955
rect 124873 1921 124907 1955
rect 127081 1921 127115 1955
rect 128185 1921 128219 1955
rect 130761 1921 130795 1955
rect 135821 1921 135855 1955
rect 138673 1921 138707 1955
rect 139501 1921 139535 1955
rect 141433 1921 141467 1955
rect 141893 1921 141927 1955
rect 144285 1921 144319 1955
rect 145941 1921 145975 1955
rect 149161 1921 149195 1955
rect 150265 1921 150299 1955
rect 152657 1921 152691 1955
rect 153669 1921 153703 1955
rect 154681 1921 154715 1955
rect 155693 1921 155727 1955
rect 156705 1921 156739 1955
rect 157165 1921 157199 1955
rect 158269 1921 158303 1955
rect 159833 1921 159867 1955
rect 160845 1921 160879 1955
rect 161949 1921 161983 1955
rect 163881 1921 163915 1955
rect 164893 1921 164927 1955
rect 166733 1921 166767 1955
rect 119537 1853 119571 1887
rect 102793 1785 102827 1819
rect 118341 1785 118375 1819
rect 125609 1853 125643 1887
rect 126621 1853 126655 1887
rect 130577 1853 130611 1887
rect 133705 1853 133739 1887
rect 134717 1853 134751 1887
rect 135361 1853 135395 1887
rect 137109 1853 137143 1887
rect 138121 1853 138155 1887
rect 143181 1853 143215 1887
rect 144193 1853 144227 1887
rect 147873 1853 147907 1887
rect 148885 1853 148919 1887
rect 165721 1853 165755 1887
rect 167101 1853 167135 1887
rect 128277 1785 128311 1819
rect 102425 1717 102459 1751
rect 111625 1717 111659 1751
rect 112269 1717 112303 1751
rect 118433 1717 118467 1751
rect 119905 1717 119939 1751
rect 120089 1717 120123 1751
rect 123953 1717 123987 1751
rect 124873 1717 124907 1751
rect 125149 1717 125183 1751
rect 129197 1717 129231 1751
rect 135913 1717 135947 1751
rect 139961 1717 139995 1751
rect 141525 1717 141559 1751
rect 156153 1717 156187 1751
rect 156797 1717 156831 1751
rect 158361 1717 158395 1751
rect 158729 1717 158763 1751
rect 159649 1717 159683 1751
rect 159925 1717 159959 1751
rect 104541 1513 104575 1547
rect 105829 1513 105863 1547
rect 117973 1513 118007 1547
rect 137569 1513 137603 1547
rect 138489 1513 138523 1547
rect 143365 1513 143399 1547
rect 158177 1513 158211 1547
rect 160109 1513 160143 1547
rect 166089 1513 166123 1547
rect 126161 1445 126195 1479
rect 102333 1377 102367 1411
rect 103529 1377 103563 1411
rect 106933 1377 106967 1411
rect 107853 1377 107887 1411
rect 110705 1377 110739 1411
rect 112637 1377 112671 1411
rect 113833 1377 113867 1411
rect 114017 1377 114051 1411
rect 116685 1377 116719 1411
rect 117421 1377 117455 1411
rect 118433 1377 118467 1411
rect 119445 1377 119479 1411
rect 121009 1377 121043 1411
rect 123953 1377 123987 1411
rect 124965 1377 124999 1411
rect 126345 1377 126379 1411
rect 129197 1377 129231 1411
rect 130209 1377 130243 1411
rect 133705 1377 133739 1411
rect 135361 1377 135395 1411
rect 136373 1377 136407 1411
rect 138673 1377 138707 1411
rect 139961 1377 139995 1411
rect 141157 1377 141191 1411
rect 142169 1377 142203 1411
rect 147873 1377 147907 1411
rect 148333 1377 148367 1411
rect 150357 1377 150391 1411
rect 156797 1377 156831 1411
rect 159281 1377 159315 1411
rect 165445 1377 165479 1411
rect 103897 1309 103931 1343
rect 105001 1309 105035 1343
rect 106013 1309 106047 1343
rect 106473 1309 106507 1343
rect 109049 1309 109083 1343
rect 109969 1309 110003 1343
rect 110613 1309 110647 1343
rect 111625 1309 111659 1343
rect 112729 1309 112763 1343
rect 113465 1309 113499 1343
rect 119905 1309 119939 1343
rect 120365 1309 120399 1343
rect 121837 1309 121871 1343
rect 122297 1309 122331 1343
rect 125517 1309 125551 1343
rect 125793 1309 125827 1343
rect 130761 1309 130795 1343
rect 131957 1309 131991 1343
rect 132233 1309 132267 1343
rect 133153 1309 133187 1343
rect 136649 1309 136683 1343
rect 137201 1309 137235 1343
rect 139777 1309 139811 1343
rect 140513 1309 140547 1343
rect 142721 1309 142755 1343
rect 142997 1309 143031 1343
rect 144929 1309 144963 1343
rect 145389 1309 145423 1343
rect 145941 1309 145975 1343
rect 146401 1309 146435 1343
rect 149897 1309 149931 1343
rect 149989 1309 150023 1343
rect 151369 1309 151403 1343
rect 152657 1309 152691 1343
rect 154405 1309 154439 1343
rect 155785 1309 155819 1343
rect 156889 1309 156923 1343
rect 157625 1309 157659 1343
rect 158269 1309 158303 1343
rect 159649 1309 159683 1343
rect 161121 1309 161155 1343
rect 161581 1309 161615 1343
rect 162409 1309 162443 1343
rect 163605 1309 163639 1343
rect 164065 1309 164099 1343
rect 164433 1309 164467 1343
rect 164985 1309 165019 1343
rect 166457 1309 166491 1343
rect 166733 1309 166767 1343
rect 167193 1309 167227 1343
rect 104265 1241 104299 1275
rect 105093 1241 105127 1275
rect 105461 1241 105495 1275
rect 108497 1241 108531 1275
rect 111073 1241 111107 1275
rect 111533 1241 111567 1275
rect 133245 1241 133279 1275
rect 145021 1241 145055 1275
rect 149161 1241 149195 1275
rect 150725 1241 150759 1275
rect 151829 1241 151863 1275
rect 160845 1241 160879 1275
rect 162961 1241 162995 1275
rect 167745 1241 167779 1275
rect 106105 1173 106139 1207
rect 107025 1173 107059 1207
rect 109509 1173 109543 1207
rect 115029 1173 115063 1207
rect 115581 1173 115615 1207
rect 116225 1173 116259 1207
rect 121929 1173 121963 1207
rect 122941 1173 122975 1207
rect 126989 1173 127023 1207
rect 128277 1173 128311 1207
rect 131129 1173 131163 1207
rect 132049 1173 132083 1207
rect 132233 1173 132267 1207
rect 132509 1173 132543 1207
rect 134349 1173 134383 1207
rect 144469 1173 144503 1207
rect 146033 1173 146067 1207
rect 146769 1173 146803 1207
rect 151461 1173 151495 1207
rect 153669 1173 153703 1207
rect 154865 1173 154899 1207
rect 161213 1173 161247 1207
rect 161949 1173 161983 1207
rect 162501 1173 162535 1207
rect 163697 1173 163731 1207
rect 166825 1173 166859 1207
rect 167561 1173 167595 1207
rect 100861 1037 100895 1071
rect 3433 969 3467 1003
rect 3617 969 3651 1003
rect 12173 969 12207 1003
rect 19349 969 19383 1003
rect 19809 969 19843 1003
rect 22201 969 22235 1003
rect 24961 969 24995 1003
rect 25881 969 25915 1003
rect 26341 969 26375 1003
rect 31861 969 31895 1003
rect 36369 969 36403 1003
rect 38485 969 38519 1003
rect 44833 969 44867 1003
rect 47685 969 47719 1003
rect 48789 969 48823 1003
rect 50077 969 50111 1003
rect 103989 969 104023 1003
rect 104633 969 104667 1003
rect 105277 969 105311 1003
rect 107853 969 107887 1003
rect 133521 969 133555 1003
rect 133705 969 133739 1003
rect 136097 969 136131 1003
rect 136373 969 136407 1003
rect 139041 969 139075 1003
rect 141065 969 141099 1003
rect 143181 969 143215 1003
rect 155233 969 155267 1003
rect 155785 969 155819 1003
rect 156613 969 156647 1003
rect 158545 969 158579 1003
rect 161305 969 161339 1003
rect 166641 969 166675 1003
rect 166825 969 166859 1003
rect 2237 901 2271 935
rect 5917 901 5951 935
rect 8769 901 8803 935
rect 3433 833 3467 867
rect 3709 833 3743 867
rect 5273 833 5307 867
rect 6193 833 6227 867
rect 7757 833 7791 867
rect 8125 833 8159 867
rect 9045 833 9079 867
rect 10609 833 10643 867
rect 12265 833 12299 867
rect 13829 833 13863 867
rect 15945 833 15979 867
rect 16681 833 16715 867
rect 16773 833 16807 867
rect 18245 833 18279 867
rect 18613 833 18647 867
rect 20729 833 20763 867
rect 21465 833 21499 867
rect 23489 833 23523 867
rect 24317 833 24351 867
rect 24869 833 24903 867
rect 26525 833 26559 867
rect 27905 833 27939 867
rect 28365 833 28399 867
rect 30389 833 30423 867
rect 30757 833 30791 867
rect 33517 833 33551 867
rect 33885 833 33919 867
rect 35449 833 35483 867
rect 36001 833 36035 867
rect 37657 833 37691 867
rect 4721 765 4755 799
rect 7205 765 7239 799
rect 10057 765 10091 799
rect 13277 765 13311 799
rect 14933 765 14967 799
rect 15761 765 15795 799
rect 16313 765 16347 799
rect 20453 765 20487 799
rect 24041 765 24075 799
rect 25421 765 25455 799
rect 27537 765 27571 799
rect 30481 765 30515 799
rect 38577 901 38611 935
rect 39129 833 39163 867
rect 41521 833 41555 867
rect 41613 833 41647 867
rect 42349 833 42383 867
rect 42717 833 42751 867
rect 43821 833 43855 867
rect 44005 833 44039 867
rect 46121 833 46155 867
rect 46305 833 46339 867
rect 47133 833 47167 867
rect 66361 901 66395 935
rect 68385 901 68419 935
rect 70593 901 70627 935
rect 70961 901 70995 935
rect 71881 901 71915 935
rect 74825 901 74859 935
rect 80529 901 80563 935
rect 84761 901 84795 935
rect 87981 901 88015 935
rect 90005 901 90039 935
rect 91845 901 91879 935
rect 92305 901 92339 935
rect 49617 833 49651 867
rect 50537 833 50571 867
rect 51641 833 51675 867
rect 51825 833 51859 867
rect 52561 833 52595 867
rect 52653 833 52687 867
rect 53481 833 53515 867
rect 54033 833 54067 867
rect 55873 833 55907 867
rect 56517 833 56551 867
rect 56885 833 56919 867
rect 58541 833 58575 867
rect 59185 833 59219 867
rect 60381 833 60415 867
rect 60473 833 60507 867
rect 61393 833 61427 867
rect 63785 833 63819 867
rect 64521 833 64555 867
rect 66453 833 66487 867
rect 68017 833 68051 867
rect 69213 833 69247 867
rect 69949 833 69983 867
rect 70501 833 70535 867
rect 71973 833 72007 867
rect 72893 833 72927 867
rect 73445 833 73479 867
rect 76481 833 76515 867
rect 76849 833 76883 867
rect 77493 833 77527 867
rect 78045 833 78079 867
rect 79333 833 79367 867
rect 79701 833 79735 867
rect 81173 833 81207 867
rect 81541 833 81575 867
rect 82093 833 82127 867
rect 83197 833 83231 867
rect 83657 833 83691 867
rect 84209 833 84243 867
rect 86049 833 86083 867
rect 86509 833 86543 867
rect 87429 833 87463 867
rect 88901 833 88935 867
rect 89913 833 89947 867
rect 90373 833 90407 867
rect 91753 833 91787 867
rect 102333 833 102367 867
rect 103897 833 103931 867
rect 41981 765 42015 799
rect 44281 765 44315 799
rect 48789 765 48823 799
rect 48973 765 49007 799
rect 110429 901 110463 935
rect 112729 901 112763 935
rect 113833 901 113867 935
rect 116225 901 116259 935
rect 105369 833 105403 867
rect 106473 833 106507 867
rect 107209 833 107243 867
rect 110889 833 110923 867
rect 111993 833 112027 867
rect 113925 833 113959 867
rect 115489 833 115523 867
rect 115857 833 115891 867
rect 116409 833 116443 867
rect 117973 833 118007 867
rect 119077 833 119111 867
rect 119261 833 119295 867
rect 120825 833 120859 867
rect 120917 833 120951 867
rect 122113 833 122147 867
rect 122665 833 122699 867
rect 123769 833 123803 867
rect 125617 833 125651 867
rect 126161 833 126195 867
rect 128277 833 128311 867
rect 128645 833 128679 867
rect 129289 833 129323 867
rect 131129 833 131163 867
rect 131405 833 131439 867
rect 132417 833 132451 867
rect 54861 765 54895 799
rect 57529 765 57563 799
rect 59645 765 59679 799
rect 61945 765 61979 799
rect 63509 765 63543 799
rect 67465 765 67499 799
rect 68937 765 68971 799
rect 75837 765 75871 799
rect 77585 765 77619 799
rect 78689 765 78723 799
rect 82645 765 82679 799
rect 89453 765 89487 799
rect 103345 765 103379 799
rect 103989 765 104023 799
rect 106381 765 106415 799
rect 109601 765 109635 799
rect 114937 765 114971 799
rect 117421 765 117455 799
rect 118341 765 118375 799
rect 5641 697 5675 731
rect 16773 697 16807 731
rect 17049 697 17083 731
rect 33333 697 33367 731
rect 38485 697 38519 731
rect 51917 697 51951 731
rect 52653 697 52687 731
rect 52929 697 52963 731
rect 68753 697 68787 731
rect 82185 697 82219 731
rect 87521 697 87555 731
rect 88993 697 89027 731
rect 112177 697 112211 731
rect 120549 697 120583 731
rect 122205 697 122239 731
rect 125701 697 125735 731
rect 131221 697 131255 731
rect 133889 833 133923 867
rect 135453 833 135487 867
rect 135821 833 135855 867
rect 167745 901 167779 935
rect 137661 833 137695 867
rect 138305 833 138339 867
rect 138857 833 138891 867
rect 140789 833 140823 867
rect 142069 833 142103 867
rect 143089 833 143123 867
rect 143549 833 143583 867
rect 146309 833 146343 867
rect 147045 833 147079 867
rect 151737 833 151771 867
rect 152473 833 152507 867
rect 158269 833 158303 867
rect 159005 833 159039 867
rect 159465 833 159499 867
rect 161029 833 161063 867
rect 161857 833 161891 867
rect 162041 833 162075 867
rect 163145 833 163179 867
rect 163881 833 163915 867
rect 164709 833 164743 867
rect 164985 833 165019 867
rect 166549 833 166583 867
rect 166641 833 166675 867
rect 134901 765 134935 799
rect 136373 765 136407 799
rect 136465 765 136499 799
rect 137753 697 137787 731
rect 10977 629 11011 663
rect 14197 629 14231 663
rect 18061 629 18095 663
rect 38025 629 38059 663
rect 53573 629 53607 663
rect 83289 629 83323 663
rect 84301 629 84335 663
rect 86141 629 86175 663
rect 104265 629 104299 663
rect 120917 629 120951 663
rect 121193 629 121227 663
rect 128369 629 128403 663
rect 128645 629 128679 663
rect 128829 629 128863 663
rect 131405 629 131439 663
rect 131681 629 131715 663
rect 132509 629 132543 663
rect 132969 629 133003 663
rect 133613 629 133647 663
rect 139225 765 139259 799
rect 140237 765 140271 799
rect 142537 765 142571 799
rect 144745 765 144779 799
rect 145205 765 145239 799
rect 147781 765 147815 799
rect 149529 765 149563 799
rect 150357 765 150391 799
rect 150633 765 150667 799
rect 156705 765 156739 799
rect 157717 765 157751 799
rect 160477 765 160511 799
rect 163053 765 163087 799
rect 165997 765 166031 799
rect 146493 697 146527 731
rect 151921 697 151955 731
rect 138857 629 138891 663
rect 142169 629 142203 663
rect 42441 425 42475 459
rect 50997 425 51031 459
rect 36461 85 36495 119
rect 36645 85 36679 119
rect 41061 85 41095 119
rect 42165 85 42199 119
rect 42257 85 42291 119
rect 111349 289 111383 323
rect 49893 17 49927 51
rect 111257 85 111291 119
rect 111349 85 111383 119
rect 111441 289 111475 323
rect 134165 289 134199 323
rect 134165 85 134199 119
<< metal1 >>
rect 23385 12971 23443 12977
rect 23385 12937 23397 12971
rect 23431 12968 23443 12971
rect 50890 12968 50896 12980
rect 23431 12940 50896 12968
rect 23431 12937 23443 12940
rect 23385 12931 23443 12937
rect 50890 12928 50896 12940
rect 50948 12928 50954 12980
rect 55217 12971 55275 12977
rect 55217 12937 55229 12971
rect 55263 12968 55275 12971
rect 56413 12971 56471 12977
rect 56413 12968 56425 12971
rect 55263 12940 56425 12968
rect 55263 12937 55275 12940
rect 55217 12931 55275 12937
rect 56413 12937 56425 12940
rect 56459 12937 56471 12971
rect 56413 12931 56471 12937
rect 56502 12928 56508 12980
rect 56560 12968 56566 12980
rect 66070 12968 66076 12980
rect 56560 12940 66076 12968
rect 56560 12928 56566 12940
rect 66070 12928 66076 12940
rect 66128 12928 66134 12980
rect 32214 12860 32220 12912
rect 32272 12900 32278 12912
rect 35894 12900 35900 12912
rect 32272 12872 35900 12900
rect 32272 12860 32278 12872
rect 35894 12860 35900 12872
rect 35952 12860 35958 12912
rect 35986 12860 35992 12912
rect 36044 12900 36050 12912
rect 36044 12872 46152 12900
rect 36044 12860 36050 12872
rect 30837 12835 30895 12841
rect 30837 12801 30849 12835
rect 30883 12832 30895 12835
rect 41322 12832 41328 12844
rect 30883 12804 41328 12832
rect 30883 12801 30895 12804
rect 30837 12795 30895 12801
rect 41322 12792 41328 12804
rect 41380 12792 41386 12844
rect 41509 12835 41567 12841
rect 41509 12801 41521 12835
rect 41555 12832 41567 12835
rect 46124 12832 46152 12872
rect 46290 12860 46296 12912
rect 46348 12900 46354 12912
rect 70854 12900 70860 12912
rect 46348 12872 70860 12900
rect 46348 12860 46354 12872
rect 70854 12860 70860 12872
rect 70912 12860 70918 12912
rect 55217 12835 55275 12841
rect 55217 12832 55229 12835
rect 41555 12804 46060 12832
rect 46124 12804 55229 12832
rect 41555 12801 41567 12804
rect 41509 12795 41567 12801
rect 22370 12724 22376 12776
rect 22428 12764 22434 12776
rect 32401 12767 32459 12773
rect 32401 12764 32413 12767
rect 22428 12736 32413 12764
rect 22428 12724 22434 12736
rect 32401 12733 32413 12736
rect 32447 12733 32459 12767
rect 32401 12727 32459 12733
rect 32493 12767 32551 12773
rect 32493 12733 32505 12767
rect 32539 12764 32551 12767
rect 39853 12767 39911 12773
rect 39853 12764 39865 12767
rect 32539 12736 39865 12764
rect 32539 12733 32551 12736
rect 32493 12727 32551 12733
rect 39853 12733 39865 12736
rect 39899 12733 39911 12767
rect 39853 12727 39911 12733
rect 40402 12724 40408 12776
rect 40460 12764 40466 12776
rect 41417 12767 41475 12773
rect 41417 12764 41429 12767
rect 40460 12736 41429 12764
rect 40460 12724 40466 12736
rect 41417 12733 41429 12736
rect 41463 12733 41475 12767
rect 45922 12764 45928 12776
rect 41417 12727 41475 12733
rect 41524 12736 45928 12764
rect 24305 12699 24363 12705
rect 24305 12665 24317 12699
rect 24351 12696 24363 12699
rect 41524 12696 41552 12736
rect 45922 12724 45928 12736
rect 45980 12724 45986 12776
rect 46032 12764 46060 12804
rect 55217 12801 55229 12804
rect 55263 12801 55275 12835
rect 55217 12795 55275 12801
rect 46293 12767 46351 12773
rect 46293 12764 46305 12767
rect 46032 12736 46305 12764
rect 46293 12733 46305 12736
rect 46339 12733 46351 12767
rect 46293 12727 46351 12733
rect 46474 12724 46480 12776
rect 46532 12764 46538 12776
rect 56413 12767 56471 12773
rect 46532 12736 55904 12764
rect 46532 12724 46538 12736
rect 24351 12668 41552 12696
rect 41601 12699 41659 12705
rect 24351 12665 24363 12668
rect 24305 12659 24363 12665
rect 41601 12665 41613 12699
rect 41647 12696 41659 12699
rect 55769 12699 55827 12705
rect 55769 12696 55781 12699
rect 41647 12668 55781 12696
rect 41647 12665 41659 12668
rect 41601 12659 41659 12665
rect 55769 12665 55781 12668
rect 55815 12665 55827 12699
rect 55876 12696 55904 12736
rect 56413 12733 56425 12767
rect 56459 12764 56471 12767
rect 57885 12767 57943 12773
rect 57885 12764 57897 12767
rect 56459 12736 57897 12764
rect 56459 12733 56471 12736
rect 56413 12727 56471 12733
rect 57885 12733 57897 12736
rect 57931 12733 57943 12767
rect 57885 12727 57943 12733
rect 58069 12767 58127 12773
rect 58069 12733 58081 12767
rect 58115 12764 58127 12767
rect 67637 12767 67695 12773
rect 67637 12764 67649 12767
rect 58115 12736 67649 12764
rect 58115 12733 58127 12736
rect 58069 12727 58127 12733
rect 67637 12733 67649 12736
rect 67683 12733 67695 12767
rect 67637 12727 67695 12733
rect 67729 12767 67787 12773
rect 67729 12733 67741 12767
rect 67775 12764 67787 12767
rect 77941 12767 77999 12773
rect 77941 12764 77953 12767
rect 67775 12736 77953 12764
rect 67775 12733 67787 12736
rect 67729 12727 67787 12733
rect 77941 12733 77953 12736
rect 77987 12733 77999 12767
rect 77941 12727 77999 12733
rect 83274 12696 83280 12708
rect 55876 12668 83280 12696
rect 55769 12659 55827 12665
rect 83274 12656 83280 12668
rect 83332 12656 83338 12708
rect 26234 12588 26240 12640
rect 26292 12628 26298 12640
rect 41690 12628 41696 12640
rect 26292 12600 41696 12628
rect 26292 12588 26298 12600
rect 41690 12588 41696 12600
rect 41748 12588 41754 12640
rect 41782 12588 41788 12640
rect 41840 12628 41846 12640
rect 50893 12631 50951 12637
rect 50893 12628 50905 12631
rect 41840 12600 50905 12628
rect 41840 12588 41846 12600
rect 50893 12597 50905 12600
rect 50939 12597 50951 12631
rect 50893 12591 50951 12597
rect 55953 12631 56011 12637
rect 55953 12597 55965 12631
rect 55999 12628 56011 12631
rect 66346 12628 66352 12640
rect 55999 12600 66352 12628
rect 55999 12597 56011 12600
rect 55953 12591 56011 12597
rect 66346 12588 66352 12600
rect 66404 12588 66410 12640
rect 98178 12588 98184 12640
rect 98236 12628 98242 12640
rect 121638 12628 121644 12640
rect 98236 12600 121644 12628
rect 98236 12588 98242 12600
rect 121638 12588 121644 12600
rect 121696 12588 121702 12640
rect 23290 12520 23296 12572
rect 23348 12560 23354 12572
rect 38010 12560 38016 12572
rect 23348 12532 38016 12560
rect 23348 12520 23354 12532
rect 38010 12520 38016 12532
rect 38068 12520 38074 12572
rect 38930 12520 38936 12572
rect 38988 12560 38994 12572
rect 40954 12560 40960 12572
rect 38988 12532 40960 12560
rect 38988 12520 38994 12532
rect 40954 12520 40960 12532
rect 41012 12520 41018 12572
rect 41046 12520 41052 12572
rect 41104 12560 41110 12572
rect 41417 12563 41475 12569
rect 41417 12560 41429 12563
rect 41104 12532 41429 12560
rect 41104 12520 41110 12532
rect 41417 12529 41429 12532
rect 41463 12529 41475 12563
rect 41417 12523 41475 12529
rect 41506 12520 41512 12572
rect 41564 12560 41570 12572
rect 55674 12560 55680 12572
rect 41564 12532 55680 12560
rect 41564 12520 41570 12532
rect 55674 12520 55680 12532
rect 55732 12520 55738 12572
rect 55769 12563 55827 12569
rect 55769 12529 55781 12563
rect 55815 12560 55827 12563
rect 61286 12560 61292 12572
rect 55815 12532 61292 12560
rect 55815 12529 55827 12532
rect 55769 12523 55827 12529
rect 61286 12520 61292 12532
rect 61344 12520 61350 12572
rect 109954 12520 109960 12572
rect 110012 12560 110018 12572
rect 123202 12560 123208 12572
rect 110012 12532 123208 12560
rect 110012 12520 110018 12532
rect 123202 12520 123208 12532
rect 123260 12520 123266 12572
rect 32401 12495 32459 12501
rect 32401 12461 32413 12495
rect 32447 12492 32459 12495
rect 36449 12495 36507 12501
rect 36449 12492 36461 12495
rect 32447 12464 36461 12492
rect 32447 12461 32459 12464
rect 32401 12455 32459 12461
rect 36449 12461 36461 12464
rect 36495 12461 36507 12495
rect 36449 12455 36507 12461
rect 36541 12495 36599 12501
rect 36541 12461 36553 12495
rect 36587 12492 36599 12495
rect 50706 12492 50712 12504
rect 36587 12464 50712 12492
rect 36587 12461 36599 12464
rect 36541 12455 36599 12461
rect 50706 12452 50712 12464
rect 50764 12452 50770 12504
rect 50893 12495 50951 12501
rect 50893 12461 50905 12495
rect 50939 12492 50951 12495
rect 56134 12492 56140 12504
rect 50939 12464 56140 12492
rect 50939 12461 50951 12464
rect 50893 12455 50951 12461
rect 56134 12452 56140 12464
rect 56192 12452 56198 12504
rect 56962 12452 56968 12504
rect 57020 12492 57026 12504
rect 58345 12495 58403 12501
rect 58345 12492 58357 12495
rect 57020 12464 58357 12492
rect 57020 12452 57026 12464
rect 58345 12461 58357 12464
rect 58391 12461 58403 12495
rect 58345 12455 58403 12461
rect 59446 12452 59452 12504
rect 59504 12492 59510 12504
rect 65705 12495 65763 12501
rect 65705 12492 65717 12495
rect 59504 12464 65717 12492
rect 59504 12452 59510 12464
rect 65705 12461 65717 12464
rect 65751 12461 65763 12495
rect 65705 12455 65763 12461
rect 96890 12452 96896 12504
rect 96948 12492 96954 12504
rect 121362 12492 121368 12504
rect 96948 12464 121368 12492
rect 96948 12452 96954 12464
rect 121362 12452 121368 12464
rect 121420 12452 121426 12504
rect 136634 12452 136640 12504
rect 136692 12492 136698 12504
rect 145098 12492 145104 12504
rect 136692 12464 145104 12492
rect 136692 12452 136698 12464
rect 145098 12452 145104 12464
rect 145156 12452 145162 12504
rect 28994 12384 29000 12436
rect 29052 12424 29058 12436
rect 32490 12424 32496 12436
rect 29052 12396 32496 12424
rect 29052 12384 29058 12396
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 32677 12427 32735 12433
rect 32677 12393 32689 12427
rect 32723 12424 32735 12427
rect 34422 12424 34428 12436
rect 32723 12396 34428 12424
rect 32723 12393 32735 12396
rect 32677 12387 32735 12393
rect 34422 12384 34428 12396
rect 34480 12384 34486 12436
rect 35618 12424 35624 12436
rect 35579 12396 35624 12424
rect 35618 12384 35624 12396
rect 35676 12384 35682 12436
rect 35713 12427 35771 12433
rect 35713 12393 35725 12427
rect 35759 12424 35771 12427
rect 82998 12424 83004 12436
rect 35759 12396 83004 12424
rect 35759 12393 35771 12396
rect 35713 12387 35771 12393
rect 82998 12384 83004 12396
rect 83056 12384 83062 12436
rect 110506 12384 110512 12436
rect 110564 12424 110570 12436
rect 123478 12424 123484 12436
rect 110564 12396 123484 12424
rect 110564 12384 110570 12396
rect 123478 12384 123484 12396
rect 123536 12384 123542 12436
rect 137002 12384 137008 12436
rect 137060 12424 137066 12436
rect 152458 12424 152464 12436
rect 137060 12396 152464 12424
rect 137060 12384 137066 12396
rect 152458 12384 152464 12396
rect 152516 12384 152522 12436
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 32309 12359 32367 12365
rect 32309 12356 32321 12359
rect 11572 12328 32321 12356
rect 11572 12316 11578 12328
rect 32309 12325 32321 12328
rect 32355 12325 32367 12359
rect 32309 12319 32367 12325
rect 32585 12359 32643 12365
rect 32585 12325 32597 12359
rect 32631 12356 32643 12359
rect 74994 12356 75000 12368
rect 32631 12328 75000 12356
rect 32631 12325 32643 12328
rect 32585 12319 32643 12325
rect 74994 12316 75000 12328
rect 75052 12316 75058 12368
rect 144730 12316 144736 12368
rect 144788 12356 144794 12368
rect 163866 12356 163872 12368
rect 144788 12328 163872 12356
rect 144788 12316 144794 12328
rect 163866 12316 163872 12328
rect 163924 12316 163930 12368
rect 24578 12248 24584 12300
rect 24636 12288 24642 12300
rect 32401 12291 32459 12297
rect 32401 12288 32413 12291
rect 24636 12260 32413 12288
rect 24636 12248 24642 12260
rect 32401 12257 32413 12260
rect 32447 12257 32459 12291
rect 32401 12251 32459 12257
rect 32490 12248 32496 12300
rect 32548 12288 32554 12300
rect 36449 12291 36507 12297
rect 32548 12260 35848 12288
rect 32548 12248 32554 12260
rect 24486 12180 24492 12232
rect 24544 12220 24550 12232
rect 28442 12220 28448 12232
rect 24544 12192 28448 12220
rect 24544 12180 24550 12192
rect 28442 12180 28448 12192
rect 28500 12180 28506 12232
rect 29178 12180 29184 12232
rect 29236 12220 29242 12232
rect 35713 12223 35771 12229
rect 35713 12220 35725 12223
rect 29236 12192 35725 12220
rect 29236 12180 29242 12192
rect 35713 12189 35725 12192
rect 35759 12189 35771 12223
rect 35820 12220 35848 12260
rect 36449 12257 36461 12291
rect 36495 12288 36507 12291
rect 38378 12288 38384 12300
rect 36495 12260 38384 12288
rect 36495 12257 36507 12260
rect 36449 12251 36507 12257
rect 38378 12248 38384 12260
rect 38436 12248 38442 12300
rect 38562 12248 38568 12300
rect 38620 12288 38626 12300
rect 55953 12291 56011 12297
rect 55953 12288 55965 12291
rect 38620 12260 55965 12288
rect 38620 12248 38626 12260
rect 55953 12257 55965 12260
rect 55999 12257 56011 12291
rect 55953 12251 56011 12257
rect 56045 12291 56103 12297
rect 56045 12257 56057 12291
rect 56091 12288 56103 12291
rect 58250 12288 58256 12300
rect 56091 12260 58256 12288
rect 56091 12257 56103 12260
rect 56045 12251 56103 12257
rect 58250 12248 58256 12260
rect 58308 12248 58314 12300
rect 58345 12291 58403 12297
rect 58345 12257 58357 12291
rect 58391 12288 58403 12291
rect 67818 12288 67824 12300
rect 58391 12260 67824 12288
rect 58391 12257 58403 12260
rect 58345 12251 58403 12257
rect 67818 12248 67824 12260
rect 67876 12248 67882 12300
rect 72418 12248 72424 12300
rect 72476 12288 72482 12300
rect 83090 12288 83096 12300
rect 72476 12260 83096 12288
rect 72476 12248 72482 12260
rect 83090 12248 83096 12260
rect 83148 12248 83154 12300
rect 108482 12248 108488 12300
rect 108540 12288 108546 12300
rect 121270 12288 121276 12300
rect 108540 12260 121276 12288
rect 108540 12248 108546 12260
rect 121270 12248 121276 12260
rect 121328 12248 121334 12300
rect 121914 12248 121920 12300
rect 121972 12288 121978 12300
rect 126882 12288 126888 12300
rect 121972 12260 126888 12288
rect 121972 12248 121978 12260
rect 126882 12248 126888 12260
rect 126940 12248 126946 12300
rect 137370 12248 137376 12300
rect 137428 12288 137434 12300
rect 162946 12288 162952 12300
rect 137428 12260 162952 12288
rect 137428 12248 137434 12260
rect 162946 12248 162952 12260
rect 163004 12248 163010 12300
rect 53098 12220 53104 12232
rect 35820 12192 53104 12220
rect 35713 12183 35771 12189
rect 53098 12180 53104 12192
rect 53156 12180 53162 12232
rect 55398 12180 55404 12232
rect 55456 12220 55462 12232
rect 65610 12220 65616 12232
rect 55456 12192 65616 12220
rect 55456 12180 55462 12192
rect 65610 12180 65616 12192
rect 65668 12180 65674 12232
rect 65705 12223 65763 12229
rect 65705 12189 65717 12223
rect 65751 12220 65763 12223
rect 79042 12220 79048 12232
rect 65751 12192 79048 12220
rect 65751 12189 65763 12192
rect 65705 12183 65763 12189
rect 79042 12180 79048 12192
rect 79100 12180 79106 12232
rect 108022 12180 108028 12232
rect 108080 12220 108086 12232
rect 125137 12223 125195 12229
rect 125137 12220 125149 12223
rect 108080 12192 113404 12220
rect 108080 12180 108086 12192
rect 113376 12164 113404 12192
rect 119632 12192 125149 12220
rect 119632 12164 119660 12192
rect 125137 12189 125149 12192
rect 125183 12189 125195 12223
rect 125137 12183 125195 12189
rect 125505 12223 125563 12229
rect 125505 12189 125517 12223
rect 125551 12220 125563 12223
rect 125594 12220 125600 12232
rect 125551 12192 125600 12220
rect 125551 12189 125563 12192
rect 125505 12183 125563 12189
rect 125594 12180 125600 12192
rect 125652 12180 125658 12232
rect 137186 12220 137192 12232
rect 132880 12192 137192 12220
rect 132880 12164 132908 12192
rect 137186 12180 137192 12192
rect 137244 12180 137250 12232
rect 137830 12180 137836 12232
rect 137888 12220 137894 12232
rect 165890 12220 165896 12232
rect 137888 12192 165896 12220
rect 137888 12180 137894 12192
rect 165890 12180 165896 12192
rect 165948 12180 165954 12232
rect 4522 12112 4528 12164
rect 4580 12152 4586 12164
rect 27614 12152 27620 12164
rect 4580 12124 27620 12152
rect 4580 12112 4586 12124
rect 27614 12112 27620 12124
rect 27672 12112 27678 12164
rect 32490 12152 32496 12164
rect 32451 12124 32496 12152
rect 32490 12112 32496 12124
rect 32548 12112 32554 12164
rect 34054 12112 34060 12164
rect 34112 12152 34118 12164
rect 46198 12152 46204 12164
rect 34112 12124 46204 12152
rect 34112 12112 34118 12124
rect 46198 12112 46204 12124
rect 46256 12112 46262 12164
rect 46293 12155 46351 12161
rect 46293 12121 46305 12155
rect 46339 12152 46351 12155
rect 61194 12152 61200 12164
rect 46339 12124 61200 12152
rect 46339 12121 46351 12124
rect 46293 12115 46351 12121
rect 61194 12112 61200 12124
rect 61252 12112 61258 12164
rect 68002 12112 68008 12164
rect 68060 12152 68066 12164
rect 80422 12152 80428 12164
rect 68060 12124 80428 12152
rect 68060 12112 68066 12124
rect 80422 12112 80428 12124
rect 80480 12112 80486 12164
rect 103146 12112 103152 12164
rect 103204 12152 103210 12164
rect 111518 12152 111524 12164
rect 103204 12124 111524 12152
rect 103204 12112 103210 12124
rect 111518 12112 111524 12124
rect 111576 12112 111582 12164
rect 113358 12112 113364 12164
rect 113416 12112 113422 12164
rect 119614 12112 119620 12164
rect 119672 12112 119678 12164
rect 119982 12112 119988 12164
rect 120040 12152 120046 12164
rect 122837 12155 122895 12161
rect 120040 12124 122788 12152
rect 120040 12112 120046 12124
rect 23382 12084 23388 12096
rect 23343 12056 23388 12084
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 24210 12044 24216 12096
rect 24268 12084 24274 12096
rect 24305 12087 24363 12093
rect 24305 12084 24317 12087
rect 24268 12056 24317 12084
rect 24268 12044 24274 12056
rect 24305 12053 24317 12056
rect 24351 12053 24363 12087
rect 24305 12047 24363 12053
rect 26878 12044 26884 12096
rect 26936 12084 26942 12096
rect 27522 12084 27528 12096
rect 26936 12056 27528 12084
rect 26936 12044 26942 12056
rect 27522 12044 27528 12056
rect 27580 12044 27586 12096
rect 27890 12044 27896 12096
rect 27948 12084 27954 12096
rect 30650 12084 30656 12096
rect 27948 12056 30656 12084
rect 27948 12044 27954 12056
rect 30650 12044 30656 12056
rect 30708 12044 30714 12096
rect 30742 12044 30748 12096
rect 30800 12084 30806 12096
rect 30837 12087 30895 12093
rect 30837 12084 30849 12087
rect 30800 12056 30849 12084
rect 30800 12044 30806 12056
rect 30837 12053 30849 12056
rect 30883 12053 30895 12087
rect 30837 12047 30895 12053
rect 31938 12044 31944 12096
rect 31996 12084 32002 12096
rect 37090 12084 37096 12096
rect 31996 12056 37096 12084
rect 31996 12044 32002 12056
rect 37090 12044 37096 12056
rect 37148 12044 37154 12096
rect 37182 12044 37188 12096
rect 37240 12084 37246 12096
rect 39574 12084 39580 12096
rect 37240 12056 39580 12084
rect 37240 12044 37246 12056
rect 39574 12044 39580 12056
rect 39632 12044 39638 12096
rect 39853 12087 39911 12093
rect 39853 12053 39865 12087
rect 39899 12084 39911 12087
rect 55769 12087 55827 12093
rect 55769 12084 55781 12087
rect 39899 12056 55781 12084
rect 39899 12053 39911 12056
rect 39853 12047 39911 12053
rect 55769 12053 55781 12056
rect 55815 12053 55827 12087
rect 55769 12047 55827 12053
rect 55858 12044 55864 12096
rect 55916 12084 55922 12096
rect 64506 12084 64512 12096
rect 55916 12056 64512 12084
rect 55916 12044 55922 12056
rect 64506 12044 64512 12056
rect 64564 12044 64570 12096
rect 73614 12044 73620 12096
rect 73672 12084 73678 12096
rect 76834 12084 76840 12096
rect 73672 12056 76840 12084
rect 73672 12044 73678 12056
rect 76834 12044 76840 12056
rect 76892 12044 76898 12096
rect 77938 12084 77944 12096
rect 77899 12056 77944 12084
rect 77938 12044 77944 12056
rect 77996 12044 78002 12096
rect 80238 12044 80244 12096
rect 80296 12084 80302 12096
rect 82906 12084 82912 12096
rect 80296 12056 82912 12084
rect 80296 12044 80302 12056
rect 82906 12044 82912 12056
rect 82964 12044 82970 12096
rect 101398 12044 101404 12096
rect 101456 12084 101462 12096
rect 118326 12084 118332 12096
rect 101456 12056 118332 12084
rect 101456 12044 101462 12056
rect 118326 12044 118332 12056
rect 118384 12044 118390 12096
rect 118694 12044 118700 12096
rect 118752 12084 118758 12096
rect 122653 12087 122711 12093
rect 122653 12084 122665 12087
rect 118752 12056 122665 12084
rect 118752 12044 118758 12056
rect 122653 12053 122665 12056
rect 122699 12053 122711 12087
rect 122760 12084 122788 12124
rect 122837 12121 122849 12155
rect 122883 12152 122895 12155
rect 127894 12152 127900 12164
rect 122883 12124 127900 12152
rect 122883 12121 122895 12124
rect 122837 12115 122895 12121
rect 127894 12112 127900 12124
rect 127952 12112 127958 12164
rect 132862 12112 132868 12164
rect 132920 12112 132926 12164
rect 134334 12112 134340 12164
rect 134392 12152 134398 12164
rect 146754 12152 146760 12164
rect 134392 12124 146760 12152
rect 134392 12112 134398 12124
rect 146754 12112 146760 12124
rect 146812 12112 146818 12164
rect 149054 12112 149060 12164
rect 149112 12152 149118 12164
rect 153286 12152 153292 12164
rect 149112 12124 153292 12152
rect 149112 12112 149118 12124
rect 153286 12112 153292 12124
rect 153344 12112 153350 12164
rect 135254 12084 135260 12096
rect 122760 12056 135260 12084
rect 122653 12047 122711 12053
rect 135254 12044 135260 12056
rect 135312 12044 135318 12096
rect 135438 12044 135444 12096
rect 135496 12084 135502 12096
rect 160370 12084 160376 12096
rect 135496 12056 160376 12084
rect 135496 12044 135502 12056
rect 160370 12044 160376 12056
rect 160428 12044 160434 12096
rect 368 11994 169556 12016
rect 368 11942 56667 11994
rect 56719 11942 56731 11994
rect 56783 11942 56795 11994
rect 56847 11942 56859 11994
rect 56911 11942 113088 11994
rect 113140 11942 113152 11994
rect 113204 11942 113216 11994
rect 113268 11942 113280 11994
rect 113332 11942 169556 11994
rect 368 11920 169556 11942
rect 29086 11880 29092 11892
rect 19260 11852 24716 11880
rect 5077 11815 5135 11821
rect 5077 11781 5089 11815
rect 5123 11812 5135 11815
rect 9674 11812 9680 11824
rect 5123 11784 9680 11812
rect 5123 11781 5135 11784
rect 5077 11775 5135 11781
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 19260 11812 19288 11852
rect 14516 11784 19288 11812
rect 14516 11772 14522 11784
rect 4798 11744 4804 11756
rect 4759 11716 4804 11744
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 8018 11744 8024 11756
rect 7791 11716 8024 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 22370 11744 22376 11756
rect 20772 11716 21864 11744
rect 22331 11716 22376 11744
rect 20772 11704 20778 11716
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 6181 11679 6239 11685
rect 6181 11676 6193 11679
rect 3375 11648 6193 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 6181 11645 6193 11648
rect 6227 11676 6239 11679
rect 6270 11676 6276 11688
rect 6227 11648 6276 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 14458 11676 14464 11688
rect 9732 11648 14464 11676
rect 9732 11636 9738 11648
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 19245 11679 19303 11685
rect 19245 11645 19257 11679
rect 19291 11676 19303 11679
rect 20162 11676 20168 11688
rect 19291 11648 20168 11676
rect 19291 11645 19303 11648
rect 19245 11639 19303 11645
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20806 11676 20812 11688
rect 20767 11648 20812 11676
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 21836 11685 21864 11716
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 24029 11747 24087 11753
rect 24029 11713 24041 11747
rect 24075 11744 24087 11747
rect 24578 11744 24584 11756
rect 24075 11716 24584 11744
rect 24075 11713 24087 11716
rect 24029 11707 24087 11713
rect 24578 11704 24584 11716
rect 24636 11704 24642 11756
rect 21821 11679 21879 11685
rect 21821 11645 21833 11679
rect 21867 11645 21879 11679
rect 21821 11639 21879 11645
rect 24121 11679 24179 11685
rect 24121 11645 24133 11679
rect 24167 11645 24179 11679
rect 24688 11676 24716 11852
rect 26896 11852 29092 11880
rect 26896 11821 26924 11852
rect 29086 11840 29092 11852
rect 29144 11840 29150 11892
rect 32030 11840 32036 11892
rect 32088 11880 32094 11892
rect 32125 11883 32183 11889
rect 32125 11880 32137 11883
rect 32088 11852 32137 11880
rect 32088 11840 32094 11852
rect 32125 11849 32137 11852
rect 32171 11849 32183 11883
rect 41138 11880 41144 11892
rect 32125 11843 32183 11849
rect 33428 11852 41144 11880
rect 26881 11815 26939 11821
rect 26881 11781 26893 11815
rect 26927 11781 26939 11815
rect 29733 11815 29791 11821
rect 26881 11775 26939 11781
rect 28184 11784 29684 11812
rect 26602 11704 26608 11756
rect 26660 11744 26666 11756
rect 26789 11747 26847 11753
rect 26789 11744 26801 11747
rect 26660 11716 26801 11744
rect 26660 11704 26666 11716
rect 26789 11713 26801 11716
rect 26835 11744 26847 11747
rect 28184 11744 28212 11784
rect 26835 11716 28212 11744
rect 26835 11713 26847 11716
rect 26789 11707 26847 11713
rect 28994 11704 29000 11756
rect 29052 11744 29058 11756
rect 29089 11747 29147 11753
rect 29089 11744 29101 11747
rect 29052 11716 29101 11744
rect 29052 11704 29058 11716
rect 29089 11713 29101 11716
rect 29135 11713 29147 11747
rect 29656 11744 29684 11784
rect 29733 11781 29745 11815
rect 29779 11812 29791 11815
rect 30926 11812 30932 11824
rect 29779 11784 30932 11812
rect 29779 11781 29791 11784
rect 29733 11775 29791 11781
rect 30926 11772 30932 11784
rect 30984 11772 30990 11824
rect 33428 11812 33456 11852
rect 41138 11840 41144 11852
rect 41196 11840 41202 11892
rect 41230 11840 41236 11892
rect 41288 11880 41294 11892
rect 42242 11880 42248 11892
rect 41288 11852 42248 11880
rect 41288 11840 41294 11852
rect 42242 11840 42248 11852
rect 42300 11840 42306 11892
rect 42426 11840 42432 11892
rect 42484 11880 42490 11892
rect 43806 11880 43812 11892
rect 42484 11852 43812 11880
rect 42484 11840 42490 11852
rect 43806 11840 43812 11852
rect 43864 11840 43870 11892
rect 46198 11840 46204 11892
rect 46256 11880 46262 11892
rect 55858 11880 55864 11892
rect 46256 11852 55864 11880
rect 46256 11840 46262 11852
rect 55858 11840 55864 11852
rect 55916 11840 55922 11892
rect 56689 11883 56747 11889
rect 56689 11849 56701 11883
rect 56735 11880 56747 11883
rect 60826 11880 60832 11892
rect 56735 11852 60832 11880
rect 56735 11849 56747 11852
rect 56689 11843 56747 11849
rect 60826 11840 60832 11852
rect 60884 11840 60890 11892
rect 63218 11880 63224 11892
rect 63179 11852 63224 11880
rect 63218 11840 63224 11852
rect 63276 11840 63282 11892
rect 70765 11883 70823 11889
rect 70765 11880 70777 11883
rect 65536 11852 70777 11880
rect 31036 11784 33456 11812
rect 31036 11744 31064 11784
rect 33502 11772 33508 11824
rect 33560 11812 33566 11824
rect 34701 11815 34759 11821
rect 34701 11812 34713 11815
rect 33560 11784 34713 11812
rect 33560 11772 33566 11784
rect 34701 11781 34713 11784
rect 34747 11781 34759 11815
rect 35805 11815 35863 11821
rect 35805 11812 35817 11815
rect 34701 11775 34759 11781
rect 35360 11784 35817 11812
rect 29656 11716 31064 11744
rect 32493 11747 32551 11753
rect 29089 11707 29147 11713
rect 32493 11713 32505 11747
rect 32539 11744 32551 11747
rect 32582 11744 32588 11756
rect 32539 11716 32588 11744
rect 32539 11713 32551 11716
rect 32493 11707 32551 11713
rect 27246 11676 27252 11688
rect 24688 11648 27252 11676
rect 24121 11639 24179 11645
rect 7653 11611 7711 11617
rect 7653 11577 7665 11611
rect 7699 11608 7711 11611
rect 17678 11608 17684 11620
rect 7699 11580 17684 11608
rect 7699 11577 7711 11580
rect 7653 11571 7711 11577
rect 17678 11568 17684 11580
rect 17736 11568 17742 11620
rect 24136 11608 24164 11639
rect 27246 11636 27252 11648
rect 27304 11636 27310 11688
rect 27338 11636 27344 11688
rect 27396 11676 27402 11688
rect 27709 11679 27767 11685
rect 27709 11676 27721 11679
rect 27396 11648 27721 11676
rect 27396 11636 27402 11648
rect 27709 11645 27721 11648
rect 27755 11645 27767 11679
rect 29104 11676 29132 11707
rect 32582 11704 32588 11716
rect 32640 11704 32646 11756
rect 35250 11744 35256 11756
rect 32692 11716 35256 11744
rect 29362 11676 29368 11688
rect 29104 11648 29368 11676
rect 27709 11639 27767 11645
rect 29362 11636 29368 11648
rect 29420 11636 29426 11688
rect 31570 11636 31576 11688
rect 31628 11676 31634 11688
rect 32692 11676 32720 11716
rect 35250 11704 35256 11716
rect 35308 11704 35314 11756
rect 35360 11753 35388 11784
rect 35805 11781 35817 11784
rect 35851 11812 35863 11815
rect 37182 11812 37188 11824
rect 35851 11784 37188 11812
rect 35851 11781 35863 11784
rect 35805 11775 35863 11781
rect 37182 11772 37188 11784
rect 37240 11772 37246 11824
rect 37553 11815 37611 11821
rect 37553 11812 37565 11815
rect 37476 11784 37565 11812
rect 35345 11747 35403 11753
rect 35345 11713 35357 11747
rect 35391 11713 35403 11747
rect 37476 11744 37504 11784
rect 37553 11781 37565 11784
rect 37599 11781 37611 11815
rect 37553 11775 37611 11781
rect 37660 11784 58204 11812
rect 37660 11744 37688 11784
rect 35345 11707 35403 11713
rect 36096 11716 37504 11744
rect 37568 11716 37688 11744
rect 38197 11747 38255 11753
rect 31628 11648 32720 11676
rect 31628 11636 31634 11648
rect 34238 11636 34244 11688
rect 34296 11676 34302 11688
rect 36096 11676 36124 11716
rect 34296 11648 36124 11676
rect 36265 11679 36323 11685
rect 34296 11636 34302 11648
rect 36265 11645 36277 11679
rect 36311 11676 36323 11679
rect 36998 11676 37004 11688
rect 36311 11648 37004 11676
rect 36311 11645 36323 11648
rect 36265 11639 36323 11645
rect 36998 11636 37004 11648
rect 37056 11636 37062 11688
rect 37182 11636 37188 11688
rect 37240 11676 37246 11688
rect 37568 11676 37596 11716
rect 38197 11713 38209 11747
rect 38243 11744 38255 11747
rect 38562 11744 38568 11756
rect 38243 11716 38568 11744
rect 38243 11713 38255 11716
rect 38197 11707 38255 11713
rect 38562 11704 38568 11716
rect 38620 11704 38626 11756
rect 39206 11704 39212 11756
rect 39264 11744 39270 11756
rect 39850 11744 39856 11756
rect 39264 11716 39856 11744
rect 39264 11704 39270 11716
rect 39850 11704 39856 11716
rect 39908 11704 39914 11756
rect 40770 11704 40776 11756
rect 40828 11744 40834 11756
rect 41046 11744 41052 11756
rect 40828 11716 41052 11744
rect 40828 11704 40834 11716
rect 41046 11704 41052 11716
rect 41104 11704 41110 11756
rect 41138 11704 41144 11756
rect 41196 11744 41202 11756
rect 41782 11744 41788 11756
rect 41196 11716 41788 11744
rect 41196 11704 41202 11716
rect 41782 11704 41788 11716
rect 41840 11704 41846 11756
rect 46109 11747 46167 11753
rect 46109 11744 46121 11747
rect 41892 11716 46121 11744
rect 37240 11648 37596 11676
rect 37240 11636 37246 11648
rect 37642 11636 37648 11688
rect 37700 11676 37706 11688
rect 41892 11676 41920 11716
rect 46109 11713 46121 11716
rect 46155 11713 46167 11747
rect 46109 11707 46167 11713
rect 46753 11747 46811 11753
rect 46753 11713 46765 11747
rect 46799 11744 46811 11747
rect 47118 11744 47124 11756
rect 46799 11716 47124 11744
rect 46799 11713 46811 11716
rect 46753 11707 46811 11713
rect 47118 11704 47124 11716
rect 47176 11704 47182 11756
rect 47673 11747 47731 11753
rect 47673 11713 47685 11747
rect 47719 11744 47731 11747
rect 48961 11747 49019 11753
rect 48961 11744 48973 11747
rect 47719 11716 48973 11744
rect 47719 11713 47731 11716
rect 47673 11707 47731 11713
rect 48961 11713 48973 11716
rect 49007 11744 49019 11747
rect 49142 11744 49148 11756
rect 49007 11716 49148 11744
rect 49007 11713 49019 11716
rect 48961 11707 49019 11713
rect 49142 11704 49148 11716
rect 49200 11704 49206 11756
rect 49602 11744 49608 11756
rect 49563 11716 49608 11744
rect 49602 11704 49608 11716
rect 49660 11704 49666 11756
rect 49786 11704 49792 11756
rect 49844 11744 49850 11756
rect 52730 11744 52736 11756
rect 49844 11716 52736 11744
rect 49844 11704 49850 11716
rect 52730 11704 52736 11716
rect 52788 11704 52794 11756
rect 53285 11747 53343 11753
rect 53285 11713 53297 11747
rect 53331 11744 53343 11747
rect 53466 11744 53472 11756
rect 53331 11716 53472 11744
rect 53331 11713 53343 11716
rect 53285 11707 53343 11713
rect 53466 11704 53472 11716
rect 53524 11704 53530 11756
rect 53745 11747 53803 11753
rect 53745 11713 53757 11747
rect 53791 11744 53803 11747
rect 54570 11744 54576 11756
rect 53791 11716 54576 11744
rect 53791 11713 53803 11716
rect 53745 11707 53803 11713
rect 54570 11704 54576 11716
rect 54628 11704 54634 11756
rect 56137 11747 56195 11753
rect 56137 11713 56149 11747
rect 56183 11744 56195 11747
rect 56318 11744 56324 11756
rect 56183 11716 56324 11744
rect 56183 11713 56195 11716
rect 56137 11707 56195 11713
rect 56318 11704 56324 11716
rect 56376 11704 56382 11756
rect 56502 11744 56508 11756
rect 56463 11716 56508 11744
rect 56502 11704 56508 11716
rect 56560 11704 56566 11756
rect 56870 11704 56876 11756
rect 56928 11744 56934 11756
rect 57422 11744 57428 11756
rect 56928 11716 57428 11744
rect 56928 11704 56934 11716
rect 57422 11704 57428 11716
rect 57480 11704 57486 11756
rect 57790 11744 57796 11756
rect 57751 11716 57796 11744
rect 57790 11704 57796 11716
rect 57848 11704 57854 11756
rect 58066 11744 58072 11756
rect 58027 11716 58072 11744
rect 58066 11704 58072 11716
rect 58124 11704 58130 11756
rect 58176 11744 58204 11784
rect 58250 11772 58256 11824
rect 58308 11812 58314 11824
rect 65536 11812 65564 11852
rect 70765 11849 70777 11852
rect 70811 11849 70823 11883
rect 70765 11843 70823 11849
rect 73893 11883 73951 11889
rect 73893 11849 73905 11883
rect 73939 11880 73951 11883
rect 74350 11880 74356 11892
rect 73939 11852 74356 11880
rect 73939 11849 73951 11852
rect 73893 11843 73951 11849
rect 58308 11784 65564 11812
rect 58308 11772 58314 11784
rect 65610 11772 65616 11824
rect 65668 11812 65674 11824
rect 73433 11815 73491 11821
rect 73433 11812 73445 11815
rect 65668 11784 73445 11812
rect 65668 11772 65674 11784
rect 73433 11781 73445 11784
rect 73479 11781 73491 11815
rect 73433 11775 73491 11781
rect 61378 11744 61384 11756
rect 58176 11716 61384 11744
rect 61378 11704 61384 11716
rect 61436 11704 61442 11756
rect 61473 11747 61531 11753
rect 61473 11713 61485 11747
rect 61519 11744 61531 11747
rect 61654 11744 61660 11756
rect 61519 11716 61660 11744
rect 61519 11713 61531 11716
rect 61473 11707 61531 11713
rect 61654 11704 61660 11716
rect 61712 11704 61718 11756
rect 61933 11747 61991 11753
rect 61933 11713 61945 11747
rect 61979 11744 61991 11747
rect 62482 11744 62488 11756
rect 61979 11716 62488 11744
rect 61979 11713 61991 11716
rect 61933 11707 61991 11713
rect 62482 11704 62488 11716
rect 62540 11704 62546 11756
rect 64690 11744 64696 11756
rect 64651 11716 64696 11744
rect 64690 11704 64696 11716
rect 64748 11704 64754 11756
rect 65150 11744 65156 11756
rect 65111 11716 65156 11744
rect 65150 11704 65156 11716
rect 65208 11704 65214 11756
rect 69201 11747 69259 11753
rect 69201 11713 69213 11747
rect 69247 11713 69259 11747
rect 69201 11707 69259 11713
rect 69661 11747 69719 11753
rect 69661 11713 69673 11747
rect 69707 11744 69719 11747
rect 70302 11744 70308 11756
rect 69707 11716 70308 11744
rect 69707 11713 69719 11716
rect 69661 11707 69719 11713
rect 37700 11648 41920 11676
rect 41969 11679 42027 11685
rect 37700 11636 37706 11648
rect 41969 11645 41981 11679
rect 42015 11676 42027 11679
rect 42058 11676 42064 11688
rect 42015 11648 42064 11676
rect 42015 11645 42027 11648
rect 41969 11639 42027 11645
rect 42058 11636 42064 11648
rect 42116 11636 42122 11688
rect 45925 11679 45983 11685
rect 45925 11645 45937 11679
rect 45971 11676 45983 11679
rect 46290 11676 46296 11688
rect 45971 11648 46296 11676
rect 45971 11645 45983 11648
rect 45925 11639 45983 11645
rect 46290 11636 46296 11648
rect 46348 11636 46354 11688
rect 46474 11636 46480 11688
rect 46532 11676 46538 11688
rect 49234 11676 49240 11688
rect 46532 11648 49240 11676
rect 46532 11636 46538 11648
rect 49234 11636 49240 11648
rect 49292 11636 49298 11688
rect 49329 11679 49387 11685
rect 49329 11645 49341 11679
rect 49375 11676 49387 11679
rect 49418 11676 49424 11688
rect 49375 11648 49424 11676
rect 49375 11645 49387 11648
rect 49329 11639 49387 11645
rect 49418 11636 49424 11648
rect 49476 11636 49482 11688
rect 49694 11636 49700 11688
rect 49752 11676 49758 11688
rect 50065 11679 50123 11685
rect 50065 11676 50077 11679
rect 49752 11648 50077 11676
rect 49752 11636 49758 11648
rect 50065 11645 50077 11648
rect 50111 11676 50123 11679
rect 50525 11679 50583 11685
rect 50525 11676 50537 11679
rect 50111 11648 50537 11676
rect 50111 11645 50123 11648
rect 50065 11639 50123 11645
rect 50525 11645 50537 11648
rect 50571 11645 50583 11679
rect 50525 11639 50583 11645
rect 50706 11636 50712 11688
rect 50764 11676 50770 11688
rect 51166 11676 51172 11688
rect 50764 11648 51172 11676
rect 50764 11636 50770 11648
rect 51166 11636 51172 11648
rect 51224 11636 51230 11688
rect 51810 11676 51816 11688
rect 51771 11648 51816 11676
rect 51810 11636 51816 11648
rect 51868 11636 51874 11688
rect 54849 11679 54907 11685
rect 54849 11645 54861 11679
rect 54895 11676 54907 11679
rect 54938 11676 54944 11688
rect 54895 11648 54944 11676
rect 54895 11645 54907 11648
rect 54849 11639 54907 11645
rect 54938 11636 54944 11648
rect 54996 11636 55002 11688
rect 55122 11636 55128 11688
rect 55180 11676 55186 11688
rect 55401 11679 55459 11685
rect 55401 11676 55413 11679
rect 55180 11648 55413 11676
rect 55180 11636 55186 11648
rect 55401 11645 55413 11648
rect 55447 11676 55459 11679
rect 56689 11679 56747 11685
rect 56689 11676 56701 11679
rect 55447 11648 56701 11676
rect 55447 11645 55459 11648
rect 55401 11639 55459 11645
rect 56689 11645 56701 11648
rect 56735 11645 56747 11679
rect 56689 11639 56747 11645
rect 56778 11636 56784 11688
rect 56836 11676 56842 11688
rect 56965 11679 57023 11685
rect 56965 11676 56977 11679
rect 56836 11648 56977 11676
rect 56836 11636 56842 11648
rect 56965 11645 56977 11648
rect 57011 11676 57023 11679
rect 59081 11679 59139 11685
rect 59081 11676 59093 11679
rect 57011 11648 59093 11676
rect 57011 11645 57023 11648
rect 56965 11639 57023 11645
rect 59081 11645 59093 11648
rect 59127 11645 59139 11679
rect 59081 11639 59139 11645
rect 60918 11636 60924 11688
rect 60976 11676 60982 11688
rect 65886 11676 65892 11688
rect 60976 11648 65892 11676
rect 60976 11636 60982 11648
rect 65886 11636 65892 11648
rect 65944 11636 65950 11688
rect 67818 11676 67824 11688
rect 67779 11648 67824 11676
rect 67818 11636 67824 11648
rect 67876 11636 67882 11688
rect 67910 11636 67916 11688
rect 67968 11676 67974 11688
rect 69216 11676 69244 11707
rect 70302 11704 70308 11716
rect 70360 11704 70366 11756
rect 71682 11704 71688 11756
rect 71740 11744 71746 11756
rect 71777 11747 71835 11753
rect 71777 11744 71789 11747
rect 71740 11716 71789 11744
rect 71740 11704 71746 11716
rect 71777 11713 71789 11716
rect 71823 11713 71835 11747
rect 71777 11707 71835 11713
rect 71866 11704 71872 11756
rect 71924 11744 71930 11756
rect 72326 11744 72332 11756
rect 71924 11716 72332 11744
rect 71924 11704 71930 11716
rect 72326 11704 72332 11716
rect 72384 11704 72390 11756
rect 73341 11747 73399 11753
rect 73341 11713 73353 11747
rect 73387 11744 73399 11747
rect 73908 11744 73936 11843
rect 74350 11840 74356 11852
rect 74408 11840 74414 11892
rect 74442 11840 74448 11892
rect 74500 11880 74506 11892
rect 79042 11880 79048 11892
rect 74500 11852 77616 11880
rect 79003 11852 79048 11880
rect 74500 11840 74506 11852
rect 75822 11772 75828 11824
rect 75880 11812 75886 11824
rect 77588 11812 77616 11852
rect 79042 11840 79048 11852
rect 79100 11840 79106 11892
rect 83274 11880 83280 11892
rect 83235 11852 83280 11880
rect 83274 11840 83280 11852
rect 83332 11840 83338 11892
rect 108206 11840 108212 11892
rect 108264 11880 108270 11892
rect 108301 11883 108359 11889
rect 108301 11880 108313 11883
rect 108264 11852 108313 11880
rect 108264 11840 108270 11852
rect 108301 11849 108313 11852
rect 108347 11880 108359 11883
rect 108482 11880 108488 11892
rect 108347 11852 108488 11880
rect 108347 11849 108359 11852
rect 108301 11843 108359 11849
rect 108482 11840 108488 11852
rect 108540 11840 108546 11892
rect 108942 11840 108948 11892
rect 109000 11880 109006 11892
rect 118694 11880 118700 11892
rect 109000 11852 118700 11880
rect 109000 11840 109006 11852
rect 118694 11840 118700 11852
rect 118752 11840 118758 11892
rect 118786 11840 118792 11892
rect 118844 11880 118850 11892
rect 124030 11880 124036 11892
rect 118844 11852 124036 11880
rect 118844 11840 118850 11852
rect 124030 11840 124036 11852
rect 124088 11840 124094 11892
rect 125594 11840 125600 11892
rect 125652 11880 125658 11892
rect 132678 11880 132684 11892
rect 125652 11852 132684 11880
rect 125652 11840 125658 11852
rect 132678 11840 132684 11852
rect 132736 11840 132742 11892
rect 134702 11840 134708 11892
rect 134760 11880 134766 11892
rect 148597 11883 148655 11889
rect 148597 11880 148609 11883
rect 134760 11852 148609 11880
rect 134760 11840 134766 11852
rect 148597 11849 148609 11852
rect 148643 11849 148655 11883
rect 148597 11843 148655 11849
rect 152458 11840 152464 11892
rect 152516 11880 152522 11892
rect 152516 11852 160140 11880
rect 152516 11840 152522 11852
rect 75880 11784 77524 11812
rect 77588 11784 79088 11812
rect 75880 11772 75886 11784
rect 74810 11744 74816 11756
rect 73387 11716 73936 11744
rect 74771 11716 74816 11744
rect 73387 11713 73399 11716
rect 73341 11707 73399 11713
rect 74810 11704 74816 11716
rect 74868 11704 74874 11756
rect 75181 11747 75239 11753
rect 75181 11713 75193 11747
rect 75227 11713 75239 11747
rect 75181 11707 75239 11713
rect 69937 11679 69995 11685
rect 69937 11676 69949 11679
rect 67968 11648 69949 11676
rect 67968 11636 67974 11648
rect 69937 11645 69949 11648
rect 69983 11645 69995 11679
rect 70486 11676 70492 11688
rect 70447 11648 70492 11676
rect 69937 11639 69995 11645
rect 70486 11636 70492 11648
rect 70544 11636 70550 11688
rect 70765 11679 70823 11685
rect 70765 11645 70777 11679
rect 70811 11676 70823 11679
rect 72145 11679 72203 11685
rect 72145 11676 72157 11679
rect 70811 11648 72157 11676
rect 70811 11645 70823 11648
rect 70765 11639 70823 11645
rect 72145 11645 72157 11648
rect 72191 11645 72203 11679
rect 72145 11639 72203 11645
rect 72878 11636 72884 11688
rect 72936 11676 72942 11688
rect 75196 11676 75224 11707
rect 75454 11704 75460 11756
rect 75512 11744 75518 11756
rect 77496 11753 77524 11784
rect 76193 11747 76251 11753
rect 76193 11744 76205 11747
rect 75512 11716 76205 11744
rect 75512 11704 75518 11716
rect 76193 11713 76205 11716
rect 76239 11744 76251 11747
rect 76653 11747 76711 11753
rect 76653 11744 76665 11747
rect 76239 11716 76665 11744
rect 76239 11713 76251 11716
rect 76193 11707 76251 11713
rect 76653 11713 76665 11716
rect 76699 11713 76711 11747
rect 76653 11707 76711 11713
rect 77481 11747 77539 11753
rect 77481 11713 77493 11747
rect 77527 11744 77539 11747
rect 77662 11744 77668 11756
rect 77527 11716 77668 11744
rect 77527 11713 77539 11716
rect 77481 11707 77539 11713
rect 77662 11704 77668 11716
rect 77720 11704 77726 11756
rect 78766 11704 78772 11756
rect 78824 11744 78830 11756
rect 78953 11747 79011 11753
rect 78953 11744 78965 11747
rect 78824 11716 78965 11744
rect 78824 11704 78830 11716
rect 78953 11713 78965 11716
rect 78999 11713 79011 11747
rect 79060 11744 79088 11784
rect 82170 11772 82176 11824
rect 82228 11812 82234 11824
rect 96890 11812 96896 11824
rect 82228 11784 84240 11812
rect 96851 11784 96896 11812
rect 82228 11772 82234 11784
rect 80974 11744 80980 11756
rect 79060 11716 80980 11744
rect 78953 11707 79011 11713
rect 80974 11704 80980 11716
rect 81032 11704 81038 11756
rect 82081 11747 82139 11753
rect 82081 11713 82093 11747
rect 82127 11713 82139 11747
rect 82081 11707 82139 11713
rect 75362 11676 75368 11688
rect 72936 11648 75368 11676
rect 72936 11636 72942 11648
rect 75362 11636 75368 11648
rect 75420 11636 75426 11688
rect 77570 11676 77576 11688
rect 77531 11648 77576 11676
rect 77570 11636 77576 11648
rect 77628 11636 77634 11688
rect 79505 11679 79563 11685
rect 79505 11645 79517 11679
rect 79551 11676 79563 11679
rect 80054 11676 80060 11688
rect 79551 11648 80060 11676
rect 79551 11645 79563 11648
rect 79505 11639 79563 11645
rect 80054 11636 80060 11648
rect 80112 11636 80118 11688
rect 80146 11636 80152 11688
rect 80204 11676 80210 11688
rect 80517 11679 80575 11685
rect 80517 11676 80529 11679
rect 80204 11648 80529 11676
rect 80204 11636 80210 11648
rect 80517 11645 80529 11648
rect 80563 11645 80575 11679
rect 80517 11639 80575 11645
rect 81529 11679 81587 11685
rect 81529 11645 81541 11679
rect 81575 11645 81587 11679
rect 81529 11639 81587 11645
rect 28350 11608 28356 11620
rect 24136 11580 28356 11608
rect 28350 11568 28356 11580
rect 28408 11568 28414 11620
rect 28442 11568 28448 11620
rect 28500 11608 28506 11620
rect 81544 11608 81572 11639
rect 81710 11636 81716 11688
rect 81768 11676 81774 11688
rect 82096 11676 82124 11707
rect 82538 11704 82544 11756
rect 82596 11744 82602 11756
rect 83185 11747 83243 11753
rect 83185 11744 83197 11747
rect 82596 11716 83197 11744
rect 82596 11704 82602 11716
rect 83185 11713 83197 11716
rect 83231 11744 83243 11747
rect 83366 11744 83372 11756
rect 83231 11716 83372 11744
rect 83231 11713 83243 11716
rect 83185 11707 83243 11713
rect 83366 11704 83372 11716
rect 83424 11704 83430 11756
rect 84212 11753 84240 11784
rect 96890 11772 96896 11784
rect 96948 11772 96954 11824
rect 112254 11812 112260 11824
rect 104636 11784 112260 11812
rect 84197 11747 84255 11753
rect 84197 11713 84209 11747
rect 84243 11744 84255 11747
rect 84746 11744 84752 11756
rect 84243 11716 84752 11744
rect 84243 11713 84255 11716
rect 84197 11707 84255 11713
rect 84746 11704 84752 11716
rect 84804 11704 84810 11756
rect 87138 11744 87144 11756
rect 87099 11716 87144 11744
rect 87138 11704 87144 11716
rect 87196 11704 87202 11756
rect 90637 11747 90695 11753
rect 90637 11713 90649 11747
rect 90683 11744 90695 11747
rect 92658 11744 92664 11756
rect 90683 11716 92664 11744
rect 90683 11713 90695 11716
rect 90637 11707 90695 11713
rect 92658 11704 92664 11716
rect 92716 11704 92722 11756
rect 93302 11744 93308 11756
rect 93263 11716 93308 11744
rect 93302 11704 93308 11716
rect 93360 11704 93366 11756
rect 96341 11747 96399 11753
rect 96341 11713 96353 11747
rect 96387 11744 96399 11747
rect 96908 11744 96936 11772
rect 98178 11744 98184 11756
rect 96387 11716 96936 11744
rect 98139 11716 98184 11744
rect 96387 11713 96399 11716
rect 96341 11707 96399 11713
rect 98178 11704 98184 11716
rect 98236 11704 98242 11756
rect 101033 11747 101091 11753
rect 101033 11713 101045 11747
rect 101079 11744 101091 11747
rect 103149 11747 103207 11753
rect 103149 11744 103161 11747
rect 101079 11716 103161 11744
rect 101079 11713 101091 11716
rect 101033 11707 101091 11713
rect 103149 11713 103161 11716
rect 103195 11744 103207 11747
rect 104066 11744 104072 11756
rect 103195 11716 104072 11744
rect 103195 11713 103207 11716
rect 103149 11707 103207 11713
rect 104066 11704 104072 11716
rect 104124 11704 104130 11756
rect 84289 11679 84347 11685
rect 84289 11676 84301 11679
rect 81768 11648 84301 11676
rect 81768 11636 81774 11648
rect 84289 11645 84301 11648
rect 84335 11645 84347 11679
rect 84289 11639 84347 11645
rect 86037 11679 86095 11685
rect 86037 11645 86049 11679
rect 86083 11676 86095 11679
rect 86954 11676 86960 11688
rect 86083 11648 86960 11676
rect 86083 11645 86095 11648
rect 86037 11639 86095 11645
rect 86954 11636 86960 11648
rect 87012 11636 87018 11688
rect 91738 11676 91744 11688
rect 91699 11648 91744 11676
rect 91738 11636 91744 11648
rect 91796 11636 91802 11688
rect 93118 11676 93124 11688
rect 93079 11648 93124 11676
rect 93118 11636 93124 11648
rect 93176 11636 93182 11688
rect 93670 11676 93676 11688
rect 93583 11648 93676 11676
rect 93670 11636 93676 11648
rect 93728 11676 93734 11688
rect 94593 11679 94651 11685
rect 94593 11676 94605 11679
rect 93728 11648 94605 11676
rect 93728 11636 93734 11648
rect 94593 11645 94605 11648
rect 94639 11645 94651 11679
rect 94593 11639 94651 11645
rect 99193 11679 99251 11685
rect 99193 11645 99205 11679
rect 99239 11676 99251 11679
rect 99466 11676 99472 11688
rect 99239 11648 99472 11676
rect 99239 11645 99251 11648
rect 99193 11639 99251 11645
rect 99466 11636 99472 11648
rect 99524 11676 99530 11688
rect 99653 11679 99711 11685
rect 99653 11676 99665 11679
rect 99524 11648 99665 11676
rect 99524 11636 99530 11648
rect 99653 11645 99665 11648
rect 99699 11645 99711 11679
rect 99653 11639 99711 11645
rect 101858 11636 101864 11688
rect 101916 11676 101922 11688
rect 104636 11685 104664 11784
rect 112254 11772 112260 11784
rect 112312 11772 112318 11824
rect 122190 11812 122196 11824
rect 112456 11784 122196 11812
rect 104713 11747 104771 11753
rect 104713 11713 104725 11747
rect 104759 11713 104771 11747
rect 104713 11707 104771 11713
rect 106645 11747 106703 11753
rect 106645 11713 106657 11747
rect 106691 11713 106703 11747
rect 107746 11744 107752 11756
rect 107707 11716 107752 11744
rect 106645 11707 106703 11713
rect 101953 11679 102011 11685
rect 101953 11676 101965 11679
rect 101916 11648 101965 11676
rect 101916 11636 101922 11648
rect 101953 11645 101965 11648
rect 101999 11676 102011 11679
rect 102045 11679 102103 11685
rect 102045 11676 102057 11679
rect 101999 11648 102057 11676
rect 101999 11645 102011 11648
rect 101953 11639 102011 11645
rect 102045 11645 102057 11648
rect 102091 11645 102103 11679
rect 102045 11639 102103 11645
rect 104621 11679 104679 11685
rect 104621 11645 104633 11679
rect 104667 11645 104679 11679
rect 104621 11639 104679 11645
rect 28500 11580 81572 11608
rect 28500 11568 28506 11580
rect 4154 11540 4160 11552
rect 4115 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 5813 11543 5871 11549
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 6086 11540 6092 11552
rect 5859 11512 6092 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 9585 11543 9643 11549
rect 9585 11509 9597 11543
rect 9631 11540 9643 11543
rect 9674 11540 9680 11552
rect 9631 11512 9680 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 17310 11540 17316 11552
rect 9824 11512 17316 11540
rect 9824 11500 9830 11512
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 20165 11543 20223 11549
rect 20165 11540 20177 11543
rect 20128 11512 20177 11540
rect 20128 11500 20134 11512
rect 20165 11509 20177 11512
rect 20211 11509 20223 11543
rect 20165 11503 20223 11509
rect 27062 11500 27068 11552
rect 27120 11540 27126 11552
rect 27249 11543 27307 11549
rect 27249 11540 27261 11543
rect 27120 11512 27261 11540
rect 27120 11500 27126 11512
rect 27249 11509 27261 11512
rect 27295 11540 27307 11543
rect 27430 11540 27436 11552
rect 27295 11512 27436 11540
rect 27295 11509 27307 11512
rect 27249 11503 27307 11509
rect 27430 11500 27436 11512
rect 27488 11500 27494 11552
rect 27522 11500 27528 11552
rect 27580 11540 27586 11552
rect 35526 11540 35532 11552
rect 27580 11512 35532 11540
rect 27580 11500 27586 11512
rect 35526 11500 35532 11512
rect 35584 11500 35590 11552
rect 35618 11500 35624 11552
rect 35676 11540 35682 11552
rect 40681 11543 40739 11549
rect 40681 11540 40693 11543
rect 35676 11512 40693 11540
rect 35676 11500 35682 11512
rect 40681 11509 40693 11512
rect 40727 11509 40739 11543
rect 40681 11503 40739 11509
rect 41322 11500 41328 11552
rect 41380 11540 41386 11552
rect 50154 11540 50160 11552
rect 41380 11512 50160 11540
rect 41380 11500 41386 11512
rect 50154 11500 50160 11512
rect 50212 11500 50218 11552
rect 50246 11500 50252 11552
rect 50304 11540 50310 11552
rect 52178 11540 52184 11552
rect 50304 11512 52184 11540
rect 50304 11500 50310 11512
rect 52178 11500 52184 11512
rect 52236 11500 52242 11552
rect 52454 11540 52460 11552
rect 52415 11512 52460 11540
rect 52454 11500 52460 11512
rect 52512 11500 52518 11552
rect 53098 11540 53104 11552
rect 53059 11512 53104 11540
rect 53098 11500 53104 11512
rect 53156 11500 53162 11552
rect 53190 11500 53196 11552
rect 53248 11540 53254 11552
rect 55953 11543 56011 11549
rect 55953 11540 55965 11543
rect 53248 11512 55965 11540
rect 53248 11500 53254 11512
rect 55953 11509 55965 11512
rect 55999 11509 56011 11543
rect 55953 11503 56011 11509
rect 56134 11500 56140 11552
rect 56192 11540 56198 11552
rect 57609 11543 57667 11549
rect 57609 11540 57621 11543
rect 56192 11512 57621 11540
rect 56192 11500 56198 11512
rect 57609 11509 57621 11512
rect 57655 11509 57667 11543
rect 59722 11540 59728 11552
rect 59635 11512 59728 11540
rect 57609 11503 57667 11509
rect 59722 11500 59728 11512
rect 59780 11540 59786 11552
rect 60642 11540 60648 11552
rect 59780 11512 60648 11540
rect 59780 11500 59786 11512
rect 60642 11500 60648 11512
rect 60700 11500 60706 11552
rect 61194 11500 61200 11552
rect 61252 11540 61258 11552
rect 61289 11543 61347 11549
rect 61289 11540 61301 11543
rect 61252 11512 61301 11540
rect 61252 11500 61258 11512
rect 61289 11509 61301 11512
rect 61335 11509 61347 11543
rect 64506 11540 64512 11552
rect 64467 11512 64512 11540
rect 61289 11503 61347 11509
rect 64506 11500 64512 11512
rect 64564 11500 64570 11552
rect 69014 11540 69020 11552
rect 68975 11512 69020 11540
rect 69014 11500 69020 11512
rect 69072 11500 69078 11552
rect 70578 11500 70584 11552
rect 70636 11540 70642 11552
rect 70949 11543 71007 11549
rect 70949 11540 70961 11543
rect 70636 11512 70961 11540
rect 70636 11500 70642 11512
rect 70949 11509 70961 11512
rect 70995 11509 71007 11543
rect 72786 11540 72792 11552
rect 72747 11512 72792 11540
rect 70949 11503 71007 11509
rect 72786 11500 72792 11512
rect 72844 11500 72850 11552
rect 74626 11500 74632 11552
rect 74684 11540 74690 11552
rect 74721 11543 74779 11549
rect 74721 11540 74733 11543
rect 74684 11512 74733 11540
rect 74684 11500 74690 11512
rect 74721 11509 74733 11512
rect 74767 11509 74779 11543
rect 76282 11540 76288 11552
rect 76243 11512 76288 11540
rect 74721 11503 74779 11509
rect 76282 11500 76288 11512
rect 76340 11500 76346 11552
rect 76742 11500 76748 11552
rect 76800 11540 76806 11552
rect 77021 11543 77079 11549
rect 77021 11540 77033 11543
rect 76800 11512 77033 11540
rect 76800 11500 76806 11512
rect 77021 11509 77033 11512
rect 77067 11509 77079 11543
rect 80146 11540 80152 11552
rect 80107 11512 80152 11540
rect 77021 11503 77079 11509
rect 80146 11500 80152 11512
rect 80204 11500 80210 11552
rect 87233 11543 87291 11549
rect 87233 11509 87245 11543
rect 87279 11540 87291 11543
rect 88334 11540 88340 11552
rect 87279 11512 88340 11540
rect 87279 11509 87291 11512
rect 87233 11503 87291 11509
rect 88334 11500 88340 11512
rect 88392 11500 88398 11552
rect 95510 11540 95516 11552
rect 95471 11512 95516 11540
rect 95510 11500 95516 11512
rect 95568 11500 95574 11552
rect 96433 11543 96491 11549
rect 96433 11509 96445 11543
rect 96479 11540 96491 11543
rect 96614 11540 96620 11552
rect 96479 11512 96620 11540
rect 96479 11509 96491 11512
rect 96433 11503 96491 11509
rect 96614 11500 96620 11512
rect 96672 11500 96678 11552
rect 98270 11540 98276 11552
rect 98231 11512 98276 11540
rect 98270 11500 98276 11512
rect 98328 11500 98334 11552
rect 104728 11540 104756 11707
rect 106550 11636 106556 11688
rect 106608 11676 106614 11688
rect 106660 11676 106688 11707
rect 107746 11704 107752 11716
rect 107804 11704 107810 11756
rect 109862 11744 109868 11756
rect 107856 11716 109868 11744
rect 107856 11676 107884 11716
rect 109862 11704 109868 11716
rect 109920 11704 109926 11756
rect 109954 11704 109960 11756
rect 110012 11744 110018 11756
rect 110049 11747 110107 11753
rect 110049 11744 110061 11747
rect 110012 11716 110061 11744
rect 110012 11704 110018 11716
rect 110049 11713 110061 11716
rect 110095 11713 110107 11747
rect 112456 11744 112484 11784
rect 122190 11772 122196 11784
rect 122248 11772 122254 11824
rect 124766 11812 124772 11824
rect 123128 11784 124772 11812
rect 123128 11756 123156 11784
rect 124766 11772 124772 11784
rect 124824 11772 124830 11824
rect 128446 11772 128452 11824
rect 128504 11812 128510 11824
rect 128504 11784 129872 11812
rect 128504 11772 128510 11784
rect 112990 11744 112996 11756
rect 110049 11707 110107 11713
rect 110156 11716 112484 11744
rect 112951 11716 112996 11744
rect 106608 11648 107884 11676
rect 108945 11679 109003 11685
rect 106608 11636 106614 11648
rect 108945 11645 108957 11679
rect 108991 11676 109003 11679
rect 109034 11676 109040 11688
rect 108991 11648 109040 11676
rect 108991 11645 109003 11648
rect 108945 11639 109003 11645
rect 109034 11636 109040 11648
rect 109092 11636 109098 11688
rect 104894 11568 104900 11620
rect 104952 11608 104958 11620
rect 110156 11608 110184 11716
rect 112990 11704 112996 11716
rect 113048 11704 113054 11756
rect 115566 11744 115572 11756
rect 113100 11716 115572 11744
rect 111702 11676 111708 11688
rect 111663 11648 111708 11676
rect 111702 11636 111708 11648
rect 111760 11636 111766 11688
rect 113100 11685 113128 11716
rect 115566 11704 115572 11716
rect 115624 11704 115630 11756
rect 116121 11747 116179 11753
rect 116121 11713 116133 11747
rect 116167 11744 116179 11747
rect 116486 11744 116492 11756
rect 116167 11716 116492 11744
rect 116167 11713 116179 11716
rect 116121 11707 116179 11713
rect 116486 11704 116492 11716
rect 116544 11704 116550 11756
rect 118237 11747 118295 11753
rect 118237 11713 118249 11747
rect 118283 11713 118295 11747
rect 118237 11707 118295 11713
rect 113085 11679 113143 11685
rect 113085 11645 113097 11679
rect 113131 11645 113143 11679
rect 113085 11639 113143 11645
rect 114557 11679 114615 11685
rect 114557 11645 114569 11679
rect 114603 11676 114615 11679
rect 114646 11676 114652 11688
rect 114603 11648 114652 11676
rect 114603 11645 114615 11648
rect 114557 11639 114615 11645
rect 114646 11636 114652 11648
rect 114704 11636 114710 11688
rect 115845 11679 115903 11685
rect 115845 11645 115857 11679
rect 115891 11676 115903 11679
rect 116302 11676 116308 11688
rect 115891 11648 116308 11676
rect 115891 11645 115903 11648
rect 115845 11639 115903 11645
rect 116302 11636 116308 11648
rect 116360 11636 116366 11688
rect 104952 11580 110184 11608
rect 110233 11611 110291 11617
rect 104952 11568 104958 11580
rect 110233 11577 110245 11611
rect 110279 11608 110291 11611
rect 114094 11608 114100 11620
rect 110279 11580 114100 11608
rect 110279 11577 110291 11580
rect 110233 11571 110291 11577
rect 114094 11568 114100 11580
rect 114152 11568 114158 11620
rect 118252 11608 118280 11707
rect 118326 11704 118332 11756
rect 118384 11744 118390 11756
rect 118384 11716 118429 11744
rect 118384 11704 118390 11716
rect 118878 11704 118884 11756
rect 118936 11744 118942 11756
rect 121825 11747 121883 11753
rect 118936 11716 121316 11744
rect 118936 11704 118942 11716
rect 120258 11676 120264 11688
rect 120219 11648 120264 11676
rect 120258 11636 120264 11648
rect 120316 11636 120322 11688
rect 121288 11685 121316 11716
rect 121825 11713 121837 11747
rect 121871 11744 121883 11747
rect 121914 11744 121920 11756
rect 121871 11716 121920 11744
rect 121871 11713 121883 11716
rect 121825 11707 121883 11713
rect 121914 11704 121920 11716
rect 121972 11704 121978 11756
rect 123110 11744 123116 11756
rect 123023 11716 123116 11744
rect 123110 11704 123116 11716
rect 123168 11704 123174 11756
rect 123202 11704 123208 11756
rect 123260 11744 123266 11756
rect 124125 11747 124183 11753
rect 123260 11716 123305 11744
rect 123260 11704 123266 11716
rect 124125 11713 124137 11747
rect 124171 11744 124183 11747
rect 124306 11744 124312 11756
rect 124171 11716 124312 11744
rect 124171 11713 124183 11716
rect 124125 11707 124183 11713
rect 124306 11704 124312 11716
rect 124364 11744 124370 11756
rect 125134 11744 125140 11756
rect 124364 11716 125140 11744
rect 124364 11704 124370 11716
rect 125134 11704 125140 11716
rect 125192 11704 125198 11756
rect 127897 11747 127955 11753
rect 127897 11713 127909 11747
rect 127943 11713 127955 11747
rect 127897 11707 127955 11713
rect 121273 11679 121331 11685
rect 121273 11645 121285 11679
rect 121319 11645 121331 11679
rect 124217 11679 124275 11685
rect 124217 11676 124229 11679
rect 121273 11639 121331 11645
rect 121472 11648 124229 11676
rect 118252 11580 118464 11608
rect 105262 11540 105268 11552
rect 104728 11512 105268 11540
rect 105262 11500 105268 11512
rect 105320 11540 105326 11552
rect 106737 11543 106795 11549
rect 106737 11540 106749 11543
rect 105320 11512 106749 11540
rect 105320 11500 105326 11512
rect 106737 11509 106749 11512
rect 106783 11509 106795 11543
rect 107102 11540 107108 11552
rect 107063 11512 107108 11540
rect 106737 11503 106795 11509
rect 107102 11500 107108 11512
rect 107160 11500 107166 11552
rect 107838 11540 107844 11552
rect 107799 11512 107844 11540
rect 107838 11500 107844 11512
rect 107896 11500 107902 11552
rect 109954 11500 109960 11552
rect 110012 11540 110018 11552
rect 110874 11540 110880 11552
rect 110012 11512 110880 11540
rect 110012 11500 110018 11512
rect 110874 11500 110880 11512
rect 110932 11500 110938 11552
rect 111242 11540 111248 11552
rect 111203 11512 111248 11540
rect 111242 11500 111248 11512
rect 111300 11500 111306 11552
rect 116486 11540 116492 11552
rect 116447 11512 116492 11540
rect 116486 11500 116492 11512
rect 116544 11500 116550 11552
rect 117958 11540 117964 11552
rect 117919 11512 117964 11540
rect 117958 11500 117964 11512
rect 118016 11500 118022 11552
rect 118436 11540 118464 11580
rect 118602 11568 118608 11620
rect 118660 11608 118666 11620
rect 121472 11608 121500 11648
rect 124217 11645 124229 11648
rect 124263 11645 124275 11679
rect 124217 11639 124275 11645
rect 126333 11679 126391 11685
rect 126333 11645 126345 11679
rect 126379 11676 126391 11679
rect 126974 11676 126980 11688
rect 126379 11648 126980 11676
rect 126379 11645 126391 11648
rect 126333 11639 126391 11645
rect 126974 11636 126980 11648
rect 127032 11636 127038 11688
rect 127345 11679 127403 11685
rect 127345 11645 127357 11679
rect 127391 11645 127403 11679
rect 127345 11639 127403 11645
rect 118660 11580 121500 11608
rect 118660 11568 118666 11580
rect 121730 11568 121736 11620
rect 121788 11608 121794 11620
rect 124398 11608 124404 11620
rect 121788 11580 124404 11608
rect 121788 11568 121794 11580
rect 124398 11568 124404 11580
rect 124456 11568 124462 11620
rect 127360 11608 127388 11639
rect 127710 11636 127716 11688
rect 127768 11676 127774 11688
rect 127912 11676 127940 11707
rect 128078 11704 128084 11756
rect 128136 11744 128142 11756
rect 129844 11753 129872 11784
rect 130654 11772 130660 11824
rect 130712 11812 130718 11824
rect 134981 11815 135039 11821
rect 134981 11812 134993 11815
rect 130712 11784 134993 11812
rect 130712 11772 130718 11784
rect 128817 11747 128875 11753
rect 128817 11744 128829 11747
rect 128136 11716 128829 11744
rect 128136 11704 128142 11716
rect 128817 11713 128829 11716
rect 128863 11744 128875 11747
rect 129277 11747 129335 11753
rect 129277 11744 129289 11747
rect 128863 11716 129289 11744
rect 128863 11713 128875 11716
rect 128817 11707 128875 11713
rect 129277 11713 129289 11716
rect 129323 11713 129335 11747
rect 129277 11707 129335 11713
rect 129829 11747 129887 11753
rect 129829 11713 129841 11747
rect 129875 11744 129887 11747
rect 130470 11744 130476 11756
rect 129875 11716 130476 11744
rect 129875 11713 129887 11716
rect 129829 11707 129887 11713
rect 130470 11704 130476 11716
rect 130528 11704 130534 11756
rect 131758 11704 131764 11756
rect 131816 11744 131822 11756
rect 133230 11744 133236 11756
rect 131816 11716 133000 11744
rect 133191 11716 133236 11744
rect 131816 11704 131822 11716
rect 129734 11676 129740 11688
rect 127768 11648 129740 11676
rect 127768 11636 127774 11648
rect 129734 11636 129740 11648
rect 129792 11636 129798 11688
rect 131669 11679 131727 11685
rect 131669 11645 131681 11679
rect 131715 11676 131727 11679
rect 132494 11676 132500 11688
rect 131715 11648 132500 11676
rect 131715 11645 131727 11648
rect 131669 11639 131727 11645
rect 132494 11636 132500 11648
rect 132552 11636 132558 11688
rect 132678 11676 132684 11688
rect 132639 11648 132684 11676
rect 132678 11636 132684 11648
rect 132736 11636 132742 11688
rect 132972 11676 133000 11716
rect 133230 11704 133236 11716
rect 133288 11704 133294 11756
rect 134536 11753 134564 11784
rect 134981 11781 134993 11784
rect 135027 11781 135039 11815
rect 134981 11775 135039 11781
rect 135070 11772 135076 11824
rect 135128 11812 135134 11824
rect 135128 11784 157380 11812
rect 135128 11772 135134 11784
rect 134521 11747 134579 11753
rect 134521 11713 134533 11747
rect 134567 11713 134579 11747
rect 134521 11707 134579 11713
rect 135533 11747 135591 11753
rect 135533 11713 135545 11747
rect 135579 11713 135591 11747
rect 135533 11707 135591 11713
rect 135548 11676 135576 11707
rect 137186 11704 137192 11756
rect 137244 11744 137250 11756
rect 137373 11747 137431 11753
rect 137373 11744 137385 11747
rect 137244 11716 137385 11744
rect 137244 11704 137250 11716
rect 137373 11713 137385 11716
rect 137419 11713 137431 11747
rect 138382 11744 138388 11756
rect 138343 11716 138388 11744
rect 137373 11707 137431 11713
rect 138382 11704 138388 11716
rect 138440 11704 138446 11756
rect 138477 11747 138535 11753
rect 138477 11713 138489 11747
rect 138523 11744 138535 11747
rect 141329 11747 141387 11753
rect 141329 11744 141341 11747
rect 138523 11716 141341 11744
rect 138523 11713 138535 11716
rect 138477 11707 138535 11713
rect 141329 11713 141341 11716
rect 141375 11744 141387 11747
rect 142065 11747 142123 11753
rect 142065 11744 142077 11747
rect 141375 11716 142077 11744
rect 141375 11713 141387 11716
rect 141329 11707 141387 11713
rect 142065 11713 142077 11716
rect 142111 11713 142123 11747
rect 142065 11707 142123 11713
rect 143350 11704 143356 11756
rect 143408 11744 143414 11756
rect 143537 11747 143595 11753
rect 143537 11744 143549 11747
rect 143408 11716 143549 11744
rect 143408 11704 143414 11716
rect 143537 11713 143549 11716
rect 143583 11713 143595 11747
rect 143537 11707 143595 11713
rect 143902 11704 143908 11756
rect 143960 11744 143966 11756
rect 144822 11744 144828 11756
rect 143960 11716 144828 11744
rect 143960 11704 143966 11716
rect 144822 11704 144828 11716
rect 144880 11704 144886 11756
rect 146754 11704 146760 11756
rect 146812 11744 146818 11756
rect 146849 11747 146907 11753
rect 146849 11744 146861 11747
rect 146812 11716 146861 11744
rect 146812 11704 146818 11716
rect 146849 11713 146861 11716
rect 146895 11744 146907 11747
rect 147309 11747 147367 11753
rect 147309 11744 147321 11747
rect 146895 11716 147321 11744
rect 146895 11713 146907 11716
rect 146849 11707 146907 11713
rect 147309 11713 147321 11716
rect 147355 11713 147367 11747
rect 147309 11707 147367 11713
rect 148597 11747 148655 11753
rect 148597 11713 148609 11747
rect 148643 11744 148655 11747
rect 150434 11744 150440 11756
rect 148643 11716 150440 11744
rect 148643 11713 148655 11716
rect 148597 11707 148655 11713
rect 150434 11704 150440 11716
rect 150492 11744 150498 11756
rect 150529 11747 150587 11753
rect 150529 11744 150541 11747
rect 150492 11716 150541 11744
rect 150492 11704 150498 11716
rect 150529 11713 150541 11716
rect 150575 11713 150587 11747
rect 150529 11707 150587 11713
rect 151446 11704 151452 11756
rect 151504 11744 151510 11756
rect 151633 11747 151691 11753
rect 151633 11744 151645 11747
rect 151504 11716 151645 11744
rect 151504 11704 151510 11716
rect 151633 11713 151645 11716
rect 151679 11713 151691 11747
rect 154482 11744 154488 11756
rect 154443 11716 154488 11744
rect 151633 11707 151691 11713
rect 154482 11704 154488 11716
rect 154540 11704 154546 11756
rect 157352 11753 157380 11784
rect 156225 11747 156283 11753
rect 156225 11744 156237 11747
rect 156156 11716 156237 11744
rect 136082 11676 136088 11688
rect 132972 11648 136088 11676
rect 136082 11636 136088 11648
rect 136140 11636 136146 11688
rect 138400 11676 138428 11704
rect 156156 11688 156184 11716
rect 156225 11713 156237 11716
rect 156271 11713 156283 11747
rect 156225 11707 156283 11713
rect 157337 11747 157395 11753
rect 157337 11713 157349 11747
rect 157383 11744 157395 11747
rect 157797 11747 157855 11753
rect 157797 11744 157809 11747
rect 157383 11716 157809 11744
rect 157383 11713 157395 11716
rect 157337 11707 157395 11713
rect 157797 11713 157809 11716
rect 157843 11713 157855 11747
rect 160112 11744 160140 11852
rect 160186 11744 160192 11756
rect 160099 11716 160192 11744
rect 157797 11707 157855 11713
rect 160186 11704 160192 11716
rect 160244 11704 160250 11756
rect 160370 11704 160376 11756
rect 160428 11744 160434 11756
rect 161937 11747 161995 11753
rect 161937 11744 161949 11747
rect 160428 11716 161949 11744
rect 160428 11704 160434 11716
rect 161937 11713 161949 11716
rect 161983 11744 161995 11747
rect 162210 11744 162216 11756
rect 161983 11716 162216 11744
rect 161983 11713 161995 11716
rect 161937 11707 161995 11713
rect 162210 11704 162216 11716
rect 162268 11704 162274 11756
rect 162946 11704 162952 11756
rect 163004 11744 163010 11756
rect 163041 11747 163099 11753
rect 163041 11744 163053 11747
rect 163004 11716 163053 11744
rect 163004 11704 163010 11716
rect 163041 11713 163053 11716
rect 163087 11744 163099 11747
rect 163501 11747 163559 11753
rect 163501 11744 163513 11747
rect 163087 11716 163513 11744
rect 163087 11713 163099 11716
rect 163041 11707 163099 11713
rect 163501 11713 163513 11716
rect 163547 11713 163559 11747
rect 165890 11744 165896 11756
rect 165851 11716 165896 11744
rect 163501 11707 163559 11713
rect 165890 11704 165896 11716
rect 165948 11704 165954 11756
rect 165985 11747 166043 11753
rect 165985 11713 165997 11747
rect 166031 11744 166043 11747
rect 167178 11744 167184 11756
rect 166031 11716 167184 11744
rect 166031 11713 166043 11716
rect 165985 11707 166043 11713
rect 167178 11704 167184 11716
rect 167236 11704 167242 11756
rect 138845 11679 138903 11685
rect 138845 11676 138857 11679
rect 138400 11648 138857 11676
rect 138845 11645 138857 11648
rect 138891 11645 138903 11679
rect 140222 11676 140228 11688
rect 140183 11648 140228 11676
rect 138845 11639 138903 11645
rect 140222 11636 140228 11648
rect 140280 11636 140286 11688
rect 140314 11636 140320 11688
rect 140372 11676 140378 11688
rect 141237 11679 141295 11685
rect 141237 11676 141249 11679
rect 140372 11648 141249 11676
rect 140372 11636 140378 11648
rect 141237 11645 141249 11648
rect 141283 11645 141295 11679
rect 144546 11676 144552 11688
rect 144507 11648 144552 11676
rect 141237 11639 141295 11645
rect 144546 11636 144552 11648
rect 144604 11636 144610 11688
rect 146478 11636 146484 11688
rect 146536 11676 146542 11688
rect 146573 11679 146631 11685
rect 146573 11676 146585 11679
rect 146536 11648 146585 11676
rect 146536 11636 146542 11648
rect 146573 11645 146585 11648
rect 146619 11676 146631 11679
rect 148781 11679 148839 11685
rect 148781 11676 148793 11679
rect 146619 11648 148793 11676
rect 146619 11645 146631 11648
rect 146573 11639 146631 11645
rect 148781 11645 148793 11648
rect 148827 11645 148839 11679
rect 156138 11676 156144 11688
rect 148781 11639 148839 11645
rect 150544 11648 156144 11676
rect 124508 11580 127388 11608
rect 129921 11611 129979 11617
rect 118786 11540 118792 11552
rect 118436 11512 118792 11540
rect 118786 11500 118792 11512
rect 118844 11500 118850 11552
rect 119246 11500 119252 11552
rect 119304 11540 119310 11552
rect 124508 11540 124536 11580
rect 129921 11577 129933 11611
rect 129967 11608 129979 11611
rect 130654 11608 130660 11620
rect 129967 11580 130660 11608
rect 129967 11577 129979 11580
rect 129921 11571 129979 11577
rect 130654 11568 130660 11580
rect 130712 11568 130718 11620
rect 134613 11611 134671 11617
rect 134613 11577 134625 11611
rect 134659 11608 134671 11611
rect 143629 11611 143687 11617
rect 134659 11580 136036 11608
rect 134659 11577 134671 11580
rect 134613 11571 134671 11577
rect 136008 11552 136036 11580
rect 143629 11577 143641 11611
rect 143675 11608 143687 11611
rect 144914 11608 144920 11620
rect 143675 11580 144920 11608
rect 143675 11577 143687 11580
rect 143629 11571 143687 11577
rect 144914 11568 144920 11580
rect 144972 11568 144978 11620
rect 145098 11568 145104 11620
rect 145156 11608 145162 11620
rect 150544 11608 150572 11648
rect 156138 11636 156144 11648
rect 156196 11636 156202 11688
rect 156874 11636 156880 11688
rect 156932 11676 156938 11688
rect 156969 11679 157027 11685
rect 156969 11676 156981 11679
rect 156932 11648 156981 11676
rect 156932 11636 156938 11648
rect 156969 11645 156981 11648
rect 157015 11676 157027 11679
rect 158349 11679 158407 11685
rect 158349 11676 158361 11679
rect 157015 11648 158361 11676
rect 157015 11645 157027 11648
rect 156969 11639 157027 11645
rect 158349 11645 158361 11648
rect 158395 11645 158407 11679
rect 158349 11639 158407 11645
rect 164789 11679 164847 11685
rect 164789 11645 164801 11679
rect 164835 11676 164847 11679
rect 166074 11676 166080 11688
rect 164835 11648 166080 11676
rect 164835 11645 164847 11648
rect 164789 11639 164847 11645
rect 166074 11636 166080 11648
rect 166132 11676 166138 11688
rect 166353 11679 166411 11685
rect 166353 11676 166365 11679
rect 166132 11648 166365 11676
rect 166132 11636 166138 11648
rect 166353 11645 166365 11648
rect 166399 11645 166411 11679
rect 166353 11639 166411 11645
rect 145156 11580 150572 11608
rect 150621 11611 150679 11617
rect 145156 11568 145162 11580
rect 150621 11577 150633 11611
rect 150667 11608 150679 11611
rect 151630 11608 151636 11620
rect 150667 11580 151636 11608
rect 150667 11577 150679 11580
rect 150621 11571 150679 11577
rect 151630 11568 151636 11580
rect 151688 11608 151694 11620
rect 152093 11611 152151 11617
rect 152093 11608 152105 11611
rect 151688 11580 152105 11608
rect 151688 11568 151694 11580
rect 152093 11577 152105 11580
rect 152139 11577 152151 11611
rect 152093 11571 152151 11577
rect 156325 11611 156383 11617
rect 156325 11577 156337 11611
rect 156371 11608 156383 11611
rect 159542 11608 159548 11620
rect 156371 11580 159548 11608
rect 156371 11577 156383 11580
rect 156325 11571 156383 11577
rect 159542 11568 159548 11580
rect 159600 11568 159606 11620
rect 160281 11611 160339 11617
rect 160281 11577 160293 11611
rect 160327 11608 160339 11611
rect 164326 11608 164332 11620
rect 160327 11580 164332 11608
rect 160327 11577 160339 11580
rect 160281 11571 160339 11577
rect 164326 11568 164332 11580
rect 164384 11568 164390 11620
rect 124674 11540 124680 11552
rect 119304 11512 124536 11540
rect 124635 11512 124680 11540
rect 119304 11500 119310 11512
rect 124674 11500 124680 11512
rect 124732 11500 124738 11552
rect 126146 11500 126152 11552
rect 126204 11540 126210 11552
rect 128909 11543 128967 11549
rect 128909 11540 128921 11543
rect 126204 11512 128921 11540
rect 126204 11500 126210 11512
rect 128909 11509 128921 11512
rect 128955 11509 128967 11543
rect 128909 11503 128967 11509
rect 130194 11500 130200 11552
rect 130252 11540 130258 11552
rect 130381 11543 130439 11549
rect 130381 11540 130393 11543
rect 130252 11512 130393 11540
rect 130252 11500 130258 11512
rect 130381 11509 130393 11512
rect 130427 11540 130439 11543
rect 131298 11540 131304 11552
rect 130427 11512 131304 11540
rect 130427 11509 130439 11512
rect 130381 11503 130439 11509
rect 131298 11500 131304 11512
rect 131356 11500 131362 11552
rect 134334 11540 134340 11552
rect 134295 11512 134340 11540
rect 134334 11500 134340 11512
rect 134392 11500 134398 11552
rect 135622 11540 135628 11552
rect 135583 11512 135628 11540
rect 135622 11500 135628 11512
rect 135680 11500 135686 11552
rect 135990 11540 135996 11552
rect 135951 11512 135996 11540
rect 135990 11500 135996 11512
rect 136048 11500 136054 11552
rect 137462 11540 137468 11552
rect 137423 11512 137468 11540
rect 137462 11500 137468 11512
rect 137520 11500 137526 11552
rect 138106 11540 138112 11552
rect 138067 11512 138112 11540
rect 138106 11500 138112 11512
rect 138164 11500 138170 11552
rect 143994 11540 144000 11552
rect 143955 11512 144000 11540
rect 143994 11500 144000 11512
rect 144052 11500 144058 11552
rect 146938 11540 146944 11552
rect 146899 11512 146944 11540
rect 146938 11500 146944 11512
rect 146996 11500 147002 11552
rect 150986 11540 150992 11552
rect 150947 11512 150992 11540
rect 150986 11500 150992 11512
rect 151044 11500 151050 11552
rect 151725 11543 151783 11549
rect 151725 11509 151737 11543
rect 151771 11540 151783 11543
rect 153194 11540 153200 11552
rect 151771 11512 153200 11540
rect 151771 11509 151783 11512
rect 151725 11503 151783 11509
rect 153194 11500 153200 11512
rect 153252 11500 153258 11552
rect 154577 11543 154635 11549
rect 154577 11509 154589 11543
rect 154623 11540 154635 11543
rect 155954 11540 155960 11552
rect 154623 11512 155960 11540
rect 154623 11509 154635 11512
rect 154577 11503 154635 11509
rect 155954 11500 155960 11512
rect 156012 11500 156018 11552
rect 157426 11540 157432 11552
rect 157387 11512 157432 11540
rect 157426 11500 157432 11512
rect 157484 11500 157490 11552
rect 162029 11543 162087 11549
rect 162029 11509 162041 11543
rect 162075 11540 162087 11543
rect 163038 11540 163044 11552
rect 162075 11512 163044 11540
rect 162075 11509 162087 11512
rect 162029 11503 162087 11509
rect 163038 11500 163044 11512
rect 163096 11500 163102 11552
rect 163133 11543 163191 11549
rect 163133 11509 163145 11543
rect 163179 11540 163191 11543
rect 166718 11540 166724 11552
rect 163179 11512 166724 11540
rect 163179 11509 163191 11512
rect 163133 11503 163191 11509
rect 166718 11500 166724 11512
rect 166776 11500 166782 11552
rect 368 11450 169556 11472
rect 368 11398 28456 11450
rect 28508 11398 28520 11450
rect 28572 11398 28584 11450
rect 28636 11398 28648 11450
rect 28700 11398 84878 11450
rect 84930 11398 84942 11450
rect 84994 11398 85006 11450
rect 85058 11398 85070 11450
rect 85122 11398 141299 11450
rect 141351 11398 141363 11450
rect 141415 11398 141427 11450
rect 141479 11398 141491 11450
rect 141543 11398 169556 11450
rect 368 11376 169556 11398
rect 4798 11336 4804 11348
rect 4759 11308 4804 11336
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 11149 11339 11207 11345
rect 11149 11305 11161 11339
rect 11195 11336 11207 11339
rect 11425 11339 11483 11345
rect 11425 11336 11437 11339
rect 11195 11308 11437 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 11425 11305 11437 11308
rect 11471 11336 11483 11339
rect 11514 11336 11520 11348
rect 11471 11308 11520 11336
rect 11471 11305 11483 11308
rect 11425 11299 11483 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 16482 11336 16488 11348
rect 16443 11308 16488 11336
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 22370 11336 22376 11348
rect 22331 11308 22376 11336
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 23569 11339 23627 11345
rect 23569 11305 23581 11339
rect 23615 11336 23627 11339
rect 27982 11336 27988 11348
rect 23615 11308 27988 11336
rect 23615 11305 23627 11308
rect 23569 11299 23627 11305
rect 27982 11296 27988 11308
rect 28040 11296 28046 11348
rect 28905 11339 28963 11345
rect 28905 11305 28917 11339
rect 28951 11336 28963 11339
rect 29178 11336 29184 11348
rect 28951 11308 29184 11336
rect 28951 11305 28963 11308
rect 28905 11299 28963 11305
rect 29178 11296 29184 11308
rect 29236 11296 29242 11348
rect 29362 11296 29368 11348
rect 29420 11336 29426 11348
rect 29457 11339 29515 11345
rect 29457 11336 29469 11339
rect 29420 11308 29469 11336
rect 29420 11296 29426 11308
rect 29457 11305 29469 11308
rect 29503 11305 29515 11339
rect 29457 11299 29515 11305
rect 30101 11339 30159 11345
rect 30101 11305 30113 11339
rect 30147 11336 30159 11339
rect 31294 11336 31300 11348
rect 30147 11308 31300 11336
rect 30147 11305 30159 11308
rect 30101 11299 30159 11305
rect 31294 11296 31300 11308
rect 31352 11296 31358 11348
rect 33134 11296 33140 11348
rect 33192 11336 33198 11348
rect 33229 11339 33287 11345
rect 33229 11336 33241 11339
rect 33192 11308 33241 11336
rect 33192 11296 33198 11308
rect 33229 11305 33241 11308
rect 33275 11305 33287 11339
rect 33229 11299 33287 11305
rect 33781 11339 33839 11345
rect 33781 11305 33793 11339
rect 33827 11336 33839 11339
rect 34054 11336 34060 11348
rect 33827 11308 34060 11336
rect 33827 11305 33839 11308
rect 33781 11299 33839 11305
rect 34054 11296 34060 11308
rect 34112 11296 34118 11348
rect 34974 11296 34980 11348
rect 35032 11336 35038 11348
rect 39669 11339 39727 11345
rect 39669 11336 39681 11339
rect 35032 11308 39681 11336
rect 35032 11296 35038 11308
rect 39669 11305 39681 11308
rect 39715 11305 39727 11339
rect 39669 11299 39727 11305
rect 39758 11296 39764 11348
rect 39816 11336 39822 11348
rect 42889 11339 42947 11345
rect 42889 11336 42901 11339
rect 39816 11308 42901 11336
rect 39816 11296 39822 11308
rect 42889 11305 42901 11308
rect 42935 11305 42947 11339
rect 42889 11299 42947 11305
rect 43441 11339 43499 11345
rect 43441 11305 43453 11339
rect 43487 11336 43499 11339
rect 43714 11336 43720 11348
rect 43487 11308 43720 11336
rect 43487 11305 43499 11308
rect 43441 11299 43499 11305
rect 43714 11296 43720 11308
rect 43772 11296 43778 11348
rect 45830 11296 45836 11348
rect 45888 11336 45894 11348
rect 46290 11336 46296 11348
rect 45888 11308 46296 11336
rect 45888 11296 45894 11308
rect 46290 11296 46296 11308
rect 46348 11296 46354 11348
rect 46566 11296 46572 11348
rect 46624 11336 46630 11348
rect 69845 11339 69903 11345
rect 69845 11336 69857 11339
rect 46624 11308 69857 11336
rect 46624 11296 46630 11308
rect 69845 11305 69857 11308
rect 69891 11305 69903 11339
rect 70762 11336 70768 11348
rect 70723 11308 70768 11336
rect 69845 11299 69903 11305
rect 70762 11296 70768 11308
rect 70820 11296 70826 11348
rect 72326 11336 72332 11348
rect 72287 11308 72332 11336
rect 72326 11296 72332 11308
rect 72384 11296 72390 11348
rect 74169 11339 74227 11345
rect 74169 11305 74181 11339
rect 74215 11336 74227 11339
rect 74442 11336 74448 11348
rect 74215 11308 74448 11336
rect 74215 11305 74227 11308
rect 74169 11299 74227 11305
rect 74442 11296 74448 11308
rect 74500 11296 74506 11348
rect 74994 11336 75000 11348
rect 74955 11308 75000 11336
rect 74994 11296 75000 11308
rect 75052 11296 75058 11348
rect 75362 11336 75368 11348
rect 75323 11308 75368 11336
rect 75362 11296 75368 11308
rect 75420 11296 75426 11348
rect 77662 11336 77668 11348
rect 77623 11308 77668 11336
rect 77662 11296 77668 11308
rect 77720 11296 77726 11348
rect 77938 11336 77944 11348
rect 77899 11308 77944 11336
rect 77938 11296 77944 11308
rect 77996 11296 78002 11348
rect 78766 11296 78772 11348
rect 78824 11336 78830 11348
rect 78953 11339 79011 11345
rect 78953 11336 78965 11339
rect 78824 11308 78965 11336
rect 78824 11296 78830 11308
rect 78953 11305 78965 11308
rect 78999 11305 79011 11339
rect 78953 11299 79011 11305
rect 80974 11296 80980 11348
rect 81032 11336 81038 11348
rect 81989 11339 82047 11345
rect 81989 11336 82001 11339
rect 81032 11308 82001 11336
rect 81032 11296 81038 11308
rect 81989 11305 82001 11308
rect 82035 11305 82047 11339
rect 82998 11336 83004 11348
rect 82959 11308 83004 11336
rect 81989 11299 82047 11305
rect 82998 11296 83004 11308
rect 83056 11296 83062 11348
rect 83366 11336 83372 11348
rect 83327 11308 83372 11336
rect 83366 11296 83372 11308
rect 83424 11296 83430 11348
rect 84746 11336 84752 11348
rect 84707 11308 84752 11336
rect 84746 11296 84752 11308
rect 84804 11296 84810 11348
rect 87138 11336 87144 11348
rect 87099 11308 87144 11336
rect 87138 11296 87144 11308
rect 87196 11296 87202 11348
rect 98178 11336 98184 11348
rect 98139 11308 98184 11336
rect 98178 11296 98184 11308
rect 98236 11296 98242 11348
rect 101125 11339 101183 11345
rect 101125 11305 101137 11339
rect 101171 11336 101183 11339
rect 101398 11336 101404 11348
rect 101171 11308 101404 11336
rect 101171 11305 101183 11308
rect 101125 11299 101183 11305
rect 101398 11296 101404 11308
rect 101456 11296 101462 11348
rect 104066 11336 104072 11348
rect 104027 11308 104072 11336
rect 104066 11296 104072 11308
rect 104124 11296 104130 11348
rect 104621 11339 104679 11345
rect 104621 11305 104633 11339
rect 104667 11336 104679 11339
rect 104894 11336 104900 11348
rect 104667 11308 104900 11336
rect 104667 11305 104679 11308
rect 104621 11299 104679 11305
rect 104894 11296 104900 11308
rect 104952 11296 104958 11348
rect 105262 11336 105268 11348
rect 105223 11308 105268 11336
rect 105262 11296 105268 11308
rect 105320 11296 105326 11348
rect 106550 11336 106556 11348
rect 106511 11308 106556 11336
rect 106550 11296 106556 11308
rect 106608 11296 106614 11348
rect 112901 11339 112959 11345
rect 108132 11308 111472 11336
rect 3694 11228 3700 11280
rect 3752 11268 3758 11280
rect 5718 11268 5724 11280
rect 3752 11240 5724 11268
rect 3752 11228 3758 11240
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 7193 11271 7251 11277
rect 7193 11237 7205 11271
rect 7239 11268 7251 11271
rect 9766 11268 9772 11280
rect 7239 11240 9772 11268
rect 7239 11237 7251 11240
rect 7193 11231 7251 11237
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 16025 11271 16083 11277
rect 16025 11237 16037 11271
rect 16071 11268 16083 11271
rect 19886 11268 19892 11280
rect 16071 11240 19892 11268
rect 16071 11237 16083 11240
rect 16025 11231 16083 11237
rect 19886 11228 19892 11240
rect 19944 11228 19950 11280
rect 22094 11228 22100 11280
rect 22152 11228 22158 11280
rect 24210 11268 24216 11280
rect 24171 11240 24216 11268
rect 24210 11228 24216 11240
rect 24268 11228 24274 11280
rect 24578 11268 24584 11280
rect 24539 11240 24584 11268
rect 24578 11228 24584 11240
rect 24636 11228 24642 11280
rect 26602 11268 26608 11280
rect 26563 11240 26608 11268
rect 26602 11228 26608 11240
rect 26660 11228 26666 11280
rect 28718 11268 28724 11280
rect 26896 11240 28724 11268
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 4338 11200 4344 11212
rect 2271 11172 4344 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 4522 11200 4528 11212
rect 4483 11172 4528 11200
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 7650 11200 7656 11212
rect 7300 11172 7656 11200
rect 4154 11132 4160 11144
rect 4115 11104 4160 11132
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 6086 11132 6092 11144
rect 5767 11104 6092 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 7300 11141 7328 11172
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11200 9551 11203
rect 9674 11200 9680 11212
rect 9539 11172 9680 11200
rect 9539 11169 9551 11172
rect 9493 11163 9551 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 16942 11200 16948 11212
rect 11011 11172 16948 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 19150 11160 19156 11212
rect 19208 11200 19214 11212
rect 21177 11203 21235 11209
rect 21177 11200 21189 11203
rect 19208 11172 21189 11200
rect 19208 11160 19214 11172
rect 21177 11169 21189 11172
rect 21223 11169 21235 11203
rect 22112 11200 22140 11228
rect 26896 11200 26924 11240
rect 28718 11228 28724 11240
rect 28776 11228 28782 11280
rect 30742 11268 30748 11280
rect 30703 11240 30748 11268
rect 30742 11228 30748 11240
rect 30800 11228 30806 11280
rect 33410 11228 33416 11280
rect 33468 11268 33474 11280
rect 37734 11268 37740 11280
rect 33468 11240 37740 11268
rect 33468 11228 33474 11240
rect 37734 11228 37740 11240
rect 37792 11228 37798 11280
rect 48774 11268 48780 11280
rect 37844 11240 48780 11268
rect 22112 11172 26924 11200
rect 21177 11163 21235 11169
rect 27062 11160 27068 11212
rect 27120 11200 27126 11212
rect 27249 11203 27307 11209
rect 27249 11200 27261 11203
rect 27120 11172 27261 11200
rect 27120 11160 27126 11172
rect 27249 11169 27261 11172
rect 27295 11169 27307 11203
rect 28258 11200 28264 11212
rect 28219 11172 28264 11200
rect 27249 11163 27307 11169
rect 28258 11160 28264 11172
rect 28316 11160 28322 11212
rect 31938 11200 31944 11212
rect 28368 11172 31944 11200
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11101 7343 11135
rect 8018 11132 8024 11144
rect 7979 11104 8024 11132
rect 7285 11095 7343 11101
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11132 11115 11135
rect 11149 11135 11207 11141
rect 11149 11132 11161 11135
rect 11103 11104 11161 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 11149 11101 11161 11104
rect 11195 11101 11207 11135
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 11149 11095 11207 11101
rect 14292 11104 14565 11132
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 8570 11064 8576 11076
rect 4120 11036 8576 11064
rect 4120 11024 4126 11036
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 11977 11067 12035 11073
rect 11977 11033 11989 11067
rect 12023 11064 12035 11067
rect 12618 11064 12624 11076
rect 12023 11036 12624 11064
rect 12023 11033 12035 11036
rect 11977 11027 12035 11033
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 14292 11073 14320 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11132 16175 11135
rect 16482 11132 16488 11144
rect 16163 11104 16488 11132
rect 16163 11101 16175 11104
rect 16117 11095 16175 11101
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 20165 11135 20223 11141
rect 20165 11132 20177 11135
rect 20128 11104 20177 11132
rect 20128 11092 20134 11104
rect 20165 11101 20177 11104
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11132 21787 11135
rect 22097 11135 22155 11141
rect 22097 11132 22109 11135
rect 21775 11104 22109 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 22097 11101 22109 11104
rect 22143 11132 22155 11135
rect 23382 11132 23388 11144
rect 22143 11104 23388 11132
rect 22143 11101 22155 11104
rect 22097 11095 22155 11101
rect 23382 11092 23388 11104
rect 23440 11092 23446 11144
rect 23753 11135 23811 11141
rect 23753 11101 23765 11135
rect 23799 11132 23811 11135
rect 24210 11132 24216 11144
rect 23799 11104 24216 11132
rect 23799 11101 23811 11104
rect 23753 11095 23811 11101
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 28368 11132 28396 11172
rect 31938 11160 31944 11172
rect 31996 11160 32002 11212
rect 32125 11203 32183 11209
rect 32125 11169 32137 11203
rect 32171 11200 32183 11203
rect 32398 11200 32404 11212
rect 32171 11172 32404 11200
rect 32171 11169 32183 11172
rect 32125 11163 32183 11169
rect 32398 11160 32404 11172
rect 32456 11160 32462 11212
rect 32582 11200 32588 11212
rect 32495 11172 32588 11200
rect 32582 11160 32588 11172
rect 32640 11200 32646 11212
rect 35526 11200 35532 11212
rect 32640 11172 34744 11200
rect 35487 11172 35532 11200
rect 32640 11160 32646 11172
rect 27264 11104 28396 11132
rect 28813 11135 28871 11141
rect 13449 11067 13507 11073
rect 13449 11033 13461 11067
rect 13495 11064 13507 11067
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 13495 11036 14289 11064
rect 13495 11033 13507 11036
rect 13449 11027 13507 11033
rect 14277 11033 14289 11036
rect 14323 11033 14335 11067
rect 14277 11027 14335 11033
rect 18877 11067 18935 11073
rect 18877 11033 18889 11067
rect 18923 11064 18935 11067
rect 19702 11064 19708 11076
rect 18923 11036 19708 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 19981 11067 20039 11073
rect 19981 11033 19993 11067
rect 20027 11064 20039 11067
rect 20806 11064 20812 11076
rect 20027 11036 20812 11064
rect 20027 11033 20039 11036
rect 19981 11027 20039 11033
rect 20806 11024 20812 11036
rect 20864 11024 20870 11076
rect 24854 11024 24860 11076
rect 24912 11064 24918 11076
rect 25777 11067 25835 11073
rect 25777 11064 25789 11067
rect 24912 11036 25789 11064
rect 24912 11024 24918 11036
rect 25777 11033 25789 11036
rect 25823 11033 25835 11067
rect 27264 11064 27292 11104
rect 28813 11101 28825 11135
rect 28859 11132 28871 11135
rect 28905 11135 28963 11141
rect 28905 11132 28917 11135
rect 28859 11104 28917 11132
rect 28859 11101 28871 11104
rect 28813 11095 28871 11101
rect 28905 11101 28917 11104
rect 28951 11101 28963 11135
rect 29638 11132 29644 11144
rect 28905 11095 28963 11101
rect 29012 11104 29644 11132
rect 25777 11027 25835 11033
rect 25884 11036 27292 11064
rect 11422 10956 11428 11008
rect 11480 10996 11486 11008
rect 24302 10996 24308 11008
rect 11480 10968 24308 10996
rect 11480 10956 11486 10968
rect 24302 10956 24308 10968
rect 24360 10956 24366 11008
rect 24670 10996 24676 11008
rect 24631 10968 24676 10996
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 24762 10956 24768 11008
rect 24820 10996 24826 11008
rect 25884 10996 25912 11036
rect 27430 11024 27436 11076
rect 27488 11064 27494 11076
rect 29012 11064 29040 11104
rect 29638 11092 29644 11104
rect 29696 11092 29702 11144
rect 30285 11135 30343 11141
rect 30285 11101 30297 11135
rect 30331 11132 30343 11135
rect 30742 11132 30748 11144
rect 30331 11104 30748 11132
rect 30331 11101 30343 11104
rect 30285 11095 30343 11101
rect 30742 11092 30748 11104
rect 30800 11092 30806 11144
rect 31205 11135 31263 11141
rect 31205 11101 31217 11135
rect 31251 11132 31263 11135
rect 32033 11135 32091 11141
rect 32033 11132 32045 11135
rect 31251 11104 32045 11132
rect 31251 11101 31263 11104
rect 31205 11095 31263 11101
rect 32033 11101 32045 11104
rect 32079 11132 32091 11135
rect 32490 11132 32496 11144
rect 32079 11104 32496 11132
rect 32079 11101 32091 11104
rect 32033 11095 32091 11101
rect 32490 11092 32496 11104
rect 32548 11092 32554 11144
rect 27488 11036 29040 11064
rect 27488 11024 27494 11036
rect 29086 11024 29092 11076
rect 29144 11064 29150 11076
rect 32122 11064 32128 11076
rect 29144 11036 32128 11064
rect 29144 11024 29150 11036
rect 32122 11024 32128 11036
rect 32180 11024 32186 11076
rect 32401 11067 32459 11073
rect 32401 11033 32413 11067
rect 32447 11064 32459 11067
rect 32600 11064 32628 11160
rect 33597 11135 33655 11141
rect 33597 11101 33609 11135
rect 33643 11132 33655 11135
rect 33781 11135 33839 11141
rect 33781 11132 33793 11135
rect 33643 11104 33793 11132
rect 33643 11101 33655 11104
rect 33597 11095 33655 11101
rect 33781 11101 33793 11104
rect 33827 11101 33839 11135
rect 33781 11095 33839 11101
rect 34517 11135 34575 11141
rect 34517 11101 34529 11135
rect 34563 11132 34575 11135
rect 34716 11132 34744 11172
rect 35526 11160 35532 11172
rect 35584 11160 35590 11212
rect 36722 11200 36728 11212
rect 35636 11172 36728 11200
rect 35636 11132 35664 11172
rect 36722 11160 36728 11172
rect 36780 11160 36786 11212
rect 36998 11200 37004 11212
rect 36959 11172 37004 11200
rect 36998 11160 37004 11172
rect 37056 11160 37062 11212
rect 37090 11160 37096 11212
rect 37148 11200 37154 11212
rect 37844 11200 37872 11240
rect 48774 11228 48780 11240
rect 48832 11228 48838 11280
rect 49142 11268 49148 11280
rect 49103 11240 49148 11268
rect 49142 11228 49148 11240
rect 49200 11228 49206 11280
rect 49234 11228 49240 11280
rect 49292 11268 49298 11280
rect 50985 11271 51043 11277
rect 50985 11268 50997 11271
rect 49292 11240 50997 11268
rect 49292 11228 49298 11240
rect 50985 11237 50997 11240
rect 51031 11237 51043 11271
rect 50985 11231 51043 11237
rect 51074 11228 51080 11280
rect 51132 11268 51138 11280
rect 51629 11271 51687 11277
rect 51629 11268 51641 11271
rect 51132 11240 51641 11268
rect 51132 11228 51138 11240
rect 51629 11237 51641 11240
rect 51675 11268 51687 11271
rect 55769 11271 55827 11277
rect 55769 11268 55781 11271
rect 51675 11240 55781 11268
rect 51675 11237 51687 11240
rect 51629 11231 51687 11237
rect 55769 11237 55781 11240
rect 55815 11237 55827 11271
rect 55769 11231 55827 11237
rect 55861 11271 55919 11277
rect 55861 11237 55873 11271
rect 55907 11268 55919 11271
rect 56962 11268 56968 11280
rect 55907 11240 56968 11268
rect 55907 11237 55919 11240
rect 55861 11231 55919 11237
rect 56962 11228 56968 11240
rect 57020 11228 57026 11280
rect 57333 11271 57391 11277
rect 57333 11237 57345 11271
rect 57379 11268 57391 11271
rect 57609 11271 57667 11277
rect 57609 11268 57621 11271
rect 57379 11240 57621 11268
rect 57379 11237 57391 11240
rect 57333 11231 57391 11237
rect 57609 11237 57621 11240
rect 57655 11268 57667 11271
rect 58894 11268 58900 11280
rect 57655 11240 58900 11268
rect 57655 11237 57667 11240
rect 57609 11231 57667 11237
rect 58894 11228 58900 11240
rect 58952 11228 58958 11280
rect 59078 11228 59084 11280
rect 59136 11268 59142 11280
rect 59541 11271 59599 11277
rect 59541 11268 59553 11271
rect 59136 11240 59553 11268
rect 59136 11228 59142 11240
rect 59541 11237 59553 11240
rect 59587 11237 59599 11271
rect 59541 11231 59599 11237
rect 60277 11271 60335 11277
rect 60277 11237 60289 11271
rect 60323 11268 60335 11271
rect 60553 11271 60611 11277
rect 60553 11268 60565 11271
rect 60323 11240 60565 11268
rect 60323 11237 60335 11240
rect 60277 11231 60335 11237
rect 60553 11237 60565 11240
rect 60599 11268 60611 11271
rect 60918 11268 60924 11280
rect 60599 11240 60924 11268
rect 60599 11237 60611 11240
rect 60553 11231 60611 11237
rect 60918 11228 60924 11240
rect 60976 11228 60982 11280
rect 61105 11271 61163 11277
rect 61105 11237 61117 11271
rect 61151 11268 61163 11271
rect 61286 11268 61292 11280
rect 61151 11240 61292 11268
rect 61151 11237 61163 11240
rect 61105 11231 61163 11237
rect 61286 11228 61292 11240
rect 61344 11228 61350 11280
rect 61378 11228 61384 11280
rect 61436 11268 61442 11280
rect 68741 11271 68799 11277
rect 68741 11268 68753 11271
rect 61436 11240 68753 11268
rect 61436 11228 61442 11240
rect 68741 11237 68753 11240
rect 68787 11237 68799 11271
rect 68741 11231 68799 11237
rect 69477 11271 69535 11277
rect 69477 11237 69489 11271
rect 69523 11268 69535 11271
rect 69753 11271 69811 11277
rect 69753 11268 69765 11271
rect 69523 11240 69765 11268
rect 69523 11237 69535 11240
rect 69477 11231 69535 11237
rect 69753 11237 69765 11240
rect 69799 11268 69811 11271
rect 69934 11268 69940 11280
rect 69799 11240 69940 11268
rect 69799 11237 69811 11240
rect 69753 11231 69811 11237
rect 69934 11228 69940 11240
rect 69992 11228 69998 11280
rect 76377 11271 76435 11277
rect 76377 11268 76389 11271
rect 72896 11240 76389 11268
rect 38010 11200 38016 11212
rect 37148 11172 37872 11200
rect 37971 11172 38016 11200
rect 37148 11160 37154 11172
rect 38010 11160 38016 11172
rect 38068 11160 38074 11212
rect 72418 11200 72424 11212
rect 38396 11172 72424 11200
rect 34563 11104 34597 11132
rect 34716 11104 35664 11132
rect 36081 11135 36139 11141
rect 34563 11101 34575 11104
rect 34517 11095 34575 11101
rect 36081 11101 36093 11135
rect 36127 11101 36139 11135
rect 36081 11095 36139 11101
rect 32447 11036 32628 11064
rect 34425 11067 34483 11073
rect 32447 11033 32459 11036
rect 32401 11027 32459 11033
rect 34425 11033 34437 11067
rect 34471 11064 34483 11067
rect 34532 11064 34560 11095
rect 34606 11064 34612 11076
rect 34471 11036 34612 11064
rect 34471 11033 34483 11036
rect 34425 11027 34483 11033
rect 34606 11024 34612 11036
rect 34664 11024 34670 11076
rect 36096 11064 36124 11095
rect 36170 11092 36176 11144
rect 36228 11132 36234 11144
rect 37642 11132 37648 11144
rect 36228 11104 37648 11132
rect 36228 11092 36234 11104
rect 37642 11092 37648 11104
rect 37700 11092 37706 11144
rect 36449 11067 36507 11073
rect 36449 11064 36461 11067
rect 36096 11036 36461 11064
rect 36449 11033 36461 11036
rect 36495 11064 36507 11067
rect 38396 11064 38424 11172
rect 72418 11160 72424 11172
rect 72476 11160 72482 11212
rect 72513 11203 72571 11209
rect 72513 11169 72525 11203
rect 72559 11200 72571 11203
rect 72786 11200 72792 11212
rect 72559 11172 72792 11200
rect 72559 11169 72571 11172
rect 72513 11163 72571 11169
rect 72786 11160 72792 11172
rect 72844 11160 72850 11212
rect 38473 11135 38531 11141
rect 38473 11101 38485 11135
rect 38519 11132 38531 11135
rect 38657 11135 38715 11141
rect 38519 11104 38608 11132
rect 38519 11101 38531 11104
rect 38473 11095 38531 11101
rect 36495 11036 38424 11064
rect 38580 11064 38608 11104
rect 38657 11101 38669 11135
rect 38703 11132 38715 11135
rect 40037 11135 40095 11141
rect 38703 11104 39528 11132
rect 38703 11101 38715 11104
rect 38657 11095 38715 11101
rect 38930 11064 38936 11076
rect 38580 11036 38936 11064
rect 36495 11033 36507 11036
rect 36449 11027 36507 11033
rect 38930 11024 38936 11036
rect 38988 11024 38994 11076
rect 24820 10968 25912 10996
rect 24820 10956 24826 10968
rect 27246 10956 27252 11008
rect 27304 10996 27310 11008
rect 27522 10996 27528 11008
rect 27304 10968 27528 10996
rect 27304 10956 27310 10968
rect 27522 10956 27528 10968
rect 27580 10956 27586 11008
rect 27614 10956 27620 11008
rect 27672 10996 27678 11008
rect 32306 10996 32312 11008
rect 27672 10968 32312 10996
rect 27672 10956 27678 10968
rect 32306 10956 32312 10968
rect 32364 10956 32370 11008
rect 32490 10956 32496 11008
rect 32548 10996 32554 11008
rect 37550 10996 37556 11008
rect 32548 10968 37556 10996
rect 32548 10956 32554 10968
rect 37550 10956 37556 10968
rect 37608 10956 37614 11008
rect 37642 10956 37648 11008
rect 37700 10996 37706 11008
rect 38657 10999 38715 11005
rect 38657 10996 38669 10999
rect 37700 10968 38669 10996
rect 37700 10956 37706 10968
rect 38657 10965 38669 10968
rect 38703 10965 38715 10999
rect 38657 10959 38715 10965
rect 38746 10956 38752 11008
rect 38804 10996 38810 11008
rect 39390 10996 39396 11008
rect 38804 10968 39396 10996
rect 38804 10956 38810 10968
rect 39390 10956 39396 10968
rect 39448 10956 39454 11008
rect 39500 10996 39528 11104
rect 40037 11101 40049 11135
rect 40083 11101 40095 11135
rect 40037 11095 40095 11101
rect 40221 11135 40279 11141
rect 40221 11101 40233 11135
rect 40267 11132 40279 11135
rect 40957 11135 41015 11141
rect 40957 11132 40969 11135
rect 40267 11104 40969 11132
rect 40267 11101 40279 11104
rect 40221 11095 40279 11101
rect 40957 11101 40969 11104
rect 41003 11101 41015 11135
rect 40957 11095 41015 11101
rect 40052 11064 40080 11095
rect 41046 11092 41052 11144
rect 41104 11132 41110 11144
rect 41601 11135 41659 11141
rect 41104 11104 41368 11132
rect 41104 11092 41110 11104
rect 40497 11067 40555 11073
rect 40497 11064 40509 11067
rect 40052 11036 40509 11064
rect 40497 11033 40509 11036
rect 40543 11064 40555 11067
rect 40586 11064 40592 11076
rect 40543 11036 40592 11064
rect 40543 11033 40555 11036
rect 40497 11027 40555 11033
rect 40586 11024 40592 11036
rect 40644 11024 40650 11076
rect 41340 11064 41368 11104
rect 41601 11101 41613 11135
rect 41647 11132 41659 11135
rect 42061 11135 42119 11141
rect 42061 11132 42073 11135
rect 41647 11104 42073 11132
rect 41647 11101 41659 11104
rect 41601 11095 41659 11101
rect 42061 11101 42073 11104
rect 42107 11132 42119 11135
rect 42794 11132 42800 11144
rect 42107 11104 42800 11132
rect 42107 11101 42119 11104
rect 42061 11095 42119 11101
rect 42794 11092 42800 11104
rect 42852 11092 42858 11144
rect 43257 11135 43315 11141
rect 43257 11101 43269 11135
rect 43303 11132 43315 11135
rect 43441 11135 43499 11141
rect 43441 11132 43453 11135
rect 43303 11104 43453 11132
rect 43303 11101 43315 11104
rect 43257 11095 43315 11101
rect 43441 11101 43453 11104
rect 43487 11101 43499 11135
rect 45646 11132 45652 11144
rect 43441 11095 43499 11101
rect 43732 11104 45652 11132
rect 43732 11064 43760 11104
rect 45646 11092 45652 11104
rect 45704 11092 45710 11144
rect 45830 11132 45836 11144
rect 45791 11104 45836 11132
rect 45830 11092 45836 11104
rect 45888 11092 45894 11144
rect 45922 11092 45928 11144
rect 45980 11132 45986 11144
rect 46017 11135 46075 11141
rect 46017 11132 46029 11135
rect 45980 11104 46029 11132
rect 45980 11092 45986 11104
rect 46017 11101 46029 11104
rect 46063 11101 46075 11135
rect 46017 11095 46075 11101
rect 46293 11135 46351 11141
rect 46293 11101 46305 11135
rect 46339 11132 46351 11135
rect 46658 11132 46664 11144
rect 46339 11104 46664 11132
rect 46339 11101 46351 11104
rect 46293 11095 46351 11101
rect 46658 11092 46664 11104
rect 46716 11092 46722 11144
rect 47118 11132 47124 11144
rect 47031 11104 47124 11132
rect 47118 11092 47124 11104
rect 47176 11132 47182 11144
rect 48682 11132 48688 11144
rect 47176 11104 48688 11132
rect 47176 11092 47182 11104
rect 48682 11092 48688 11104
rect 48740 11092 48746 11144
rect 48774 11092 48780 11144
rect 48832 11132 48838 11144
rect 49418 11132 49424 11144
rect 48832 11104 49424 11132
rect 48832 11092 48838 11104
rect 49418 11092 49424 11104
rect 49476 11092 49482 11144
rect 49694 11132 49700 11144
rect 49655 11104 49700 11132
rect 49694 11092 49700 11104
rect 49752 11092 49758 11144
rect 50246 11132 50252 11144
rect 50080 11104 50252 11132
rect 41340 11036 43760 11064
rect 44637 11067 44695 11073
rect 44637 11033 44649 11067
rect 44683 11064 44695 11067
rect 46382 11064 46388 11076
rect 44683 11036 46388 11064
rect 44683 11033 44695 11036
rect 44637 11027 44695 11033
rect 46382 11024 46388 11036
rect 46440 11024 46446 11076
rect 49602 11064 49608 11076
rect 46584 11036 47164 11064
rect 40221 10999 40279 11005
rect 40221 10996 40233 10999
rect 39500 10968 40233 10996
rect 40221 10965 40233 10968
rect 40267 10965 40279 10999
rect 40770 10996 40776 11008
rect 40731 10968 40776 10996
rect 40221 10959 40279 10965
rect 40770 10956 40776 10968
rect 40828 10956 40834 11008
rect 40954 10956 40960 11008
rect 41012 10996 41018 11008
rect 41782 10996 41788 11008
rect 41012 10968 41788 10996
rect 41012 10956 41018 10968
rect 41782 10956 41788 10968
rect 41840 10956 41846 11008
rect 42058 10956 42064 11008
rect 42116 10996 42122 11008
rect 46584 10996 46612 11036
rect 42116 10968 46612 10996
rect 42116 10956 42122 10968
rect 46658 10956 46664 11008
rect 46716 10996 46722 11008
rect 46753 10999 46811 11005
rect 46753 10996 46765 10999
rect 46716 10968 46765 10996
rect 46716 10956 46722 10968
rect 46753 10965 46765 10968
rect 46799 10996 46811 10999
rect 47026 10996 47032 11008
rect 46799 10968 47032 10996
rect 46799 10965 46811 10968
rect 46753 10959 46811 10965
rect 47026 10956 47032 10968
rect 47084 10956 47090 11008
rect 47136 10996 47164 11036
rect 48056 11036 48360 11064
rect 49515 11036 49608 11064
rect 48056 10996 48084 11036
rect 48222 10996 48228 11008
rect 47136 10968 48084 10996
rect 48183 10968 48228 10996
rect 48222 10956 48228 10968
rect 48280 10956 48286 11008
rect 48332 10996 48360 11036
rect 49602 11024 49608 11036
rect 49660 11064 49666 11076
rect 50080 11064 50108 11104
rect 50246 11092 50252 11104
rect 50304 11092 50310 11144
rect 50522 11092 50528 11144
rect 50580 11132 50586 11144
rect 50706 11132 50712 11144
rect 50580 11104 50712 11132
rect 50580 11092 50586 11104
rect 50706 11092 50712 11104
rect 50764 11092 50770 11144
rect 50982 11132 50988 11144
rect 50943 11104 50988 11132
rect 50982 11092 50988 11104
rect 51040 11092 51046 11144
rect 52454 11132 52460 11144
rect 52415 11104 52460 11132
rect 52454 11092 52460 11104
rect 52512 11092 52518 11144
rect 52549 11135 52607 11141
rect 52549 11101 52561 11135
rect 52595 11101 52607 11135
rect 52549 11095 52607 11101
rect 52917 11135 52975 11141
rect 52917 11101 52929 11135
rect 52963 11132 52975 11135
rect 53285 11135 53343 11141
rect 53285 11132 53297 11135
rect 52963 11104 53297 11132
rect 52963 11101 52975 11104
rect 52917 11095 52975 11101
rect 53285 11101 53297 11104
rect 53331 11132 53343 11135
rect 55122 11132 55128 11144
rect 53331 11104 54984 11132
rect 55083 11104 55128 11132
rect 53331 11101 53343 11104
rect 53285 11095 53343 11101
rect 49660 11036 50108 11064
rect 49660 11024 49666 11036
rect 50154 11024 50160 11076
rect 50212 11064 50218 11076
rect 52564 11064 52592 11095
rect 53558 11064 53564 11076
rect 50212 11036 52592 11064
rect 53519 11036 53564 11064
rect 50212 11024 50218 11036
rect 53558 11024 53564 11036
rect 53616 11024 53622 11076
rect 53929 11067 53987 11073
rect 53929 11033 53941 11067
rect 53975 11064 53987 11067
rect 54662 11064 54668 11076
rect 53975 11036 54668 11064
rect 53975 11033 53987 11036
rect 53929 11027 53987 11033
rect 54662 11024 54668 11036
rect 54720 11024 54726 11076
rect 54956 11064 54984 11104
rect 55122 11092 55128 11104
rect 55180 11092 55186 11144
rect 55306 11132 55312 11144
rect 55267 11104 55312 11132
rect 55306 11092 55312 11104
rect 55364 11092 55370 11144
rect 55490 11132 55496 11144
rect 55451 11104 55496 11132
rect 55490 11092 55496 11104
rect 55548 11092 55554 11144
rect 55861 11135 55919 11141
rect 55861 11132 55873 11135
rect 55600 11104 55873 11132
rect 55600 11064 55628 11104
rect 55861 11101 55873 11104
rect 55907 11101 55919 11135
rect 56042 11132 56048 11144
rect 56003 11104 56048 11132
rect 55861 11095 55919 11101
rect 56042 11092 56048 11104
rect 56100 11092 56106 11144
rect 56413 11135 56471 11141
rect 56413 11101 56425 11135
rect 56459 11132 56471 11135
rect 56502 11132 56508 11144
rect 56459 11104 56508 11132
rect 56459 11101 56471 11104
rect 56413 11095 56471 11101
rect 56502 11092 56508 11104
rect 56560 11092 56566 11144
rect 56778 11132 56784 11144
rect 56739 11104 56784 11132
rect 56778 11092 56784 11104
rect 56836 11092 56842 11144
rect 56873 11135 56931 11141
rect 56873 11101 56885 11135
rect 56919 11132 56931 11135
rect 57146 11132 57152 11144
rect 56919 11104 57152 11132
rect 56919 11101 56931 11104
rect 56873 11095 56931 11101
rect 57146 11092 57152 11104
rect 57204 11092 57210 11144
rect 57241 11135 57299 11141
rect 57241 11101 57253 11135
rect 57287 11132 57299 11135
rect 57333 11135 57391 11141
rect 57333 11132 57345 11135
rect 57287 11104 57345 11132
rect 57287 11101 57299 11104
rect 57241 11095 57299 11101
rect 57333 11101 57345 11104
rect 57379 11101 57391 11135
rect 59538 11132 59544 11144
rect 57333 11095 57391 11101
rect 57440 11104 59544 11132
rect 54956 11036 55628 11064
rect 55769 11067 55827 11073
rect 55769 11033 55781 11067
rect 55815 11064 55827 11067
rect 57440 11064 57468 11104
rect 59538 11092 59544 11104
rect 59596 11092 59602 11144
rect 59722 11132 59728 11144
rect 59683 11104 59728 11132
rect 59722 11092 59728 11104
rect 59780 11092 59786 11144
rect 60185 11135 60243 11141
rect 60185 11101 60197 11135
rect 60231 11132 60243 11135
rect 60277 11135 60335 11141
rect 60277 11132 60289 11135
rect 60231 11104 60289 11132
rect 60231 11101 60243 11104
rect 60185 11095 60243 11101
rect 60277 11101 60289 11104
rect 60323 11101 60335 11135
rect 60277 11095 60335 11101
rect 60921 11135 60979 11141
rect 60921 11101 60933 11135
rect 60967 11132 60979 11135
rect 61286 11132 61292 11144
rect 60967 11104 61292 11132
rect 60967 11101 60979 11104
rect 60921 11095 60979 11101
rect 61286 11092 61292 11104
rect 61344 11092 61350 11144
rect 61749 11135 61807 11141
rect 61749 11101 61761 11135
rect 61795 11132 61807 11135
rect 62117 11135 62175 11141
rect 62117 11132 62129 11135
rect 61795 11104 62129 11132
rect 61795 11101 61807 11104
rect 61749 11095 61807 11101
rect 62117 11101 62129 11104
rect 62163 11132 62175 11135
rect 63402 11132 63408 11144
rect 62163 11104 63408 11132
rect 62163 11101 62175 11104
rect 62117 11095 62175 11101
rect 63402 11092 63408 11104
rect 63460 11092 63466 11144
rect 63586 11132 63592 11144
rect 63547 11104 63592 11132
rect 63586 11092 63592 11104
rect 63644 11092 63650 11144
rect 64690 11132 64696 11144
rect 64603 11104 64696 11132
rect 64690 11092 64696 11104
rect 64748 11132 64754 11144
rect 66073 11135 66131 11141
rect 66073 11132 66085 11135
rect 64748 11104 66085 11132
rect 64748 11092 64754 11104
rect 66073 11101 66085 11104
rect 66119 11101 66131 11135
rect 66073 11095 66131 11101
rect 67637 11135 67695 11141
rect 67637 11101 67649 11135
rect 67683 11132 67695 11135
rect 67910 11132 67916 11144
rect 67683 11104 67916 11132
rect 67683 11101 67695 11104
rect 67637 11095 67695 11101
rect 67910 11092 67916 11104
rect 67968 11092 67974 11144
rect 68557 11135 68615 11141
rect 68557 11101 68569 11135
rect 68603 11132 68615 11135
rect 68922 11132 68928 11144
rect 68603 11104 68928 11132
rect 68603 11101 68615 11104
rect 68557 11095 68615 11101
rect 68922 11092 68928 11104
rect 68980 11092 68986 11144
rect 69385 11135 69443 11141
rect 69385 11101 69397 11135
rect 69431 11132 69443 11135
rect 69477 11135 69535 11141
rect 69477 11132 69489 11135
rect 69431 11104 69489 11132
rect 69431 11101 69443 11104
rect 69385 11095 69443 11101
rect 69477 11101 69489 11104
rect 69523 11101 69535 11135
rect 69477 11095 69535 11101
rect 70121 11135 70179 11141
rect 70121 11101 70133 11135
rect 70167 11132 70179 11135
rect 70302 11132 70308 11144
rect 70167 11104 70308 11132
rect 70167 11101 70179 11104
rect 70121 11095 70179 11101
rect 70302 11092 70308 11104
rect 70360 11092 70366 11144
rect 70578 11092 70584 11144
rect 70636 11132 70642 11144
rect 70673 11135 70731 11141
rect 70673 11132 70685 11135
rect 70636 11104 70685 11132
rect 70636 11092 70642 11104
rect 70673 11101 70685 11104
rect 70719 11101 70731 11135
rect 70673 11095 70731 11101
rect 71130 11092 71136 11144
rect 71188 11132 71194 11144
rect 71225 11135 71283 11141
rect 71225 11132 71237 11135
rect 71188 11104 71237 11132
rect 71188 11092 71194 11104
rect 71225 11101 71237 11104
rect 71271 11132 71283 11135
rect 71685 11135 71743 11141
rect 71685 11132 71697 11135
rect 71271 11104 71697 11132
rect 71271 11101 71283 11104
rect 71225 11095 71283 11101
rect 71685 11101 71697 11104
rect 71731 11101 71743 11135
rect 71685 11095 71743 11101
rect 55815 11036 57468 11064
rect 55815 11033 55827 11036
rect 55769 11027 55827 11033
rect 57790 11024 57796 11076
rect 57848 11064 57854 11076
rect 57977 11067 58035 11073
rect 57977 11064 57989 11067
rect 57848 11036 57989 11064
rect 57848 11024 57854 11036
rect 57977 11033 57989 11036
rect 58023 11064 58035 11067
rect 62577 11067 62635 11073
rect 62577 11064 62589 11067
rect 58023 11036 62589 11064
rect 58023 11033 58035 11036
rect 57977 11027 58035 11033
rect 62577 11033 62589 11036
rect 62623 11033 62635 11067
rect 62577 11027 62635 11033
rect 65150 11024 65156 11076
rect 65208 11064 65214 11076
rect 65613 11067 65671 11073
rect 65613 11064 65625 11067
rect 65208 11036 65625 11064
rect 65208 11024 65214 11036
rect 65613 11033 65625 11036
rect 65659 11064 65671 11067
rect 69566 11064 69572 11076
rect 65659 11036 69572 11064
rect 65659 11033 65671 11036
rect 65613 11027 65671 11033
rect 69566 11024 69572 11036
rect 69624 11024 69630 11076
rect 69845 11067 69903 11073
rect 69845 11033 69857 11067
rect 69891 11064 69903 11067
rect 72896 11064 72924 11240
rect 76377 11237 76389 11240
rect 76423 11237 76435 11271
rect 76377 11231 76435 11237
rect 79134 11228 79140 11280
rect 79192 11268 79198 11280
rect 79192 11240 81940 11268
rect 79192 11228 79198 11240
rect 73522 11200 73528 11212
rect 73483 11172 73528 11200
rect 73522 11160 73528 11172
rect 73580 11160 73586 11212
rect 76190 11160 76196 11212
rect 76248 11200 76254 11212
rect 78309 11203 78367 11209
rect 78309 11200 78321 11203
rect 76248 11172 78321 11200
rect 76248 11160 76254 11172
rect 74077 11135 74135 11141
rect 74077 11101 74089 11135
rect 74123 11132 74135 11135
rect 74169 11135 74227 11141
rect 74169 11132 74181 11135
rect 74123 11104 74181 11132
rect 74123 11101 74135 11104
rect 74077 11095 74135 11101
rect 74169 11101 74181 11104
rect 74215 11101 74227 11135
rect 74169 11095 74227 11101
rect 74718 11092 74724 11144
rect 74776 11132 74782 11144
rect 74905 11135 74963 11141
rect 74905 11132 74917 11135
rect 74776 11104 74917 11132
rect 74776 11092 74782 11104
rect 74905 11101 74917 11104
rect 74951 11132 74963 11135
rect 75733 11135 75791 11141
rect 75733 11132 75745 11135
rect 74951 11104 75745 11132
rect 74951 11101 74963 11104
rect 74905 11095 74963 11101
rect 75733 11101 75745 11104
rect 75779 11101 75791 11135
rect 75733 11095 75791 11101
rect 76006 11092 76012 11144
rect 76064 11132 76070 11144
rect 76285 11135 76343 11141
rect 76285 11132 76297 11135
rect 76064 11104 76297 11132
rect 76064 11092 76070 11104
rect 76285 11101 76297 11104
rect 76331 11132 76343 11135
rect 76742 11132 76748 11144
rect 76331 11104 76748 11132
rect 76331 11101 76343 11104
rect 76285 11095 76343 11101
rect 76742 11092 76748 11104
rect 76800 11092 76806 11144
rect 76834 11092 76840 11144
rect 76892 11132 76898 11144
rect 77864 11141 77892 11172
rect 78309 11169 78321 11172
rect 78355 11169 78367 11203
rect 80422 11200 80428 11212
rect 80383 11172 80428 11200
rect 78309 11163 78367 11169
rect 80422 11160 80428 11172
rect 80480 11160 80486 11212
rect 81710 11200 81716 11212
rect 81671 11172 81716 11200
rect 81710 11160 81716 11172
rect 81768 11160 81774 11212
rect 77297 11135 77355 11141
rect 77297 11132 77309 11135
rect 76892 11104 77309 11132
rect 76892 11092 76898 11104
rect 77297 11101 77309 11104
rect 77343 11101 77355 11135
rect 77297 11095 77355 11101
rect 77849 11135 77907 11141
rect 77849 11101 77861 11135
rect 77895 11101 77907 11135
rect 77849 11095 77907 11101
rect 79413 11135 79471 11141
rect 79413 11101 79425 11135
rect 79459 11132 79471 11135
rect 80054 11132 80060 11144
rect 79459 11104 80060 11132
rect 79459 11101 79471 11104
rect 79413 11095 79471 11101
rect 80054 11092 80060 11104
rect 80112 11092 80118 11144
rect 81912 11141 81940 11240
rect 82446 11228 82452 11280
rect 82504 11268 82510 11280
rect 85393 11271 85451 11277
rect 85393 11268 85405 11271
rect 82504 11240 85405 11268
rect 82504 11228 82510 11240
rect 81986 11160 81992 11212
rect 82044 11200 82050 11212
rect 84381 11203 84439 11209
rect 84381 11200 84393 11203
rect 82044 11172 84393 11200
rect 82044 11160 82050 11172
rect 80977 11135 81035 11141
rect 80977 11101 80989 11135
rect 81023 11101 81035 11135
rect 80977 11095 81035 11101
rect 81897 11135 81955 11141
rect 81897 11101 81909 11135
rect 81943 11132 81955 11135
rect 82357 11135 82415 11141
rect 82357 11132 82369 11135
rect 81943 11104 82369 11132
rect 81943 11101 81955 11104
rect 81897 11095 81955 11101
rect 82357 11101 82369 11104
rect 82403 11101 82415 11135
rect 82906 11132 82912 11144
rect 82867 11104 82912 11132
rect 82357 11095 82415 11101
rect 74810 11064 74816 11076
rect 69891 11036 72924 11064
rect 74771 11036 74816 11064
rect 69891 11033 69903 11036
rect 69845 11027 69903 11033
rect 74810 11024 74816 11036
rect 74868 11024 74874 11076
rect 80992 11064 81020 11095
rect 82906 11092 82912 11104
rect 82964 11132 82970 11144
rect 83936 11141 83964 11172
rect 84381 11169 84393 11172
rect 84427 11169 84439 11203
rect 84381 11163 84439 11169
rect 84948 11141 84976 11240
rect 85393 11237 85405 11240
rect 85439 11237 85451 11271
rect 85393 11231 85451 11237
rect 92937 11271 92995 11277
rect 92937 11237 92949 11271
rect 92983 11268 92995 11271
rect 93302 11268 93308 11280
rect 92983 11240 93308 11268
rect 92983 11237 92995 11240
rect 92937 11231 92995 11237
rect 93302 11228 93308 11240
rect 93360 11268 93366 11280
rect 96798 11268 96804 11280
rect 93360 11240 96804 11268
rect 93360 11228 93366 11240
rect 96798 11228 96804 11240
rect 96856 11228 96862 11280
rect 96985 11271 97043 11277
rect 96985 11237 96997 11271
rect 97031 11268 97043 11271
rect 100941 11271 100999 11277
rect 97031 11240 100892 11268
rect 97031 11237 97043 11240
rect 96985 11231 97043 11237
rect 93121 11203 93179 11209
rect 93121 11169 93133 11203
rect 93167 11200 93179 11203
rect 93670 11200 93676 11212
rect 93167 11172 93676 11200
rect 93167 11169 93179 11172
rect 93121 11163 93179 11169
rect 93670 11160 93676 11172
rect 93728 11160 93734 11212
rect 93854 11160 93860 11212
rect 93912 11200 93918 11212
rect 94133 11203 94191 11209
rect 94133 11200 94145 11203
rect 93912 11172 94145 11200
rect 93912 11160 93918 11172
rect 94133 11169 94145 11172
rect 94179 11169 94191 11203
rect 95510 11200 95516 11212
rect 95471 11172 95516 11200
rect 94133 11163 94191 11169
rect 95510 11160 95516 11172
rect 95568 11160 95574 11212
rect 99466 11200 99472 11212
rect 99427 11172 99472 11200
rect 99466 11160 99472 11172
rect 99524 11160 99530 11212
rect 83737 11135 83795 11141
rect 83737 11132 83749 11135
rect 82964 11104 83749 11132
rect 82964 11092 82970 11104
rect 83737 11101 83749 11104
rect 83783 11101 83795 11135
rect 83737 11095 83795 11101
rect 83921 11135 83979 11141
rect 83921 11101 83933 11135
rect 83967 11101 83979 11135
rect 83921 11095 83979 11101
rect 84933 11135 84991 11141
rect 84933 11101 84945 11135
rect 84979 11101 84991 11135
rect 84933 11095 84991 11101
rect 94685 11135 94743 11141
rect 94685 11101 94697 11135
rect 94731 11101 94743 11135
rect 96614 11132 96620 11144
rect 96575 11104 96620 11132
rect 94685 11095 94743 11101
rect 81345 11067 81403 11073
rect 81345 11064 81357 11067
rect 77864 11036 78076 11064
rect 80992 11036 81357 11064
rect 51442 10996 51448 11008
rect 48332 10968 51448 10996
rect 51442 10956 51448 10968
rect 51500 10956 51506 11008
rect 51534 10956 51540 11008
rect 51592 10996 51598 11008
rect 53006 10996 53012 11008
rect 51592 10968 53012 10996
rect 51592 10956 51598 10968
rect 53006 10956 53012 10968
rect 53064 10956 53070 11008
rect 54481 10999 54539 11005
rect 54481 10965 54493 10999
rect 54527 10996 54539 10999
rect 54570 10996 54576 11008
rect 54527 10968 54576 10996
rect 54527 10965 54539 10968
rect 54481 10959 54539 10965
rect 54570 10956 54576 10968
rect 54628 10956 54634 11008
rect 55122 10956 55128 11008
rect 55180 10996 55186 11008
rect 57146 10996 57152 11008
rect 55180 10968 57152 10996
rect 55180 10956 55186 10968
rect 57146 10956 57152 10968
rect 57204 10956 57210 11008
rect 58066 10996 58072 11008
rect 58027 10968 58072 10996
rect 58066 10956 58072 10968
rect 58124 10956 58130 11008
rect 58434 10956 58440 11008
rect 58492 10996 58498 11008
rect 58529 10999 58587 11005
rect 58529 10996 58541 10999
rect 58492 10968 58541 10996
rect 58492 10956 58498 10968
rect 58529 10965 58541 10968
rect 58575 10965 58587 10999
rect 58529 10959 58587 10965
rect 60458 10956 60464 11008
rect 60516 10996 60522 11008
rect 61930 10996 61936 11008
rect 60516 10968 61936 10996
rect 60516 10956 60522 10968
rect 61930 10956 61936 10968
rect 61988 10956 61994 11008
rect 62482 10996 62488 11008
rect 62443 10968 62488 10996
rect 62482 10956 62488 10968
rect 62540 10956 62546 11008
rect 65061 10999 65119 11005
rect 65061 10965 65073 10999
rect 65107 10996 65119 10999
rect 65242 10996 65248 11008
rect 65107 10968 65248 10996
rect 65107 10965 65119 10968
rect 65061 10959 65119 10965
rect 65242 10956 65248 10968
rect 65300 10956 65306 11008
rect 65334 10956 65340 11008
rect 65392 10996 65398 11008
rect 77864 10996 77892 11036
rect 65392 10968 77892 10996
rect 78048 10996 78076 11036
rect 81345 11033 81357 11036
rect 81391 11064 81403 11067
rect 84013 11067 84071 11073
rect 84013 11064 84025 11067
rect 81391 11036 84025 11064
rect 81391 11033 81403 11036
rect 81345 11027 81403 11033
rect 84013 11033 84025 11036
rect 84059 11033 84071 11067
rect 84013 11027 84071 11033
rect 85025 11067 85083 11073
rect 85025 11033 85037 11067
rect 85071 11064 85083 11067
rect 85758 11064 85764 11076
rect 85071 11036 85764 11064
rect 85071 11033 85083 11036
rect 85025 11027 85083 11033
rect 85758 11024 85764 11036
rect 85816 11024 85822 11076
rect 87506 11064 87512 11076
rect 87467 11036 87512 11064
rect 87506 11024 87512 11036
rect 87564 11024 87570 11076
rect 91738 11064 91744 11076
rect 91699 11036 91744 11064
rect 91738 11024 91744 11036
rect 91796 11024 91802 11076
rect 92014 11064 92020 11076
rect 91975 11036 92020 11064
rect 92014 11024 92020 11036
rect 92072 11024 92078 11076
rect 94700 11064 94728 11095
rect 96614 11092 96620 11104
rect 96672 11132 96678 11144
rect 97353 11135 97411 11141
rect 97353 11132 97365 11135
rect 96672 11104 97365 11132
rect 96672 11092 96678 11104
rect 97353 11101 97365 11104
rect 97399 11101 97411 11135
rect 97353 11095 97411 11101
rect 100757 11135 100815 11141
rect 100757 11101 100769 11135
rect 100803 11101 100815 11135
rect 100864 11132 100892 11240
rect 100941 11237 100953 11271
rect 100987 11268 100999 11271
rect 108022 11268 108028 11280
rect 100987 11240 108028 11268
rect 100987 11237 100999 11240
rect 100941 11231 100999 11237
rect 108022 11228 108028 11240
rect 108080 11228 108086 11280
rect 108132 11277 108160 11308
rect 108117 11271 108175 11277
rect 108117 11237 108129 11271
rect 108163 11237 108175 11271
rect 108117 11231 108175 11237
rect 101858 11200 101864 11212
rect 101819 11172 101864 11200
rect 101858 11160 101864 11172
rect 101916 11160 101922 11212
rect 103146 11200 103152 11212
rect 103107 11172 103152 11200
rect 103146 11160 103152 11172
rect 103204 11160 103210 11212
rect 105633 11203 105691 11209
rect 103256 11172 104756 11200
rect 103256 11132 103284 11172
rect 100864 11104 103284 11132
rect 103425 11135 103483 11141
rect 100757 11095 100815 11101
rect 103425 11101 103437 11135
rect 103471 11101 103483 11135
rect 103425 11095 103483 11101
rect 104345 11135 104403 11141
rect 104345 11101 104357 11135
rect 104391 11132 104403 11135
rect 104621 11135 104679 11141
rect 104621 11132 104633 11135
rect 104391 11104 104633 11132
rect 104391 11101 104403 11104
rect 104345 11095 104403 11101
rect 104621 11101 104633 11104
rect 104667 11101 104679 11135
rect 104621 11095 104679 11101
rect 95053 11067 95111 11073
rect 95053 11064 95065 11067
rect 94700 11036 95065 11064
rect 95053 11033 95065 11036
rect 95099 11064 95111 11067
rect 100662 11064 100668 11076
rect 95099 11036 100668 11064
rect 95099 11033 95111 11036
rect 95053 11027 95111 11033
rect 100662 11024 100668 11036
rect 100720 11024 100726 11076
rect 100772 11064 100800 11095
rect 101125 11067 101183 11073
rect 101125 11064 101137 11067
rect 100772 11036 101137 11064
rect 101125 11033 101137 11036
rect 101171 11033 101183 11067
rect 103440 11064 103468 11095
rect 103793 11067 103851 11073
rect 103793 11064 103805 11067
rect 103440 11036 103805 11064
rect 101125 11027 101183 11033
rect 103793 11033 103805 11036
rect 103839 11064 103851 11067
rect 104437 11067 104495 11073
rect 104437 11064 104449 11067
rect 103839 11036 104449 11064
rect 103839 11033 103851 11036
rect 103793 11027 103851 11033
rect 104437 11033 104449 11036
rect 104483 11033 104495 11067
rect 104728 11064 104756 11172
rect 105633 11169 105645 11203
rect 105679 11200 105691 11203
rect 106645 11203 106703 11209
rect 106645 11200 106657 11203
rect 105679 11172 106657 11200
rect 105679 11169 105691 11172
rect 105633 11163 105691 11169
rect 106645 11169 106657 11172
rect 106691 11200 106703 11203
rect 107102 11200 107108 11212
rect 106691 11172 107108 11200
rect 106691 11169 106703 11172
rect 106645 11163 106703 11169
rect 107102 11160 107108 11172
rect 107160 11160 107166 11212
rect 110874 11160 110880 11212
rect 110932 11200 110938 11212
rect 111242 11200 111248 11212
rect 110932 11172 110977 11200
rect 111203 11172 111248 11200
rect 110932 11160 110938 11172
rect 111242 11160 111248 11172
rect 111300 11160 111306 11212
rect 108206 11132 108212 11144
rect 108167 11104 108212 11132
rect 108206 11092 108212 11104
rect 108264 11092 108270 11144
rect 108574 11132 108580 11144
rect 108535 11104 108580 11132
rect 108574 11092 108580 11104
rect 108632 11092 108638 11144
rect 109957 11135 110015 11141
rect 109957 11101 109969 11135
rect 110003 11132 110015 11135
rect 110506 11132 110512 11144
rect 110003 11104 110512 11132
rect 110003 11101 110015 11104
rect 109957 11095 110015 11101
rect 110506 11092 110512 11104
rect 110564 11092 110570 11144
rect 110049 11067 110107 11073
rect 104728 11036 110000 11064
rect 104437 11027 104495 11033
rect 78306 10996 78312 11008
rect 78048 10968 78312 10996
rect 65392 10956 65398 10968
rect 78306 10956 78312 10968
rect 78364 10956 78370 11008
rect 85942 10996 85948 11008
rect 85903 10968 85948 10996
rect 85942 10956 85948 10968
rect 86000 10956 86006 11008
rect 90358 10996 90364 11008
rect 90319 10968 90364 10996
rect 90358 10956 90364 10968
rect 90416 10956 90422 11008
rect 107746 10956 107752 11008
rect 107804 10996 107810 11008
rect 108574 10996 108580 11008
rect 107804 10968 108580 10996
rect 107804 10956 107810 10968
rect 108574 10956 108580 10968
rect 108632 10956 108638 11008
rect 109034 10956 109040 11008
rect 109092 10996 109098 11008
rect 109972 10996 110000 11036
rect 110049 11033 110061 11067
rect 110095 11064 110107 11067
rect 110966 11064 110972 11076
rect 110095 11036 110972 11064
rect 110095 11033 110107 11036
rect 110049 11027 110107 11033
rect 110966 11024 110972 11036
rect 111024 11024 111030 11076
rect 111444 11064 111472 11308
rect 112901 11305 112913 11339
rect 112947 11336 112959 11339
rect 113177 11339 113235 11345
rect 113177 11336 113189 11339
rect 112947 11308 113189 11336
rect 112947 11305 112959 11308
rect 112901 11299 112959 11305
rect 113177 11305 113189 11308
rect 113223 11336 113235 11339
rect 118602 11336 118608 11348
rect 113223 11308 118608 11336
rect 113223 11305 113235 11308
rect 113177 11299 113235 11305
rect 118602 11296 118608 11308
rect 118660 11296 118666 11348
rect 121270 11336 121276 11348
rect 121231 11308 121276 11336
rect 121270 11296 121276 11308
rect 121328 11296 121334 11348
rect 121457 11339 121515 11345
rect 121457 11305 121469 11339
rect 121503 11336 121515 11339
rect 121730 11336 121736 11348
rect 121503 11308 121736 11336
rect 121503 11305 121515 11308
rect 121457 11299 121515 11305
rect 121730 11296 121736 11308
rect 121788 11296 121794 11348
rect 121914 11296 121920 11348
rect 121972 11336 121978 11348
rect 122009 11339 122067 11345
rect 122009 11336 122021 11339
rect 121972 11308 122021 11336
rect 121972 11296 121978 11308
rect 122009 11305 122021 11308
rect 122055 11305 122067 11339
rect 123110 11336 123116 11348
rect 123071 11308 123116 11336
rect 122009 11299 122067 11305
rect 123110 11296 123116 11308
rect 123168 11296 123174 11348
rect 124217 11339 124275 11345
rect 124217 11305 124229 11339
rect 124263 11336 124275 11339
rect 124306 11336 124312 11348
rect 124263 11308 124312 11336
rect 124263 11305 124275 11308
rect 124217 11299 124275 11305
rect 124306 11296 124312 11308
rect 124364 11296 124370 11348
rect 127158 11336 127164 11348
rect 125612 11308 127164 11336
rect 112717 11271 112775 11277
rect 112717 11237 112729 11271
rect 112763 11268 112775 11271
rect 114462 11268 114468 11280
rect 112763 11240 114468 11268
rect 112763 11237 112775 11240
rect 112717 11231 112775 11237
rect 114462 11228 114468 11240
rect 114520 11228 114526 11280
rect 123021 11271 123079 11277
rect 123021 11268 123033 11271
rect 114848 11240 123033 11268
rect 112990 11160 112996 11212
rect 113048 11200 113054 11212
rect 113545 11203 113603 11209
rect 113545 11200 113557 11203
rect 113048 11172 113557 11200
rect 113048 11160 113054 11172
rect 113545 11169 113557 11172
rect 113591 11200 113603 11203
rect 114848 11200 114876 11240
rect 123021 11237 123033 11240
rect 123067 11237 123079 11271
rect 123386 11268 123392 11280
rect 123347 11240 123392 11268
rect 123021 11231 123079 11237
rect 123386 11228 123392 11240
rect 123444 11228 123450 11280
rect 123573 11271 123631 11277
rect 123573 11237 123585 11271
rect 123619 11268 123631 11271
rect 123849 11271 123907 11277
rect 123849 11268 123861 11271
rect 123619 11240 123861 11268
rect 123619 11237 123631 11240
rect 123573 11231 123631 11237
rect 123849 11237 123861 11240
rect 123895 11268 123907 11271
rect 125502 11268 125508 11280
rect 123895 11240 125508 11268
rect 123895 11237 123907 11240
rect 123849 11231 123907 11237
rect 125502 11228 125508 11240
rect 125560 11228 125566 11280
rect 115014 11200 115020 11212
rect 113591 11172 114876 11200
rect 114975 11172 115020 11200
rect 113591 11169 113603 11172
rect 113545 11163 113603 11169
rect 115014 11160 115020 11172
rect 115072 11160 115078 11212
rect 115198 11160 115204 11212
rect 115256 11200 115262 11212
rect 116581 11203 116639 11209
rect 116581 11200 116593 11203
rect 115256 11172 116593 11200
rect 115256 11160 115262 11172
rect 116581 11169 116593 11172
rect 116627 11169 116639 11203
rect 117958 11200 117964 11212
rect 117919 11172 117964 11200
rect 116581 11163 116639 11169
rect 117958 11160 117964 11172
rect 118016 11160 118022 11212
rect 118694 11160 118700 11212
rect 118752 11200 118758 11212
rect 118973 11203 119031 11209
rect 118973 11200 118985 11203
rect 118752 11172 118985 11200
rect 118752 11160 118758 11172
rect 118973 11169 118985 11172
rect 119019 11169 119031 11203
rect 122926 11200 122932 11212
rect 118973 11163 119031 11169
rect 119448 11172 122932 11200
rect 112809 11135 112867 11141
rect 112809 11101 112821 11135
rect 112855 11132 112867 11135
rect 112901 11135 112959 11141
rect 112901 11132 112913 11135
rect 112855 11104 112913 11132
rect 112855 11101 112867 11104
rect 112809 11095 112867 11101
rect 112901 11101 112913 11104
rect 112947 11101 112959 11135
rect 112901 11095 112959 11101
rect 114465 11135 114523 11141
rect 114465 11101 114477 11135
rect 114511 11132 114523 11135
rect 115032 11132 115060 11160
rect 114511 11104 115060 11132
rect 115385 11135 115443 11141
rect 114511 11101 114523 11104
rect 114465 11095 114523 11101
rect 115385 11101 115397 11135
rect 115431 11132 115443 11135
rect 115566 11132 115572 11144
rect 115431 11104 115572 11132
rect 115431 11101 115443 11104
rect 115385 11095 115443 11101
rect 115566 11092 115572 11104
rect 115624 11092 115630 11144
rect 117133 11135 117191 11141
rect 117133 11101 117145 11135
rect 117179 11101 117191 11135
rect 117133 11095 117191 11101
rect 113726 11064 113732 11076
rect 111444 11036 113732 11064
rect 113726 11024 113732 11036
rect 113784 11024 113790 11076
rect 114373 11067 114431 11073
rect 114373 11033 114385 11067
rect 114419 11064 114431 11067
rect 114646 11064 114652 11076
rect 114419 11036 114652 11064
rect 114419 11033 114431 11036
rect 114373 11027 114431 11033
rect 114646 11024 114652 11036
rect 114704 11064 114710 11076
rect 116578 11064 116584 11076
rect 114704 11036 116584 11064
rect 114704 11024 114710 11036
rect 116578 11024 116584 11036
rect 116636 11024 116642 11076
rect 117148 11064 117176 11095
rect 117501 11067 117559 11073
rect 117501 11064 117513 11067
rect 117148 11036 117513 11064
rect 117501 11033 117513 11036
rect 117547 11064 117559 11067
rect 119448 11064 119476 11172
rect 122926 11160 122932 11172
rect 122984 11160 122990 11212
rect 125318 11200 125324 11212
rect 123036 11172 124812 11200
rect 125279 11172 125324 11200
rect 119525 11135 119583 11141
rect 119525 11101 119537 11135
rect 119571 11132 119583 11135
rect 119893 11135 119951 11141
rect 119893 11132 119905 11135
rect 119571 11104 119905 11132
rect 119571 11101 119583 11104
rect 119525 11095 119583 11101
rect 119893 11101 119905 11104
rect 119939 11132 119951 11135
rect 121181 11135 121239 11141
rect 119939 11104 121132 11132
rect 119939 11101 119951 11104
rect 119893 11095 119951 11101
rect 120258 11064 120264 11076
rect 117547 11036 119476 11064
rect 120219 11036 120264 11064
rect 117547 11033 117559 11036
rect 117501 11027 117559 11033
rect 120258 11024 120264 11036
rect 120316 11024 120322 11076
rect 121104 11064 121132 11104
rect 121181 11101 121193 11135
rect 121227 11132 121239 11135
rect 121457 11135 121515 11141
rect 121457 11132 121469 11135
rect 121227 11104 121469 11132
rect 121227 11101 121239 11104
rect 121181 11095 121239 11101
rect 121457 11101 121469 11104
rect 121503 11101 121515 11135
rect 123036 11132 123064 11172
rect 121457 11095 121515 11101
rect 122024 11104 123064 11132
rect 123297 11135 123355 11141
rect 122024 11064 122052 11104
rect 123297 11101 123309 11135
rect 123343 11132 123355 11135
rect 123573 11135 123631 11141
rect 123573 11132 123585 11135
rect 123343 11104 123585 11132
rect 123343 11101 123355 11104
rect 123297 11095 123355 11101
rect 123573 11101 123585 11104
rect 123619 11101 123631 11135
rect 123573 11095 123631 11101
rect 124309 11135 124367 11141
rect 124309 11101 124321 11135
rect 124355 11132 124367 11135
rect 124674 11132 124680 11144
rect 124355 11104 124680 11132
rect 124355 11101 124367 11104
rect 124309 11095 124367 11101
rect 124674 11092 124680 11104
rect 124732 11092 124738 11144
rect 124784 11132 124812 11172
rect 125318 11160 125324 11172
rect 125376 11160 125382 11212
rect 125612 11132 125640 11308
rect 127158 11296 127164 11308
rect 127216 11296 127222 11348
rect 127710 11336 127716 11348
rect 127671 11308 127716 11336
rect 127710 11296 127716 11308
rect 127768 11296 127774 11348
rect 130470 11336 130476 11348
rect 130431 11308 130476 11336
rect 130470 11296 130476 11308
rect 130528 11296 130534 11348
rect 132497 11339 132555 11345
rect 132497 11305 132509 11339
rect 132543 11336 132555 11339
rect 133230 11336 133236 11348
rect 132543 11308 133236 11336
rect 132543 11305 132555 11308
rect 132497 11299 132555 11305
rect 133230 11296 133236 11308
rect 133288 11296 133294 11348
rect 136082 11336 136088 11348
rect 136043 11308 136088 11336
rect 136082 11296 136088 11308
rect 136140 11296 136146 11348
rect 137186 11296 137192 11348
rect 137244 11336 137250 11348
rect 137465 11339 137523 11345
rect 137465 11336 137477 11339
rect 137244 11308 137477 11336
rect 137244 11296 137250 11308
rect 137465 11305 137477 11308
rect 137511 11305 137523 11339
rect 137465 11299 137523 11305
rect 141053 11339 141111 11345
rect 141053 11305 141065 11339
rect 141099 11336 141111 11339
rect 144546 11336 144552 11348
rect 141099 11308 144552 11336
rect 141099 11305 141111 11308
rect 141053 11299 141111 11305
rect 126146 11268 126152 11280
rect 126107 11240 126152 11268
rect 126146 11228 126152 11240
rect 126204 11228 126210 11280
rect 128541 11271 128599 11277
rect 128541 11237 128553 11271
rect 128587 11268 128599 11271
rect 131942 11268 131948 11280
rect 128587 11240 131948 11268
rect 128587 11237 128599 11240
rect 128541 11231 128599 11237
rect 124784 11104 125640 11132
rect 125873 11135 125931 11141
rect 125873 11101 125885 11135
rect 125919 11132 125931 11135
rect 126164 11132 126192 11228
rect 126333 11203 126391 11209
rect 126333 11169 126345 11203
rect 126379 11200 126391 11203
rect 126885 11203 126943 11209
rect 126885 11200 126897 11203
rect 126379 11172 126897 11200
rect 126379 11169 126391 11172
rect 126333 11163 126391 11169
rect 126885 11169 126897 11172
rect 126931 11169 126943 11203
rect 126885 11163 126943 11169
rect 125919 11104 126192 11132
rect 125919 11101 125931 11104
rect 125873 11095 125931 11101
rect 126238 11092 126244 11144
rect 126296 11132 126302 11144
rect 126793 11135 126851 11141
rect 126793 11132 126805 11135
rect 126296 11104 126805 11132
rect 126296 11092 126302 11104
rect 126793 11101 126805 11104
rect 126839 11132 126851 11135
rect 127253 11135 127311 11141
rect 127253 11132 127265 11135
rect 126839 11104 127265 11132
rect 126839 11101 126851 11104
rect 126793 11095 126851 11101
rect 127253 11101 127265 11104
rect 127299 11101 127311 11135
rect 128556 11132 128584 11231
rect 131942 11228 131948 11240
rect 132000 11228 132006 11280
rect 135622 11228 135628 11280
rect 135680 11268 135686 11280
rect 139305 11271 139363 11277
rect 135680 11240 139256 11268
rect 135680 11228 135686 11240
rect 129645 11203 129703 11209
rect 129645 11200 129657 11203
rect 128740 11172 129657 11200
rect 128633 11135 128691 11141
rect 128633 11132 128645 11135
rect 128556 11104 128645 11132
rect 127253 11095 127311 11101
rect 128633 11101 128645 11104
rect 128679 11101 128691 11135
rect 128633 11095 128691 11101
rect 122190 11064 122196 11076
rect 121104 11036 122052 11064
rect 122151 11036 122196 11064
rect 122190 11024 122196 11036
rect 122248 11024 122254 11076
rect 123021 11067 123079 11073
rect 123021 11033 123033 11067
rect 123067 11064 123079 11067
rect 126333 11067 126391 11073
rect 126333 11064 126345 11067
rect 123067 11036 126345 11064
rect 123067 11033 123079 11036
rect 123021 11027 123079 11033
rect 126333 11033 126345 11036
rect 126379 11033 126391 11067
rect 126333 11027 126391 11033
rect 126609 11067 126667 11073
rect 126609 11033 126621 11067
rect 126655 11064 126667 11067
rect 126974 11064 126980 11076
rect 126655 11036 126980 11064
rect 126655 11033 126667 11036
rect 126609 11027 126667 11033
rect 126974 11024 126980 11036
rect 127032 11064 127038 11076
rect 127802 11064 127808 11076
rect 127032 11036 127808 11064
rect 127032 11024 127038 11036
rect 127802 11024 127808 11036
rect 127860 11024 127866 11076
rect 127894 11024 127900 11076
rect 127952 11064 127958 11076
rect 128740 11064 128768 11172
rect 129645 11169 129657 11172
rect 129691 11169 129703 11203
rect 129645 11163 129703 11169
rect 130286 11160 130292 11212
rect 130344 11200 130350 11212
rect 132865 11203 132923 11209
rect 132865 11200 132877 11203
rect 130344 11172 132877 11200
rect 130344 11160 130350 11172
rect 130194 11132 130200 11144
rect 130155 11104 130200 11132
rect 130194 11092 130200 11104
rect 130252 11092 130258 11144
rect 132420 11141 132448 11172
rect 132865 11169 132877 11172
rect 132911 11169 132923 11203
rect 135254 11200 135260 11212
rect 135215 11172 135260 11200
rect 132865 11163 132923 11169
rect 135254 11160 135260 11172
rect 135312 11160 135318 11212
rect 137462 11160 137468 11212
rect 137520 11200 137526 11212
rect 139228 11200 139256 11240
rect 139305 11237 139317 11271
rect 139351 11268 139363 11271
rect 139486 11268 139492 11280
rect 139351 11240 139492 11268
rect 139351 11237 139363 11240
rect 139305 11231 139363 11237
rect 139486 11228 139492 11240
rect 139544 11228 139550 11280
rect 140866 11200 140872 11212
rect 137520 11172 139164 11200
rect 139228 11172 140872 11200
rect 137520 11160 137526 11172
rect 131025 11135 131083 11141
rect 131025 11132 131037 11135
rect 130488 11104 131037 11132
rect 127952 11036 128768 11064
rect 127952 11024 127958 11036
rect 128814 11024 128820 11076
rect 128872 11064 128878 11076
rect 130488 11064 130516 11104
rect 131025 11101 131037 11104
rect 131071 11132 131083 11135
rect 131485 11135 131543 11141
rect 131485 11132 131497 11135
rect 131071 11104 131497 11132
rect 131071 11101 131083 11104
rect 131025 11095 131083 11101
rect 131485 11101 131497 11104
rect 131531 11101 131543 11135
rect 131485 11095 131543 11101
rect 132405 11135 132463 11141
rect 132405 11101 132417 11135
rect 132451 11101 132463 11135
rect 132405 11095 132463 11101
rect 134245 11135 134303 11141
rect 134245 11101 134257 11135
rect 134291 11132 134303 11135
rect 134334 11132 134340 11144
rect 134291 11104 134340 11132
rect 134291 11101 134303 11104
rect 134245 11095 134303 11101
rect 134334 11092 134340 11104
rect 134392 11132 134398 11144
rect 135162 11132 135168 11144
rect 134392 11104 135168 11132
rect 134392 11092 134398 11104
rect 135162 11092 135168 11104
rect 135220 11092 135226 11144
rect 135809 11135 135867 11141
rect 135809 11101 135821 11135
rect 135855 11132 135867 11135
rect 135990 11132 135996 11144
rect 135855 11104 135996 11132
rect 135855 11101 135867 11104
rect 135809 11095 135867 11101
rect 135990 11092 135996 11104
rect 136048 11092 136054 11144
rect 136634 11132 136640 11144
rect 136595 11104 136640 11132
rect 136634 11092 136640 11104
rect 136692 11132 136698 11144
rect 137097 11135 137155 11141
rect 137097 11132 137109 11135
rect 136692 11104 137109 11132
rect 136692 11092 136698 11104
rect 137097 11101 137109 11104
rect 137143 11101 137155 11135
rect 137097 11095 137155 11101
rect 138017 11135 138075 11141
rect 138017 11101 138029 11135
rect 138063 11132 138075 11135
rect 138106 11132 138112 11144
rect 138063 11104 138112 11132
rect 138063 11101 138075 11104
rect 138017 11095 138075 11101
rect 138106 11092 138112 11104
rect 138164 11092 138170 11144
rect 139136 11141 139164 11172
rect 140866 11160 140872 11172
rect 140924 11160 140930 11212
rect 141160 11209 141188 11308
rect 144546 11296 144552 11308
rect 144604 11296 144610 11348
rect 144822 11296 144828 11348
rect 144880 11336 144886 11348
rect 144880 11308 152412 11336
rect 144880 11296 144886 11308
rect 141234 11228 141240 11280
rect 141292 11268 141298 11280
rect 150434 11268 150440 11280
rect 141292 11240 144684 11268
rect 150395 11240 150440 11268
rect 141292 11228 141298 11240
rect 141145 11203 141203 11209
rect 141145 11169 141157 11203
rect 141191 11169 141203 11203
rect 141145 11163 141203 11169
rect 142338 11160 142344 11212
rect 142396 11200 142402 11212
rect 144656 11209 144684 11240
rect 150434 11228 150440 11240
rect 150492 11228 150498 11280
rect 144641 11203 144699 11209
rect 142396 11172 142441 11200
rect 142396 11160 142402 11172
rect 144641 11169 144653 11203
rect 144687 11169 144699 11203
rect 146478 11200 146484 11212
rect 146439 11172 146484 11200
rect 144641 11163 144699 11169
rect 146478 11160 146484 11172
rect 146536 11160 146542 11212
rect 147490 11200 147496 11212
rect 147451 11172 147496 11200
rect 147490 11160 147496 11172
rect 147548 11160 147554 11212
rect 149517 11203 149575 11209
rect 149517 11169 149529 11203
rect 149563 11200 149575 11203
rect 150529 11203 150587 11209
rect 150529 11200 150541 11203
rect 149563 11172 150541 11200
rect 149563 11169 149575 11172
rect 149517 11163 149575 11169
rect 150529 11169 150541 11172
rect 150575 11200 150587 11203
rect 150986 11200 150992 11212
rect 150575 11172 150992 11200
rect 150575 11169 150587 11172
rect 150529 11163 150587 11169
rect 150986 11160 150992 11172
rect 151044 11160 151050 11212
rect 151538 11200 151544 11212
rect 151499 11172 151544 11200
rect 151538 11160 151544 11172
rect 151596 11160 151602 11212
rect 152384 11200 152412 11308
rect 156138 11296 156144 11348
rect 156196 11336 156202 11348
rect 156233 11339 156291 11345
rect 156233 11336 156245 11339
rect 156196 11308 156245 11336
rect 156196 11296 156202 11308
rect 156233 11305 156245 11308
rect 156279 11305 156291 11339
rect 160186 11336 160192 11348
rect 160147 11308 160192 11336
rect 156233 11299 156291 11305
rect 160186 11296 160192 11308
rect 160244 11296 160250 11348
rect 162210 11296 162216 11348
rect 162268 11336 162274 11348
rect 162305 11339 162363 11345
rect 162305 11336 162317 11339
rect 162268 11308 162317 11336
rect 162268 11296 162274 11308
rect 162305 11305 162317 11308
rect 162351 11305 162363 11339
rect 165890 11336 165896 11348
rect 165851 11308 165896 11336
rect 162305 11299 162363 11305
rect 165890 11296 165896 11308
rect 165948 11296 165954 11348
rect 153286 11228 153292 11280
rect 153344 11268 153350 11280
rect 153344 11240 167132 11268
rect 153344 11228 153350 11240
rect 157889 11203 157947 11209
rect 157889 11200 157901 11203
rect 152384 11172 157901 11200
rect 157889 11169 157901 11172
rect 157935 11169 157947 11203
rect 163866 11200 163872 11212
rect 163827 11172 163872 11200
rect 157889 11163 157947 11169
rect 163866 11160 163872 11172
rect 163924 11160 163930 11212
rect 166074 11200 166080 11212
rect 166035 11172 166080 11200
rect 166074 11160 166080 11172
rect 166132 11160 166138 11212
rect 167104 11209 167132 11240
rect 167089 11203 167147 11209
rect 167089 11169 167101 11203
rect 167135 11169 167147 11203
rect 167089 11163 167147 11169
rect 139121 11135 139179 11141
rect 139121 11101 139133 11135
rect 139167 11132 139179 11135
rect 139857 11135 139915 11141
rect 139857 11132 139869 11135
rect 139167 11104 139869 11132
rect 139167 11101 139179 11104
rect 139121 11095 139179 11101
rect 139857 11101 139869 11104
rect 139903 11101 139915 11135
rect 142249 11135 142307 11141
rect 142249 11132 142261 11135
rect 139857 11095 139915 11101
rect 140056 11104 142261 11132
rect 131114 11064 131120 11076
rect 128872 11036 130516 11064
rect 131075 11036 131120 11064
rect 128872 11024 128878 11036
rect 131114 11024 131120 11036
rect 131172 11024 131178 11076
rect 131945 11067 132003 11073
rect 131945 11033 131957 11067
rect 131991 11064 132003 11067
rect 132494 11064 132500 11076
rect 131991 11036 132500 11064
rect 131991 11033 132003 11036
rect 131945 11027 132003 11033
rect 132494 11024 132500 11036
rect 132552 11064 132558 11076
rect 133138 11064 133144 11076
rect 132552 11036 133144 11064
rect 132552 11024 132558 11036
rect 133138 11024 133144 11036
rect 133196 11024 133202 11076
rect 136729 11067 136787 11073
rect 136729 11033 136741 11067
rect 136775 11064 136787 11067
rect 140056 11064 140084 11104
rect 142249 11101 142261 11104
rect 142295 11132 142307 11135
rect 142985 11135 143043 11141
rect 142985 11132 142997 11135
rect 142295 11104 142997 11132
rect 142295 11101 142307 11104
rect 142249 11095 142307 11101
rect 142985 11101 142997 11104
rect 143031 11101 143043 11135
rect 143350 11132 143356 11144
rect 143311 11104 143356 11132
rect 142985 11095 143043 11101
rect 143350 11092 143356 11104
rect 143408 11092 143414 11144
rect 143629 11135 143687 11141
rect 143629 11101 143641 11135
rect 143675 11132 143687 11135
rect 143994 11132 144000 11144
rect 143675 11104 144000 11132
rect 143675 11101 143687 11104
rect 143629 11095 143687 11101
rect 140222 11064 140228 11076
rect 136775 11036 140084 11064
rect 140183 11036 140228 11064
rect 136775 11033 136787 11036
rect 136729 11027 136787 11033
rect 140222 11024 140228 11036
rect 140280 11024 140286 11076
rect 140682 11024 140688 11076
rect 140740 11064 140746 11076
rect 143644 11064 143672 11095
rect 143994 11092 144000 11104
rect 144052 11092 144058 11144
rect 145006 11132 145012 11144
rect 144967 11104 145012 11132
rect 145006 11092 145012 11104
rect 145064 11132 145070 11144
rect 145469 11135 145527 11141
rect 145469 11132 145481 11135
rect 145064 11104 145481 11132
rect 145064 11092 145070 11104
rect 145469 11101 145481 11104
rect 145515 11101 145527 11135
rect 145469 11095 145527 11101
rect 146938 11092 146944 11144
rect 146996 11132 147002 11144
rect 147585 11135 147643 11141
rect 147585 11132 147597 11135
rect 146996 11104 147597 11132
rect 146996 11092 147002 11104
rect 147585 11101 147597 11104
rect 147631 11132 147643 11135
rect 148321 11135 148379 11141
rect 148321 11132 148333 11135
rect 147631 11104 148333 11132
rect 147631 11101 147643 11104
rect 147585 11095 147643 11101
rect 148321 11101 148333 11104
rect 148367 11101 148379 11135
rect 151630 11132 151636 11144
rect 151591 11104 151636 11132
rect 148321 11095 148379 11101
rect 151630 11092 151636 11104
rect 151688 11092 151694 11144
rect 152369 11135 152427 11141
rect 152369 11132 152381 11135
rect 151740 11104 152381 11132
rect 140740 11036 143672 11064
rect 140740 11024 140746 11036
rect 150710 11024 150716 11076
rect 150768 11064 150774 11076
rect 151446 11064 151452 11076
rect 150768 11036 151452 11064
rect 150768 11024 150774 11036
rect 151446 11024 151452 11036
rect 151504 11064 151510 11076
rect 151740 11064 151768 11104
rect 152369 11101 152381 11104
rect 152415 11101 152427 11135
rect 156874 11132 156880 11144
rect 156835 11104 156880 11132
rect 152369 11095 152427 11101
rect 156874 11092 156880 11104
rect 156932 11092 156938 11144
rect 157426 11092 157432 11144
rect 157484 11132 157490 11144
rect 157981 11135 158039 11141
rect 157981 11132 157993 11135
rect 157484 11104 157993 11132
rect 157484 11092 157490 11104
rect 157981 11101 157993 11104
rect 158027 11132 158039 11135
rect 158717 11135 158775 11141
rect 158717 11132 158729 11135
rect 158027 11104 158729 11132
rect 158027 11101 158039 11104
rect 157981 11095 158039 11101
rect 158717 11101 158729 11104
rect 158763 11101 158775 11135
rect 162857 11135 162915 11141
rect 162857 11132 162869 11135
rect 158717 11095 158775 11101
rect 162688 11104 162869 11132
rect 151504 11036 151768 11064
rect 151504 11024 151510 11036
rect 151814 11024 151820 11076
rect 151872 11064 151878 11076
rect 152921 11067 152979 11073
rect 152921 11064 152933 11067
rect 151872 11036 152933 11064
rect 151872 11024 151878 11036
rect 152921 11033 152933 11036
rect 152967 11033 152979 11067
rect 152921 11027 152979 11033
rect 154114 11024 154120 11076
rect 154172 11064 154178 11076
rect 154482 11064 154488 11076
rect 154172 11036 154488 11064
rect 154172 11024 154178 11036
rect 154482 11024 154488 11036
rect 154540 11024 154546 11076
rect 162688 11073 162716 11104
rect 162857 11101 162869 11104
rect 162903 11101 162915 11135
rect 162857 11095 162915 11101
rect 163038 11092 163044 11144
rect 163096 11132 163102 11144
rect 163961 11135 164019 11141
rect 163961 11132 163973 11135
rect 163096 11104 163973 11132
rect 163096 11092 163102 11104
rect 163961 11101 163973 11104
rect 164007 11132 164019 11135
rect 164697 11135 164755 11141
rect 164697 11132 164709 11135
rect 164007 11104 164709 11132
rect 164007 11101 164019 11104
rect 163961 11095 164019 11101
rect 164697 11101 164709 11104
rect 164743 11101 164755 11135
rect 167178 11132 167184 11144
rect 167139 11104 167184 11132
rect 164697 11095 164755 11101
rect 167178 11092 167184 11104
rect 167236 11132 167242 11144
rect 167917 11135 167975 11141
rect 167917 11132 167929 11135
rect 167236 11104 167929 11132
rect 167236 11092 167242 11104
rect 167917 11101 167929 11104
rect 167963 11101 167975 11135
rect 167917 11095 167975 11101
rect 161845 11067 161903 11073
rect 161845 11033 161857 11067
rect 161891 11064 161903 11067
rect 162673 11067 162731 11073
rect 162673 11064 162685 11067
rect 161891 11036 162685 11064
rect 161891 11033 161903 11036
rect 161845 11027 161903 11033
rect 162673 11033 162685 11036
rect 162719 11033 162731 11067
rect 162673 11027 162731 11033
rect 110782 10996 110788 11008
rect 109092 10968 109137 10996
rect 109972 10968 110788 10996
rect 109092 10956 109098 10968
rect 110782 10956 110788 10968
rect 110840 10956 110846 11008
rect 110874 10956 110880 11008
rect 110932 10996 110938 11008
rect 111886 10996 111892 11008
rect 110932 10968 111892 10996
rect 110932 10956 110938 10968
rect 111886 10956 111892 10968
rect 111944 10956 111950 11008
rect 114554 10996 114560 11008
rect 114515 10968 114560 10996
rect 114554 10956 114560 10968
rect 114612 10956 114618 11008
rect 117774 10956 117780 11008
rect 117832 10996 117838 11008
rect 119706 10996 119712 11008
rect 117832 10968 119712 10996
rect 117832 10956 117838 10968
rect 119706 10956 119712 10968
rect 119764 10956 119770 11008
rect 120442 10956 120448 11008
rect 120500 10996 120506 11008
rect 128262 10996 128268 11008
rect 120500 10968 128268 10996
rect 120500 10956 120506 10968
rect 128262 10956 128268 10968
rect 128320 10956 128326 11008
rect 155129 10999 155187 11005
rect 155129 10965 155141 10999
rect 155175 10996 155187 10999
rect 155310 10996 155316 11008
rect 155175 10968 155316 10996
rect 155175 10965 155187 10968
rect 155129 10959 155187 10965
rect 155310 10956 155316 10968
rect 155368 10956 155374 11008
rect 159266 10996 159272 11008
rect 159227 10968 159272 10996
rect 159266 10956 159272 10968
rect 159324 10956 159330 11008
rect 368 10906 169556 10928
rect 368 10854 56667 10906
rect 56719 10854 56731 10906
rect 56783 10854 56795 10906
rect 56847 10854 56859 10906
rect 56911 10854 113088 10906
rect 113140 10854 113152 10906
rect 113204 10854 113216 10906
rect 113268 10854 113280 10906
rect 113332 10854 169556 10906
rect 368 10832 169556 10854
rect 6270 10792 6276 10804
rect 6231 10764 6276 10792
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 9732 10764 10149 10792
rect 9732 10752 9738 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 23566 10792 23572 10804
rect 23479 10764 23572 10792
rect 10137 10755 10195 10761
rect 23566 10752 23572 10764
rect 23624 10792 23630 10804
rect 24670 10792 24676 10804
rect 23624 10764 24676 10792
rect 23624 10752 23630 10764
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 25792 10764 26004 10792
rect 24489 10727 24547 10733
rect 14200 10696 19840 10724
rect 3694 10616 3700 10668
rect 3752 10656 3758 10668
rect 3970 10656 3976 10668
rect 3752 10628 3976 10656
rect 3752 10616 3758 10628
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4338 10656 4344 10668
rect 4299 10628 4344 10656
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 4798 10656 4804 10668
rect 4755 10628 4804 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 5074 10656 5080 10668
rect 5035 10628 5080 10656
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 12618 10656 12624 10668
rect 12579 10628 12624 10656
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14200 10665 14228 10696
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 14056 10628 14197 10656
rect 14056 10616 14062 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10625 18751 10659
rect 19702 10656 19708 10668
rect 19663 10628 19708 10656
rect 18693 10619 18751 10625
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 6733 10591 6791 10597
rect 3375 10560 4016 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3988 10464 4016 10560
rect 6733 10557 6745 10591
rect 6779 10588 6791 10591
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 6779 10560 7757 10588
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 7745 10557 7757 10560
rect 7791 10588 7803 10591
rect 8294 10588 8300 10600
rect 7791 10560 8300 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10588 16267 10591
rect 17310 10588 17316 10600
rect 16255 10560 17316 10588
rect 16255 10557 16267 10560
rect 16209 10551 16267 10557
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 9217 10523 9275 10529
rect 9217 10489 9229 10523
rect 9263 10520 9275 10523
rect 14093 10523 14151 10529
rect 9263 10492 13124 10520
rect 9263 10489 9275 10492
rect 9217 10483 9275 10489
rect 3970 10452 3976 10464
rect 3931 10424 3976 10452
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 13096 10452 13124 10492
rect 14093 10489 14105 10523
rect 14139 10520 14151 10523
rect 18046 10520 18052 10532
rect 14139 10492 18052 10520
rect 14139 10489 14151 10492
rect 14093 10483 14151 10489
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 18414 10480 18420 10532
rect 18472 10520 18478 10532
rect 18601 10523 18659 10529
rect 18601 10520 18613 10523
rect 18472 10492 18613 10520
rect 18472 10480 18478 10492
rect 18601 10489 18613 10492
rect 18647 10489 18659 10523
rect 18601 10483 18659 10489
rect 18708 10464 18736 10619
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 19812 10656 19840 10696
rect 24489 10693 24501 10727
rect 24535 10724 24547 10727
rect 25792 10724 25820 10764
rect 24535 10696 25820 10724
rect 25976 10724 26004 10764
rect 26050 10752 26056 10804
rect 26108 10792 26114 10804
rect 51166 10792 51172 10804
rect 26108 10764 51172 10792
rect 26108 10752 26114 10764
rect 51166 10752 51172 10764
rect 51224 10752 51230 10804
rect 51258 10752 51264 10804
rect 51316 10792 51322 10804
rect 60458 10792 60464 10804
rect 51316 10764 60464 10792
rect 51316 10752 51322 10764
rect 60458 10752 60464 10764
rect 60516 10752 60522 10804
rect 60645 10795 60703 10801
rect 60645 10761 60657 10795
rect 60691 10792 60703 10795
rect 60734 10792 60740 10804
rect 60691 10764 60740 10792
rect 60691 10761 60703 10764
rect 60645 10755 60703 10761
rect 28810 10724 28816 10736
rect 25976 10696 28816 10724
rect 24535 10693 24547 10696
rect 24489 10687 24547 10693
rect 28810 10684 28816 10696
rect 28868 10684 28874 10736
rect 29086 10724 29092 10736
rect 28920 10696 29092 10724
rect 21269 10659 21327 10665
rect 19812 10628 20852 10656
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 18840 10560 20729 10588
rect 18840 10548 18846 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20824 10588 20852 10628
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 21634 10656 21640 10668
rect 21315 10628 21640 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 21634 10616 21640 10628
rect 21692 10616 21698 10668
rect 24397 10659 24455 10665
rect 24397 10625 24409 10659
rect 24443 10656 24455 10659
rect 24762 10656 24768 10668
rect 24443 10628 24768 10656
rect 24443 10625 24455 10628
rect 24397 10619 24455 10625
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 25866 10656 25872 10668
rect 25827 10628 25872 10656
rect 25866 10616 25872 10628
rect 25924 10616 25930 10668
rect 26053 10659 26111 10665
rect 26053 10625 26065 10659
rect 26099 10656 26111 10659
rect 27246 10656 27252 10668
rect 26099 10628 27252 10656
rect 26099 10625 26111 10628
rect 26053 10619 26111 10625
rect 27246 10616 27252 10628
rect 27304 10616 27310 10668
rect 27430 10656 27436 10668
rect 27391 10628 27436 10656
rect 27430 10616 27436 10628
rect 27488 10616 27494 10668
rect 27709 10659 27767 10665
rect 27709 10625 27721 10659
rect 27755 10656 27767 10659
rect 28920 10656 28948 10696
rect 29086 10684 29092 10696
rect 29144 10684 29150 10736
rect 30558 10724 30564 10736
rect 29380 10696 30564 10724
rect 27755 10628 28948 10656
rect 27755 10625 27767 10628
rect 27709 10619 27767 10625
rect 28994 10616 29000 10668
rect 29052 10656 29058 10668
rect 29273 10659 29331 10665
rect 29052 10628 29097 10656
rect 29052 10616 29058 10628
rect 29273 10625 29285 10659
rect 29319 10656 29331 10659
rect 29380 10656 29408 10696
rect 30558 10684 30564 10696
rect 30616 10684 30622 10736
rect 30837 10727 30895 10733
rect 30837 10693 30849 10727
rect 30883 10724 30895 10727
rect 31662 10724 31668 10736
rect 30883 10696 31668 10724
rect 30883 10693 30895 10696
rect 30837 10687 30895 10693
rect 31662 10684 31668 10696
rect 31720 10684 31726 10736
rect 32401 10727 32459 10733
rect 32401 10693 32413 10727
rect 32447 10724 32459 10727
rect 32766 10724 32772 10736
rect 32447 10696 32772 10724
rect 32447 10693 32459 10696
rect 32401 10687 32459 10693
rect 32766 10684 32772 10696
rect 32824 10684 32830 10736
rect 33870 10684 33876 10736
rect 33928 10724 33934 10736
rect 34517 10727 34575 10733
rect 34517 10724 34529 10727
rect 33928 10696 34529 10724
rect 33928 10684 33934 10696
rect 34517 10693 34529 10696
rect 34563 10693 34575 10727
rect 41966 10724 41972 10736
rect 34517 10687 34575 10693
rect 34624 10696 41972 10724
rect 30742 10656 30748 10668
rect 29319 10628 29408 10656
rect 30703 10628 30748 10656
rect 29319 10625 29331 10628
rect 29273 10619 29331 10625
rect 30742 10616 30748 10628
rect 30800 10616 30806 10668
rect 31386 10616 31392 10668
rect 31444 10656 31450 10668
rect 32214 10656 32220 10668
rect 31444 10628 31800 10656
rect 32175 10628 32220 10656
rect 31444 10616 31450 10628
rect 20824 10560 24256 10588
rect 20717 10551 20775 10557
rect 16574 10452 16580 10464
rect 13096 10424 16580 10452
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 18690 10452 18696 10464
rect 18603 10424 18696 10452
rect 18690 10412 18696 10424
rect 18748 10452 18754 10464
rect 24118 10452 24124 10464
rect 18748 10424 24124 10452
rect 18748 10412 18754 10424
rect 24118 10412 24124 10424
rect 24176 10412 24182 10464
rect 24228 10452 24256 10560
rect 27798 10548 27804 10600
rect 27856 10588 27862 10600
rect 29454 10588 29460 10600
rect 27856 10560 29460 10588
rect 27856 10548 27862 10560
rect 29454 10548 29460 10560
rect 29512 10548 29518 10600
rect 29546 10548 29552 10600
rect 29604 10588 29610 10600
rect 31772 10588 31800 10628
rect 32214 10616 32220 10628
rect 32272 10616 32278 10668
rect 32306 10616 32312 10668
rect 32364 10656 32370 10668
rect 34624 10656 34652 10696
rect 41966 10684 41972 10696
rect 42024 10684 42030 10736
rect 42058 10684 42064 10736
rect 42116 10724 42122 10736
rect 42334 10724 42340 10736
rect 42116 10696 42340 10724
rect 42116 10684 42122 10696
rect 42334 10684 42340 10696
rect 42392 10684 42398 10736
rect 42426 10684 42432 10736
rect 42484 10684 42490 10736
rect 45373 10727 45431 10733
rect 45373 10693 45385 10727
rect 45419 10724 45431 10727
rect 45830 10724 45836 10736
rect 45419 10696 45836 10724
rect 45419 10693 45431 10696
rect 45373 10687 45431 10693
rect 45830 10684 45836 10696
rect 45888 10684 45894 10736
rect 47397 10727 47455 10733
rect 47397 10724 47409 10727
rect 46400 10696 47409 10724
rect 35158 10656 35164 10668
rect 32364 10628 34652 10656
rect 35119 10628 35164 10656
rect 32364 10616 32370 10628
rect 35158 10616 35164 10628
rect 35216 10616 35222 10668
rect 35342 10616 35348 10668
rect 35400 10656 35406 10668
rect 37458 10656 37464 10668
rect 35400 10628 37228 10656
rect 37419 10628 37464 10656
rect 35400 10616 35406 10628
rect 35618 10588 35624 10600
rect 29604 10560 31708 10588
rect 31772 10560 35624 10588
rect 29604 10548 29610 10560
rect 24302 10480 24308 10532
rect 24360 10520 24366 10532
rect 31570 10520 31576 10532
rect 24360 10492 31576 10520
rect 24360 10480 24366 10492
rect 31570 10480 31576 10492
rect 31628 10480 31634 10532
rect 31680 10520 31708 10560
rect 35618 10548 35624 10560
rect 35676 10548 35682 10600
rect 36078 10588 36084 10600
rect 36039 10560 36084 10588
rect 36078 10548 36084 10560
rect 36136 10548 36142 10600
rect 36354 10548 36360 10600
rect 36412 10588 36418 10600
rect 36998 10588 37004 10600
rect 36412 10560 37004 10588
rect 36412 10548 36418 10560
rect 36998 10548 37004 10560
rect 37056 10548 37062 10600
rect 37093 10591 37151 10597
rect 37093 10557 37105 10591
rect 37139 10557 37151 10591
rect 37093 10551 37151 10557
rect 37108 10520 37136 10551
rect 31680 10492 37136 10520
rect 37200 10520 37228 10628
rect 37458 10616 37464 10628
rect 37516 10616 37522 10668
rect 37550 10616 37556 10668
rect 37608 10656 37614 10668
rect 41046 10656 41052 10668
rect 37608 10628 41052 10656
rect 37608 10616 37614 10628
rect 41046 10616 41052 10628
rect 41104 10616 41110 10668
rect 41141 10659 41199 10665
rect 41141 10625 41153 10659
rect 41187 10656 41199 10659
rect 41598 10656 41604 10668
rect 41187 10628 41604 10656
rect 41187 10625 41199 10628
rect 41141 10619 41199 10625
rect 41598 10616 41604 10628
rect 41656 10616 41662 10668
rect 41690 10616 41696 10668
rect 41748 10656 41754 10668
rect 41748 10628 42288 10656
rect 41748 10616 41754 10628
rect 37642 10548 37648 10600
rect 37700 10588 37706 10600
rect 38013 10591 38071 10597
rect 38013 10588 38025 10591
rect 37700 10560 38025 10588
rect 37700 10548 37706 10560
rect 38013 10557 38025 10560
rect 38059 10588 38071 10591
rect 38473 10591 38531 10597
rect 38473 10588 38485 10591
rect 38059 10560 38485 10588
rect 38059 10557 38071 10560
rect 38013 10551 38071 10557
rect 38473 10557 38485 10560
rect 38519 10557 38531 10591
rect 38473 10551 38531 10557
rect 38580 10560 42196 10588
rect 38580 10520 38608 10560
rect 37200 10492 38608 10520
rect 38654 10480 38660 10532
rect 38712 10520 38718 10532
rect 41690 10520 41696 10532
rect 38712 10492 41696 10520
rect 38712 10480 38718 10492
rect 41690 10480 41696 10492
rect 41748 10480 41754 10532
rect 41782 10480 41788 10532
rect 41840 10520 41846 10532
rect 41966 10520 41972 10532
rect 41840 10492 41972 10520
rect 41840 10480 41846 10492
rect 41966 10480 41972 10492
rect 42024 10480 42030 10532
rect 26142 10452 26148 10464
rect 24228 10424 26148 10452
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 27341 10455 27399 10461
rect 27341 10421 27353 10455
rect 27387 10452 27399 10455
rect 27430 10452 27436 10464
rect 27387 10424 27436 10452
rect 27387 10421 27399 10424
rect 27341 10415 27399 10421
rect 27430 10412 27436 10424
rect 27488 10412 27494 10464
rect 27522 10412 27528 10464
rect 27580 10452 27586 10464
rect 27709 10455 27767 10461
rect 27709 10452 27721 10455
rect 27580 10424 27721 10452
rect 27580 10412 27586 10424
rect 27709 10421 27721 10424
rect 27755 10421 27767 10455
rect 27709 10415 27767 10421
rect 27798 10412 27804 10464
rect 27856 10452 27862 10464
rect 27893 10455 27951 10461
rect 27893 10452 27905 10455
rect 27856 10424 27905 10452
rect 27856 10412 27862 10424
rect 27893 10421 27905 10424
rect 27939 10421 27951 10455
rect 27893 10415 27951 10421
rect 27982 10412 27988 10464
rect 28040 10452 28046 10464
rect 31478 10452 31484 10464
rect 28040 10424 31484 10452
rect 28040 10412 28046 10424
rect 31478 10412 31484 10424
rect 31536 10412 31542 10464
rect 32582 10412 32588 10464
rect 32640 10452 32646 10464
rect 32677 10455 32735 10461
rect 32677 10452 32689 10455
rect 32640 10424 32689 10452
rect 32640 10412 32646 10424
rect 32677 10421 32689 10424
rect 32723 10421 32735 10455
rect 32677 10415 32735 10421
rect 35066 10412 35072 10464
rect 35124 10452 35130 10464
rect 35529 10455 35587 10461
rect 35529 10452 35541 10455
rect 35124 10424 35541 10452
rect 35124 10412 35130 10424
rect 35529 10421 35541 10424
rect 35575 10421 35587 10455
rect 35529 10415 35587 10421
rect 35618 10412 35624 10464
rect 35676 10452 35682 10464
rect 42058 10452 42064 10464
rect 35676 10424 42064 10452
rect 35676 10412 35682 10424
rect 42058 10412 42064 10424
rect 42116 10412 42122 10464
rect 42168 10452 42196 10560
rect 42260 10520 42288 10628
rect 42444 10597 42472 10684
rect 46400 10668 46428 10696
rect 47397 10693 47409 10696
rect 47443 10693 47455 10727
rect 47397 10687 47455 10693
rect 47504 10696 51396 10724
rect 42705 10659 42763 10665
rect 42705 10625 42717 10659
rect 42751 10625 42763 10659
rect 42705 10619 42763 10625
rect 42429 10591 42487 10597
rect 42429 10557 42441 10591
rect 42475 10557 42487 10591
rect 42720 10588 42748 10619
rect 43346 10616 43352 10668
rect 43404 10656 43410 10668
rect 46382 10656 46388 10668
rect 43404 10628 46152 10656
rect 46343 10628 46388 10656
rect 43404 10616 43410 10628
rect 43162 10588 43168 10600
rect 42720 10560 43168 10588
rect 42429 10551 42487 10557
rect 43162 10548 43168 10560
rect 43220 10548 43226 10600
rect 44269 10591 44327 10597
rect 44269 10557 44281 10591
rect 44315 10588 44327 10591
rect 45830 10588 45836 10600
rect 44315 10560 45836 10588
rect 44315 10557 44327 10560
rect 44269 10551 44327 10557
rect 45830 10548 45836 10560
rect 45888 10588 45894 10600
rect 46017 10591 46075 10597
rect 46017 10588 46029 10591
rect 45888 10560 46029 10588
rect 45888 10548 45894 10560
rect 46017 10557 46029 10560
rect 46063 10557 46075 10591
rect 46124 10588 46152 10628
rect 46382 10616 46388 10628
rect 46440 10616 46446 10668
rect 47118 10656 47124 10668
rect 47079 10628 47124 10656
rect 47118 10616 47124 10628
rect 47176 10616 47182 10668
rect 47504 10588 47532 10696
rect 47949 10659 48007 10665
rect 47949 10625 47961 10659
rect 47995 10656 48007 10659
rect 48222 10656 48228 10668
rect 47995 10628 48228 10656
rect 47995 10625 48007 10628
rect 47949 10619 48007 10625
rect 48222 10616 48228 10628
rect 48280 10616 48286 10668
rect 49513 10659 49571 10665
rect 49513 10625 49525 10659
rect 49559 10656 49571 10659
rect 49694 10656 49700 10668
rect 49559 10628 49700 10656
rect 49559 10625 49571 10628
rect 49513 10619 49571 10625
rect 49694 10616 49700 10628
rect 49752 10656 49758 10668
rect 50614 10656 50620 10668
rect 49752 10628 50620 10656
rect 49752 10616 49758 10628
rect 50614 10616 50620 10628
rect 50672 10616 50678 10668
rect 50706 10616 50712 10668
rect 50764 10656 50770 10668
rect 51077 10659 51135 10665
rect 51077 10656 51089 10659
rect 50764 10628 51089 10656
rect 50764 10616 50770 10628
rect 51077 10625 51089 10628
rect 51123 10625 51135 10659
rect 51368 10656 51396 10696
rect 51442 10684 51448 10736
rect 51500 10724 51506 10736
rect 55306 10724 55312 10736
rect 51500 10696 55312 10724
rect 51500 10684 51506 10696
rect 55306 10684 55312 10696
rect 55364 10684 55370 10736
rect 55769 10727 55827 10733
rect 55769 10724 55781 10727
rect 55508 10696 55781 10724
rect 51718 10656 51724 10668
rect 51368 10628 51488 10656
rect 51679 10628 51724 10656
rect 51077 10619 51135 10625
rect 48958 10588 48964 10600
rect 46124 10560 47532 10588
rect 48919 10560 48964 10588
rect 46017 10551 46075 10557
rect 48958 10548 48964 10560
rect 49016 10548 49022 10600
rect 49050 10548 49056 10600
rect 49108 10588 49114 10600
rect 51353 10591 51411 10597
rect 51353 10588 51365 10591
rect 49108 10560 51365 10588
rect 49108 10548 49114 10560
rect 51353 10557 51365 10560
rect 51399 10557 51411 10591
rect 51460 10588 51488 10628
rect 51718 10616 51724 10628
rect 51776 10616 51782 10668
rect 51810 10616 51816 10668
rect 51868 10656 51874 10668
rect 52362 10656 52368 10668
rect 51868 10628 52368 10656
rect 51868 10616 51874 10628
rect 52362 10616 52368 10628
rect 52420 10656 52426 10668
rect 52549 10659 52607 10665
rect 52549 10656 52561 10659
rect 52420 10628 52561 10656
rect 52420 10616 52426 10628
rect 52549 10625 52561 10628
rect 52595 10625 52607 10659
rect 52549 10619 52607 10625
rect 53285 10659 53343 10665
rect 53285 10625 53297 10659
rect 53331 10656 53343 10659
rect 53466 10656 53472 10668
rect 53331 10628 53472 10656
rect 53331 10625 53343 10628
rect 53285 10619 53343 10625
rect 53466 10616 53472 10628
rect 53524 10616 53530 10668
rect 54938 10656 54944 10668
rect 54899 10628 54944 10656
rect 54938 10616 54944 10628
rect 54996 10616 55002 10668
rect 55508 10665 55536 10696
rect 55769 10693 55781 10696
rect 55815 10693 55827 10727
rect 55769 10687 55827 10693
rect 55858 10684 55864 10736
rect 55916 10724 55922 10736
rect 56045 10727 56103 10733
rect 56045 10724 56057 10727
rect 55916 10696 56057 10724
rect 55916 10684 55922 10696
rect 56045 10693 56057 10696
rect 56091 10724 56103 10727
rect 58066 10724 58072 10736
rect 56091 10696 58072 10724
rect 56091 10693 56103 10696
rect 56045 10687 56103 10693
rect 58066 10684 58072 10696
rect 58124 10684 58130 10736
rect 60660 10724 60688 10755
rect 60734 10752 60740 10764
rect 60792 10752 60798 10804
rect 60918 10752 60924 10804
rect 60976 10792 60982 10804
rect 61746 10792 61752 10804
rect 60976 10764 61752 10792
rect 60976 10752 60982 10764
rect 61746 10752 61752 10764
rect 61804 10752 61810 10804
rect 63770 10752 63776 10804
rect 63828 10792 63834 10804
rect 71682 10792 71688 10804
rect 63828 10764 71688 10792
rect 63828 10752 63834 10764
rect 71682 10752 71688 10764
rect 71740 10752 71746 10804
rect 71774 10752 71780 10804
rect 71832 10792 71838 10804
rect 72053 10795 72111 10801
rect 72053 10792 72065 10795
rect 71832 10764 72065 10792
rect 71832 10752 71838 10764
rect 72053 10761 72065 10764
rect 72099 10761 72111 10795
rect 72053 10755 72111 10761
rect 73246 10752 73252 10804
rect 73304 10792 73310 10804
rect 74350 10792 74356 10804
rect 73304 10764 74356 10792
rect 73304 10752 73310 10764
rect 74350 10752 74356 10764
rect 74408 10752 74414 10804
rect 74534 10752 74540 10804
rect 74592 10792 74598 10804
rect 75089 10795 75147 10801
rect 75089 10792 75101 10795
rect 74592 10764 75101 10792
rect 74592 10752 74598 10764
rect 75089 10761 75101 10764
rect 75135 10761 75147 10795
rect 75089 10755 75147 10761
rect 78030 10752 78036 10804
rect 78088 10792 78094 10804
rect 78309 10795 78367 10801
rect 78309 10792 78321 10795
rect 78088 10764 78321 10792
rect 78088 10752 78094 10764
rect 78309 10761 78321 10764
rect 78355 10761 78367 10795
rect 78309 10755 78367 10761
rect 82906 10752 82912 10804
rect 82964 10792 82970 10804
rect 83093 10795 83151 10801
rect 83093 10792 83105 10795
rect 82964 10764 83105 10792
rect 82964 10752 82970 10764
rect 83093 10761 83105 10764
rect 83139 10792 83151 10795
rect 83918 10792 83924 10804
rect 83139 10764 83924 10792
rect 83139 10761 83151 10764
rect 83093 10755 83151 10761
rect 83918 10752 83924 10764
rect 83976 10752 83982 10804
rect 86954 10792 86960 10804
rect 86915 10764 86960 10792
rect 86954 10752 86960 10764
rect 87012 10792 87018 10804
rect 87012 10764 87092 10792
rect 87012 10752 87018 10764
rect 70670 10724 70676 10736
rect 60200 10696 60688 10724
rect 69400 10696 70676 10724
rect 55493 10659 55551 10665
rect 55493 10625 55505 10659
rect 55539 10625 55551 10659
rect 56226 10656 56232 10668
rect 55493 10619 55551 10625
rect 55692 10628 56232 10656
rect 55692 10588 55720 10628
rect 56226 10616 56232 10628
rect 56284 10616 56290 10668
rect 56410 10616 56416 10668
rect 56468 10656 56474 10668
rect 57149 10659 57207 10665
rect 56468 10628 57100 10656
rect 56468 10616 56474 10628
rect 51460 10560 55720 10588
rect 55769 10591 55827 10597
rect 51353 10551 51411 10557
rect 55769 10557 55781 10591
rect 55815 10588 55827 10591
rect 56962 10588 56968 10600
rect 55815 10560 56968 10588
rect 55815 10557 55827 10560
rect 55769 10551 55827 10557
rect 56962 10548 56968 10560
rect 57020 10548 57026 10600
rect 57072 10588 57100 10628
rect 57149 10625 57161 10659
rect 57195 10656 57207 10659
rect 57882 10656 57888 10668
rect 57195 10628 57888 10656
rect 57195 10625 57207 10628
rect 57149 10619 57207 10625
rect 57882 10616 57888 10628
rect 57940 10616 57946 10668
rect 58713 10659 58771 10665
rect 58713 10625 58725 10659
rect 58759 10656 58771 10659
rect 59446 10656 59452 10668
rect 58759 10628 59452 10656
rect 58759 10625 58771 10628
rect 58713 10619 58771 10625
rect 59446 10616 59452 10628
rect 59504 10616 59510 10668
rect 59817 10659 59875 10665
rect 59817 10625 59829 10659
rect 59863 10656 59875 10659
rect 60200 10656 60228 10696
rect 69400 10668 69428 10696
rect 70670 10684 70676 10696
rect 70728 10684 70734 10736
rect 72510 10684 72516 10736
rect 72568 10724 72574 10736
rect 80422 10724 80428 10736
rect 72568 10696 74028 10724
rect 72568 10684 72574 10696
rect 59863 10628 60228 10656
rect 60277 10659 60335 10665
rect 59863 10625 59875 10628
rect 59817 10619 59875 10625
rect 60277 10625 60289 10659
rect 60323 10625 60335 10659
rect 60277 10619 60335 10625
rect 57072 10560 57560 10588
rect 46477 10523 46535 10529
rect 46477 10520 46489 10523
rect 42260 10492 46489 10520
rect 46477 10489 46489 10492
rect 46523 10489 46535 10523
rect 46477 10483 46535 10489
rect 46566 10480 46572 10532
rect 46624 10520 46630 10532
rect 46624 10492 56456 10520
rect 46624 10480 46630 10492
rect 43346 10452 43352 10464
rect 42168 10424 43352 10452
rect 43346 10412 43352 10424
rect 43404 10412 43410 10464
rect 45554 10412 45560 10464
rect 45612 10452 45618 10464
rect 49786 10452 49792 10464
rect 45612 10424 49792 10452
rect 45612 10412 45618 10424
rect 49786 10412 49792 10424
rect 49844 10412 49850 10464
rect 49970 10412 49976 10464
rect 50028 10452 50034 10464
rect 50028 10424 50073 10452
rect 50028 10412 50034 10424
rect 50154 10412 50160 10464
rect 50212 10452 50218 10464
rect 51442 10452 51448 10464
rect 50212 10424 51448 10452
rect 50212 10412 50218 10424
rect 51442 10412 51448 10424
rect 51500 10412 51506 10464
rect 51626 10412 51632 10464
rect 51684 10452 51690 10464
rect 51997 10455 52055 10461
rect 51997 10452 52009 10455
rect 51684 10424 52009 10452
rect 51684 10412 51690 10424
rect 51997 10421 52009 10424
rect 52043 10421 52055 10455
rect 51997 10415 52055 10421
rect 52641 10455 52699 10461
rect 52641 10421 52653 10455
rect 52687 10452 52699 10455
rect 52822 10452 52828 10464
rect 52687 10424 52828 10452
rect 52687 10421 52699 10424
rect 52641 10415 52699 10421
rect 52822 10412 52828 10424
rect 52880 10412 52886 10464
rect 55033 10455 55091 10461
rect 55033 10421 55045 10455
rect 55079 10452 55091 10455
rect 55214 10452 55220 10464
rect 55079 10424 55220 10452
rect 55079 10421 55091 10424
rect 55033 10415 55091 10421
rect 55214 10412 55220 10424
rect 55272 10412 55278 10464
rect 55490 10412 55496 10464
rect 55548 10452 55554 10464
rect 56042 10452 56048 10464
rect 55548 10424 56048 10452
rect 55548 10412 55554 10424
rect 56042 10412 56048 10424
rect 56100 10412 56106 10464
rect 56318 10452 56324 10464
rect 56279 10424 56324 10452
rect 56318 10412 56324 10424
rect 56376 10412 56382 10464
rect 56428 10452 56456 10492
rect 56502 10480 56508 10532
rect 56560 10520 56566 10532
rect 57422 10520 57428 10532
rect 56560 10492 57428 10520
rect 56560 10480 56566 10492
rect 57422 10480 57428 10492
rect 57480 10480 57486 10532
rect 57532 10520 57560 10560
rect 57974 10548 57980 10600
rect 58032 10588 58038 10600
rect 59909 10591 59967 10597
rect 59909 10588 59921 10591
rect 58032 10560 59921 10588
rect 58032 10548 58038 10560
rect 59909 10557 59921 10560
rect 59955 10557 59967 10591
rect 60292 10588 60320 10619
rect 60642 10616 60648 10668
rect 60700 10656 60706 10668
rect 62209 10659 62267 10665
rect 62209 10656 62221 10659
rect 60700 10628 62221 10656
rect 60700 10616 60706 10628
rect 62209 10625 62221 10628
rect 62255 10625 62267 10659
rect 62209 10619 62267 10625
rect 62298 10616 62304 10668
rect 62356 10656 62362 10668
rect 65334 10656 65340 10668
rect 62356 10628 65340 10656
rect 62356 10616 62362 10628
rect 65334 10616 65340 10628
rect 65392 10616 65398 10668
rect 66254 10656 66260 10668
rect 66215 10628 66260 10656
rect 66254 10616 66260 10628
rect 66312 10616 66318 10668
rect 67818 10616 67824 10668
rect 67876 10656 67882 10668
rect 68649 10659 68707 10665
rect 68649 10656 68661 10659
rect 67876 10628 68661 10656
rect 67876 10616 67882 10628
rect 68649 10625 68661 10628
rect 68695 10656 68707 10659
rect 68738 10656 68744 10668
rect 68695 10628 68744 10656
rect 68695 10625 68707 10628
rect 68649 10619 68707 10625
rect 68738 10616 68744 10628
rect 68796 10616 68802 10668
rect 69382 10656 69388 10668
rect 69295 10628 69388 10656
rect 69382 10616 69388 10628
rect 69440 10616 69446 10668
rect 70213 10659 70271 10665
rect 70213 10625 70225 10659
rect 70259 10656 70271 10659
rect 70486 10656 70492 10668
rect 70259 10628 70492 10656
rect 70259 10625 70271 10628
rect 70213 10619 70271 10625
rect 70486 10616 70492 10628
rect 70544 10616 70550 10668
rect 71777 10659 71835 10665
rect 71777 10625 71789 10659
rect 71823 10656 71835 10659
rect 71869 10659 71927 10665
rect 71869 10656 71881 10659
rect 71823 10628 71881 10656
rect 71823 10625 71835 10628
rect 71777 10619 71835 10625
rect 71869 10625 71881 10628
rect 71915 10625 71927 10659
rect 73614 10656 73620 10668
rect 73575 10628 73620 10656
rect 71869 10619 71927 10625
rect 73614 10616 73620 10628
rect 73672 10616 73678 10668
rect 74000 10665 74028 10696
rect 74552 10696 80428 10724
rect 73985 10659 74043 10665
rect 73985 10625 73997 10659
rect 74031 10656 74043 10659
rect 74442 10656 74448 10668
rect 74031 10628 74448 10656
rect 74031 10625 74043 10628
rect 73985 10619 74043 10625
rect 74442 10616 74448 10628
rect 74500 10616 74506 10668
rect 60734 10588 60740 10600
rect 60292 10560 60740 10588
rect 59909 10551 59967 10557
rect 60734 10548 60740 10560
rect 60792 10588 60798 10600
rect 60918 10588 60924 10600
rect 60792 10560 60924 10588
rect 60792 10548 60798 10560
rect 60918 10548 60924 10560
rect 60976 10548 60982 10600
rect 61105 10591 61163 10597
rect 61105 10557 61117 10591
rect 61151 10557 61163 10591
rect 61105 10551 61163 10557
rect 58437 10523 58495 10529
rect 58437 10520 58449 10523
rect 57532 10492 58449 10520
rect 58437 10489 58449 10492
rect 58483 10489 58495 10523
rect 58437 10483 58495 10489
rect 58544 10492 60320 10520
rect 58544 10452 58572 10492
rect 56428 10424 58572 10452
rect 58618 10412 58624 10464
rect 58676 10452 58682 10464
rect 60182 10452 60188 10464
rect 58676 10424 60188 10452
rect 58676 10412 58682 10424
rect 60182 10412 60188 10424
rect 60240 10412 60246 10464
rect 60292 10452 60320 10492
rect 60366 10480 60372 10532
rect 60424 10520 60430 10532
rect 61120 10520 61148 10551
rect 61930 10548 61936 10600
rect 61988 10588 61994 10600
rect 63221 10591 63279 10597
rect 63221 10588 63233 10591
rect 61988 10560 63233 10588
rect 61988 10548 61994 10560
rect 63221 10557 63233 10560
rect 63267 10557 63279 10591
rect 63221 10551 63279 10557
rect 64877 10591 64935 10597
rect 64877 10557 64889 10591
rect 64923 10588 64935 10591
rect 65242 10588 65248 10600
rect 64923 10560 65248 10588
rect 64923 10557 64935 10560
rect 64877 10551 64935 10557
rect 65242 10548 65248 10560
rect 65300 10548 65306 10600
rect 74552 10588 74580 10696
rect 80422 10684 80428 10696
rect 80480 10684 80486 10736
rect 82633 10727 82691 10733
rect 82633 10724 82645 10727
rect 81728 10696 82645 10724
rect 74997 10659 75055 10665
rect 74997 10625 75009 10659
rect 75043 10656 75055 10659
rect 75086 10656 75092 10668
rect 75043 10628 75092 10656
rect 75043 10625 75055 10628
rect 74997 10619 75055 10625
rect 75086 10616 75092 10628
rect 75144 10616 75150 10668
rect 77665 10659 77723 10665
rect 77665 10625 77677 10659
rect 77711 10625 77723 10659
rect 77665 10619 77723 10625
rect 65352 10560 73568 10588
rect 65352 10520 65380 10560
rect 66162 10520 66168 10532
rect 60424 10492 61148 10520
rect 61488 10492 65380 10520
rect 66123 10492 66168 10520
rect 60424 10480 60430 10492
rect 61488 10452 61516 10492
rect 66162 10480 66168 10492
rect 66220 10480 66226 10532
rect 66346 10480 66352 10532
rect 66404 10520 66410 10532
rect 68741 10523 68799 10529
rect 68741 10520 68753 10523
rect 66404 10492 68753 10520
rect 66404 10480 66410 10492
rect 68741 10489 68753 10492
rect 68787 10489 68799 10523
rect 71498 10520 71504 10532
rect 71459 10492 71504 10520
rect 68741 10483 68799 10489
rect 71498 10480 71504 10492
rect 71556 10480 71562 10532
rect 71869 10523 71927 10529
rect 71869 10489 71881 10523
rect 71915 10520 71927 10523
rect 72050 10520 72056 10532
rect 71915 10492 72056 10520
rect 71915 10489 71927 10492
rect 71869 10483 71927 10489
rect 72050 10480 72056 10492
rect 72108 10520 72114 10532
rect 73540 10529 73568 10560
rect 73632 10560 74580 10588
rect 76193 10591 76251 10597
rect 73525 10523 73583 10529
rect 72108 10492 72556 10520
rect 72108 10480 72114 10492
rect 61654 10452 61660 10464
rect 60292 10424 61516 10452
rect 61615 10424 61660 10452
rect 61654 10412 61660 10424
rect 61712 10412 61718 10464
rect 72418 10452 72424 10464
rect 72379 10424 72424 10452
rect 72418 10412 72424 10424
rect 72476 10412 72482 10464
rect 72528 10452 72556 10492
rect 73525 10489 73537 10523
rect 73571 10489 73583 10523
rect 73525 10483 73583 10489
rect 73632 10452 73660 10560
rect 76193 10557 76205 10591
rect 76239 10588 76251 10591
rect 76282 10588 76288 10600
rect 76239 10560 76288 10588
rect 76239 10557 76251 10560
rect 76193 10551 76251 10557
rect 76282 10548 76288 10560
rect 76340 10548 76346 10600
rect 77386 10588 77392 10600
rect 77347 10560 77392 10588
rect 77386 10548 77392 10560
rect 77444 10548 77450 10600
rect 77680 10588 77708 10619
rect 77754 10616 77760 10668
rect 77812 10656 77818 10668
rect 79042 10656 79048 10668
rect 77812 10628 79048 10656
rect 77812 10616 77818 10628
rect 79042 10616 79048 10628
rect 79100 10616 79106 10668
rect 81526 10616 81532 10668
rect 81584 10656 81590 10668
rect 81728 10665 81756 10696
rect 82633 10693 82645 10696
rect 82679 10693 82691 10727
rect 82633 10687 82691 10693
rect 81713 10659 81771 10665
rect 81713 10656 81725 10659
rect 81584 10628 81725 10656
rect 81584 10616 81590 10628
rect 81713 10625 81725 10628
rect 81759 10625 81771 10659
rect 81713 10619 81771 10625
rect 82541 10659 82599 10665
rect 82541 10625 82553 10659
rect 82587 10625 82599 10659
rect 82541 10619 82599 10625
rect 80149 10591 80207 10597
rect 77680 10560 78260 10588
rect 78232 10532 78260 10560
rect 80149 10557 80161 10591
rect 80195 10588 80207 10591
rect 80238 10588 80244 10600
rect 80195 10560 80244 10588
rect 80195 10557 80207 10560
rect 80149 10551 80207 10557
rect 80238 10548 80244 10560
rect 80296 10548 80302 10600
rect 81158 10588 81164 10600
rect 81119 10560 81164 10588
rect 81158 10548 81164 10560
rect 81216 10548 81222 10600
rect 81434 10548 81440 10600
rect 81492 10588 81498 10600
rect 82556 10588 82584 10619
rect 83182 10616 83188 10668
rect 83240 10656 83246 10668
rect 83550 10656 83556 10668
rect 83240 10628 83556 10656
rect 83240 10616 83246 10628
rect 83550 10616 83556 10628
rect 83608 10616 83614 10668
rect 85758 10656 85764 10668
rect 85719 10628 85764 10656
rect 85758 10616 85764 10628
rect 85816 10656 85822 10668
rect 87064 10665 87092 10764
rect 90358 10752 90364 10804
rect 90416 10792 90422 10804
rect 90453 10795 90511 10801
rect 90453 10792 90465 10795
rect 90416 10764 90465 10792
rect 90416 10752 90422 10764
rect 90453 10761 90465 10764
rect 90499 10761 90511 10795
rect 90453 10755 90511 10761
rect 91005 10795 91063 10801
rect 91005 10761 91017 10795
rect 91051 10792 91063 10795
rect 91738 10792 91744 10804
rect 91051 10764 91744 10792
rect 91051 10761 91063 10764
rect 91005 10755 91063 10761
rect 91738 10752 91744 10764
rect 91796 10752 91802 10804
rect 94593 10795 94651 10801
rect 94593 10761 94605 10795
rect 94639 10792 94651 10795
rect 95510 10792 95516 10804
rect 94639 10764 95516 10792
rect 94639 10761 94651 10764
rect 94593 10755 94651 10761
rect 95510 10752 95516 10764
rect 95568 10752 95574 10804
rect 106182 10752 106188 10804
rect 106240 10792 106246 10804
rect 111058 10792 111064 10804
rect 106240 10764 111064 10792
rect 106240 10752 106246 10764
rect 111058 10752 111064 10764
rect 111116 10752 111122 10804
rect 118513 10795 118571 10801
rect 118513 10761 118525 10795
rect 118559 10792 118571 10795
rect 120258 10792 120264 10804
rect 118559 10764 120264 10792
rect 118559 10761 118571 10764
rect 118513 10755 118571 10761
rect 120258 10752 120264 10764
rect 120316 10752 120322 10804
rect 120718 10752 120724 10804
rect 120776 10792 120782 10804
rect 123754 10792 123760 10804
rect 120776 10764 123760 10792
rect 120776 10752 120782 10764
rect 123754 10752 123760 10764
rect 123812 10752 123818 10804
rect 124766 10792 124772 10804
rect 124727 10764 124772 10792
rect 124766 10752 124772 10764
rect 124824 10752 124830 10804
rect 127158 10752 127164 10804
rect 127216 10792 127222 10804
rect 128173 10795 128231 10801
rect 128173 10792 128185 10795
rect 127216 10764 128185 10792
rect 127216 10752 127222 10764
rect 128173 10761 128185 10764
rect 128219 10761 128231 10795
rect 128173 10755 128231 10761
rect 128262 10752 128268 10804
rect 128320 10792 128326 10804
rect 131942 10792 131948 10804
rect 128320 10764 131436 10792
rect 131903 10764 131948 10792
rect 128320 10752 128326 10764
rect 110874 10724 110880 10736
rect 107488 10696 110880 10724
rect 86497 10659 86555 10665
rect 86497 10656 86509 10659
rect 85816 10628 86509 10656
rect 85816 10616 85822 10628
rect 86497 10625 86509 10628
rect 86543 10625 86555 10659
rect 86497 10619 86555 10625
rect 87049 10659 87107 10665
rect 87049 10625 87061 10659
rect 87095 10625 87107 10659
rect 88334 10656 88340 10668
rect 88295 10628 88340 10656
rect 87049 10619 87107 10625
rect 88334 10616 88340 10628
rect 88392 10656 88398 10668
rect 88889 10659 88947 10665
rect 88889 10656 88901 10659
rect 88392 10628 88901 10656
rect 88392 10616 88398 10628
rect 88889 10625 88901 10628
rect 88935 10625 88947 10659
rect 88889 10619 88947 10625
rect 90910 10616 90916 10668
rect 90968 10656 90974 10668
rect 93765 10659 93823 10665
rect 90968 10628 93256 10656
rect 90968 10616 90974 10628
rect 82722 10588 82728 10600
rect 81492 10560 82728 10588
rect 81492 10548 81498 10560
rect 82722 10548 82728 10560
rect 82780 10548 82786 10600
rect 84654 10588 84660 10600
rect 84615 10560 84660 10588
rect 84654 10548 84660 10560
rect 84712 10548 84718 10600
rect 85666 10588 85672 10600
rect 85627 10560 85672 10588
rect 85666 10548 85672 10560
rect 85724 10548 85730 10600
rect 88058 10588 88064 10600
rect 88019 10560 88064 10588
rect 88058 10548 88064 10560
rect 88116 10548 88122 10600
rect 92201 10591 92259 10597
rect 92201 10557 92213 10591
rect 92247 10588 92259 10591
rect 93118 10588 93124 10600
rect 92247 10560 93124 10588
rect 92247 10557 92259 10560
rect 92201 10551 92259 10557
rect 93118 10548 93124 10560
rect 93176 10548 93182 10600
rect 93228 10597 93256 10628
rect 93765 10625 93777 10659
rect 93811 10656 93823 10659
rect 93811 10628 94176 10656
rect 93811 10625 93823 10628
rect 93765 10619 93823 10625
rect 93213 10591 93271 10597
rect 93213 10557 93225 10591
rect 93259 10557 93271 10591
rect 93213 10551 93271 10557
rect 73890 10480 73896 10532
rect 73948 10520 73954 10532
rect 73948 10492 74764 10520
rect 73948 10480 73954 10492
rect 72528 10424 73660 10452
rect 74074 10412 74080 10464
rect 74132 10452 74138 10464
rect 74445 10455 74503 10461
rect 74445 10452 74457 10455
rect 74132 10424 74457 10452
rect 74132 10412 74138 10424
rect 74445 10421 74457 10424
rect 74491 10421 74503 10455
rect 74736 10452 74764 10492
rect 78214 10480 78220 10532
rect 78272 10520 78278 10532
rect 83645 10523 83703 10529
rect 83645 10520 83657 10523
rect 78272 10492 83657 10520
rect 78272 10480 78278 10492
rect 83645 10489 83657 10492
rect 83691 10489 83703 10523
rect 83645 10483 83703 10489
rect 94148 10461 94176 10628
rect 96062 10616 96068 10668
rect 96120 10656 96126 10668
rect 98914 10656 98920 10668
rect 96120 10628 98500 10656
rect 98827 10628 98920 10656
rect 96120 10616 96126 10628
rect 95878 10588 95884 10600
rect 95839 10560 95884 10588
rect 95878 10548 95884 10560
rect 95936 10548 95942 10600
rect 97353 10591 97411 10597
rect 97353 10557 97365 10591
rect 97399 10588 97411 10591
rect 98362 10588 98368 10600
rect 97399 10560 98368 10588
rect 97399 10557 97411 10560
rect 97353 10551 97411 10557
rect 98362 10548 98368 10560
rect 98420 10548 98426 10600
rect 98472 10597 98500 10628
rect 98914 10616 98920 10628
rect 98972 10656 98978 10668
rect 101766 10656 101772 10668
rect 98972 10628 101772 10656
rect 98972 10616 98978 10628
rect 101766 10616 101772 10628
rect 101824 10616 101830 10668
rect 103793 10659 103851 10665
rect 103793 10625 103805 10659
rect 103839 10656 103851 10659
rect 104250 10656 104256 10668
rect 103839 10628 104256 10656
rect 103839 10625 103851 10628
rect 103793 10619 103851 10625
rect 104250 10616 104256 10628
rect 104308 10616 104314 10668
rect 106182 10656 106188 10668
rect 106143 10628 106188 10656
rect 106182 10616 106188 10628
rect 106240 10616 106246 10668
rect 98457 10591 98515 10597
rect 98457 10557 98469 10591
rect 98503 10557 98515 10591
rect 98457 10551 98515 10557
rect 99558 10548 99564 10600
rect 99616 10588 99622 10600
rect 99745 10591 99803 10597
rect 99745 10588 99757 10591
rect 99616 10560 99757 10588
rect 99616 10548 99622 10560
rect 99745 10557 99757 10560
rect 99791 10557 99803 10591
rect 102226 10588 102232 10600
rect 102187 10560 102232 10588
rect 99745 10551 99803 10557
rect 102226 10548 102232 10560
rect 102284 10548 102290 10600
rect 103238 10588 103244 10600
rect 103199 10560 103244 10588
rect 103238 10548 103244 10560
rect 103296 10548 103302 10600
rect 104618 10588 104624 10600
rect 104579 10560 104624 10588
rect 104618 10548 104624 10560
rect 104676 10548 104682 10600
rect 106093 10591 106151 10597
rect 106093 10557 106105 10591
rect 106139 10588 106151 10591
rect 107488 10588 107516 10696
rect 110874 10684 110880 10696
rect 110932 10684 110938 10736
rect 119614 10724 119620 10736
rect 117240 10696 119620 10724
rect 107838 10616 107844 10668
rect 107896 10656 107902 10668
rect 108761 10659 108819 10665
rect 108761 10656 108773 10659
rect 107896 10628 108773 10656
rect 107896 10616 107902 10628
rect 108761 10625 108773 10628
rect 108807 10656 108819 10659
rect 108942 10656 108948 10668
rect 108807 10628 108948 10656
rect 108807 10625 108819 10628
rect 108761 10619 108819 10625
rect 108942 10616 108948 10628
rect 109000 10616 109006 10668
rect 111334 10656 111340 10668
rect 111295 10628 111340 10656
rect 111334 10616 111340 10628
rect 111392 10616 111398 10668
rect 112622 10656 112628 10668
rect 111536 10628 112628 10656
rect 107654 10588 107660 10600
rect 106139 10560 107516 10588
rect 107615 10560 107660 10588
rect 106139 10557 106151 10560
rect 106093 10551 106151 10557
rect 107654 10548 107660 10560
rect 107712 10548 107718 10600
rect 110046 10588 110052 10600
rect 110007 10560 110052 10588
rect 110046 10548 110052 10560
rect 110104 10548 110110 10600
rect 111536 10588 111564 10628
rect 112622 10616 112628 10628
rect 112680 10616 112686 10668
rect 114649 10659 114707 10665
rect 114649 10625 114661 10659
rect 114695 10625 114707 10659
rect 114649 10619 114707 10625
rect 110800 10560 111564 10588
rect 105630 10480 105636 10532
rect 105688 10520 105694 10532
rect 108850 10520 108856 10532
rect 105688 10492 108856 10520
rect 105688 10480 105694 10492
rect 108850 10480 108856 10492
rect 108908 10480 108914 10532
rect 108945 10523 109003 10529
rect 108945 10489 108957 10523
rect 108991 10520 109003 10523
rect 110800 10520 110828 10560
rect 112898 10548 112904 10600
rect 112956 10548 112962 10600
rect 113269 10591 113327 10597
rect 113269 10557 113281 10591
rect 113315 10588 113327 10591
rect 113450 10588 113456 10600
rect 113315 10560 113456 10588
rect 113315 10557 113327 10560
rect 113269 10551 113327 10557
rect 113450 10548 113456 10560
rect 113508 10548 113514 10600
rect 108991 10492 110828 10520
rect 108991 10489 109003 10492
rect 108945 10483 109003 10489
rect 110966 10480 110972 10532
rect 111024 10520 111030 10532
rect 111334 10520 111340 10532
rect 111024 10492 111340 10520
rect 111024 10480 111030 10492
rect 111334 10480 111340 10492
rect 111392 10480 111398 10532
rect 111521 10523 111579 10529
rect 111521 10489 111533 10523
rect 111567 10520 111579 10523
rect 112916 10520 112944 10548
rect 114664 10532 114692 10619
rect 117130 10616 117136 10668
rect 117188 10656 117194 10668
rect 117240 10665 117268 10696
rect 119614 10684 119620 10696
rect 119672 10684 119678 10736
rect 119706 10684 119712 10736
rect 119764 10724 119770 10736
rect 119764 10696 129688 10724
rect 119764 10684 119770 10696
rect 117225 10659 117283 10665
rect 117225 10656 117237 10659
rect 117188 10628 117237 10656
rect 117188 10616 117194 10628
rect 117225 10625 117237 10628
rect 117271 10625 117283 10659
rect 121086 10656 121092 10668
rect 121047 10628 121092 10656
rect 117225 10619 117283 10625
rect 121086 10616 121092 10628
rect 121144 10616 121150 10668
rect 122837 10659 122895 10665
rect 122837 10625 122849 10659
rect 122883 10656 122895 10659
rect 123110 10656 123116 10668
rect 122883 10628 123116 10656
rect 122883 10625 122895 10628
rect 122837 10619 122895 10625
rect 123110 10616 123116 10628
rect 123168 10656 123174 10668
rect 124677 10659 124735 10665
rect 123168 10628 123708 10656
rect 123168 10616 123174 10628
rect 114741 10591 114799 10597
rect 114741 10557 114753 10591
rect 114787 10588 114799 10591
rect 114830 10588 114836 10600
rect 114787 10560 114836 10588
rect 114787 10557 114799 10560
rect 114741 10551 114799 10557
rect 114830 10548 114836 10560
rect 114888 10548 114894 10600
rect 115661 10591 115719 10597
rect 115661 10557 115673 10591
rect 115707 10588 115719 10591
rect 115842 10588 115848 10600
rect 115707 10560 115848 10588
rect 115707 10557 115719 10560
rect 115661 10551 115719 10557
rect 115842 10548 115848 10560
rect 115900 10548 115906 10600
rect 116670 10588 116676 10600
rect 116631 10560 116676 10588
rect 116670 10548 116676 10560
rect 116728 10548 116734 10600
rect 119522 10588 119528 10600
rect 119483 10560 119528 10588
rect 119522 10548 119528 10560
rect 119580 10548 119586 10600
rect 120534 10588 120540 10600
rect 120495 10560 120540 10588
rect 120534 10548 120540 10560
rect 120592 10548 120598 10600
rect 123386 10588 123392 10600
rect 121012 10560 123392 10588
rect 114646 10520 114652 10532
rect 111567 10492 112944 10520
rect 114559 10492 114652 10520
rect 111567 10489 111579 10492
rect 111521 10483 111579 10489
rect 114646 10480 114652 10492
rect 114704 10520 114710 10532
rect 121012 10520 121040 10560
rect 123386 10548 123392 10560
rect 123444 10548 123450 10600
rect 123680 10588 123708 10628
rect 124677 10625 124689 10659
rect 124723 10656 124735 10659
rect 124950 10656 124956 10668
rect 124723 10628 124956 10656
rect 124723 10625 124735 10628
rect 124677 10619 124735 10625
rect 124950 10616 124956 10628
rect 125008 10656 125014 10668
rect 127066 10656 127072 10668
rect 125008 10628 127072 10656
rect 125008 10616 125014 10628
rect 127066 10616 127072 10628
rect 127124 10616 127130 10668
rect 127253 10659 127311 10665
rect 127253 10625 127265 10659
rect 127299 10656 127311 10659
rect 127618 10656 127624 10668
rect 127299 10628 127624 10656
rect 127299 10625 127311 10628
rect 127253 10619 127311 10625
rect 127618 10616 127624 10628
rect 127676 10616 127682 10668
rect 128081 10659 128139 10665
rect 128081 10625 128093 10659
rect 128127 10656 128139 10659
rect 128354 10656 128360 10668
rect 128127 10628 128360 10656
rect 128127 10625 128139 10628
rect 128081 10619 128139 10625
rect 128354 10616 128360 10628
rect 128412 10656 128418 10668
rect 129182 10656 129188 10668
rect 128412 10628 129188 10656
rect 128412 10616 128418 10628
rect 129182 10616 129188 10628
rect 129240 10616 129246 10668
rect 125594 10588 125600 10600
rect 123680 10560 125600 10588
rect 125594 10548 125600 10560
rect 125652 10548 125658 10600
rect 125689 10591 125747 10597
rect 125689 10557 125701 10591
rect 125735 10588 125747 10591
rect 126238 10588 126244 10600
rect 125735 10560 126244 10588
rect 125735 10557 125747 10560
rect 125689 10551 125747 10557
rect 126238 10548 126244 10560
rect 126296 10548 126302 10600
rect 126701 10591 126759 10597
rect 126701 10557 126713 10591
rect 126747 10557 126759 10591
rect 129550 10588 129556 10600
rect 129511 10560 129556 10588
rect 126701 10551 126759 10557
rect 126716 10520 126744 10551
rect 129550 10548 129556 10560
rect 129608 10548 129614 10600
rect 129660 10588 129688 10696
rect 130654 10656 130660 10668
rect 130615 10628 130660 10656
rect 130654 10616 130660 10628
rect 130712 10616 130718 10668
rect 130565 10591 130623 10597
rect 130565 10588 130577 10591
rect 129660 10560 130577 10588
rect 130565 10557 130577 10560
rect 130611 10557 130623 10591
rect 130565 10551 130623 10557
rect 114704 10492 121040 10520
rect 121104 10492 126744 10520
rect 131408 10520 131436 10764
rect 131942 10752 131948 10764
rect 132000 10752 132006 10804
rect 148318 10752 148324 10804
rect 148376 10792 148382 10804
rect 148376 10764 165752 10792
rect 148376 10752 148382 10764
rect 131574 10684 131580 10736
rect 131632 10724 131638 10736
rect 135070 10724 135076 10736
rect 131632 10696 135076 10724
rect 131632 10684 131638 10696
rect 135070 10684 135076 10696
rect 135128 10724 135134 10736
rect 135257 10727 135315 10733
rect 135128 10696 135208 10724
rect 135128 10684 135134 10696
rect 134058 10656 134064 10668
rect 134019 10628 134064 10656
rect 134058 10616 134064 10628
rect 134116 10616 134122 10668
rect 135180 10665 135208 10696
rect 135257 10693 135269 10727
rect 135303 10724 135315 10727
rect 139118 10724 139124 10736
rect 135303 10696 139124 10724
rect 135303 10693 135315 10696
rect 135257 10687 135315 10693
rect 139118 10684 139124 10696
rect 139176 10724 139182 10736
rect 139489 10727 139547 10733
rect 139489 10724 139501 10727
rect 139176 10696 139501 10724
rect 139176 10684 139182 10696
rect 139489 10693 139501 10696
rect 139535 10693 139547 10727
rect 145006 10724 145012 10736
rect 139489 10687 139547 10693
rect 141988 10696 145012 10724
rect 135165 10659 135223 10665
rect 135165 10625 135177 10659
rect 135211 10625 135223 10659
rect 137281 10659 137339 10665
rect 137281 10656 137293 10659
rect 135165 10619 135223 10625
rect 136100 10628 137293 10656
rect 132954 10588 132960 10600
rect 132915 10560 132960 10588
rect 132954 10548 132960 10560
rect 133012 10548 133018 10600
rect 134153 10591 134211 10597
rect 134153 10557 134165 10591
rect 134199 10588 134211 10591
rect 136100 10588 136128 10628
rect 137281 10625 137293 10628
rect 137327 10656 137339 10659
rect 137462 10656 137468 10668
rect 137327 10628 137468 10656
rect 137327 10625 137339 10628
rect 137281 10619 137339 10625
rect 137462 10616 137468 10628
rect 137520 10616 137526 10668
rect 139026 10656 139032 10668
rect 138987 10628 139032 10656
rect 139026 10616 139032 10628
rect 139084 10616 139090 10668
rect 141988 10656 142016 10696
rect 145006 10684 145012 10696
rect 145064 10684 145070 10736
rect 146846 10684 146852 10736
rect 146904 10724 146910 10736
rect 146904 10696 159496 10724
rect 146904 10684 146910 10696
rect 142154 10656 142160 10668
rect 139136 10628 142016 10656
rect 142115 10628 142160 10656
rect 134199 10560 136128 10588
rect 136177 10591 136235 10597
rect 134199 10557 134211 10560
rect 134153 10551 134211 10557
rect 136177 10557 136189 10591
rect 136223 10588 136235 10591
rect 136266 10588 136272 10600
rect 136223 10560 136272 10588
rect 136223 10557 136235 10560
rect 136177 10551 136235 10557
rect 136266 10548 136272 10560
rect 136324 10548 136330 10600
rect 139136 10597 139164 10628
rect 142154 10616 142160 10628
rect 142212 10616 142218 10668
rect 144914 10656 144920 10668
rect 144875 10628 144920 10656
rect 144914 10616 144920 10628
rect 144972 10656 144978 10668
rect 145653 10659 145711 10665
rect 145653 10656 145665 10659
rect 144972 10628 145665 10656
rect 144972 10616 144978 10628
rect 145653 10625 145665 10628
rect 145699 10625 145711 10659
rect 147858 10656 147864 10668
rect 147819 10628 147864 10656
rect 145653 10619 145711 10625
rect 147858 10616 147864 10628
rect 147916 10616 147922 10668
rect 150897 10659 150955 10665
rect 150897 10625 150909 10659
rect 150943 10656 150955 10659
rect 151630 10656 151636 10668
rect 150943 10628 151636 10656
rect 150943 10625 150955 10628
rect 150897 10619 150955 10625
rect 151630 10616 151636 10628
rect 151688 10616 151694 10668
rect 153194 10656 153200 10668
rect 153155 10628 153200 10656
rect 153194 10616 153200 10628
rect 153252 10616 153258 10668
rect 155954 10656 155960 10668
rect 155915 10628 155960 10656
rect 155954 10616 155960 10628
rect 156012 10616 156018 10668
rect 158441 10659 158499 10665
rect 158441 10625 158453 10659
rect 158487 10656 158499 10659
rect 158714 10656 158720 10668
rect 158487 10628 158720 10656
rect 158487 10625 158499 10628
rect 158441 10619 158499 10625
rect 158714 10616 158720 10628
rect 158772 10656 158778 10668
rect 159266 10656 159272 10668
rect 158772 10628 159272 10656
rect 158772 10616 158778 10628
rect 159266 10616 159272 10628
rect 159324 10616 159330 10668
rect 137189 10591 137247 10597
rect 137189 10557 137201 10591
rect 137235 10557 137247 10591
rect 137189 10551 137247 10557
rect 139121 10591 139179 10597
rect 139121 10557 139133 10591
rect 139167 10557 139179 10591
rect 139121 10551 139179 10557
rect 140961 10591 141019 10597
rect 140961 10557 140973 10591
rect 141007 10588 141019 10591
rect 141050 10588 141056 10600
rect 141007 10560 141056 10588
rect 141007 10557 141019 10560
rect 140961 10551 141019 10557
rect 137204 10520 137232 10551
rect 141050 10548 141056 10560
rect 141108 10548 141114 10600
rect 143813 10591 143871 10597
rect 143813 10557 143825 10591
rect 143859 10588 143871 10591
rect 144178 10588 144184 10600
rect 143859 10560 144184 10588
rect 143859 10557 143871 10560
rect 143813 10551 143871 10557
rect 144178 10548 144184 10560
rect 144236 10548 144242 10600
rect 146389 10591 146447 10597
rect 146389 10557 146401 10591
rect 146435 10588 146447 10591
rect 146938 10588 146944 10600
rect 146435 10560 146944 10588
rect 146435 10557 146447 10560
rect 146389 10551 146447 10557
rect 146938 10548 146944 10560
rect 146996 10548 147002 10600
rect 148778 10548 148784 10600
rect 148836 10588 148842 10600
rect 149333 10591 149391 10597
rect 149333 10588 149345 10591
rect 148836 10560 149345 10588
rect 148836 10548 148842 10560
rect 149333 10557 149345 10560
rect 149379 10557 149391 10591
rect 149333 10551 149391 10557
rect 152001 10591 152059 10597
rect 152001 10557 152013 10591
rect 152047 10588 152059 10591
rect 152090 10588 152096 10600
rect 152047 10560 152096 10588
rect 152047 10557 152059 10560
rect 152001 10551 152059 10557
rect 152090 10548 152096 10560
rect 152148 10548 152154 10600
rect 154761 10591 154819 10597
rect 154761 10557 154773 10591
rect 154807 10588 154819 10591
rect 155310 10588 155316 10600
rect 154807 10560 155316 10588
rect 154807 10557 154819 10560
rect 154761 10551 154819 10557
rect 155310 10548 155316 10560
rect 155368 10548 155374 10600
rect 156138 10588 156144 10600
rect 156099 10560 156144 10588
rect 156138 10548 156144 10560
rect 156196 10548 156202 10600
rect 157242 10548 157248 10600
rect 157300 10588 157306 10600
rect 159468 10597 159496 10696
rect 159542 10616 159548 10668
rect 159600 10656 159606 10668
rect 161109 10659 161167 10665
rect 159600 10628 159645 10656
rect 159600 10616 159606 10628
rect 161109 10625 161121 10659
rect 161155 10656 161167 10659
rect 162854 10656 162860 10668
rect 161155 10628 162860 10656
rect 161155 10625 161167 10628
rect 161109 10619 161167 10625
rect 162854 10616 162860 10628
rect 162912 10616 162918 10668
rect 164326 10656 164332 10668
rect 164287 10628 164332 10656
rect 164326 10616 164332 10628
rect 164384 10616 164390 10668
rect 159453 10591 159511 10597
rect 157300 10560 157380 10588
rect 157300 10548 157306 10560
rect 142246 10520 142252 10532
rect 131408 10492 137232 10520
rect 142207 10492 142252 10520
rect 114704 10480 114710 10492
rect 79137 10455 79195 10461
rect 79137 10452 79149 10455
rect 74736 10424 79149 10452
rect 74445 10415 74503 10421
rect 79137 10421 79149 10424
rect 79183 10421 79195 10455
rect 79137 10415 79195 10421
rect 94133 10455 94191 10461
rect 94133 10421 94145 10455
rect 94179 10452 94191 10455
rect 109678 10452 109684 10464
rect 94179 10424 109684 10452
rect 94179 10421 94191 10424
rect 94133 10415 94191 10421
rect 109678 10412 109684 10424
rect 109736 10412 109742 10464
rect 111150 10412 111156 10464
rect 111208 10452 111214 10464
rect 111702 10452 111708 10464
rect 111208 10424 111708 10452
rect 111208 10412 111214 10424
rect 111702 10412 111708 10424
rect 111760 10452 111766 10464
rect 111889 10455 111947 10461
rect 111889 10452 111901 10455
rect 111760 10424 111901 10452
rect 111760 10412 111766 10424
rect 111889 10421 111901 10424
rect 111935 10421 111947 10455
rect 112898 10452 112904 10464
rect 112859 10424 112904 10452
rect 111889 10415 111947 10421
rect 112898 10412 112904 10424
rect 112956 10412 112962 10464
rect 112990 10412 112996 10464
rect 113048 10452 113054 10464
rect 121104 10452 121132 10492
rect 142246 10480 142252 10492
rect 142304 10480 142310 10532
rect 145098 10520 145104 10532
rect 145059 10492 145104 10520
rect 145098 10480 145104 10492
rect 145156 10480 145162 10532
rect 147861 10523 147919 10529
rect 147861 10489 147873 10523
rect 147907 10520 147919 10523
rect 149790 10520 149796 10532
rect 147907 10492 149796 10520
rect 147907 10489 147919 10492
rect 147861 10483 147919 10489
rect 149790 10480 149796 10492
rect 149848 10480 149854 10532
rect 150805 10523 150863 10529
rect 150805 10489 150817 10523
rect 150851 10520 150863 10523
rect 152366 10520 152372 10532
rect 150851 10492 152372 10520
rect 150851 10489 150863 10492
rect 150805 10483 150863 10489
rect 152366 10480 152372 10492
rect 152424 10480 152430 10532
rect 153286 10520 153292 10532
rect 153247 10492 153292 10520
rect 153286 10480 153292 10492
rect 153344 10480 153350 10532
rect 157352 10520 157380 10560
rect 159453 10557 159465 10591
rect 159499 10557 159511 10591
rect 159453 10551 159511 10557
rect 162121 10591 162179 10597
rect 162121 10557 162133 10591
rect 162167 10588 162179 10591
rect 162670 10588 162676 10600
rect 162167 10560 162676 10588
rect 162167 10557 162179 10560
rect 162121 10551 162179 10557
rect 162670 10548 162676 10560
rect 162728 10588 162734 10600
rect 163225 10591 163283 10597
rect 163225 10588 163237 10591
rect 162728 10560 163237 10588
rect 162728 10548 162734 10560
rect 163225 10557 163237 10560
rect 163271 10557 163283 10591
rect 163225 10551 163283 10557
rect 164237 10591 164295 10597
rect 164237 10557 164249 10591
rect 164283 10557 164295 10591
rect 165614 10588 165620 10600
rect 165575 10560 165620 10588
rect 164237 10551 164295 10557
rect 164252 10520 164280 10551
rect 165614 10548 165620 10560
rect 165672 10548 165678 10600
rect 165724 10588 165752 10764
rect 166718 10656 166724 10668
rect 166679 10628 166724 10656
rect 166718 10616 166724 10628
rect 166776 10616 166782 10668
rect 166629 10591 166687 10597
rect 166629 10588 166641 10591
rect 165724 10560 166641 10588
rect 166629 10557 166641 10560
rect 166675 10557 166687 10591
rect 166629 10551 166687 10557
rect 157352 10492 164280 10520
rect 113048 10424 121132 10452
rect 113048 10412 113054 10424
rect 121178 10412 121184 10464
rect 121236 10452 121242 10464
rect 121365 10455 121423 10461
rect 121365 10452 121377 10455
rect 121236 10424 121377 10452
rect 121236 10412 121242 10424
rect 121365 10421 121377 10424
rect 121411 10421 121423 10455
rect 121365 10415 121423 10421
rect 122561 10455 122619 10461
rect 122561 10421 122573 10455
rect 122607 10452 122619 10455
rect 122742 10452 122748 10464
rect 122607 10424 122748 10452
rect 122607 10421 122619 10424
rect 122561 10415 122619 10421
rect 122742 10412 122748 10424
rect 122800 10412 122806 10464
rect 122926 10452 122932 10464
rect 122887 10424 122932 10452
rect 122926 10412 122932 10424
rect 122984 10412 122990 10464
rect 123754 10412 123760 10464
rect 123812 10452 123818 10464
rect 127434 10452 127440 10464
rect 123812 10424 127440 10452
rect 123812 10412 123818 10424
rect 127434 10412 127440 10424
rect 127492 10412 127498 10464
rect 127618 10452 127624 10464
rect 127579 10424 127624 10452
rect 127618 10412 127624 10424
rect 127676 10412 127682 10464
rect 128078 10412 128084 10464
rect 128136 10452 128142 10464
rect 128541 10455 128599 10461
rect 128541 10452 128553 10455
rect 128136 10424 128553 10452
rect 128136 10412 128142 10424
rect 128541 10421 128553 10424
rect 128587 10421 128599 10455
rect 132402 10452 132408 10464
rect 132363 10424 132408 10452
rect 128541 10415 128599 10421
rect 132402 10412 132408 10424
rect 132460 10412 132466 10464
rect 133506 10412 133512 10464
rect 133564 10452 133570 10464
rect 133693 10455 133751 10461
rect 133693 10452 133705 10455
rect 133564 10424 133705 10452
rect 133564 10412 133570 10424
rect 133693 10421 133705 10424
rect 133739 10421 133751 10455
rect 133693 10415 133751 10421
rect 138014 10412 138020 10464
rect 138072 10452 138078 10464
rect 140406 10452 140412 10464
rect 138072 10424 138117 10452
rect 140367 10424 140412 10452
rect 138072 10412 138078 10424
rect 140406 10412 140412 10424
rect 140464 10412 140470 10464
rect 147582 10412 147588 10464
rect 147640 10452 147646 10464
rect 157242 10452 157248 10464
rect 147640 10424 157248 10452
rect 147640 10412 147646 10424
rect 157242 10412 157248 10424
rect 157300 10412 157306 10464
rect 157978 10452 157984 10464
rect 157939 10424 157984 10452
rect 157978 10412 157984 10424
rect 158036 10412 158042 10464
rect 160462 10452 160468 10464
rect 160423 10424 160468 10452
rect 160462 10412 160468 10424
rect 160520 10412 160526 10464
rect 368 10362 169556 10384
rect 368 10310 28456 10362
rect 28508 10310 28520 10362
rect 28572 10310 28584 10362
rect 28636 10310 28648 10362
rect 28700 10310 84878 10362
rect 84930 10310 84942 10362
rect 84994 10310 85006 10362
rect 85058 10310 85070 10362
rect 85122 10310 141299 10362
rect 141351 10310 141363 10362
rect 141415 10310 141427 10362
rect 141479 10310 141491 10362
rect 141543 10310 169556 10362
rect 368 10288 169556 10310
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 5353 10251 5411 10257
rect 5353 10248 5365 10251
rect 4396 10220 5365 10248
rect 4396 10208 4402 10220
rect 5353 10217 5365 10220
rect 5399 10217 5411 10251
rect 8294 10248 8300 10260
rect 8255 10220 8300 10248
rect 5353 10211 5411 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 9217 10251 9275 10257
rect 9217 10217 9229 10251
rect 9263 10248 9275 10251
rect 9306 10248 9312 10260
rect 9263 10220 9312 10248
rect 9263 10217 9275 10220
rect 9217 10211 9275 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13998 10248 14004 10260
rect 13959 10220 14004 10248
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 17310 10248 17316 10260
rect 17271 10220 17316 10248
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18690 10248 18696 10260
rect 18651 10220 18696 10248
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 19702 10248 19708 10260
rect 19663 10220 19708 10248
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 24121 10251 24179 10257
rect 24121 10217 24133 10251
rect 24167 10248 24179 10251
rect 24397 10251 24455 10257
rect 24397 10248 24409 10251
rect 24167 10220 24409 10248
rect 24167 10217 24179 10220
rect 24121 10211 24179 10217
rect 24397 10217 24409 10220
rect 24443 10248 24455 10251
rect 29086 10248 29092 10260
rect 24443 10220 29092 10248
rect 24443 10217 24455 10220
rect 24397 10211 24455 10217
rect 29086 10208 29092 10220
rect 29144 10208 29150 10260
rect 30742 10208 30748 10260
rect 30800 10248 30806 10260
rect 30837 10251 30895 10257
rect 30837 10248 30849 10251
rect 30800 10220 30849 10248
rect 30800 10208 30806 10220
rect 30837 10217 30849 10220
rect 30883 10248 30895 10251
rect 33870 10248 33876 10260
rect 30883 10220 33876 10248
rect 30883 10217 30895 10220
rect 30837 10211 30895 10217
rect 33870 10208 33876 10220
rect 33928 10208 33934 10260
rect 34701 10251 34759 10257
rect 34701 10217 34713 10251
rect 34747 10248 34759 10251
rect 35158 10248 35164 10260
rect 34747 10220 35164 10248
rect 34747 10217 34759 10220
rect 34701 10211 34759 10217
rect 35158 10208 35164 10220
rect 35216 10208 35222 10260
rect 35621 10251 35679 10257
rect 35621 10217 35633 10251
rect 35667 10248 35679 10251
rect 35897 10251 35955 10257
rect 35897 10248 35909 10251
rect 35667 10220 35909 10248
rect 35667 10217 35679 10220
rect 35621 10211 35679 10217
rect 35897 10217 35909 10220
rect 35943 10248 35955 10251
rect 35943 10220 36676 10248
rect 35943 10217 35955 10220
rect 35897 10211 35955 10217
rect 2866 10140 2872 10192
rect 2924 10180 2930 10192
rect 9674 10180 9680 10192
rect 2924 10152 9680 10180
rect 2924 10140 2930 10152
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 19518 10140 19524 10192
rect 19576 10180 19582 10192
rect 19576 10152 21220 10180
rect 19576 10140 19582 10152
rect 4154 10112 4160 10124
rect 4115 10084 4160 10112
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 4264 10084 6224 10112
rect 3970 10044 3976 10056
rect 3931 10016 3976 10044
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4264 10044 4292 10084
rect 4120 10016 4292 10044
rect 4525 10047 4583 10053
rect 4120 10004 4126 10016
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 4706 10044 4712 10056
rect 4571 10016 4712 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10013 6147 10047
rect 6196 10044 6224 10084
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 7064 10084 7113 10112
rect 7064 10072 7070 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 19061 10115 19119 10121
rect 7101 10075 7159 10081
rect 7484 10084 8156 10112
rect 7484 10044 7512 10084
rect 6196 10016 7512 10044
rect 7653 10047 7711 10053
rect 6089 10007 6147 10013
rect 7653 10013 7665 10047
rect 7699 10044 7711 10047
rect 7699 10016 8064 10044
rect 7699 10013 7711 10016
rect 7653 10007 7711 10013
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 4430 9908 4436 9920
rect 3660 9880 4436 9908
rect 3660 9868 3666 9880
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 5074 9908 5080 9920
rect 5035 9880 5080 9908
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5997 9911 6055 9917
rect 5997 9877 6009 9911
rect 6043 9908 6055 9911
rect 6104 9908 6132 10007
rect 8036 9920 8064 10016
rect 8128 9976 8156 10084
rect 19061 10081 19073 10115
rect 19107 10112 19119 10115
rect 20070 10112 20076 10124
rect 19107 10084 20076 10112
rect 19107 10081 19119 10084
rect 19061 10075 19119 10081
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 20162 10072 20168 10124
rect 20220 10112 20226 10124
rect 20714 10112 20720 10124
rect 20220 10084 20720 10112
rect 20220 10072 20226 10084
rect 20714 10072 20720 10084
rect 20772 10072 20778 10124
rect 21192 10121 21220 10152
rect 24026 10140 24032 10192
rect 24084 10180 24090 10192
rect 25130 10180 25136 10192
rect 24084 10152 25136 10180
rect 24084 10140 24090 10152
rect 25130 10140 25136 10152
rect 25188 10140 25194 10192
rect 25593 10183 25651 10189
rect 25593 10149 25605 10183
rect 25639 10180 25651 10183
rect 25866 10180 25872 10192
rect 25639 10152 25872 10180
rect 25639 10149 25651 10152
rect 25593 10143 25651 10149
rect 25866 10140 25872 10152
rect 25924 10140 25930 10192
rect 26970 10180 26976 10192
rect 25976 10152 26976 10180
rect 21177 10115 21235 10121
rect 21177 10081 21189 10115
rect 21223 10081 21235 10115
rect 24762 10112 24768 10124
rect 21177 10075 21235 10081
rect 21652 10084 24256 10112
rect 24723 10084 24768 10112
rect 17310 10004 17316 10056
rect 17368 10044 17374 10056
rect 19889 10047 19947 10053
rect 19889 10044 19901 10047
rect 17368 10016 19901 10044
rect 17368 10004 17374 10016
rect 19889 10013 19901 10016
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 21652 9976 21680 10084
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10044 21787 10047
rect 22097 10047 22155 10053
rect 22097 10044 22109 10047
rect 21775 10016 22109 10044
rect 21775 10013 21787 10016
rect 21729 10007 21787 10013
rect 22097 10013 22109 10016
rect 22143 10044 22155 10047
rect 23382 10044 23388 10056
rect 22143 10016 23388 10044
rect 22143 10013 22155 10016
rect 22097 10007 22155 10013
rect 23382 10004 23388 10016
rect 23440 10004 23446 10056
rect 23566 10044 23572 10056
rect 23527 10016 23572 10044
rect 23566 10004 23572 10016
rect 23624 10004 23630 10056
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10044 23719 10047
rect 23934 10044 23940 10056
rect 23707 10016 23940 10044
rect 23707 10013 23719 10016
rect 23661 10007 23719 10013
rect 23934 10004 23940 10016
rect 23992 10004 23998 10056
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10044 24087 10047
rect 24121 10047 24179 10053
rect 24121 10044 24133 10047
rect 24075 10016 24133 10044
rect 24075 10013 24087 10016
rect 24029 10007 24087 10013
rect 24121 10013 24133 10016
rect 24167 10013 24179 10047
rect 24228 10044 24256 10084
rect 24762 10072 24768 10084
rect 24820 10072 24826 10124
rect 25976 10044 26004 10152
rect 26970 10140 26976 10152
rect 27028 10140 27034 10192
rect 27065 10183 27123 10189
rect 27065 10149 27077 10183
rect 27111 10180 27123 10183
rect 27890 10180 27896 10192
rect 27111 10152 27896 10180
rect 27111 10149 27123 10152
rect 27065 10143 27123 10149
rect 27080 10112 27108 10143
rect 27890 10140 27896 10152
rect 27948 10140 27954 10192
rect 28905 10183 28963 10189
rect 28905 10149 28917 10183
rect 28951 10180 28963 10183
rect 28994 10180 29000 10192
rect 28951 10152 29000 10180
rect 28951 10149 28963 10152
rect 28905 10143 28963 10149
rect 28994 10140 29000 10152
rect 29052 10140 29058 10192
rect 30653 10183 30711 10189
rect 30653 10149 30665 10183
rect 30699 10180 30711 10183
rect 34330 10180 34336 10192
rect 30699 10152 34336 10180
rect 30699 10149 30711 10152
rect 30653 10143 30711 10149
rect 34330 10140 34336 10152
rect 34388 10140 34394 10192
rect 34514 10140 34520 10192
rect 34572 10180 34578 10192
rect 34885 10183 34943 10189
rect 34885 10180 34897 10183
rect 34572 10152 34897 10180
rect 34572 10140 34578 10152
rect 34885 10149 34897 10152
rect 34931 10149 34943 10183
rect 34885 10143 34943 10149
rect 35434 10140 35440 10192
rect 35492 10180 35498 10192
rect 36648 10180 36676 10220
rect 36814 10208 36820 10260
rect 36872 10248 36878 10260
rect 40313 10251 40371 10257
rect 40313 10248 40325 10251
rect 36872 10220 40325 10248
rect 36872 10208 36878 10220
rect 40313 10217 40325 10220
rect 40359 10217 40371 10251
rect 40313 10211 40371 10217
rect 40957 10251 41015 10257
rect 40957 10217 40969 10251
rect 41003 10248 41015 10251
rect 41049 10251 41107 10257
rect 41049 10248 41061 10251
rect 41003 10220 41061 10248
rect 41003 10217 41015 10220
rect 40957 10211 41015 10217
rect 41049 10217 41061 10220
rect 41095 10248 41107 10251
rect 41233 10251 41291 10257
rect 41233 10248 41245 10251
rect 41095 10220 41245 10248
rect 41095 10217 41107 10220
rect 41049 10211 41107 10217
rect 41233 10217 41245 10220
rect 41279 10217 41291 10251
rect 41233 10211 41291 10217
rect 41509 10251 41567 10257
rect 41509 10217 41521 10251
rect 41555 10248 41567 10251
rect 41598 10248 41604 10260
rect 41555 10220 41604 10248
rect 41555 10217 41567 10220
rect 41509 10211 41567 10217
rect 41598 10208 41604 10220
rect 41656 10248 41662 10260
rect 41874 10248 41880 10260
rect 41656 10220 41880 10248
rect 41656 10208 41662 10220
rect 41874 10208 41880 10220
rect 41932 10208 41938 10260
rect 42058 10208 42064 10260
rect 42116 10248 42122 10260
rect 42426 10248 42432 10260
rect 42116 10220 42432 10248
rect 42116 10208 42122 10220
rect 42426 10208 42432 10220
rect 42484 10208 42490 10260
rect 42794 10208 42800 10260
rect 42852 10248 42858 10260
rect 46566 10248 46572 10260
rect 42852 10220 46572 10248
rect 42852 10208 42858 10220
rect 46566 10208 46572 10220
rect 46624 10208 46630 10260
rect 48041 10251 48099 10257
rect 48041 10217 48053 10251
rect 48087 10248 48099 10251
rect 48222 10248 48228 10260
rect 48087 10220 48228 10248
rect 48087 10217 48099 10220
rect 48041 10211 48099 10217
rect 48222 10208 48228 10220
rect 48280 10208 48286 10260
rect 48317 10251 48375 10257
rect 48317 10217 48329 10251
rect 48363 10248 48375 10251
rect 48590 10248 48596 10260
rect 48363 10220 48596 10248
rect 48363 10217 48375 10220
rect 48317 10211 48375 10217
rect 48590 10208 48596 10220
rect 48648 10208 48654 10260
rect 49053 10251 49111 10257
rect 49053 10217 49065 10251
rect 49099 10248 49111 10251
rect 49329 10251 49387 10257
rect 49329 10248 49341 10251
rect 49099 10220 49341 10248
rect 49099 10217 49111 10220
rect 49053 10211 49111 10217
rect 49329 10217 49341 10220
rect 49375 10248 49387 10251
rect 50798 10248 50804 10260
rect 49375 10220 50804 10248
rect 49375 10217 49387 10220
rect 49329 10211 49387 10217
rect 50798 10208 50804 10220
rect 50856 10208 50862 10260
rect 50893 10251 50951 10257
rect 50893 10217 50905 10251
rect 50939 10248 50951 10251
rect 50982 10248 50988 10260
rect 50939 10220 50988 10248
rect 50939 10217 50951 10220
rect 50893 10211 50951 10217
rect 50982 10208 50988 10220
rect 51040 10248 51046 10260
rect 51534 10248 51540 10260
rect 51040 10220 51540 10248
rect 51040 10208 51046 10220
rect 51534 10208 51540 10220
rect 51592 10208 51598 10260
rect 51718 10208 51724 10260
rect 51776 10248 51782 10260
rect 52181 10251 52239 10257
rect 52181 10248 52193 10251
rect 51776 10220 52193 10248
rect 51776 10208 51782 10220
rect 52181 10217 52193 10220
rect 52227 10217 52239 10251
rect 52181 10211 52239 10217
rect 52362 10208 52368 10260
rect 52420 10248 52426 10260
rect 53561 10251 53619 10257
rect 53561 10248 53573 10251
rect 52420 10220 53573 10248
rect 52420 10208 52426 10220
rect 53561 10217 53573 10220
rect 53607 10217 53619 10251
rect 53561 10211 53619 10217
rect 54938 10208 54944 10260
rect 54996 10248 55002 10260
rect 55125 10251 55183 10257
rect 55125 10248 55137 10251
rect 54996 10220 55137 10248
rect 54996 10208 55002 10220
rect 55125 10217 55137 10220
rect 55171 10217 55183 10251
rect 55398 10248 55404 10260
rect 55359 10220 55404 10248
rect 55125 10211 55183 10217
rect 55398 10208 55404 10220
rect 55456 10208 55462 10260
rect 55490 10208 55496 10260
rect 55548 10248 55554 10260
rect 60369 10251 60427 10257
rect 60369 10248 60381 10251
rect 55548 10220 60381 10248
rect 55548 10208 55554 10220
rect 60369 10217 60381 10220
rect 60415 10217 60427 10251
rect 60369 10211 60427 10217
rect 60734 10208 60740 10260
rect 60792 10248 60798 10260
rect 60829 10251 60887 10257
rect 60829 10248 60841 10251
rect 60792 10220 60841 10248
rect 60792 10208 60798 10220
rect 60829 10217 60841 10220
rect 60875 10217 60887 10251
rect 60829 10211 60887 10217
rect 60918 10208 60924 10260
rect 60976 10248 60982 10260
rect 64230 10248 64236 10260
rect 60976 10220 64236 10248
rect 60976 10208 60982 10220
rect 64230 10208 64236 10220
rect 64288 10208 64294 10260
rect 65242 10248 65248 10260
rect 65203 10220 65248 10248
rect 65242 10208 65248 10220
rect 65300 10208 65306 10260
rect 68738 10248 68744 10260
rect 68699 10220 68744 10248
rect 68738 10208 68744 10220
rect 68796 10208 68802 10260
rect 69382 10248 69388 10260
rect 69343 10220 69388 10248
rect 69382 10208 69388 10220
rect 69440 10208 69446 10260
rect 70305 10251 70363 10257
rect 70305 10217 70317 10251
rect 70351 10248 70363 10251
rect 70486 10248 70492 10260
rect 70351 10220 70492 10248
rect 70351 10217 70363 10220
rect 70305 10211 70363 10217
rect 70486 10208 70492 10220
rect 70544 10208 70550 10260
rect 70765 10251 70823 10257
rect 70765 10217 70777 10251
rect 70811 10248 70823 10251
rect 70854 10248 70860 10260
rect 70811 10220 70860 10248
rect 70811 10217 70823 10220
rect 70765 10211 70823 10217
rect 70854 10208 70860 10220
rect 70912 10208 70918 10260
rect 74442 10208 74448 10260
rect 74500 10248 74506 10260
rect 74813 10251 74871 10257
rect 74813 10248 74825 10251
rect 74500 10220 74825 10248
rect 74500 10208 74506 10220
rect 74813 10217 74825 10220
rect 74859 10217 74871 10251
rect 74813 10211 74871 10217
rect 75086 10208 75092 10260
rect 75144 10248 75150 10260
rect 75549 10251 75607 10257
rect 75549 10248 75561 10251
rect 75144 10220 75561 10248
rect 75144 10208 75150 10220
rect 75549 10217 75561 10220
rect 75595 10217 75607 10251
rect 76374 10248 76380 10260
rect 76335 10220 76380 10248
rect 75549 10211 75607 10217
rect 76374 10208 76380 10220
rect 76432 10208 76438 10260
rect 76558 10208 76564 10260
rect 76616 10248 76622 10260
rect 76745 10251 76803 10257
rect 76745 10248 76757 10251
rect 76616 10220 76757 10248
rect 76616 10208 76622 10220
rect 76745 10217 76757 10220
rect 76791 10217 76803 10251
rect 78214 10248 78220 10260
rect 78175 10220 78220 10248
rect 76745 10211 76803 10217
rect 78214 10208 78220 10220
rect 78272 10208 78278 10260
rect 78306 10208 78312 10260
rect 78364 10248 78370 10260
rect 78401 10251 78459 10257
rect 78401 10248 78413 10251
rect 78364 10220 78413 10248
rect 78364 10208 78370 10220
rect 78401 10217 78413 10220
rect 78447 10217 78459 10251
rect 79042 10248 79048 10260
rect 79003 10220 79048 10248
rect 78401 10211 78459 10217
rect 79042 10208 79048 10220
rect 79100 10208 79106 10260
rect 80238 10248 80244 10260
rect 80199 10220 80244 10248
rect 80238 10208 80244 10220
rect 80296 10208 80302 10260
rect 80422 10248 80428 10260
rect 80383 10220 80428 10248
rect 80422 10208 80428 10220
rect 80480 10208 80486 10260
rect 81526 10248 81532 10260
rect 81487 10220 81532 10248
rect 81526 10208 81532 10220
rect 81584 10208 81590 10260
rect 82722 10248 82728 10260
rect 82683 10220 82728 10248
rect 82722 10208 82728 10220
rect 82780 10208 82786 10260
rect 83550 10248 83556 10260
rect 83511 10220 83556 10248
rect 83550 10208 83556 10220
rect 83608 10208 83614 10260
rect 84654 10248 84660 10260
rect 84615 10220 84660 10248
rect 84654 10208 84660 10220
rect 84712 10208 84718 10260
rect 89441 10251 89499 10257
rect 89441 10217 89453 10251
rect 89487 10248 89499 10251
rect 93486 10248 93492 10260
rect 89487 10220 93492 10248
rect 89487 10217 89499 10220
rect 89441 10211 89499 10217
rect 41966 10180 41972 10192
rect 35492 10152 36124 10180
rect 36648 10152 41972 10180
rect 35492 10140 35498 10152
rect 26620 10084 27108 10112
rect 27433 10115 27491 10121
rect 26620 10053 26648 10084
rect 27433 10081 27445 10115
rect 27479 10112 27491 10115
rect 27614 10112 27620 10124
rect 27479 10084 27620 10112
rect 27479 10081 27491 10084
rect 27433 10075 27491 10081
rect 27614 10072 27620 10084
rect 27672 10072 27678 10124
rect 29362 10072 29368 10124
rect 29420 10112 29426 10124
rect 35989 10115 36047 10121
rect 35989 10112 36001 10115
rect 29420 10084 36001 10112
rect 29420 10072 29426 10084
rect 35989 10081 36001 10084
rect 36035 10081 36047 10115
rect 36096 10112 36124 10152
rect 41966 10140 41972 10152
rect 42024 10140 42030 10192
rect 42337 10183 42395 10189
rect 42337 10149 42349 10183
rect 42383 10180 42395 10183
rect 44542 10180 44548 10192
rect 42383 10152 44548 10180
rect 42383 10149 42395 10152
rect 42337 10143 42395 10149
rect 44542 10140 44548 10152
rect 44600 10140 44606 10192
rect 48958 10180 48964 10192
rect 45204 10152 48964 10180
rect 37090 10112 37096 10124
rect 36096 10084 37096 10112
rect 35989 10075 36047 10081
rect 37090 10072 37096 10084
rect 37148 10072 37154 10124
rect 37458 10112 37464 10124
rect 37419 10084 37464 10112
rect 37458 10072 37464 10084
rect 37516 10072 37522 10124
rect 37642 10112 37648 10124
rect 37603 10084 37648 10112
rect 37642 10072 37648 10084
rect 37700 10072 37706 10124
rect 37734 10072 37740 10124
rect 37792 10112 37798 10124
rect 38657 10115 38715 10121
rect 38657 10112 38669 10115
rect 37792 10084 38669 10112
rect 37792 10072 37798 10084
rect 38657 10081 38669 10084
rect 38703 10081 38715 10115
rect 38657 10075 38715 10081
rect 38838 10072 38844 10124
rect 38896 10112 38902 10124
rect 41233 10115 41291 10121
rect 38896 10084 41092 10112
rect 38896 10072 38902 10084
rect 24228 10016 26004 10044
rect 26605 10047 26663 10053
rect 24121 10007 24179 10013
rect 26605 10013 26617 10047
rect 26651 10013 26663 10047
rect 26605 10007 26663 10013
rect 26697 10047 26755 10053
rect 26697 10013 26709 10047
rect 26743 10044 26755 10047
rect 27154 10044 27160 10056
rect 26743 10016 27160 10044
rect 26743 10013 26755 10016
rect 26697 10007 26755 10013
rect 27154 10004 27160 10016
rect 27212 10004 27218 10056
rect 27798 10044 27804 10056
rect 27759 10016 27804 10044
rect 27798 10004 27804 10016
rect 27856 10004 27862 10056
rect 27890 10004 27896 10056
rect 27948 10044 27954 10056
rect 28261 10047 28319 10053
rect 27948 10016 27993 10044
rect 27948 10004 27954 10016
rect 28261 10013 28273 10047
rect 28307 10044 28319 10047
rect 28629 10047 28687 10053
rect 28629 10044 28641 10047
rect 28307 10016 28641 10044
rect 28307 10013 28319 10016
rect 28261 10007 28319 10013
rect 28629 10013 28641 10016
rect 28675 10044 28687 10047
rect 32398 10044 32404 10056
rect 28675 10016 32404 10044
rect 28675 10013 28687 10016
rect 28629 10007 28687 10013
rect 32398 10004 32404 10016
rect 32456 10004 32462 10056
rect 32582 10044 32588 10056
rect 32543 10016 32588 10044
rect 32582 10004 32588 10016
rect 32640 10004 32646 10056
rect 32674 10004 32680 10056
rect 32732 10044 32738 10056
rect 33045 10047 33103 10053
rect 32732 10016 32777 10044
rect 32732 10004 32738 10016
rect 33045 10013 33057 10047
rect 33091 10044 33103 10047
rect 33410 10044 33416 10056
rect 33091 10016 33416 10044
rect 33091 10013 33103 10016
rect 33045 10007 33103 10013
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 35066 10044 35072 10056
rect 35027 10016 35072 10044
rect 35066 10004 35072 10016
rect 35124 10004 35130 10056
rect 35529 10047 35587 10053
rect 35529 10013 35541 10047
rect 35575 10044 35587 10047
rect 35621 10047 35679 10053
rect 35621 10044 35633 10047
rect 35575 10016 35633 10044
rect 35575 10013 35587 10016
rect 35529 10007 35587 10013
rect 35621 10013 35633 10016
rect 35667 10013 35679 10047
rect 39114 10044 39120 10056
rect 35621 10007 35679 10013
rect 35728 10016 39120 10044
rect 8128 9948 21680 9976
rect 24210 9936 24216 9988
rect 24268 9976 24274 9988
rect 27522 9976 27528 9988
rect 24268 9948 27528 9976
rect 24268 9936 24274 9948
rect 27522 9936 27528 9948
rect 27580 9936 27586 9988
rect 27706 9936 27712 9988
rect 27764 9976 27770 9988
rect 30653 9979 30711 9985
rect 30653 9976 30665 9979
rect 27764 9948 30665 9976
rect 27764 9936 27770 9948
rect 30653 9945 30665 9948
rect 30699 9945 30711 9979
rect 30653 9939 30711 9945
rect 30742 9936 30748 9988
rect 30800 9976 30806 9988
rect 30800 9948 33548 9976
rect 30800 9936 30806 9948
rect 7098 9908 7104 9920
rect 6043 9880 7104 9908
rect 6043 9877 6055 9880
rect 5997 9871 6055 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 16393 9911 16451 9917
rect 16393 9877 16405 9911
rect 16439 9908 16451 9911
rect 17310 9908 17316 9920
rect 16439 9880 17316 9908
rect 16439 9877 16451 9880
rect 16393 9871 16451 9877
rect 17310 9868 17316 9880
rect 17368 9868 17374 9920
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 24026 9908 24032 9920
rect 19935 9880 24032 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 24026 9868 24032 9880
rect 24084 9868 24090 9920
rect 24118 9868 24124 9920
rect 24176 9908 24182 9920
rect 27982 9908 27988 9920
rect 24176 9880 27988 9908
rect 24176 9868 24182 9880
rect 27982 9868 27988 9880
rect 28040 9868 28046 9920
rect 28074 9868 28080 9920
rect 28132 9908 28138 9920
rect 28994 9908 29000 9920
rect 28132 9880 29000 9908
rect 28132 9868 28138 9880
rect 28994 9868 29000 9880
rect 29052 9868 29058 9920
rect 29089 9911 29147 9917
rect 29089 9877 29101 9911
rect 29135 9908 29147 9911
rect 29638 9908 29644 9920
rect 29135 9880 29644 9908
rect 29135 9877 29147 9880
rect 29089 9871 29147 9877
rect 29638 9868 29644 9880
rect 29696 9868 29702 9920
rect 30282 9908 30288 9920
rect 30243 9880 30288 9908
rect 30282 9868 30288 9880
rect 30340 9868 30346 9920
rect 32125 9911 32183 9917
rect 32125 9877 32137 9911
rect 32171 9908 32183 9911
rect 32214 9908 32220 9920
rect 32171 9880 32220 9908
rect 32171 9877 32183 9880
rect 32125 9871 32183 9877
rect 32214 9868 32220 9880
rect 32272 9868 32278 9920
rect 33410 9908 33416 9920
rect 33371 9880 33416 9908
rect 33410 9868 33416 9880
rect 33468 9868 33474 9920
rect 33520 9908 33548 9948
rect 33870 9936 33876 9988
rect 33928 9976 33934 9988
rect 35728 9976 35756 10016
rect 39114 10004 39120 10016
rect 39172 10004 39178 10056
rect 39209 10047 39267 10053
rect 39209 10013 39221 10047
rect 39255 10044 39267 10047
rect 39301 10047 39359 10053
rect 39301 10044 39313 10047
rect 39255 10016 39313 10044
rect 39255 10013 39267 10016
rect 39209 10007 39267 10013
rect 39301 10013 39313 10016
rect 39347 10013 39359 10047
rect 39301 10007 39359 10013
rect 40681 10047 40739 10053
rect 40681 10013 40693 10047
rect 40727 10044 40739 10047
rect 40957 10047 41015 10053
rect 40957 10044 40969 10047
rect 40727 10016 40969 10044
rect 40727 10013 40739 10016
rect 40681 10007 40739 10013
rect 40957 10013 40969 10016
rect 41003 10013 41015 10047
rect 41064 10044 41092 10084
rect 41233 10081 41245 10115
rect 41279 10112 41291 10115
rect 45094 10112 45100 10124
rect 41279 10084 45100 10112
rect 41279 10081 41291 10084
rect 41233 10075 41291 10081
rect 45094 10072 45100 10084
rect 45152 10072 45158 10124
rect 45204 10044 45232 10152
rect 48958 10140 48964 10152
rect 49016 10140 49022 10192
rect 49694 10180 49700 10192
rect 49655 10152 49700 10180
rect 49694 10140 49700 10152
rect 49752 10140 49758 10192
rect 49878 10180 49884 10192
rect 49839 10152 49884 10180
rect 49878 10140 49884 10152
rect 49936 10140 49942 10192
rect 50816 10152 51028 10180
rect 45278 10072 45284 10124
rect 45336 10112 45342 10124
rect 50816 10112 50844 10152
rect 45336 10084 50844 10112
rect 51000 10112 51028 10152
rect 51258 10140 51264 10192
rect 51316 10180 51322 10192
rect 73157 10183 73215 10189
rect 73157 10180 73169 10183
rect 51316 10152 73169 10180
rect 51316 10140 51322 10152
rect 73157 10149 73169 10152
rect 73203 10149 73215 10183
rect 73157 10143 73215 10149
rect 73433 10183 73491 10189
rect 73433 10149 73445 10183
rect 73479 10180 73491 10183
rect 79410 10180 79416 10192
rect 73479 10152 77892 10180
rect 79371 10152 79416 10180
rect 73479 10149 73491 10152
rect 73433 10143 73491 10149
rect 55490 10112 55496 10124
rect 51000 10084 55496 10112
rect 45336 10072 45342 10084
rect 55490 10072 55496 10084
rect 55548 10072 55554 10124
rect 56134 10112 56140 10124
rect 56095 10084 56140 10112
rect 56134 10072 56140 10084
rect 56192 10072 56198 10124
rect 56229 10115 56287 10121
rect 56229 10081 56241 10115
rect 56275 10112 56287 10115
rect 56502 10112 56508 10124
rect 56275 10084 56508 10112
rect 56275 10081 56287 10084
rect 56229 10075 56287 10081
rect 56502 10072 56508 10084
rect 56560 10072 56566 10124
rect 57164 10084 57652 10112
rect 45830 10044 45836 10056
rect 41064 10016 45232 10044
rect 45791 10016 45836 10044
rect 40957 10007 41015 10013
rect 45830 10004 45836 10016
rect 45888 10004 45894 10056
rect 46201 10047 46259 10053
rect 46201 10013 46213 10047
rect 46247 10013 46259 10047
rect 46201 10007 46259 10013
rect 46569 10047 46627 10053
rect 46569 10013 46581 10047
rect 46615 10044 46627 10047
rect 46937 10047 46995 10053
rect 46937 10044 46949 10047
rect 46615 10016 46949 10044
rect 46615 10013 46627 10016
rect 46569 10007 46627 10013
rect 46937 10013 46949 10016
rect 46983 10044 46995 10047
rect 48222 10044 48228 10056
rect 46983 10016 48228 10044
rect 46983 10013 46995 10016
rect 46937 10007 46995 10013
rect 33928 9948 35756 9976
rect 35989 9979 36047 9985
rect 33928 9936 33934 9948
rect 35989 9945 36001 9979
rect 36035 9976 36047 9979
rect 42337 9979 42395 9985
rect 42337 9976 42349 9979
rect 36035 9948 42349 9976
rect 36035 9945 36047 9948
rect 35989 9939 36047 9945
rect 42337 9945 42349 9948
rect 42383 9945 42395 9979
rect 46216 9976 46244 10007
rect 48222 10004 48228 10016
rect 48280 10004 48286 10056
rect 48406 10044 48412 10056
rect 48367 10016 48412 10044
rect 48406 10004 48412 10016
rect 48464 10004 48470 10056
rect 48961 10047 49019 10053
rect 48961 10013 48973 10047
rect 49007 10044 49019 10047
rect 49053 10047 49111 10053
rect 49053 10044 49065 10047
rect 49007 10016 49065 10044
rect 49007 10013 49019 10016
rect 48961 10007 49019 10013
rect 49053 10013 49065 10016
rect 49099 10013 49111 10047
rect 49970 10044 49976 10056
rect 49931 10016 49976 10044
rect 49053 10007 49111 10013
rect 49970 10004 49976 10016
rect 50028 10004 50034 10056
rect 50525 10047 50583 10053
rect 50525 10013 50537 10047
rect 50571 10044 50583 10047
rect 50890 10044 50896 10056
rect 50571 10016 50896 10044
rect 50571 10013 50583 10016
rect 50525 10007 50583 10013
rect 50890 10004 50896 10016
rect 50948 10004 50954 10056
rect 51626 10044 51632 10056
rect 51587 10016 51632 10044
rect 51626 10004 51632 10016
rect 51684 10004 51690 10056
rect 51721 10047 51779 10053
rect 51721 10013 51733 10047
rect 51767 10013 51779 10047
rect 51721 10007 51779 10013
rect 52089 10047 52147 10053
rect 52089 10013 52101 10047
rect 52135 10013 52147 10047
rect 52089 10007 52147 10013
rect 52181 10047 52239 10053
rect 52181 10013 52193 10047
rect 52227 10044 52239 10047
rect 52457 10047 52515 10053
rect 52457 10044 52469 10047
rect 52227 10016 52469 10044
rect 52227 10013 52239 10016
rect 52181 10007 52239 10013
rect 52457 10013 52469 10016
rect 52503 10044 52515 10047
rect 53374 10044 53380 10056
rect 52503 10016 53380 10044
rect 52503 10013 52515 10016
rect 52457 10007 52515 10013
rect 42337 9939 42395 9945
rect 42444 9948 46244 9976
rect 35342 9908 35348 9920
rect 33520 9880 35348 9908
rect 35342 9868 35348 9880
rect 35400 9868 35406 9920
rect 36078 9868 36084 9920
rect 36136 9908 36142 9920
rect 36265 9911 36323 9917
rect 36265 9908 36277 9911
rect 36136 9880 36277 9908
rect 36136 9868 36142 9880
rect 36265 9877 36277 9880
rect 36311 9908 36323 9911
rect 36998 9908 37004 9920
rect 36311 9880 37004 9908
rect 36311 9877 36323 9880
rect 36265 9871 36323 9877
rect 36998 9868 37004 9880
rect 37056 9868 37062 9920
rect 37090 9868 37096 9920
rect 37148 9908 37154 9920
rect 39206 9908 39212 9920
rect 37148 9880 39212 9908
rect 37148 9868 37154 9880
rect 39206 9868 39212 9880
rect 39264 9868 39270 9920
rect 39301 9911 39359 9917
rect 39301 9877 39313 9911
rect 39347 9908 39359 9911
rect 39577 9911 39635 9917
rect 39577 9908 39589 9911
rect 39347 9880 39589 9908
rect 39347 9877 39359 9880
rect 39301 9871 39359 9877
rect 39577 9877 39589 9880
rect 39623 9908 39635 9911
rect 40034 9908 40040 9920
rect 39623 9880 40040 9908
rect 39623 9877 39635 9880
rect 39577 9871 39635 9877
rect 40034 9868 40040 9880
rect 40092 9868 40098 9920
rect 40402 9868 40408 9920
rect 40460 9908 40466 9920
rect 42444 9908 42472 9948
rect 47118 9936 47124 9988
rect 47176 9976 47182 9988
rect 47305 9979 47363 9985
rect 47305 9976 47317 9979
rect 47176 9948 47317 9976
rect 47176 9936 47182 9948
rect 47305 9945 47317 9948
rect 47351 9976 47363 9979
rect 50246 9976 50252 9988
rect 47351 9948 50252 9976
rect 47351 9945 47363 9948
rect 47305 9939 47363 9945
rect 50246 9936 50252 9948
rect 50304 9936 50310 9988
rect 50338 9936 50344 9988
rect 50396 9976 50402 9988
rect 51736 9976 51764 10007
rect 50396 9948 51764 9976
rect 50396 9936 50402 9948
rect 42610 9908 42616 9920
rect 40460 9880 42472 9908
rect 42571 9880 42616 9908
rect 40460 9868 40466 9880
rect 42610 9868 42616 9880
rect 42668 9868 42674 9920
rect 43162 9908 43168 9920
rect 43123 9880 43168 9908
rect 43162 9868 43168 9880
rect 43220 9868 43226 9920
rect 44082 9868 44088 9920
rect 44140 9908 44146 9920
rect 50614 9908 50620 9920
rect 44140 9880 50620 9908
rect 44140 9868 44146 9880
rect 50614 9868 50620 9880
rect 50672 9868 50678 9920
rect 50706 9868 50712 9920
rect 50764 9908 50770 9920
rect 51169 9911 51227 9917
rect 51169 9908 51181 9911
rect 50764 9880 51181 9908
rect 50764 9868 50770 9880
rect 51169 9877 51181 9880
rect 51215 9877 51227 9911
rect 52104 9908 52132 10007
rect 53374 10004 53380 10016
rect 53432 10004 53438 10056
rect 55585 10047 55643 10053
rect 55585 10013 55597 10047
rect 55631 10044 55643 10047
rect 55858 10044 55864 10056
rect 55631 10016 55864 10044
rect 55631 10013 55643 10016
rect 55585 10007 55643 10013
rect 55858 10004 55864 10016
rect 55916 10004 55922 10056
rect 56045 10047 56103 10053
rect 56045 10013 56057 10047
rect 56091 10013 56103 10047
rect 56045 10007 56103 10013
rect 56413 10047 56471 10053
rect 56413 10013 56425 10047
rect 56459 10044 56471 10047
rect 56778 10044 56784 10056
rect 56459 10016 56784 10044
rect 56459 10013 56471 10016
rect 56413 10007 56471 10013
rect 53285 9979 53343 9985
rect 53285 9945 53297 9979
rect 53331 9976 53343 9979
rect 53466 9976 53472 9988
rect 53331 9948 53472 9976
rect 53331 9945 53343 9948
rect 53285 9939 53343 9945
rect 53466 9936 53472 9948
rect 53524 9936 53530 9988
rect 54478 9976 54484 9988
rect 53576 9948 54484 9976
rect 52825 9911 52883 9917
rect 52825 9908 52837 9911
rect 52104 9880 52837 9908
rect 51169 9871 51227 9877
rect 52825 9877 52837 9880
rect 52871 9908 52883 9911
rect 53576 9908 53604 9948
rect 54478 9936 54484 9948
rect 54536 9936 54542 9988
rect 54570 9936 54576 9988
rect 54628 9976 54634 9988
rect 54628 9948 55904 9976
rect 54628 9936 54634 9948
rect 55876 9920 55904 9948
rect 52871 9880 53604 9908
rect 54297 9911 54355 9917
rect 52871 9877 52883 9880
rect 52825 9871 52883 9877
rect 54297 9877 54309 9911
rect 54343 9908 54355 9911
rect 55122 9908 55128 9920
rect 54343 9880 55128 9908
rect 54343 9877 54355 9880
rect 54297 9871 54355 9877
rect 55122 9868 55128 9880
rect 55180 9868 55186 9920
rect 55858 9868 55864 9920
rect 55916 9868 55922 9920
rect 56060 9908 56088 10007
rect 56778 10004 56784 10016
rect 56836 10004 56842 10056
rect 57164 10053 57192 10084
rect 57149 10047 57207 10053
rect 57149 10013 57161 10047
rect 57195 10013 57207 10047
rect 57149 10007 57207 10013
rect 57241 10047 57299 10053
rect 57241 10013 57253 10047
rect 57287 10044 57299 10047
rect 57517 10047 57575 10053
rect 57287 10016 57468 10044
rect 57287 10013 57299 10016
rect 57241 10007 57299 10013
rect 57440 9988 57468 10016
rect 57517 10013 57529 10047
rect 57563 10013 57575 10047
rect 57624 10044 57652 10084
rect 57698 10072 57704 10124
rect 57756 10112 57762 10124
rect 57756 10084 57801 10112
rect 57756 10072 57762 10084
rect 57882 10072 57888 10124
rect 57940 10112 57946 10124
rect 58989 10115 59047 10121
rect 58989 10112 59001 10115
rect 57940 10084 59001 10112
rect 57940 10072 57946 10084
rect 58989 10081 59001 10084
rect 59035 10081 59047 10115
rect 59446 10112 59452 10124
rect 58989 10075 59047 10081
rect 59096 10084 59452 10112
rect 57790 10044 57796 10056
rect 57624 10016 57796 10044
rect 57517 10007 57575 10013
rect 56594 9936 56600 9988
rect 56652 9976 56658 9988
rect 57054 9976 57060 9988
rect 56652 9948 57060 9976
rect 56652 9936 56658 9948
rect 57054 9936 57060 9948
rect 57112 9936 57118 9988
rect 57422 9936 57428 9988
rect 57480 9936 57486 9988
rect 57532 9976 57560 10007
rect 57790 10004 57796 10016
rect 57848 10044 57854 10056
rect 58618 10044 58624 10056
rect 57848 10016 58624 10044
rect 57848 10004 57854 10016
rect 58618 10004 58624 10016
rect 58676 10004 58682 10056
rect 58713 10047 58771 10053
rect 58713 10013 58725 10047
rect 58759 10044 58771 10047
rect 59096 10044 59124 10084
rect 59446 10072 59452 10084
rect 59504 10072 59510 10124
rect 60734 10112 60740 10124
rect 59648 10084 60740 10112
rect 59648 10053 59676 10084
rect 60734 10072 60740 10084
rect 60792 10072 60798 10124
rect 68922 10112 68928 10124
rect 68883 10084 68928 10112
rect 68922 10072 68928 10084
rect 68980 10072 68986 10124
rect 72050 10072 72056 10124
rect 72108 10112 72114 10124
rect 72108 10084 72153 10112
rect 72108 10072 72114 10084
rect 72234 10072 72240 10124
rect 72292 10112 72298 10124
rect 73249 10115 73307 10121
rect 73249 10112 73261 10115
rect 72292 10084 73261 10112
rect 72292 10072 72298 10084
rect 58759 10016 59124 10044
rect 59265 10047 59323 10053
rect 58759 10013 58771 10016
rect 58713 10007 58771 10013
rect 59265 10013 59277 10047
rect 59311 10044 59323 10047
rect 59633 10047 59691 10053
rect 59633 10044 59645 10047
rect 59311 10016 59645 10044
rect 59311 10013 59323 10016
rect 59265 10007 59323 10013
rect 59633 10013 59645 10016
rect 59679 10013 59691 10047
rect 59814 10044 59820 10056
rect 59775 10016 59820 10044
rect 59633 10007 59691 10013
rect 59814 10004 59820 10016
rect 59872 10004 59878 10056
rect 60185 10047 60243 10053
rect 60185 10013 60197 10047
rect 60231 10044 60243 10047
rect 60458 10044 60464 10056
rect 60231 10016 60464 10044
rect 60231 10013 60243 10016
rect 60185 10007 60243 10013
rect 60458 10004 60464 10016
rect 60516 10004 60522 10056
rect 60550 10004 60556 10056
rect 60608 10044 60614 10056
rect 61013 10047 61071 10053
rect 61013 10044 61025 10047
rect 60608 10016 61025 10044
rect 60608 10004 60614 10016
rect 61013 10013 61025 10016
rect 61059 10013 61071 10047
rect 62022 10044 62028 10056
rect 61983 10016 62028 10044
rect 61013 10007 61071 10013
rect 62022 10004 62028 10016
rect 62080 10004 62086 10056
rect 62758 10004 62764 10056
rect 62816 10044 62822 10056
rect 70121 10047 70179 10053
rect 70121 10044 70133 10047
rect 62816 10016 70133 10044
rect 62816 10004 62822 10016
rect 70121 10013 70133 10016
rect 70167 10013 70179 10047
rect 70854 10044 70860 10056
rect 70815 10016 70860 10044
rect 70121 10007 70179 10013
rect 70854 10004 70860 10016
rect 70912 10004 70918 10056
rect 71406 10044 71412 10056
rect 71367 10016 71412 10044
rect 71406 10004 71412 10016
rect 71464 10044 71470 10056
rect 71685 10047 71743 10053
rect 71685 10044 71697 10047
rect 71464 10016 71697 10044
rect 71464 10004 71470 10016
rect 71685 10013 71697 10016
rect 71731 10013 71743 10047
rect 72418 10044 72424 10056
rect 72379 10016 72424 10044
rect 71685 10007 71743 10013
rect 72418 10004 72424 10016
rect 72476 10004 72482 10056
rect 72602 10044 72608 10056
rect 72563 10016 72608 10044
rect 72602 10004 72608 10016
rect 72660 10004 72666 10056
rect 72804 10053 72832 10084
rect 73249 10081 73261 10084
rect 73295 10081 73307 10115
rect 73249 10075 73307 10081
rect 72789 10047 72847 10053
rect 72789 10013 72801 10047
rect 72835 10013 72847 10047
rect 72789 10007 72847 10013
rect 73157 10047 73215 10053
rect 73157 10013 73169 10047
rect 73203 10044 73215 10047
rect 73890 10044 73896 10056
rect 73203 10016 73896 10044
rect 73203 10013 73215 10016
rect 73157 10007 73215 10013
rect 73890 10004 73896 10016
rect 73948 10004 73954 10056
rect 74074 10044 74080 10056
rect 74035 10016 74080 10044
rect 74074 10004 74080 10016
rect 74132 10004 74138 10056
rect 74169 10047 74227 10053
rect 74169 10013 74181 10047
rect 74215 10013 74227 10047
rect 74350 10044 74356 10056
rect 74311 10016 74356 10044
rect 74169 10007 74227 10013
rect 57977 9979 58035 9985
rect 57977 9976 57989 9979
rect 57532 9948 57989 9976
rect 57977 9945 57989 9948
rect 58023 9976 58035 9979
rect 60274 9976 60280 9988
rect 58023 9948 60280 9976
rect 58023 9945 58035 9948
rect 57977 9939 58035 9945
rect 60274 9936 60280 9948
rect 60332 9936 60338 9988
rect 60369 9979 60427 9985
rect 60369 9945 60381 9979
rect 60415 9976 60427 9979
rect 74184 9976 74212 10007
rect 74350 10004 74356 10016
rect 74408 10044 74414 10056
rect 75181 10047 75239 10053
rect 75181 10044 75193 10047
rect 74408 10016 75193 10044
rect 74408 10004 74414 10016
rect 75181 10013 75193 10016
rect 75227 10013 75239 10047
rect 75181 10007 75239 10013
rect 76285 10047 76343 10053
rect 76285 10013 76297 10047
rect 76331 10044 76343 10047
rect 76558 10044 76564 10056
rect 76331 10016 76564 10044
rect 76331 10013 76343 10016
rect 76285 10007 76343 10013
rect 76558 10004 76564 10016
rect 76616 10004 76622 10056
rect 77294 10044 77300 10056
rect 77255 10016 77300 10044
rect 77294 10004 77300 10016
rect 77352 10044 77358 10056
rect 77757 10047 77815 10053
rect 77757 10044 77769 10047
rect 77352 10016 77769 10044
rect 77352 10004 77358 10016
rect 77757 10013 77769 10016
rect 77803 10013 77815 10047
rect 77757 10007 77815 10013
rect 77386 9976 77392 9988
rect 60415 9948 74212 9976
rect 77347 9948 77392 9976
rect 60415 9945 60427 9948
rect 60369 9939 60427 9945
rect 77386 9936 77392 9948
rect 77444 9936 77450 9988
rect 77864 9976 77892 10152
rect 79410 10140 79416 10152
rect 79468 10140 79474 10192
rect 79781 10115 79839 10121
rect 79781 10112 79793 10115
rect 79336 10084 79793 10112
rect 78030 10004 78036 10056
rect 78088 10044 78094 10056
rect 78309 10047 78367 10053
rect 78309 10044 78321 10047
rect 78088 10016 78321 10044
rect 78088 10004 78094 10016
rect 78309 10013 78321 10016
rect 78355 10013 78367 10047
rect 78309 10007 78367 10013
rect 78398 10004 78404 10056
rect 78456 10044 78462 10056
rect 79336 10053 79364 10084
rect 79781 10081 79793 10084
rect 79827 10081 79839 10115
rect 79781 10075 79839 10081
rect 80057 10115 80115 10121
rect 80057 10081 80069 10115
rect 80103 10112 80115 10115
rect 83001 10115 83059 10121
rect 83001 10112 83013 10115
rect 80103 10084 83013 10112
rect 80103 10081 80115 10084
rect 80057 10075 80115 10081
rect 83001 10081 83013 10084
rect 83047 10081 83059 10115
rect 83001 10075 83059 10081
rect 83921 10115 83979 10121
rect 83921 10081 83933 10115
rect 83967 10112 83979 10115
rect 84672 10112 84700 10208
rect 85206 10140 85212 10192
rect 85264 10180 85270 10192
rect 85264 10152 86080 10180
rect 85264 10140 85270 10152
rect 83967 10084 84700 10112
rect 85025 10115 85083 10121
rect 83967 10081 83979 10084
rect 83921 10075 83979 10081
rect 85025 10081 85037 10115
rect 85071 10112 85083 10115
rect 85114 10112 85120 10124
rect 85071 10084 85120 10112
rect 85071 10081 85083 10084
rect 85025 10075 85083 10081
rect 85114 10072 85120 10084
rect 85172 10112 85178 10124
rect 85942 10112 85948 10124
rect 85172 10084 85948 10112
rect 85172 10072 85178 10084
rect 85942 10072 85948 10084
rect 86000 10072 86006 10124
rect 86052 10121 86080 10152
rect 86037 10115 86095 10121
rect 86037 10081 86049 10115
rect 86083 10081 86095 10115
rect 86037 10075 86095 10081
rect 87230 10072 87236 10124
rect 87288 10112 87294 10124
rect 88521 10115 88579 10121
rect 88521 10112 88533 10115
rect 87288 10084 88533 10112
rect 87288 10072 87294 10084
rect 88521 10081 88533 10084
rect 88567 10081 88579 10115
rect 89456 10112 89484 10211
rect 93486 10208 93492 10220
rect 93544 10208 93550 10260
rect 95878 10248 95884 10260
rect 95839 10220 95884 10248
rect 95878 10208 95884 10220
rect 95936 10208 95942 10260
rect 97997 10251 98055 10257
rect 97997 10217 98009 10251
rect 98043 10248 98055 10251
rect 98270 10248 98276 10260
rect 98043 10220 98276 10248
rect 98043 10217 98055 10220
rect 97997 10211 98055 10217
rect 91925 10183 91983 10189
rect 91925 10149 91937 10183
rect 91971 10180 91983 10183
rect 92382 10180 92388 10192
rect 91971 10152 92388 10180
rect 91971 10149 91983 10152
rect 91925 10143 91983 10149
rect 92382 10140 92388 10152
rect 92440 10140 92446 10192
rect 88521 10075 88579 10081
rect 88996 10084 89484 10112
rect 79321 10047 79379 10053
rect 79321 10044 79333 10047
rect 78456 10016 79333 10044
rect 78456 10004 78462 10016
rect 79321 10013 79333 10016
rect 79367 10013 79379 10047
rect 79321 10007 79379 10013
rect 79502 10004 79508 10056
rect 79560 10044 79566 10056
rect 80333 10047 80391 10053
rect 80333 10044 80345 10047
rect 79560 10016 80345 10044
rect 79560 10004 79566 10016
rect 80333 10013 80345 10016
rect 80379 10044 80391 10047
rect 80793 10047 80851 10053
rect 80793 10044 80805 10047
rect 80379 10016 80805 10044
rect 80379 10013 80391 10016
rect 80333 10007 80391 10013
rect 80793 10013 80805 10016
rect 80839 10013 80851 10047
rect 80793 10007 80851 10013
rect 81066 10004 81072 10056
rect 81124 10044 81130 10056
rect 81897 10047 81955 10053
rect 81897 10044 81909 10047
rect 81124 10016 81909 10044
rect 81124 10004 81130 10016
rect 81897 10013 81909 10016
rect 81943 10044 81955 10047
rect 82357 10047 82415 10053
rect 82357 10044 82369 10047
rect 81943 10016 82369 10044
rect 81943 10013 81955 10016
rect 81897 10007 81955 10013
rect 82357 10013 82369 10016
rect 82403 10013 82415 10047
rect 82906 10044 82912 10056
rect 82867 10016 82912 10044
rect 82357 10007 82415 10013
rect 82906 10004 82912 10016
rect 82964 10004 82970 10056
rect 88996 10053 89024 10084
rect 90358 10072 90364 10124
rect 90416 10112 90422 10124
rect 90453 10115 90511 10121
rect 90453 10112 90465 10115
rect 90416 10084 90465 10112
rect 90416 10072 90422 10084
rect 90453 10081 90465 10084
rect 90499 10081 90511 10115
rect 90453 10075 90511 10081
rect 92750 10072 92756 10124
rect 92808 10112 92814 10124
rect 94133 10115 94191 10121
rect 94133 10112 94145 10115
rect 92808 10084 94145 10112
rect 92808 10072 92814 10084
rect 94133 10081 94145 10084
rect 94179 10081 94191 10115
rect 95896 10112 95924 10208
rect 97534 10180 97540 10192
rect 97495 10152 97540 10180
rect 97534 10140 97540 10152
rect 97592 10140 97598 10192
rect 96065 10115 96123 10121
rect 96065 10112 96077 10115
rect 95896 10084 96077 10112
rect 94133 10075 94191 10081
rect 96065 10081 96077 10084
rect 96111 10081 96123 10115
rect 96065 10075 96123 10081
rect 86589 10047 86647 10053
rect 86589 10013 86601 10047
rect 86635 10044 86647 10047
rect 87509 10047 87567 10053
rect 86635 10016 87000 10044
rect 86635 10013 86647 10016
rect 86589 10007 86647 10013
rect 81989 9979 82047 9985
rect 81989 9976 82001 9979
rect 77864 9948 82001 9976
rect 81989 9945 82001 9948
rect 82035 9945 82047 9979
rect 81989 9939 82047 9945
rect 86972 9920 87000 10016
rect 87509 10013 87521 10047
rect 87555 10013 87567 10047
rect 87509 10007 87567 10013
rect 88981 10047 89039 10053
rect 88981 10013 88993 10047
rect 89027 10013 89039 10047
rect 91922 10044 91928 10056
rect 91883 10016 91928 10044
rect 88981 10007 89039 10013
rect 56781 9911 56839 9917
rect 56781 9908 56793 9911
rect 56060 9880 56793 9908
rect 56781 9877 56793 9880
rect 56827 9908 56839 9911
rect 57701 9911 57759 9917
rect 57701 9908 57713 9911
rect 56827 9880 57713 9908
rect 56827 9877 56839 9880
rect 56781 9871 56839 9877
rect 57701 9877 57713 9880
rect 57747 9877 57759 9911
rect 57701 9871 57759 9877
rect 58529 9911 58587 9917
rect 58529 9877 58541 9911
rect 58575 9908 58587 9911
rect 58713 9911 58771 9917
rect 58713 9908 58725 9911
rect 58575 9880 58725 9908
rect 58575 9877 58587 9880
rect 58529 9871 58587 9877
rect 58713 9877 58725 9880
rect 58759 9877 58771 9911
rect 58713 9871 58771 9877
rect 58897 9911 58955 9917
rect 58897 9877 58909 9911
rect 58943 9908 58955 9911
rect 58989 9911 59047 9917
rect 58989 9908 59001 9911
rect 58943 9880 59001 9908
rect 58943 9877 58955 9880
rect 58897 9871 58955 9877
rect 58989 9877 59001 9880
rect 59035 9908 59047 9911
rect 60918 9908 60924 9920
rect 59035 9880 60924 9908
rect 59035 9877 59047 9880
rect 58989 9871 59047 9877
rect 60918 9868 60924 9880
rect 60976 9868 60982 9920
rect 61286 9868 61292 9920
rect 61344 9908 61350 9920
rect 63037 9911 63095 9917
rect 63037 9908 63049 9911
rect 61344 9880 63049 9908
rect 61344 9868 61350 9880
rect 63037 9877 63049 9880
rect 63083 9877 63095 9911
rect 66254 9908 66260 9920
rect 66215 9880 66260 9908
rect 63037 9871 63095 9877
rect 66254 9868 66260 9880
rect 66312 9868 66318 9920
rect 70121 9911 70179 9917
rect 70121 9877 70133 9911
rect 70167 9908 70179 9911
rect 73433 9911 73491 9917
rect 73433 9908 73445 9911
rect 70167 9880 73445 9908
rect 70167 9877 70179 9880
rect 70121 9871 70179 9877
rect 73433 9877 73445 9880
rect 73479 9877 73491 9911
rect 73614 9908 73620 9920
rect 73575 9880 73620 9908
rect 73433 9871 73491 9877
rect 73614 9868 73620 9880
rect 73672 9868 73678 9920
rect 76101 9911 76159 9917
rect 76101 9877 76113 9911
rect 76147 9908 76159 9911
rect 76282 9908 76288 9920
rect 76147 9880 76288 9908
rect 76147 9877 76159 9880
rect 76101 9871 76159 9877
rect 76282 9868 76288 9880
rect 76340 9868 76346 9920
rect 78490 9868 78496 9920
rect 78548 9908 78554 9920
rect 80057 9911 80115 9917
rect 80057 9908 80069 9911
rect 78548 9880 80069 9908
rect 78548 9868 78554 9880
rect 80057 9877 80069 9880
rect 80103 9877 80115 9911
rect 86954 9908 86960 9920
rect 86915 9880 86960 9908
rect 80057 9871 80115 9877
rect 86954 9868 86960 9880
rect 87012 9868 87018 9920
rect 87230 9908 87236 9920
rect 87191 9880 87236 9908
rect 87230 9868 87236 9880
rect 87288 9908 87294 9920
rect 87524 9908 87552 10007
rect 91922 10004 91928 10016
rect 91980 10044 91986 10056
rect 92293 10047 92351 10053
rect 92293 10044 92305 10047
rect 91980 10016 92305 10044
rect 91980 10004 91986 10016
rect 92293 10013 92305 10016
rect 92339 10013 92351 10047
rect 92293 10007 92351 10013
rect 92658 10004 92664 10056
rect 92716 10044 92722 10056
rect 93121 10047 93179 10053
rect 93121 10044 93133 10047
rect 92716 10016 93133 10044
rect 92716 10004 92722 10016
rect 93121 10013 93133 10016
rect 93167 10044 93179 10047
rect 93302 10044 93308 10056
rect 93167 10016 93308 10044
rect 93167 10013 93179 10016
rect 93121 10007 93179 10013
rect 93302 10004 93308 10016
rect 93360 10004 93366 10056
rect 94222 10044 94228 10056
rect 94183 10016 94228 10044
rect 94222 10004 94228 10016
rect 94280 10044 94286 10056
rect 94961 10047 95019 10053
rect 94961 10044 94973 10047
rect 94280 10016 94973 10044
rect 94280 10004 94286 10016
rect 94961 10013 94973 10016
rect 95007 10013 95019 10047
rect 94961 10007 95019 10013
rect 97629 10047 97687 10053
rect 97629 10013 97641 10047
rect 97675 10044 97687 10047
rect 98012 10044 98040 10211
rect 98270 10208 98276 10220
rect 98328 10208 98334 10260
rect 98362 10208 98368 10260
rect 98420 10248 98426 10260
rect 98457 10251 98515 10257
rect 98457 10248 98469 10251
rect 98420 10220 98469 10248
rect 98420 10208 98426 10220
rect 98457 10217 98469 10220
rect 98503 10217 98515 10251
rect 99558 10248 99564 10260
rect 99519 10220 99564 10248
rect 98457 10211 98515 10217
rect 99558 10208 99564 10220
rect 99616 10248 99622 10260
rect 107654 10248 107660 10260
rect 99616 10220 99696 10248
rect 107615 10220 107660 10248
rect 99616 10208 99622 10220
rect 98914 10112 98920 10124
rect 98875 10084 98920 10112
rect 98914 10072 98920 10084
rect 98972 10072 98978 10124
rect 99668 10121 99696 10220
rect 107654 10208 107660 10220
rect 107712 10208 107718 10260
rect 108942 10248 108948 10260
rect 108903 10220 108948 10248
rect 108942 10208 108948 10220
rect 109000 10208 109006 10260
rect 109678 10208 109684 10260
rect 109736 10248 109742 10260
rect 110966 10248 110972 10260
rect 109736 10220 110972 10248
rect 109736 10208 109742 10220
rect 110966 10208 110972 10220
rect 111024 10208 111030 10260
rect 111334 10208 111340 10260
rect 111392 10248 111398 10260
rect 111429 10251 111487 10257
rect 111429 10248 111441 10251
rect 111392 10220 111441 10248
rect 111392 10208 111398 10220
rect 111429 10217 111441 10220
rect 111475 10217 111487 10251
rect 111429 10211 111487 10217
rect 112809 10251 112867 10257
rect 112809 10217 112821 10251
rect 112855 10248 112867 10251
rect 116946 10248 116952 10260
rect 112855 10220 116952 10248
rect 112855 10217 112867 10220
rect 112809 10211 112867 10217
rect 116946 10208 116952 10220
rect 117004 10208 117010 10260
rect 117130 10248 117136 10260
rect 117091 10220 117136 10248
rect 117130 10208 117136 10220
rect 117188 10208 117194 10260
rect 119433 10251 119491 10257
rect 119433 10217 119445 10251
rect 119479 10248 119491 10251
rect 119522 10248 119528 10260
rect 119479 10220 119528 10248
rect 119479 10217 119491 10220
rect 119433 10211 119491 10217
rect 119522 10208 119528 10220
rect 119580 10208 119586 10260
rect 119614 10208 119620 10260
rect 119672 10248 119678 10260
rect 122098 10248 122104 10260
rect 119672 10220 122104 10248
rect 119672 10208 119678 10220
rect 122098 10208 122104 10220
rect 122156 10208 122162 10260
rect 123110 10248 123116 10260
rect 123071 10220 123116 10248
rect 123110 10208 123116 10220
rect 123168 10208 123174 10260
rect 124950 10248 124956 10260
rect 124911 10220 124956 10248
rect 124950 10208 124956 10220
rect 125008 10208 125014 10260
rect 125781 10251 125839 10257
rect 125781 10217 125793 10251
rect 125827 10248 125839 10251
rect 125965 10251 126023 10257
rect 125965 10248 125977 10251
rect 125827 10220 125977 10248
rect 125827 10217 125839 10220
rect 125781 10211 125839 10217
rect 125965 10217 125977 10220
rect 126011 10248 126023 10251
rect 126606 10248 126612 10260
rect 126011 10220 126612 10248
rect 126011 10217 126023 10220
rect 125965 10211 126023 10217
rect 126606 10208 126612 10220
rect 126664 10208 126670 10260
rect 127342 10248 127348 10260
rect 127303 10220 127348 10248
rect 127342 10208 127348 10220
rect 127400 10208 127406 10260
rect 127434 10208 127440 10260
rect 127492 10248 127498 10260
rect 127897 10251 127955 10257
rect 127492 10220 127664 10248
rect 127492 10208 127498 10220
rect 106734 10140 106740 10192
rect 106792 10180 106798 10192
rect 124677 10183 124735 10189
rect 106792 10152 116164 10180
rect 106792 10140 106798 10152
rect 99653 10115 99711 10121
rect 99653 10081 99665 10115
rect 99699 10081 99711 10115
rect 100846 10112 100852 10124
rect 100807 10084 100852 10112
rect 99653 10075 99711 10081
rect 100846 10072 100852 10084
rect 100904 10072 100910 10124
rect 102226 10112 102232 10124
rect 102187 10084 102232 10112
rect 102226 10072 102232 10084
rect 102284 10112 102290 10124
rect 102689 10115 102747 10121
rect 102689 10112 102701 10115
rect 102284 10084 102701 10112
rect 102284 10072 102290 10084
rect 102689 10081 102701 10084
rect 102735 10081 102747 10115
rect 102689 10075 102747 10081
rect 107013 10115 107071 10121
rect 107013 10081 107025 10115
rect 107059 10112 107071 10115
rect 107654 10112 107660 10124
rect 107059 10084 107660 10112
rect 107059 10081 107071 10084
rect 107013 10075 107071 10081
rect 107654 10072 107660 10084
rect 107712 10072 107718 10124
rect 108117 10115 108175 10121
rect 108117 10081 108129 10115
rect 108163 10112 108175 10115
rect 110046 10112 110052 10124
rect 108163 10084 110052 10112
rect 108163 10081 108175 10084
rect 108117 10075 108175 10081
rect 110046 10072 110052 10084
rect 110104 10112 110110 10124
rect 110417 10115 110475 10121
rect 110417 10112 110429 10115
rect 110104 10084 110429 10112
rect 110104 10072 110110 10084
rect 110417 10081 110429 10084
rect 110463 10081 110475 10115
rect 110417 10075 110475 10081
rect 110969 10115 111027 10121
rect 110969 10081 110981 10115
rect 111015 10112 111027 10115
rect 111242 10112 111248 10124
rect 111015 10084 111248 10112
rect 111015 10081 111027 10084
rect 110969 10075 111027 10081
rect 111242 10072 111248 10084
rect 111300 10072 111306 10124
rect 112530 10112 112536 10124
rect 111352 10084 112536 10112
rect 97675 10016 98040 10044
rect 101217 10047 101275 10053
rect 97675 10013 97687 10016
rect 97629 10007 97687 10013
rect 101217 10013 101229 10047
rect 101263 10044 101275 10047
rect 101582 10044 101588 10056
rect 101263 10016 101588 10044
rect 101263 10013 101275 10016
rect 101217 10007 101275 10013
rect 101582 10004 101588 10016
rect 101640 10004 101646 10056
rect 101766 10004 101772 10056
rect 101824 10044 101830 10056
rect 111352 10044 111380 10084
rect 112530 10072 112536 10084
rect 112588 10072 112594 10124
rect 114281 10115 114339 10121
rect 114281 10081 114293 10115
rect 114327 10112 114339 10115
rect 115566 10112 115572 10124
rect 114327 10084 114968 10112
rect 115527 10084 115572 10112
rect 114327 10081 114339 10084
rect 114281 10075 114339 10081
rect 101824 10016 111380 10044
rect 101824 10004 101830 10016
rect 112254 10004 112260 10056
rect 112312 10044 112318 10056
rect 112898 10044 112904 10056
rect 112312 10016 112904 10044
rect 112312 10004 112318 10016
rect 112898 10004 112904 10016
rect 112956 10004 112962 10056
rect 114373 10047 114431 10053
rect 114373 10013 114385 10047
rect 114419 10013 114431 10047
rect 114373 10007 114431 10013
rect 109034 9936 109040 9988
rect 109092 9976 109098 9988
rect 109957 9979 110015 9985
rect 109957 9976 109969 9979
rect 109092 9948 109969 9976
rect 109092 9936 109098 9948
rect 109957 9945 109969 9948
rect 110003 9945 110015 9979
rect 109957 9939 110015 9945
rect 110046 9936 110052 9988
rect 110104 9976 110110 9988
rect 112809 9979 112867 9985
rect 112809 9976 112821 9979
rect 110104 9948 112821 9976
rect 110104 9936 110110 9948
rect 112809 9945 112821 9948
rect 112855 9945 112867 9979
rect 114388 9976 114416 10007
rect 114646 10004 114652 10056
rect 114704 10044 114710 10056
rect 114741 10047 114799 10053
rect 114741 10044 114753 10047
rect 114704 10016 114753 10044
rect 114704 10004 114710 10016
rect 114741 10013 114753 10016
rect 114787 10013 114799 10047
rect 114940 10044 114968 10084
rect 115566 10072 115572 10084
rect 115624 10072 115630 10124
rect 115934 10044 115940 10056
rect 114940 10016 115940 10044
rect 114741 10007 114799 10013
rect 115934 10004 115940 10016
rect 115992 10004 115998 10056
rect 116136 10044 116164 10152
rect 124677 10149 124689 10183
rect 124723 10180 124735 10183
rect 125321 10183 125379 10189
rect 125321 10180 125333 10183
rect 124723 10152 125333 10180
rect 124723 10149 124735 10152
rect 124677 10143 124735 10149
rect 125321 10149 125333 10152
rect 125367 10180 125379 10183
rect 127526 10180 127532 10192
rect 125367 10152 127532 10180
rect 125367 10149 125379 10152
rect 125321 10143 125379 10149
rect 127526 10140 127532 10152
rect 127584 10140 127590 10192
rect 127636 10180 127664 10220
rect 127897 10217 127909 10251
rect 127943 10248 127955 10251
rect 128354 10248 128360 10260
rect 127943 10220 128360 10248
rect 127943 10217 127955 10220
rect 127897 10211 127955 10217
rect 128354 10208 128360 10220
rect 128412 10208 128418 10260
rect 129550 10208 129556 10260
rect 129608 10248 129614 10260
rect 130289 10251 130347 10257
rect 130289 10248 130301 10251
rect 129608 10220 130301 10248
rect 129608 10208 129614 10220
rect 130289 10217 130301 10220
rect 130335 10248 130347 10251
rect 132954 10248 132960 10260
rect 130335 10220 132960 10248
rect 130335 10217 130347 10220
rect 130289 10211 130347 10217
rect 132954 10208 132960 10220
rect 133012 10208 133018 10260
rect 134058 10208 134064 10260
rect 134116 10248 134122 10260
rect 134245 10251 134303 10257
rect 134245 10248 134257 10251
rect 134116 10220 134257 10248
rect 134116 10208 134122 10220
rect 134245 10217 134257 10220
rect 134291 10217 134303 10251
rect 134245 10211 134303 10217
rect 135070 10208 135076 10260
rect 135128 10248 135134 10260
rect 135257 10251 135315 10257
rect 135257 10248 135269 10251
rect 135128 10220 135269 10248
rect 135128 10208 135134 10220
rect 135257 10217 135269 10220
rect 135303 10217 135315 10251
rect 137462 10248 137468 10260
rect 137423 10220 137468 10248
rect 135257 10211 135315 10217
rect 137462 10208 137468 10220
rect 137520 10208 137526 10260
rect 149057 10251 149115 10257
rect 137572 10220 139072 10248
rect 137572 10180 137600 10220
rect 127636 10152 137600 10180
rect 116578 10112 116584 10124
rect 116539 10084 116584 10112
rect 116578 10072 116584 10084
rect 116636 10072 116642 10124
rect 117593 10115 117651 10121
rect 117593 10081 117605 10115
rect 117639 10112 117651 10115
rect 117958 10112 117964 10124
rect 117639 10084 117964 10112
rect 117639 10081 117651 10084
rect 117593 10075 117651 10081
rect 117958 10072 117964 10084
rect 118016 10072 118022 10124
rect 122193 10115 122251 10121
rect 122193 10112 122205 10115
rect 118988 10084 122205 10112
rect 118988 10044 119016 10084
rect 122193 10081 122205 10084
rect 122239 10081 122251 10115
rect 126885 10115 126943 10121
rect 126885 10112 126897 10115
rect 122193 10075 122251 10081
rect 122300 10084 126897 10112
rect 116136 10016 119016 10044
rect 119065 10047 119123 10053
rect 119065 10013 119077 10047
rect 119111 10044 119123 10047
rect 119433 10047 119491 10053
rect 119433 10044 119445 10047
rect 119111 10016 119445 10044
rect 119111 10013 119123 10016
rect 119065 10007 119123 10013
rect 119433 10013 119445 10016
rect 119479 10013 119491 10047
rect 119433 10007 119491 10013
rect 120077 10047 120135 10053
rect 120077 10013 120089 10047
rect 120123 10044 120135 10047
rect 121178 10044 121184 10056
rect 120123 10016 121184 10044
rect 120123 10013 120135 10016
rect 120077 10007 120135 10013
rect 121178 10004 121184 10016
rect 121236 10004 121242 10056
rect 122098 10004 122104 10056
rect 122156 10044 122162 10056
rect 122300 10044 122328 10084
rect 126885 10081 126897 10084
rect 126931 10081 126943 10115
rect 128998 10112 129004 10124
rect 128959 10084 129004 10112
rect 126885 10075 126943 10081
rect 128998 10072 129004 10084
rect 129056 10072 129062 10124
rect 129734 10072 129740 10124
rect 129792 10112 129798 10124
rect 130473 10115 130531 10121
rect 130473 10112 130485 10115
rect 129792 10084 130485 10112
rect 129792 10072 129798 10084
rect 130473 10081 130485 10084
rect 130519 10081 130531 10115
rect 130473 10075 130531 10081
rect 130654 10072 130660 10124
rect 130712 10112 130718 10124
rect 131209 10115 131267 10121
rect 131209 10112 131221 10115
rect 130712 10084 131221 10112
rect 130712 10072 130718 10084
rect 131209 10081 131221 10084
rect 131255 10081 131267 10115
rect 132402 10112 132408 10124
rect 132363 10084 132408 10112
rect 131209 10075 131267 10081
rect 132402 10072 132408 10084
rect 132460 10072 132466 10124
rect 133414 10112 133420 10124
rect 133375 10084 133420 10112
rect 133414 10072 133420 10084
rect 133472 10072 133478 10124
rect 136266 10112 136272 10124
rect 136227 10084 136272 10112
rect 136266 10072 136272 10084
rect 136324 10112 136330 10124
rect 139044 10121 139072 10220
rect 149057 10217 149069 10251
rect 149103 10248 149115 10251
rect 151909 10251 151967 10257
rect 151909 10248 151921 10251
rect 149103 10220 151921 10248
rect 149103 10217 149115 10220
rect 149057 10211 149115 10217
rect 146205 10183 146263 10189
rect 146205 10149 146217 10183
rect 146251 10180 146263 10183
rect 147214 10180 147220 10192
rect 146251 10152 147220 10180
rect 146251 10149 146263 10152
rect 146205 10143 146263 10149
rect 147214 10140 147220 10152
rect 147272 10140 147278 10192
rect 136729 10115 136787 10121
rect 136729 10112 136741 10115
rect 136324 10084 136741 10112
rect 136324 10072 136330 10084
rect 136729 10081 136741 10084
rect 136775 10081 136787 10115
rect 136729 10075 136787 10081
rect 139029 10115 139087 10121
rect 139029 10081 139041 10115
rect 139075 10081 139087 10115
rect 139029 10075 139087 10081
rect 140774 10072 140780 10124
rect 140832 10112 140838 10124
rect 141421 10115 141479 10121
rect 141421 10112 141433 10115
rect 140832 10084 141433 10112
rect 140832 10072 140838 10084
rect 141421 10081 141433 10084
rect 141467 10081 141479 10115
rect 141421 10075 141479 10081
rect 142154 10072 142160 10124
rect 142212 10112 142218 10124
rect 142249 10115 142307 10121
rect 142249 10112 142261 10115
rect 142212 10084 142261 10112
rect 142212 10072 142218 10084
rect 142249 10081 142261 10084
rect 142295 10081 142307 10115
rect 142249 10075 142307 10081
rect 122742 10044 122748 10056
rect 122156 10016 122328 10044
rect 122703 10016 122748 10044
rect 122156 10004 122162 10016
rect 122742 10004 122748 10016
rect 122800 10004 122806 10056
rect 124401 10047 124459 10053
rect 124401 10013 124413 10047
rect 124447 10044 124459 10047
rect 124677 10047 124735 10053
rect 124677 10044 124689 10047
rect 124447 10016 124689 10044
rect 124447 10013 124459 10016
rect 124401 10007 124459 10013
rect 124677 10013 124689 10016
rect 124723 10013 124735 10047
rect 124677 10007 124735 10013
rect 125413 10047 125471 10053
rect 125413 10013 125425 10047
rect 125459 10044 125471 10047
rect 125781 10047 125839 10053
rect 125781 10044 125793 10047
rect 125459 10016 125793 10044
rect 125459 10013 125471 10016
rect 125413 10007 125471 10013
rect 125781 10013 125793 10016
rect 125827 10013 125839 10047
rect 125781 10007 125839 10013
rect 126793 10047 126851 10053
rect 126793 10013 126805 10047
rect 126839 10044 126851 10047
rect 127342 10044 127348 10056
rect 126839 10016 127348 10044
rect 126839 10013 126851 10016
rect 126793 10007 126851 10013
rect 127342 10004 127348 10016
rect 127400 10004 127406 10056
rect 127989 10047 128047 10053
rect 127989 10013 128001 10047
rect 128035 10044 128047 10047
rect 128078 10044 128084 10056
rect 128035 10016 128084 10044
rect 128035 10013 128047 10016
rect 127989 10007 128047 10013
rect 128078 10004 128084 10016
rect 128136 10004 128142 10056
rect 129553 10047 129611 10053
rect 129553 10013 129565 10047
rect 129599 10013 129611 10047
rect 129553 10007 129611 10013
rect 115201 9979 115259 9985
rect 115201 9976 115213 9979
rect 114388 9948 115213 9976
rect 112809 9939 112867 9945
rect 115201 9945 115213 9948
rect 115247 9976 115259 9979
rect 115247 9948 116164 9976
rect 115247 9945 115259 9948
rect 115201 9939 115259 9945
rect 87288 9880 87552 9908
rect 92753 9911 92811 9917
rect 87288 9868 87294 9880
rect 92753 9877 92765 9911
rect 92799 9908 92811 9911
rect 93118 9908 93124 9920
rect 92799 9880 93124 9908
rect 92799 9877 92811 9880
rect 92753 9871 92811 9877
rect 93118 9868 93124 9880
rect 93176 9868 93182 9920
rect 93394 9868 93400 9920
rect 93452 9908 93458 9920
rect 98362 9908 98368 9920
rect 93452 9880 98368 9908
rect 93452 9868 93458 9880
rect 98362 9868 98368 9880
rect 98420 9868 98426 9920
rect 98457 9911 98515 9917
rect 98457 9877 98469 9911
rect 98503 9908 98515 9911
rect 102134 9908 102140 9920
rect 98503 9880 102140 9908
rect 98503 9877 98515 9880
rect 98457 9871 98515 9877
rect 102134 9868 102140 9880
rect 102192 9868 102198 9920
rect 103241 9911 103299 9917
rect 103241 9877 103253 9911
rect 103287 9908 103299 9911
rect 103330 9908 103336 9920
rect 103287 9880 103336 9908
rect 103287 9877 103299 9880
rect 103241 9871 103299 9877
rect 103330 9868 103336 9880
rect 103388 9868 103394 9920
rect 103793 9911 103851 9917
rect 103793 9877 103805 9911
rect 103839 9908 103851 9911
rect 104250 9908 104256 9920
rect 103839 9880 104256 9908
rect 103839 9877 103851 9880
rect 103793 9871 103851 9877
rect 104250 9868 104256 9880
rect 104308 9868 104314 9920
rect 104618 9908 104624 9920
rect 104579 9880 104624 9908
rect 104618 9868 104624 9880
rect 104676 9868 104682 9920
rect 106001 9911 106059 9917
rect 106001 9877 106013 9911
rect 106047 9908 106059 9911
rect 106182 9908 106188 9920
rect 106047 9880 106188 9908
rect 106047 9877 106059 9880
rect 106001 9871 106059 9877
rect 106182 9868 106188 9880
rect 106240 9908 106246 9920
rect 114554 9908 114560 9920
rect 106240 9880 114560 9908
rect 106240 9868 106246 9880
rect 114554 9868 114560 9880
rect 114612 9868 114618 9920
rect 115842 9868 115848 9920
rect 115900 9908 115906 9920
rect 116029 9911 116087 9917
rect 116029 9908 116041 9911
rect 115900 9880 116041 9908
rect 115900 9868 115906 9880
rect 116029 9877 116041 9880
rect 116075 9877 116087 9911
rect 116136 9908 116164 9948
rect 120902 9936 120908 9988
rect 120960 9976 120966 9988
rect 125505 9979 125563 9985
rect 125505 9976 125517 9979
rect 120960 9948 125517 9976
rect 120960 9936 120966 9948
rect 125505 9945 125517 9948
rect 125551 9945 125563 9979
rect 129568 9976 129596 10007
rect 129918 10004 129924 10056
rect 129976 10044 129982 10056
rect 130381 10047 130439 10053
rect 130381 10044 130393 10047
rect 129976 10016 130393 10044
rect 129976 10004 129982 10016
rect 130381 10013 130393 10016
rect 130427 10044 130439 10047
rect 130841 10047 130899 10053
rect 130841 10044 130853 10047
rect 130427 10016 130853 10044
rect 130427 10013 130439 10016
rect 130381 10007 130439 10013
rect 130841 10013 130853 10016
rect 130887 10013 130899 10047
rect 133506 10044 133512 10056
rect 133467 10016 133512 10044
rect 130841 10007 130899 10013
rect 133506 10004 133512 10016
rect 133564 10004 133570 10056
rect 134794 10044 134800 10056
rect 134755 10016 134800 10044
rect 134794 10004 134800 10016
rect 134852 10044 134858 10056
rect 135625 10047 135683 10053
rect 135625 10044 135637 10047
rect 134852 10016 135637 10044
rect 134852 10004 134858 10016
rect 135625 10013 135637 10016
rect 135671 10013 135683 10047
rect 135625 10007 135683 10013
rect 138014 10004 138020 10056
rect 138072 10044 138078 10056
rect 139118 10044 139124 10056
rect 138072 10016 138117 10044
rect 139079 10016 139124 10044
rect 138072 10004 138078 10016
rect 139118 10004 139124 10016
rect 139176 10004 139182 10056
rect 140406 10044 140412 10056
rect 140367 10016 140412 10044
rect 140406 10004 140412 10016
rect 140464 10004 140470 10056
rect 140866 10004 140872 10056
rect 140924 10044 140930 10056
rect 149256 10053 149284 10220
rect 151909 10217 151921 10220
rect 151955 10217 151967 10251
rect 152090 10248 152096 10260
rect 152051 10220 152096 10248
rect 151909 10211 151967 10217
rect 152090 10208 152096 10220
rect 152148 10208 152154 10260
rect 153194 10208 153200 10260
rect 153252 10248 153258 10260
rect 153289 10251 153347 10257
rect 153289 10248 153301 10251
rect 153252 10220 153301 10248
rect 153252 10208 153258 10220
rect 153289 10217 153301 10220
rect 153335 10217 153347 10251
rect 155310 10248 155316 10260
rect 155271 10220 155316 10248
rect 153289 10211 153347 10217
rect 155310 10208 155316 10220
rect 155368 10208 155374 10260
rect 155954 10208 155960 10260
rect 156012 10248 156018 10260
rect 156325 10251 156383 10257
rect 156325 10248 156337 10251
rect 156012 10220 156337 10248
rect 156012 10208 156018 10220
rect 156325 10217 156337 10220
rect 156371 10217 156383 10251
rect 156325 10211 156383 10217
rect 157889 10251 157947 10257
rect 157889 10217 157901 10251
rect 157935 10248 157947 10251
rect 158714 10248 158720 10260
rect 157935 10220 158720 10248
rect 157935 10217 157947 10220
rect 157889 10211 157947 10217
rect 158714 10208 158720 10220
rect 158772 10208 158778 10260
rect 159542 10208 159548 10260
rect 159600 10248 159606 10260
rect 159821 10251 159879 10257
rect 159821 10248 159833 10251
rect 159600 10220 159833 10248
rect 159600 10208 159606 10220
rect 159821 10217 159833 10220
rect 159867 10217 159879 10251
rect 162670 10248 162676 10260
rect 162631 10220 162676 10248
rect 159821 10211 159879 10217
rect 162670 10208 162676 10220
rect 162728 10208 162734 10260
rect 164326 10208 164332 10260
rect 164384 10248 164390 10260
rect 165065 10251 165123 10257
rect 165065 10248 165077 10251
rect 164384 10220 165077 10248
rect 164384 10208 164390 10220
rect 165065 10217 165077 10220
rect 165111 10217 165123 10251
rect 165614 10248 165620 10260
rect 165575 10220 165620 10248
rect 165065 10211 165123 10217
rect 165614 10208 165620 10220
rect 165672 10208 165678 10260
rect 166718 10208 166724 10260
rect 166776 10248 166782 10260
rect 166905 10251 166963 10257
rect 166905 10248 166917 10251
rect 166776 10220 166917 10248
rect 166776 10208 166782 10220
rect 166905 10217 166917 10220
rect 166951 10217 166963 10251
rect 166905 10211 166963 10217
rect 150713 10183 150771 10189
rect 150713 10149 150725 10183
rect 150759 10180 150771 10183
rect 151262 10180 151268 10192
rect 150759 10152 151268 10180
rect 150759 10149 150771 10152
rect 150713 10143 150771 10149
rect 151262 10140 151268 10152
rect 151320 10140 151326 10192
rect 151633 10115 151691 10121
rect 151633 10081 151645 10115
rect 151679 10112 151691 10115
rect 152108 10112 152136 10208
rect 162302 10140 162308 10192
rect 162360 10180 162366 10192
rect 162360 10152 163912 10180
rect 162360 10140 162366 10152
rect 151679 10084 152136 10112
rect 156969 10115 157027 10121
rect 151679 10081 151691 10084
rect 151633 10075 151691 10081
rect 156969 10081 156981 10115
rect 157015 10112 157027 10115
rect 157978 10112 157984 10124
rect 157015 10084 157984 10112
rect 157015 10081 157027 10084
rect 156969 10075 157027 10081
rect 157978 10072 157984 10084
rect 158036 10072 158042 10124
rect 159358 10112 159364 10124
rect 159319 10084 159364 10112
rect 159358 10072 159364 10084
rect 159416 10072 159422 10124
rect 160462 10112 160468 10124
rect 160423 10084 160468 10112
rect 160462 10072 160468 10084
rect 160520 10072 160526 10124
rect 160554 10072 160560 10124
rect 160612 10112 160618 10124
rect 161477 10115 161535 10121
rect 161477 10112 161489 10115
rect 160612 10084 161489 10112
rect 160612 10072 160618 10084
rect 161477 10081 161489 10084
rect 161523 10081 161535 10115
rect 162854 10112 162860 10124
rect 162815 10084 162860 10112
rect 161477 10075 161535 10081
rect 162854 10072 162860 10084
rect 162912 10072 162918 10124
rect 163884 10121 163912 10152
rect 163869 10115 163927 10121
rect 163869 10081 163881 10115
rect 163915 10081 163927 10115
rect 165632 10112 165660 10208
rect 166077 10115 166135 10121
rect 166077 10112 166089 10115
rect 165632 10084 166089 10112
rect 163869 10075 163927 10081
rect 166077 10081 166089 10084
rect 166123 10081 166135 10115
rect 166077 10075 166135 10081
rect 141513 10047 141571 10053
rect 141513 10044 141525 10047
rect 140924 10016 141525 10044
rect 140924 10004 140930 10016
rect 141513 10013 141525 10016
rect 141559 10044 141571 10047
rect 142617 10047 142675 10053
rect 142617 10044 142629 10047
rect 141559 10016 142629 10044
rect 141559 10013 141571 10016
rect 141513 10007 141571 10013
rect 142617 10013 142629 10016
rect 142663 10013 142675 10047
rect 142617 10007 142675 10013
rect 144733 10047 144791 10053
rect 144733 10013 144745 10047
rect 144779 10013 144791 10047
rect 144733 10007 144791 10013
rect 146297 10047 146355 10053
rect 146297 10013 146309 10047
rect 146343 10013 146355 10047
rect 146297 10007 146355 10013
rect 149241 10047 149299 10053
rect 149241 10013 149253 10047
rect 149287 10013 149299 10047
rect 149241 10007 149299 10013
rect 150345 10047 150403 10053
rect 150345 10013 150357 10047
rect 150391 10013 150403 10047
rect 159542 10044 159548 10056
rect 159503 10016 159548 10044
rect 150345 10007 150403 10013
rect 134889 9979 134947 9985
rect 129568 9948 129964 9976
rect 125505 9939 125563 9945
rect 120718 9908 120724 9920
rect 116136 9880 120724 9908
rect 116029 9871 116087 9877
rect 120718 9868 120724 9880
rect 120776 9868 120782 9920
rect 120813 9911 120871 9917
rect 120813 9877 120825 9911
rect 120859 9908 120871 9911
rect 121086 9908 121092 9920
rect 120859 9880 121092 9908
rect 120859 9877 120871 9880
rect 120813 9871 120871 9877
rect 121086 9868 121092 9880
rect 121144 9908 121150 9920
rect 124493 9911 124551 9917
rect 124493 9908 124505 9911
rect 121144 9880 124505 9908
rect 121144 9868 121150 9880
rect 124493 9877 124505 9880
rect 124539 9877 124551 9911
rect 126238 9908 126244 9920
rect 126199 9880 126244 9908
rect 124493 9871 124551 9877
rect 126238 9868 126244 9880
rect 126296 9868 126302 9920
rect 129936 9917 129964 9948
rect 134889 9945 134901 9979
rect 134935 9976 134947 9979
rect 137830 9976 137836 9988
rect 134935 9948 137836 9976
rect 134935 9945 134947 9948
rect 134889 9939 134947 9945
rect 137830 9936 137836 9948
rect 137888 9936 137894 9988
rect 139026 9936 139032 9988
rect 139084 9976 139090 9988
rect 139857 9979 139915 9985
rect 139857 9976 139869 9979
rect 139084 9948 139869 9976
rect 139084 9936 139090 9948
rect 139857 9945 139869 9948
rect 139903 9945 139915 9979
rect 139857 9939 139915 9945
rect 141050 9936 141056 9988
rect 141108 9976 141114 9988
rect 143629 9979 143687 9985
rect 143629 9976 143641 9979
rect 141108 9948 143641 9976
rect 141108 9936 141114 9948
rect 143629 9945 143641 9948
rect 143675 9945 143687 9979
rect 143629 9939 143687 9945
rect 129921 9911 129979 9917
rect 129921 9877 129933 9911
rect 129967 9908 129979 9911
rect 130194 9908 130200 9920
rect 129967 9880 130200 9908
rect 129967 9877 129979 9880
rect 129921 9871 129979 9877
rect 130194 9868 130200 9880
rect 130252 9868 130258 9920
rect 144178 9908 144184 9920
rect 144139 9880 144184 9908
rect 144178 9868 144184 9880
rect 144236 9868 144242 9920
rect 144546 9908 144552 9920
rect 144507 9880 144552 9908
rect 144546 9868 144552 9880
rect 144604 9908 144610 9920
rect 144748 9908 144776 10007
rect 144604 9880 144776 9908
rect 146312 9908 146340 10007
rect 147769 9979 147827 9985
rect 147769 9945 147781 9979
rect 147815 9976 147827 9979
rect 147858 9976 147864 9988
rect 147815 9948 147864 9976
rect 147815 9945 147827 9948
rect 147769 9939 147827 9945
rect 147858 9936 147864 9948
rect 147916 9976 147922 9988
rect 148689 9979 148747 9985
rect 147916 9948 148456 9976
rect 147916 9936 147922 9948
rect 146662 9908 146668 9920
rect 146312 9880 146668 9908
rect 144604 9868 144610 9880
rect 146662 9868 146668 9880
rect 146720 9868 146726 9920
rect 146938 9908 146944 9920
rect 146899 9880 146944 9908
rect 146938 9868 146944 9880
rect 146996 9868 147002 9920
rect 147122 9908 147128 9920
rect 147083 9880 147128 9908
rect 147122 9868 147128 9880
rect 147180 9868 147186 9920
rect 148134 9908 148140 9920
rect 148095 9880 148140 9908
rect 148134 9868 148140 9880
rect 148192 9868 148198 9920
rect 148428 9908 148456 9948
rect 148689 9945 148701 9979
rect 148735 9976 148747 9979
rect 148778 9976 148784 9988
rect 148735 9948 148784 9976
rect 148735 9945 148747 9948
rect 148689 9939 148747 9945
rect 148778 9936 148784 9948
rect 148836 9936 148842 9988
rect 150360 9976 150388 10007
rect 159542 10004 159548 10016
rect 159600 10004 159606 10056
rect 161566 10044 161572 10056
rect 161527 10016 161572 10044
rect 161566 10004 161572 10016
rect 161624 10044 161630 10056
rect 162305 10047 162363 10053
rect 162305 10044 162317 10047
rect 161624 10016 162317 10044
rect 161624 10004 161630 10016
rect 162305 10013 162317 10016
rect 162351 10013 162363 10047
rect 163958 10044 163964 10056
rect 163919 10016 163964 10044
rect 162305 10007 162363 10013
rect 163958 10004 163964 10016
rect 164016 10044 164022 10056
rect 164697 10047 164755 10053
rect 164697 10044 164709 10047
rect 164016 10016 164709 10044
rect 164016 10004 164022 10016
rect 164697 10013 164709 10016
rect 164743 10013 164755 10047
rect 164697 10007 164755 10013
rect 151909 9979 151967 9985
rect 150360 9948 151124 9976
rect 151096 9920 151124 9948
rect 151909 9945 151921 9979
rect 151955 9976 151967 9979
rect 152645 9979 152703 9985
rect 152645 9976 152657 9979
rect 151955 9948 152657 9976
rect 151955 9945 151967 9948
rect 151909 9939 151967 9945
rect 152645 9945 152657 9948
rect 152691 9945 152703 9979
rect 152645 9939 152703 9945
rect 149974 9908 149980 9920
rect 148428 9880 149980 9908
rect 149974 9868 149980 9880
rect 150032 9868 150038 9920
rect 151078 9908 151084 9920
rect 151039 9880 151084 9908
rect 151078 9868 151084 9880
rect 151136 9868 151142 9920
rect 151541 9911 151599 9917
rect 151541 9877 151553 9911
rect 151587 9908 151599 9911
rect 151630 9908 151636 9920
rect 151587 9880 151636 9908
rect 151587 9877 151599 9880
rect 151541 9871 151599 9877
rect 151630 9868 151636 9880
rect 151688 9868 151694 9920
rect 153194 9868 153200 9920
rect 153252 9908 153258 9920
rect 153657 9911 153715 9917
rect 153657 9908 153669 9911
rect 153252 9880 153669 9908
rect 153252 9868 153258 9880
rect 153657 9877 153669 9880
rect 153703 9877 153715 9911
rect 154850 9908 154856 9920
rect 154811 9880 154856 9908
rect 153657 9871 153715 9877
rect 154850 9868 154856 9880
rect 154908 9868 154914 9920
rect 154942 9868 154948 9920
rect 155000 9908 155006 9920
rect 155865 9911 155923 9917
rect 155865 9908 155877 9911
rect 155000 9880 155877 9908
rect 155000 9868 155006 9880
rect 155865 9877 155877 9880
rect 155911 9877 155923 9911
rect 155865 9871 155923 9877
rect 368 9818 169556 9840
rect 368 9766 56667 9818
rect 56719 9766 56731 9818
rect 56783 9766 56795 9818
rect 56847 9766 56859 9818
rect 56911 9766 113088 9818
rect 113140 9766 113152 9818
rect 113204 9766 113216 9818
rect 113268 9766 113280 9818
rect 113332 9766 169556 9818
rect 368 9744 169556 9766
rect 7098 9704 7104 9716
rect 7059 9676 7104 9704
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 24210 9704 24216 9716
rect 8076 9676 24216 9704
rect 8076 9664 8082 9676
rect 24210 9664 24216 9676
rect 24268 9664 24274 9716
rect 25130 9664 25136 9716
rect 25188 9704 25194 9716
rect 26786 9704 26792 9716
rect 25188 9676 26792 9704
rect 25188 9664 25194 9676
rect 26786 9664 26792 9676
rect 26844 9664 26850 9716
rect 27614 9704 27620 9716
rect 27575 9676 27620 9704
rect 27614 9664 27620 9676
rect 27672 9664 27678 9716
rect 27798 9664 27804 9716
rect 27856 9704 27862 9716
rect 28537 9707 28595 9713
rect 28537 9704 28549 9707
rect 27856 9676 28549 9704
rect 27856 9664 27862 9676
rect 28537 9673 28549 9676
rect 28583 9673 28595 9707
rect 28537 9667 28595 9673
rect 28810 9664 28816 9716
rect 28868 9704 28874 9716
rect 31386 9704 31392 9716
rect 28868 9676 31392 9704
rect 28868 9664 28874 9676
rect 31386 9664 31392 9676
rect 31444 9664 31450 9716
rect 32309 9707 32367 9713
rect 31588 9676 31892 9704
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 6086 9636 6092 9648
rect 3016 9608 5948 9636
rect 6047 9608 6092 9636
rect 3016 9596 3022 9608
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 4522 9568 4528 9580
rect 3384 9540 4528 9568
rect 3384 9528 3390 9540
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 5920 9568 5948 9608
rect 6086 9596 6092 9608
rect 6144 9596 6150 9648
rect 15286 9636 15292 9648
rect 15247 9608 15292 9636
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 15620 9608 20760 9636
rect 15620 9596 15626 9608
rect 7006 9568 7012 9580
rect 5920 9540 7012 9568
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 14366 9528 14372 9580
rect 14424 9568 14430 9580
rect 18785 9571 18843 9577
rect 14424 9540 18736 9568
rect 14424 9528 14430 9540
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3936 9472 3985 9500
rect 3936 9460 3942 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 5960 9472 8800 9500
rect 5960 9460 5966 9472
rect 2590 9392 2596 9444
rect 2648 9432 2654 9444
rect 6914 9432 6920 9444
rect 2648 9404 6920 9432
rect 2648 9392 2654 9404
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 1118 9324 1124 9376
rect 1176 9364 1182 9376
rect 4062 9364 4068 9376
rect 1176 9336 4068 9364
rect 1176 9324 1182 9336
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4706 9364 4712 9376
rect 4571 9336 4712 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6420 9336 6561 9364
rect 6420 9324 6426 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 8772 9364 8800 9472
rect 10318 9460 10324 9512
rect 10376 9500 10382 9512
rect 15565 9503 15623 9509
rect 10376 9472 15516 9500
rect 10376 9460 10382 9472
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 15488 9432 15516 9472
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 17494 9500 17500 9512
rect 15611 9472 17500 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 17773 9503 17831 9509
rect 17773 9469 17785 9503
rect 17819 9500 17831 9503
rect 18598 9500 18604 9512
rect 17819 9472 18604 9500
rect 17819 9469 17831 9472
rect 17773 9463 17831 9469
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 18708 9500 18736 9540
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 19797 9571 19855 9577
rect 19797 9568 19809 9571
rect 18831 9540 19809 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 19797 9537 19809 9540
rect 19843 9568 19855 9571
rect 19886 9568 19892 9580
rect 19843 9540 19892 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 20530 9568 20536 9580
rect 20491 9540 20536 9568
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 20732 9568 20760 9608
rect 20806 9596 20812 9648
rect 20864 9636 20870 9648
rect 21361 9639 21419 9645
rect 21361 9636 21373 9639
rect 20864 9608 21373 9636
rect 20864 9596 20870 9608
rect 21361 9605 21373 9608
rect 21407 9605 21419 9639
rect 21361 9599 21419 9605
rect 21450 9596 21456 9648
rect 21508 9636 21514 9648
rect 22738 9636 22744 9648
rect 21508 9608 22744 9636
rect 21508 9596 21514 9608
rect 22738 9596 22744 9608
rect 22796 9596 22802 9648
rect 31588 9636 31616 9676
rect 24688 9608 31616 9636
rect 31864 9636 31892 9676
rect 32309 9673 32321 9707
rect 32355 9704 32367 9707
rect 32582 9704 32588 9716
rect 32355 9676 32588 9704
rect 32355 9673 32367 9676
rect 32309 9667 32367 9673
rect 32582 9664 32588 9676
rect 32640 9664 32646 9716
rect 33410 9664 33416 9716
rect 33468 9704 33474 9716
rect 41782 9704 41788 9716
rect 33468 9676 41788 9704
rect 33468 9664 33474 9676
rect 41782 9664 41788 9676
rect 41840 9664 41846 9716
rect 41966 9664 41972 9716
rect 42024 9704 42030 9716
rect 46750 9704 46756 9716
rect 42024 9676 46756 9704
rect 42024 9664 42030 9676
rect 46750 9664 46756 9676
rect 46808 9664 46814 9716
rect 48314 9664 48320 9716
rect 48372 9704 48378 9716
rect 49789 9707 49847 9713
rect 48372 9676 48636 9704
rect 48372 9664 48378 9676
rect 33318 9636 33324 9648
rect 31864 9608 33324 9636
rect 24688 9568 24716 9608
rect 33318 9596 33324 9608
rect 33376 9596 33382 9648
rect 33502 9596 33508 9648
rect 33560 9636 33566 9648
rect 34422 9636 34428 9648
rect 33560 9608 34428 9636
rect 33560 9596 33566 9608
rect 34422 9596 34428 9608
rect 34480 9596 34486 9648
rect 34606 9596 34612 9648
rect 34664 9636 34670 9648
rect 34701 9639 34759 9645
rect 34701 9636 34713 9639
rect 34664 9608 34713 9636
rect 34664 9596 34670 9608
rect 34701 9605 34713 9608
rect 34747 9605 34759 9639
rect 35618 9636 35624 9648
rect 34701 9599 34759 9605
rect 34900 9608 35624 9636
rect 24854 9568 24860 9580
rect 20732 9540 24716 9568
rect 24815 9540 24860 9568
rect 24854 9528 24860 9540
rect 24912 9528 24918 9580
rect 24949 9571 25007 9577
rect 24949 9537 24961 9571
rect 24995 9568 25007 9571
rect 25130 9568 25136 9580
rect 24995 9540 25136 9568
rect 24995 9537 25007 9540
rect 24949 9531 25007 9537
rect 25130 9528 25136 9540
rect 25188 9528 25194 9580
rect 25314 9568 25320 9580
rect 25275 9540 25320 9568
rect 25314 9528 25320 9540
rect 25372 9528 25378 9580
rect 26421 9571 26479 9577
rect 26421 9537 26433 9571
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 26881 9571 26939 9577
rect 26881 9537 26893 9571
rect 26927 9568 26939 9571
rect 26970 9568 26976 9580
rect 26927 9540 26976 9568
rect 26927 9537 26939 9540
rect 26881 9531 26939 9537
rect 20622 9500 20628 9512
rect 18708 9472 20628 9500
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 20809 9503 20867 9509
rect 20809 9500 20821 9503
rect 20772 9472 20821 9500
rect 20772 9460 20778 9472
rect 20809 9469 20821 9472
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 21358 9460 21364 9512
rect 21416 9500 21422 9512
rect 21818 9500 21824 9512
rect 21416 9472 21824 9500
rect 21416 9460 21422 9472
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23106 9500 23112 9512
rect 22971 9472 23112 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23106 9460 23112 9472
rect 23164 9460 23170 9512
rect 23198 9460 23204 9512
rect 23256 9500 23262 9512
rect 26326 9500 26332 9512
rect 23256 9472 26332 9500
rect 23256 9460 23262 9472
rect 26326 9460 26332 9472
rect 26384 9460 26390 9512
rect 26436 9500 26464 9531
rect 26970 9528 26976 9540
rect 27028 9528 27034 9580
rect 27249 9571 27307 9577
rect 27249 9537 27261 9571
rect 27295 9568 27307 9571
rect 27338 9568 27344 9580
rect 27295 9540 27344 9568
rect 27295 9537 27307 9540
rect 27249 9531 27307 9537
rect 27264 9500 27292 9531
rect 27338 9528 27344 9540
rect 27396 9528 27402 9580
rect 27430 9528 27436 9580
rect 27488 9568 27494 9580
rect 30190 9568 30196 9580
rect 27488 9540 30196 9568
rect 27488 9528 27494 9540
rect 30190 9528 30196 9540
rect 30248 9528 30254 9580
rect 30282 9528 30288 9580
rect 30340 9568 30346 9580
rect 30745 9571 30803 9577
rect 30745 9568 30757 9571
rect 30340 9540 30757 9568
rect 30340 9528 30346 9540
rect 30745 9537 30757 9540
rect 30791 9537 30803 9571
rect 31478 9568 31484 9580
rect 31439 9540 31484 9568
rect 30745 9531 30803 9537
rect 31478 9528 31484 9540
rect 31536 9528 31542 9580
rect 31938 9528 31944 9580
rect 31996 9568 32002 9580
rect 34900 9568 34928 9608
rect 35618 9596 35624 9608
rect 35676 9596 35682 9648
rect 35710 9596 35716 9648
rect 35768 9636 35774 9648
rect 37921 9639 37979 9645
rect 37921 9636 37933 9639
rect 35768 9608 37933 9636
rect 35768 9596 35774 9608
rect 37921 9605 37933 9608
rect 37967 9605 37979 9639
rect 37921 9599 37979 9605
rect 39114 9596 39120 9648
rect 39172 9636 39178 9648
rect 41233 9639 41291 9645
rect 39172 9608 41184 9636
rect 39172 9596 39178 9608
rect 31996 9540 34928 9568
rect 31996 9528 32002 9540
rect 34974 9528 34980 9580
rect 35032 9568 35038 9580
rect 36357 9571 36415 9577
rect 36357 9568 36369 9571
rect 35032 9540 36369 9568
rect 35032 9528 35038 9540
rect 36357 9537 36369 9540
rect 36403 9537 36415 9571
rect 36814 9568 36820 9580
rect 36775 9540 36820 9568
rect 36357 9531 36415 9537
rect 36814 9528 36820 9540
rect 36872 9528 36878 9580
rect 36906 9528 36912 9580
rect 36964 9568 36970 9580
rect 38470 9568 38476 9580
rect 36964 9540 38476 9568
rect 36964 9528 36970 9540
rect 38470 9528 38476 9540
rect 38528 9528 38534 9580
rect 38565 9571 38623 9577
rect 38565 9537 38577 9571
rect 38611 9568 38623 9571
rect 39206 9568 39212 9580
rect 38611 9540 39212 9568
rect 38611 9537 38623 9540
rect 38565 9531 38623 9537
rect 39206 9528 39212 9540
rect 39264 9528 39270 9580
rect 39298 9528 39304 9580
rect 39356 9568 39362 9580
rect 40218 9568 40224 9580
rect 39356 9540 40224 9568
rect 39356 9528 39362 9540
rect 40218 9528 40224 9540
rect 40276 9528 40282 9580
rect 40405 9571 40463 9577
rect 40405 9537 40417 9571
rect 40451 9568 40463 9571
rect 40865 9571 40923 9577
rect 40451 9540 40816 9568
rect 40451 9537 40463 9540
rect 40405 9531 40463 9537
rect 34606 9500 34612 9512
rect 26436 9472 27292 9500
rect 27356 9472 34612 9500
rect 22830 9432 22836 9444
rect 8904 9404 15424 9432
rect 15488 9404 22836 9432
rect 8904 9392 8910 9404
rect 15194 9364 15200 9376
rect 8772 9336 15200 9364
rect 6549 9327 6607 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 15396 9364 15424 9404
rect 22830 9392 22836 9404
rect 22888 9392 22894 9444
rect 27356 9432 27384 9472
rect 34606 9460 34612 9472
rect 34664 9460 34670 9512
rect 35526 9460 35532 9512
rect 35584 9500 35590 9512
rect 40586 9500 40592 9512
rect 35584 9472 40592 9500
rect 35584 9460 35590 9472
rect 40586 9460 40592 9472
rect 40644 9460 40650 9512
rect 40788 9500 40816 9540
rect 40865 9537 40877 9571
rect 40911 9568 40923 9571
rect 41046 9568 41052 9580
rect 40911 9540 41052 9568
rect 40911 9537 40923 9540
rect 40865 9531 40923 9537
rect 41046 9528 41052 9540
rect 41104 9528 41110 9580
rect 41156 9568 41184 9608
rect 41233 9605 41245 9639
rect 41279 9636 41291 9639
rect 41322 9636 41328 9648
rect 41279 9608 41328 9636
rect 41279 9605 41291 9608
rect 41233 9599 41291 9605
rect 41322 9596 41328 9608
rect 41380 9636 41386 9648
rect 42610 9636 42616 9648
rect 41380 9608 42616 9636
rect 41380 9596 41386 9608
rect 42610 9596 42616 9608
rect 42668 9596 42674 9648
rect 42978 9596 42984 9648
rect 43036 9636 43042 9648
rect 43898 9636 43904 9648
rect 43036 9608 43904 9636
rect 43036 9596 43042 9608
rect 43898 9596 43904 9608
rect 43956 9596 43962 9648
rect 48041 9639 48099 9645
rect 44008 9608 46704 9636
rect 41874 9568 41880 9580
rect 41156 9540 41736 9568
rect 41835 9540 41880 9568
rect 41322 9500 41328 9512
rect 40788 9472 41328 9500
rect 41322 9460 41328 9472
rect 41380 9460 41386 9512
rect 22940 9404 27384 9432
rect 19242 9364 19248 9376
rect 15396 9336 19248 9364
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 19889 9367 19947 9373
rect 19889 9364 19901 9367
rect 19392 9336 19901 9364
rect 19392 9324 19398 9336
rect 19889 9333 19901 9336
rect 19935 9333 19947 9367
rect 19889 9327 19947 9333
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 21140 9336 21833 9364
rect 21140 9324 21146 9336
rect 21821 9333 21833 9336
rect 21867 9364 21879 9367
rect 21910 9364 21916 9376
rect 21867 9336 21916 9364
rect 21867 9333 21879 9336
rect 21821 9327 21879 9333
rect 21910 9324 21916 9336
rect 21968 9324 21974 9376
rect 22002 9324 22008 9376
rect 22060 9364 22066 9376
rect 22940 9364 22968 9404
rect 27430 9392 27436 9444
rect 27488 9432 27494 9444
rect 29822 9432 29828 9444
rect 27488 9404 29828 9432
rect 27488 9392 27494 9404
rect 29822 9392 29828 9404
rect 29880 9392 29886 9444
rect 31938 9432 31944 9444
rect 29932 9404 31944 9432
rect 22060 9336 22968 9364
rect 22060 9324 22066 9336
rect 23014 9324 23020 9376
rect 23072 9364 23078 9376
rect 25866 9364 25872 9376
rect 23072 9336 25872 9364
rect 23072 9324 23078 9336
rect 25866 9324 25872 9336
rect 25924 9324 25930 9376
rect 26050 9364 26056 9376
rect 26011 9336 26056 9364
rect 26050 9324 26056 9336
rect 26108 9324 26114 9376
rect 26237 9367 26295 9373
rect 26237 9333 26249 9367
rect 26283 9364 26295 9367
rect 26326 9364 26332 9376
rect 26283 9336 26332 9364
rect 26283 9333 26295 9336
rect 26237 9327 26295 9333
rect 26326 9324 26332 9336
rect 26384 9324 26390 9376
rect 26418 9324 26424 9376
rect 26476 9364 26482 9376
rect 29270 9364 29276 9376
rect 26476 9336 29276 9364
rect 26476 9324 26482 9336
rect 29270 9324 29276 9336
rect 29328 9324 29334 9376
rect 29362 9324 29368 9376
rect 29420 9364 29426 9376
rect 29932 9364 29960 9404
rect 31938 9392 31944 9404
rect 31996 9392 32002 9444
rect 41708 9432 41736 9540
rect 41874 9528 41880 9540
rect 41932 9528 41938 9580
rect 41966 9528 41972 9580
rect 42024 9568 42030 9580
rect 42061 9571 42119 9577
rect 42061 9568 42073 9571
rect 42024 9540 42073 9568
rect 42024 9528 42030 9540
rect 42061 9537 42073 9540
rect 42107 9537 42119 9571
rect 42426 9568 42432 9580
rect 42339 9540 42432 9568
rect 42061 9531 42119 9537
rect 42426 9528 42432 9540
rect 42484 9568 42490 9580
rect 44008 9568 44036 9608
rect 46566 9568 46572 9580
rect 42484 9540 44036 9568
rect 46527 9540 46572 9568
rect 42484 9528 42490 9540
rect 46566 9528 46572 9540
rect 46624 9528 46630 9580
rect 46676 9568 46704 9608
rect 48041 9605 48053 9639
rect 48087 9636 48099 9639
rect 48406 9636 48412 9648
rect 48087 9608 48412 9636
rect 48087 9605 48099 9608
rect 48041 9599 48099 9605
rect 48406 9596 48412 9608
rect 48464 9636 48470 9648
rect 48501 9639 48559 9645
rect 48501 9636 48513 9639
rect 48464 9608 48513 9636
rect 48464 9596 48470 9608
rect 48501 9605 48513 9608
rect 48547 9605 48559 9639
rect 48608 9636 48636 9676
rect 49789 9673 49801 9707
rect 49835 9704 49847 9707
rect 49970 9704 49976 9716
rect 49835 9676 49976 9704
rect 49835 9673 49847 9676
rect 49789 9667 49847 9673
rect 49970 9664 49976 9676
rect 50028 9664 50034 9716
rect 50246 9664 50252 9716
rect 50304 9704 50310 9716
rect 51350 9704 51356 9716
rect 50304 9676 51356 9704
rect 50304 9664 50310 9676
rect 51350 9664 51356 9676
rect 51408 9664 51414 9716
rect 51460 9676 57836 9704
rect 50154 9636 50160 9648
rect 48608 9608 50160 9636
rect 48501 9599 48559 9605
rect 50154 9596 50160 9608
rect 50212 9596 50218 9648
rect 51166 9596 51172 9648
rect 51224 9636 51230 9648
rect 51460 9636 51488 9676
rect 52086 9636 52092 9648
rect 51224 9608 51488 9636
rect 51736 9608 52092 9636
rect 51224 9596 51230 9608
rect 47118 9568 47124 9580
rect 46676 9540 46980 9568
rect 47031 9540 47124 9568
rect 41782 9460 41788 9512
rect 41840 9500 41846 9512
rect 46290 9500 46296 9512
rect 41840 9472 46296 9500
rect 41840 9460 41846 9472
rect 46290 9460 46296 9472
rect 46348 9460 46354 9512
rect 46952 9500 46980 9540
rect 47118 9528 47124 9540
rect 47176 9568 47182 9580
rect 50522 9568 50528 9580
rect 47176 9540 50528 9568
rect 47176 9528 47182 9540
rect 50522 9528 50528 9540
rect 50580 9528 50586 9580
rect 51074 9528 51080 9580
rect 51132 9568 51138 9580
rect 51132 9540 51177 9568
rect 51132 9528 51138 9540
rect 51258 9528 51264 9580
rect 51316 9528 51322 9580
rect 51736 9577 51764 9608
rect 52086 9596 52092 9608
rect 52144 9596 52150 9648
rect 52178 9596 52184 9648
rect 52236 9636 52242 9648
rect 54662 9636 54668 9648
rect 52236 9608 54340 9636
rect 54623 9608 54668 9636
rect 52236 9596 52242 9608
rect 51721 9571 51779 9577
rect 51721 9537 51733 9571
rect 51767 9537 51779 9571
rect 51721 9531 51779 9537
rect 53190 9528 53196 9580
rect 53248 9568 53254 9580
rect 53285 9571 53343 9577
rect 53285 9568 53297 9571
rect 53248 9540 53297 9568
rect 53248 9528 53254 9540
rect 53285 9537 53297 9540
rect 53331 9537 53343 9571
rect 53834 9568 53840 9580
rect 53285 9531 53343 9537
rect 53392 9540 53840 9568
rect 49510 9500 49516 9512
rect 46952 9472 49516 9500
rect 49510 9460 49516 9472
rect 49568 9460 49574 9512
rect 50614 9460 50620 9512
rect 50672 9500 50678 9512
rect 51276 9500 51304 9528
rect 50672 9472 51304 9500
rect 50672 9460 50678 9472
rect 51626 9460 51632 9512
rect 51684 9500 51690 9512
rect 53392 9500 53420 9540
rect 53834 9528 53840 9540
rect 53892 9528 53898 9580
rect 54021 9571 54079 9577
rect 54021 9537 54033 9571
rect 54067 9568 54079 9571
rect 54113 9571 54171 9577
rect 54113 9568 54125 9571
rect 54067 9540 54125 9568
rect 54067 9537 54079 9540
rect 54021 9531 54079 9537
rect 54113 9537 54125 9540
rect 54159 9537 54171 9571
rect 54312 9568 54340 9608
rect 54662 9596 54668 9608
rect 54720 9596 54726 9648
rect 54846 9596 54852 9648
rect 54904 9636 54910 9648
rect 55674 9636 55680 9648
rect 54904 9608 55680 9636
rect 54904 9596 54910 9608
rect 55674 9596 55680 9608
rect 55732 9596 55738 9648
rect 56134 9596 56140 9648
rect 56192 9636 56198 9648
rect 57241 9639 57299 9645
rect 56192 9608 56916 9636
rect 56192 9596 56198 9608
rect 54938 9568 54944 9580
rect 54312 9540 54944 9568
rect 54113 9531 54171 9537
rect 54938 9528 54944 9540
rect 54996 9528 55002 9580
rect 55122 9568 55128 9580
rect 55083 9540 55128 9568
rect 55122 9528 55128 9540
rect 55180 9528 55186 9580
rect 55493 9571 55551 9577
rect 55493 9537 55505 9571
rect 55539 9568 55551 9571
rect 55858 9568 55864 9580
rect 55539 9540 55864 9568
rect 55539 9537 55551 9540
rect 55493 9531 55551 9537
rect 55858 9528 55864 9540
rect 55916 9568 55922 9580
rect 56778 9568 56784 9580
rect 55916 9540 56784 9568
rect 55916 9528 55922 9540
rect 56778 9528 56784 9540
rect 56836 9528 56842 9580
rect 51684 9472 53420 9500
rect 51684 9460 51690 9472
rect 53466 9460 53472 9512
rect 53524 9500 53530 9512
rect 55582 9500 55588 9512
rect 53524 9472 55588 9500
rect 53524 9460 53530 9472
rect 55582 9460 55588 9472
rect 55640 9460 55646 9512
rect 56888 9500 56916 9608
rect 57241 9605 57253 9639
rect 57287 9636 57299 9639
rect 57698 9636 57704 9648
rect 57287 9608 57704 9636
rect 57287 9605 57299 9608
rect 57241 9599 57299 9605
rect 57698 9596 57704 9608
rect 57756 9596 57762 9648
rect 57808 9636 57836 9676
rect 57882 9664 57888 9716
rect 57940 9704 57946 9716
rect 57940 9676 59216 9704
rect 57940 9664 57946 9676
rect 59078 9636 59084 9648
rect 57808 9608 59084 9636
rect 59078 9596 59084 9608
rect 59136 9596 59142 9648
rect 59188 9636 59216 9676
rect 59354 9664 59360 9716
rect 59412 9704 59418 9716
rect 60550 9704 60556 9716
rect 59412 9676 60556 9704
rect 59412 9664 59418 9676
rect 60550 9664 60556 9676
rect 60608 9664 60614 9716
rect 60734 9664 60740 9716
rect 60792 9704 60798 9716
rect 62022 9704 62028 9716
rect 60792 9676 62028 9704
rect 60792 9664 60798 9676
rect 62022 9664 62028 9676
rect 62080 9664 62086 9716
rect 64230 9704 64236 9716
rect 64191 9676 64236 9704
rect 64230 9664 64236 9676
rect 64288 9664 64294 9716
rect 71682 9664 71688 9716
rect 71740 9704 71746 9716
rect 78490 9704 78496 9716
rect 71740 9676 78496 9704
rect 71740 9664 71746 9676
rect 78490 9664 78496 9676
rect 78548 9664 78554 9716
rect 85114 9704 85120 9716
rect 85075 9676 85120 9704
rect 85114 9664 85120 9676
rect 85172 9664 85178 9716
rect 86954 9664 86960 9716
rect 87012 9704 87018 9716
rect 93302 9704 93308 9716
rect 87012 9676 93164 9704
rect 93263 9676 93308 9704
rect 87012 9664 87018 9676
rect 60645 9639 60703 9645
rect 60645 9636 60657 9639
rect 59188 9608 60657 9636
rect 60645 9605 60657 9608
rect 60691 9605 60703 9639
rect 60645 9599 60703 9605
rect 61654 9596 61660 9648
rect 61712 9636 61718 9648
rect 63221 9639 63279 9645
rect 63221 9636 63233 9639
rect 61712 9608 63233 9636
rect 61712 9596 61718 9608
rect 63221 9605 63233 9608
rect 63267 9605 63279 9639
rect 63221 9599 63279 9605
rect 63494 9596 63500 9648
rect 63552 9636 63558 9648
rect 68830 9636 68836 9648
rect 63552 9608 68836 9636
rect 63552 9596 63558 9608
rect 68830 9596 68836 9608
rect 68888 9596 68894 9648
rect 70213 9639 70271 9645
rect 70213 9605 70225 9639
rect 70259 9636 70271 9639
rect 70854 9636 70860 9648
rect 70259 9608 70860 9636
rect 70259 9605 70271 9608
rect 70213 9599 70271 9605
rect 70854 9596 70860 9608
rect 70912 9596 70918 9648
rect 71225 9639 71283 9645
rect 71225 9605 71237 9639
rect 71271 9636 71283 9639
rect 71774 9636 71780 9648
rect 71271 9608 71780 9636
rect 71271 9605 71283 9608
rect 71225 9599 71283 9605
rect 71774 9596 71780 9608
rect 71832 9596 71838 9648
rect 72329 9639 72387 9645
rect 72329 9605 72341 9639
rect 72375 9636 72387 9639
rect 72786 9636 72792 9648
rect 72375 9608 72792 9636
rect 72375 9605 72387 9608
rect 72329 9599 72387 9605
rect 72786 9596 72792 9608
rect 72844 9596 72850 9648
rect 73982 9596 73988 9648
rect 74040 9636 74046 9648
rect 74442 9636 74448 9648
rect 74040 9608 74448 9636
rect 74040 9596 74046 9608
rect 74442 9596 74448 9608
rect 74500 9636 74506 9648
rect 79689 9639 79747 9645
rect 74500 9608 74764 9636
rect 74500 9596 74506 9608
rect 57793 9571 57851 9577
rect 57793 9537 57805 9571
rect 57839 9568 57851 9571
rect 57882 9568 57888 9580
rect 57839 9540 57888 9568
rect 57839 9537 57851 9540
rect 57793 9531 57851 9537
rect 57882 9528 57888 9540
rect 57940 9528 57946 9580
rect 58253 9571 58311 9577
rect 58253 9537 58265 9571
rect 58299 9568 58311 9571
rect 58621 9571 58679 9577
rect 58621 9568 58633 9571
rect 58299 9540 58633 9568
rect 58299 9537 58311 9540
rect 58253 9531 58311 9537
rect 58621 9537 58633 9540
rect 58667 9568 58679 9571
rect 58802 9568 58808 9580
rect 58667 9540 58808 9568
rect 58667 9537 58679 9540
rect 58621 9531 58679 9537
rect 58802 9528 58808 9540
rect 58860 9528 58866 9580
rect 59354 9568 59360 9580
rect 59315 9540 59360 9568
rect 59354 9528 59360 9540
rect 59412 9528 59418 9580
rect 59817 9571 59875 9577
rect 59817 9537 59829 9571
rect 59863 9568 59875 9571
rect 59906 9568 59912 9580
rect 59863 9540 59912 9568
rect 59863 9537 59875 9540
rect 59817 9531 59875 9537
rect 59906 9528 59912 9540
rect 59964 9568 59970 9580
rect 59964 9540 60688 9568
rect 59964 9528 59970 9540
rect 57974 9500 57980 9512
rect 56888 9472 57980 9500
rect 57974 9460 57980 9472
rect 58032 9460 58038 9512
rect 47302 9432 47308 9444
rect 34348 9404 41644 9432
rect 41708 9404 47308 9432
rect 30834 9364 30840 9376
rect 29420 9336 29960 9364
rect 30795 9336 30840 9364
rect 29420 9324 29426 9336
rect 30834 9324 30840 9336
rect 30892 9324 30898 9376
rect 31478 9324 31484 9376
rect 31536 9364 31542 9376
rect 31662 9364 31668 9376
rect 31536 9336 31668 9364
rect 31536 9324 31542 9336
rect 31662 9324 31668 9336
rect 31720 9364 31726 9376
rect 34348 9364 34376 9404
rect 31720 9336 34376 9364
rect 31720 9324 31726 9336
rect 34422 9324 34428 9376
rect 34480 9364 34486 9376
rect 37918 9364 37924 9376
rect 34480 9336 37924 9364
rect 34480 9324 34486 9336
rect 37918 9324 37924 9336
rect 37976 9324 37982 9376
rect 39022 9364 39028 9376
rect 38983 9336 39028 9364
rect 39022 9324 39028 9336
rect 39080 9324 39086 9376
rect 40218 9364 40224 9376
rect 40179 9336 40224 9364
rect 40218 9324 40224 9336
rect 40276 9324 40282 9376
rect 40310 9324 40316 9376
rect 40368 9364 40374 9376
rect 41506 9364 41512 9376
rect 40368 9336 41512 9364
rect 40368 9324 40374 9336
rect 41506 9324 41512 9336
rect 41564 9324 41570 9376
rect 41616 9364 41644 9404
rect 47302 9392 47308 9404
rect 47360 9392 47366 9444
rect 48314 9392 48320 9444
rect 48372 9432 48378 9444
rect 51077 9435 51135 9441
rect 48372 9404 50568 9432
rect 48372 9392 48378 9404
rect 42610 9364 42616 9376
rect 41616 9336 42616 9364
rect 42610 9324 42616 9336
rect 42668 9324 42674 9376
rect 42794 9364 42800 9376
rect 42755 9336 42800 9364
rect 42794 9324 42800 9336
rect 42852 9324 42858 9376
rect 44450 9324 44456 9376
rect 44508 9364 44514 9376
rect 46569 9367 46627 9373
rect 46569 9364 46581 9367
rect 44508 9336 46581 9364
rect 44508 9324 44514 9336
rect 46569 9333 46581 9336
rect 46615 9333 46627 9367
rect 46569 9327 46627 9333
rect 46658 9324 46664 9376
rect 46716 9364 46722 9376
rect 50430 9364 50436 9376
rect 46716 9336 50436 9364
rect 46716 9324 46722 9336
rect 50430 9324 50436 9336
rect 50488 9324 50494 9376
rect 50540 9364 50568 9404
rect 51077 9401 51089 9435
rect 51123 9432 51135 9435
rect 51350 9432 51356 9444
rect 51123 9404 51356 9432
rect 51123 9401 51135 9404
rect 51077 9395 51135 9401
rect 51350 9392 51356 9404
rect 51408 9392 51414 9444
rect 53742 9432 53748 9444
rect 51460 9404 53748 9432
rect 51460 9364 51488 9404
rect 53742 9392 53748 9404
rect 53800 9392 53806 9444
rect 54294 9392 54300 9444
rect 54352 9432 54358 9444
rect 54941 9435 54999 9441
rect 54941 9432 54953 9435
rect 54352 9404 54953 9432
rect 54352 9392 54358 9404
rect 54941 9401 54953 9404
rect 54987 9401 54999 9435
rect 54941 9395 54999 9401
rect 55030 9392 55036 9444
rect 55088 9432 55094 9444
rect 56134 9432 56140 9444
rect 55088 9404 56140 9432
rect 55088 9392 55094 9404
rect 56134 9392 56140 9404
rect 56192 9392 56198 9444
rect 56428 9404 57744 9432
rect 50540 9336 51488 9364
rect 51626 9324 51632 9376
rect 51684 9364 51690 9376
rect 52270 9364 52276 9376
rect 51684 9336 52276 9364
rect 51684 9324 51690 9336
rect 52270 9324 52276 9336
rect 52328 9324 52334 9376
rect 52454 9324 52460 9376
rect 52512 9364 52518 9376
rect 53377 9367 53435 9373
rect 53377 9364 53389 9367
rect 52512 9336 53389 9364
rect 52512 9324 52518 9336
rect 53377 9333 53389 9336
rect 53423 9333 53435 9367
rect 53377 9327 53435 9333
rect 54113 9367 54171 9373
rect 54113 9333 54125 9367
rect 54159 9364 54171 9367
rect 54389 9367 54447 9373
rect 54389 9364 54401 9367
rect 54159 9336 54401 9364
rect 54159 9333 54171 9336
rect 54113 9327 54171 9333
rect 54389 9333 54401 9336
rect 54435 9364 54447 9367
rect 56428 9364 56456 9404
rect 54435 9336 56456 9364
rect 54435 9333 54447 9336
rect 54389 9327 54447 9333
rect 56502 9324 56508 9376
rect 56560 9364 56566 9376
rect 56781 9367 56839 9373
rect 56781 9364 56793 9367
rect 56560 9336 56793 9364
rect 56560 9324 56566 9336
rect 56781 9333 56793 9336
rect 56827 9333 56839 9367
rect 56781 9327 56839 9333
rect 56870 9324 56876 9376
rect 56928 9364 56934 9376
rect 57330 9364 57336 9376
rect 56928 9336 57336 9364
rect 56928 9324 56934 9336
rect 57330 9324 57336 9336
rect 57388 9324 57394 9376
rect 57514 9324 57520 9376
rect 57572 9364 57578 9376
rect 57609 9367 57667 9373
rect 57609 9364 57621 9367
rect 57572 9336 57621 9364
rect 57572 9324 57578 9336
rect 57609 9333 57621 9336
rect 57655 9333 57667 9367
rect 57716 9364 57744 9404
rect 57790 9392 57796 9444
rect 57848 9432 57854 9444
rect 60366 9432 60372 9444
rect 57848 9404 60372 9432
rect 57848 9392 57854 9404
rect 60366 9392 60372 9404
rect 60424 9392 60430 9444
rect 60660 9432 60688 9540
rect 60826 9528 60832 9580
rect 60884 9568 60890 9580
rect 62209 9571 62267 9577
rect 62209 9568 62221 9571
rect 60884 9540 62221 9568
rect 60884 9528 60890 9540
rect 62209 9537 62221 9540
rect 62255 9537 62267 9571
rect 62209 9531 62267 9537
rect 62482 9528 62488 9580
rect 62540 9568 62546 9580
rect 69106 9568 69112 9580
rect 62540 9540 69112 9568
rect 62540 9528 62546 9540
rect 69106 9528 69112 9540
rect 69164 9528 69170 9580
rect 69201 9571 69259 9577
rect 69201 9537 69213 9571
rect 69247 9568 69259 9571
rect 70578 9568 70584 9580
rect 69247 9540 70584 9568
rect 69247 9537 69259 9540
rect 69201 9531 69259 9537
rect 70578 9528 70584 9540
rect 70636 9528 70642 9580
rect 74350 9568 74356 9580
rect 74311 9540 74356 9568
rect 74350 9528 74356 9540
rect 74408 9528 74414 9580
rect 74736 9577 74764 9608
rect 79689 9605 79701 9639
rect 79735 9636 79747 9639
rect 80238 9636 80244 9648
rect 79735 9608 80244 9636
rect 79735 9605 79747 9608
rect 79689 9599 79747 9605
rect 80238 9596 80244 9608
rect 80296 9596 80302 9648
rect 82814 9596 82820 9648
rect 82872 9636 82878 9648
rect 87138 9636 87144 9648
rect 82872 9608 87144 9636
rect 82872 9596 82878 9608
rect 87138 9596 87144 9608
rect 87196 9596 87202 9648
rect 93136 9636 93164 9676
rect 93302 9664 93308 9676
rect 93360 9664 93366 9716
rect 93394 9664 93400 9716
rect 93452 9664 93458 9716
rect 93486 9664 93492 9716
rect 93544 9704 93550 9716
rect 106182 9704 106188 9716
rect 93544 9676 106188 9704
rect 93544 9664 93550 9676
rect 106182 9664 106188 9676
rect 106240 9664 106246 9716
rect 108574 9664 108580 9716
rect 108632 9704 108638 9716
rect 120994 9704 121000 9716
rect 108632 9676 121000 9704
rect 108632 9664 108638 9676
rect 120994 9664 121000 9676
rect 121052 9664 121058 9716
rect 121196 9676 122604 9704
rect 93412 9636 93440 9664
rect 93136 9608 93440 9636
rect 97626 9596 97632 9648
rect 97684 9636 97690 9648
rect 100846 9636 100852 9648
rect 97684 9608 100852 9636
rect 97684 9596 97690 9608
rect 100846 9596 100852 9608
rect 100904 9596 100910 9648
rect 101585 9639 101643 9645
rect 101585 9605 101597 9639
rect 101631 9636 101643 9639
rect 104618 9636 104624 9648
rect 101631 9608 104624 9636
rect 101631 9605 101643 9608
rect 101585 9599 101643 9605
rect 104618 9596 104624 9608
rect 104676 9596 104682 9648
rect 104986 9596 104992 9648
rect 105044 9636 105050 9648
rect 111150 9636 111156 9648
rect 105044 9608 111012 9636
rect 111111 9608 111156 9636
rect 105044 9596 105050 9608
rect 74721 9571 74779 9577
rect 74721 9537 74733 9571
rect 74767 9537 74779 9571
rect 74721 9531 74779 9537
rect 76377 9571 76435 9577
rect 76377 9537 76389 9571
rect 76423 9568 76435 9571
rect 76926 9568 76932 9580
rect 76423 9540 76932 9568
rect 76423 9537 76435 9540
rect 76377 9531 76435 9537
rect 76926 9528 76932 9540
rect 76984 9528 76990 9580
rect 80606 9528 80612 9580
rect 80664 9568 80670 9580
rect 80701 9571 80759 9577
rect 80701 9568 80713 9571
rect 80664 9540 80713 9568
rect 80664 9528 80670 9540
rect 80701 9537 80713 9540
rect 80747 9537 80759 9571
rect 80701 9531 80759 9537
rect 81897 9571 81955 9577
rect 81897 9537 81909 9571
rect 81943 9537 81955 9571
rect 81897 9531 81955 9537
rect 82909 9571 82967 9577
rect 82909 9537 82921 9571
rect 82955 9568 82967 9571
rect 83182 9568 83188 9580
rect 82955 9540 83188 9568
rect 82955 9537 82967 9540
rect 82909 9531 82967 9537
rect 61930 9460 61936 9512
rect 61988 9500 61994 9512
rect 66990 9500 66996 9512
rect 61988 9472 66996 9500
rect 61988 9460 61994 9472
rect 66990 9460 66996 9472
rect 67048 9460 67054 9512
rect 74534 9500 74540 9512
rect 74495 9472 74540 9500
rect 74534 9460 74540 9472
rect 74592 9460 74598 9512
rect 80790 9500 80796 9512
rect 80751 9472 80796 9500
rect 80790 9460 80796 9472
rect 80848 9460 80854 9512
rect 81912 9500 81940 9531
rect 83182 9528 83188 9540
rect 83240 9568 83246 9580
rect 84562 9568 84568 9580
rect 83240 9540 84568 9568
rect 83240 9528 83246 9540
rect 84562 9528 84568 9540
rect 84620 9528 84626 9580
rect 86589 9571 86647 9577
rect 86589 9537 86601 9571
rect 86635 9568 86647 9571
rect 86954 9568 86960 9580
rect 86635 9540 86960 9568
rect 86635 9537 86647 9540
rect 86589 9531 86647 9537
rect 86954 9528 86960 9540
rect 87012 9568 87018 9580
rect 87506 9568 87512 9580
rect 87012 9540 87512 9568
rect 87012 9528 87018 9540
rect 87506 9528 87512 9540
rect 87564 9528 87570 9580
rect 88153 9571 88211 9577
rect 88153 9537 88165 9571
rect 88199 9568 88211 9571
rect 88518 9568 88524 9580
rect 88199 9540 88524 9568
rect 88199 9537 88211 9540
rect 88153 9531 88211 9537
rect 88518 9528 88524 9540
rect 88576 9528 88582 9580
rect 91465 9571 91523 9577
rect 91465 9537 91477 9571
rect 91511 9568 91523 9571
rect 92014 9568 92020 9580
rect 91511 9540 92020 9568
rect 91511 9537 91523 9540
rect 91465 9531 91523 9537
rect 92014 9528 92020 9540
rect 92072 9528 92078 9580
rect 92750 9568 92756 9580
rect 92711 9540 92756 9568
rect 92750 9528 92756 9540
rect 92808 9528 92814 9580
rect 94314 9528 94320 9580
rect 94372 9568 94378 9580
rect 97902 9568 97908 9580
rect 94372 9540 97488 9568
rect 97863 9540 97908 9568
rect 94372 9528 94378 9540
rect 83458 9500 83464 9512
rect 81912 9472 83464 9500
rect 83458 9460 83464 9472
rect 83516 9460 83522 9512
rect 86494 9460 86500 9512
rect 86552 9500 86558 9512
rect 87601 9503 87659 9509
rect 87601 9500 87613 9503
rect 86552 9472 87613 9500
rect 86552 9460 86558 9472
rect 87601 9469 87613 9472
rect 87647 9469 87659 9503
rect 87601 9463 87659 9469
rect 88981 9503 89039 9509
rect 88981 9469 88993 9503
rect 89027 9500 89039 9503
rect 89898 9500 89904 9512
rect 89027 9472 89904 9500
rect 89027 9469 89039 9472
rect 88981 9463 89039 9469
rect 89898 9460 89904 9472
rect 89956 9460 89962 9512
rect 90266 9500 90272 9512
rect 90227 9472 90272 9500
rect 90266 9460 90272 9472
rect 90324 9460 90330 9512
rect 91646 9460 91652 9512
rect 91704 9500 91710 9512
rect 92477 9503 92535 9509
rect 92477 9500 92489 9503
rect 91704 9472 92489 9500
rect 91704 9460 91710 9472
rect 92477 9469 92489 9472
rect 92523 9469 92535 9503
rect 92477 9463 92535 9469
rect 92842 9460 92848 9512
rect 92900 9500 92906 9512
rect 93857 9503 93915 9509
rect 93857 9500 93869 9503
rect 92900 9472 93869 9500
rect 92900 9460 92906 9472
rect 93857 9469 93869 9472
rect 93903 9469 93915 9503
rect 93857 9463 93915 9469
rect 96433 9503 96491 9509
rect 96433 9469 96445 9503
rect 96479 9500 96491 9503
rect 96614 9500 96620 9512
rect 96479 9472 96620 9500
rect 96479 9469 96491 9472
rect 96433 9463 96491 9469
rect 96614 9460 96620 9472
rect 96672 9460 96678 9512
rect 97460 9509 97488 9540
rect 97902 9528 97908 9540
rect 97960 9528 97966 9580
rect 100389 9571 100447 9577
rect 100389 9537 100401 9571
rect 100435 9568 100447 9571
rect 101030 9568 101036 9580
rect 100435 9540 101036 9568
rect 100435 9537 100447 9540
rect 100389 9531 100447 9537
rect 101030 9528 101036 9540
rect 101088 9528 101094 9580
rect 104710 9568 104716 9580
rect 104084 9540 104572 9568
rect 104671 9540 104716 9568
rect 97445 9503 97503 9509
rect 97445 9469 97457 9503
rect 97491 9469 97503 9503
rect 97445 9463 97503 9469
rect 98178 9460 98184 9512
rect 98236 9500 98242 9512
rect 98825 9503 98883 9509
rect 98825 9500 98837 9503
rect 98236 9472 98837 9500
rect 98236 9460 98242 9472
rect 98825 9469 98837 9472
rect 98871 9500 98883 9503
rect 99742 9500 99748 9512
rect 98871 9472 99748 9500
rect 98871 9469 98883 9472
rect 98825 9463 98883 9469
rect 99742 9460 99748 9472
rect 99800 9460 99806 9512
rect 99837 9503 99895 9509
rect 99837 9469 99849 9503
rect 99883 9469 99895 9503
rect 99837 9463 99895 9469
rect 103149 9503 103207 9509
rect 103149 9469 103161 9503
rect 103195 9500 103207 9503
rect 103330 9500 103336 9512
rect 103195 9472 103336 9500
rect 103195 9469 103207 9472
rect 103149 9463 103207 9469
rect 62206 9432 62212 9444
rect 60660 9404 62212 9432
rect 62206 9392 62212 9404
rect 62264 9392 62270 9444
rect 83001 9435 83059 9441
rect 83001 9401 83013 9435
rect 83047 9432 83059 9435
rect 83090 9432 83096 9444
rect 83047 9404 83096 9432
rect 83047 9401 83059 9404
rect 83001 9395 83059 9401
rect 83090 9392 83096 9404
rect 83148 9392 83154 9444
rect 95694 9392 95700 9444
rect 95752 9432 95758 9444
rect 99852 9432 99880 9463
rect 103330 9460 103336 9472
rect 103388 9460 103394 9512
rect 95752 9404 99880 9432
rect 95752 9392 95758 9404
rect 100938 9392 100944 9444
rect 100996 9432 101002 9444
rect 104084 9432 104112 9540
rect 104161 9503 104219 9509
rect 104161 9469 104173 9503
rect 104207 9469 104219 9503
rect 104161 9463 104219 9469
rect 100996 9404 104112 9432
rect 100996 9392 101002 9404
rect 59078 9364 59084 9376
rect 57716 9336 59084 9364
rect 57609 9327 57667 9333
rect 59078 9324 59084 9336
rect 59136 9324 59142 9376
rect 59173 9367 59231 9373
rect 59173 9333 59185 9367
rect 59219 9364 59231 9367
rect 59538 9364 59544 9376
rect 59219 9336 59544 9364
rect 59219 9333 59231 9336
rect 59173 9327 59231 9333
rect 59538 9324 59544 9336
rect 59596 9324 59602 9376
rect 60458 9324 60464 9376
rect 60516 9364 60522 9376
rect 62942 9364 62948 9376
rect 60516 9336 62948 9364
rect 60516 9324 60522 9336
rect 62942 9324 62948 9336
rect 63000 9324 63006 9376
rect 63034 9324 63040 9376
rect 63092 9364 63098 9376
rect 68462 9364 68468 9376
rect 63092 9336 68468 9364
rect 63092 9324 63098 9336
rect 68462 9324 68468 9336
rect 68520 9324 68526 9376
rect 76466 9364 76472 9376
rect 76427 9336 76472 9364
rect 76466 9324 76472 9336
rect 76524 9324 76530 9376
rect 76558 9324 76564 9376
rect 76616 9364 76622 9376
rect 81989 9367 82047 9373
rect 81989 9364 82001 9367
rect 76616 9336 82001 9364
rect 76616 9324 76622 9336
rect 81989 9333 82001 9336
rect 82035 9333 82047 9367
rect 88518 9364 88524 9376
rect 88479 9336 88524 9364
rect 81989 9327 82047 9333
rect 88518 9324 88524 9336
rect 88576 9324 88582 9376
rect 90174 9324 90180 9376
rect 90232 9364 90238 9376
rect 91186 9364 91192 9376
rect 90232 9336 91192 9364
rect 90232 9324 90238 9336
rect 91186 9324 91192 9336
rect 91244 9324 91250 9376
rect 94314 9364 94320 9376
rect 94275 9336 94320 9364
rect 94314 9324 94320 9336
rect 94372 9324 94378 9376
rect 99650 9324 99656 9376
rect 99708 9364 99714 9376
rect 104176 9364 104204 9463
rect 99708 9336 104204 9364
rect 104544 9364 104572 9540
rect 104710 9528 104716 9540
rect 104768 9528 104774 9580
rect 105998 9528 106004 9580
rect 106056 9568 106062 9580
rect 108206 9568 108212 9580
rect 106056 9540 108212 9568
rect 106056 9528 106062 9540
rect 108206 9528 108212 9540
rect 108264 9528 108270 9580
rect 109586 9568 109592 9580
rect 109547 9540 109592 9568
rect 109586 9528 109592 9540
rect 109644 9528 109650 9580
rect 110984 9568 111012 9608
rect 111150 9596 111156 9608
rect 111208 9596 111214 9648
rect 112809 9639 112867 9645
rect 112809 9605 112821 9639
rect 112855 9636 112867 9639
rect 113361 9639 113419 9645
rect 113361 9636 113373 9639
rect 112855 9608 113373 9636
rect 112855 9605 112867 9608
rect 112809 9599 112867 9605
rect 113361 9605 113373 9608
rect 113407 9636 113419 9639
rect 113450 9636 113456 9648
rect 113407 9608 113456 9636
rect 113407 9605 113419 9608
rect 113361 9599 113419 9605
rect 113450 9596 113456 9608
rect 113508 9596 113514 9648
rect 113542 9596 113548 9648
rect 113600 9636 113606 9648
rect 119246 9636 119252 9648
rect 113600 9608 119252 9636
rect 113600 9596 113606 9608
rect 119246 9596 119252 9608
rect 119304 9596 119310 9648
rect 121196 9636 121224 9676
rect 119356 9608 121224 9636
rect 122576 9636 122604 9676
rect 122742 9664 122748 9716
rect 122800 9704 122806 9716
rect 129182 9704 129188 9716
rect 122800 9676 129188 9704
rect 122800 9664 122806 9676
rect 129182 9664 129188 9676
rect 129240 9664 129246 9716
rect 132129 9707 132187 9713
rect 132129 9673 132141 9707
rect 132175 9704 132187 9707
rect 132402 9704 132408 9716
rect 132175 9676 132408 9704
rect 132175 9673 132187 9676
rect 132129 9667 132187 9673
rect 132402 9664 132408 9676
rect 132460 9664 132466 9716
rect 141050 9704 141056 9716
rect 134996 9676 135300 9704
rect 141011 9676 141056 9704
rect 125318 9636 125324 9648
rect 122576 9608 125324 9636
rect 112533 9571 112591 9577
rect 112533 9568 112545 9571
rect 110984 9540 112545 9568
rect 112533 9537 112545 9540
rect 112579 9537 112591 9571
rect 115198 9568 115204 9580
rect 115159 9540 115204 9568
rect 112533 9531 112591 9537
rect 115198 9528 115204 9540
rect 115256 9528 115262 9580
rect 117406 9528 117412 9580
rect 117464 9568 117470 9580
rect 119356 9568 119384 9608
rect 125318 9596 125324 9608
rect 125376 9596 125382 9648
rect 126882 9636 126888 9648
rect 126843 9608 126888 9636
rect 126882 9596 126888 9608
rect 126940 9596 126946 9648
rect 127802 9636 127808 9648
rect 127763 9608 127808 9636
rect 127802 9596 127808 9608
rect 127860 9596 127866 9648
rect 133138 9636 133144 9648
rect 133099 9608 133144 9636
rect 133138 9596 133144 9608
rect 133196 9596 133202 9648
rect 133322 9596 133328 9648
rect 133380 9636 133386 9648
rect 134996 9636 135024 9676
rect 135162 9636 135168 9648
rect 133380 9608 135024 9636
rect 135123 9608 135168 9636
rect 133380 9596 133386 9608
rect 135162 9596 135168 9608
rect 135220 9596 135226 9648
rect 135272 9636 135300 9676
rect 141050 9664 141056 9676
rect 141108 9664 141114 9716
rect 143997 9707 144055 9713
rect 143997 9673 144009 9707
rect 144043 9704 144055 9707
rect 144546 9704 144552 9716
rect 144043 9676 144552 9704
rect 144043 9673 144055 9676
rect 143997 9667 144055 9673
rect 144546 9664 144552 9676
rect 144604 9664 144610 9716
rect 148226 9704 148232 9716
rect 148187 9676 148232 9704
rect 148226 9664 148232 9676
rect 148284 9664 148290 9716
rect 148778 9664 148784 9716
rect 148836 9704 148842 9716
rect 153013 9707 153071 9713
rect 153013 9704 153025 9707
rect 148836 9676 153025 9704
rect 148836 9664 148842 9676
rect 153013 9673 153025 9676
rect 153059 9673 153071 9707
rect 153013 9667 153071 9673
rect 137741 9639 137799 9645
rect 135272 9608 136772 9636
rect 120442 9568 120448 9580
rect 117464 9540 119384 9568
rect 120403 9540 120448 9568
rect 117464 9528 117470 9540
rect 120442 9528 120448 9540
rect 120500 9528 120506 9580
rect 121454 9568 121460 9580
rect 121367 9540 121460 9568
rect 121454 9528 121460 9540
rect 121512 9568 121518 9580
rect 122190 9568 122196 9580
rect 121512 9540 122196 9568
rect 121512 9528 121518 9540
rect 122190 9528 122196 9540
rect 122248 9528 122254 9580
rect 123021 9571 123079 9577
rect 123021 9537 123033 9571
rect 123067 9568 123079 9571
rect 123570 9568 123576 9580
rect 123067 9540 123576 9568
rect 123067 9537 123079 9540
rect 123021 9531 123079 9537
rect 123570 9528 123576 9540
rect 123628 9528 123634 9580
rect 125965 9571 126023 9577
rect 125965 9537 125977 9571
rect 126011 9537 126023 9571
rect 125965 9531 126023 9537
rect 126793 9571 126851 9577
rect 126793 9537 126805 9571
rect 126839 9568 126851 9571
rect 127066 9568 127072 9580
rect 126839 9540 127072 9568
rect 126839 9537 126851 9540
rect 126793 9531 126851 9537
rect 108117 9503 108175 9509
rect 108117 9469 108129 9503
rect 108163 9500 108175 9503
rect 108298 9500 108304 9512
rect 108163 9472 108304 9500
rect 108163 9469 108175 9472
rect 108117 9463 108175 9469
rect 108298 9460 108304 9472
rect 108356 9460 108362 9512
rect 108482 9460 108488 9512
rect 108540 9500 108546 9512
rect 109129 9503 109187 9509
rect 109129 9500 109141 9503
rect 108540 9472 109141 9500
rect 108540 9460 108546 9472
rect 109129 9469 109141 9472
rect 109175 9469 109187 9503
rect 109129 9463 109187 9469
rect 113910 9460 113916 9512
rect 113968 9500 113974 9512
rect 114005 9503 114063 9509
rect 114005 9500 114017 9503
rect 113968 9472 114017 9500
rect 113968 9460 113974 9472
rect 114005 9469 114017 9472
rect 114051 9469 114063 9503
rect 114005 9463 114063 9469
rect 114112 9472 115428 9500
rect 107930 9392 107936 9444
rect 107988 9432 107994 9444
rect 114112 9432 114140 9472
rect 115290 9432 115296 9444
rect 107988 9404 114140 9432
rect 115251 9404 115296 9432
rect 107988 9392 107994 9404
rect 115290 9392 115296 9404
rect 115348 9392 115354 9444
rect 115400 9432 115428 9472
rect 115566 9460 115572 9512
rect 115624 9500 115630 9512
rect 115937 9503 115995 9509
rect 115937 9500 115949 9503
rect 115624 9472 115949 9500
rect 115624 9460 115630 9472
rect 115937 9469 115949 9472
rect 115983 9500 115995 9503
rect 116397 9503 116455 9509
rect 116397 9500 116409 9503
rect 115983 9472 116409 9500
rect 115983 9469 115995 9472
rect 115937 9463 115995 9469
rect 116397 9469 116409 9472
rect 116443 9469 116455 9503
rect 116397 9463 116455 9469
rect 118786 9460 118792 9512
rect 118844 9500 118850 9512
rect 118881 9503 118939 9509
rect 118881 9500 118893 9503
rect 118844 9472 118893 9500
rect 118844 9460 118850 9472
rect 118881 9469 118893 9472
rect 118927 9469 118939 9503
rect 119890 9500 119896 9512
rect 119851 9472 119896 9500
rect 118881 9463 118939 9469
rect 119890 9460 119896 9472
rect 119948 9460 119954 9512
rect 120994 9460 121000 9512
rect 121052 9500 121058 9512
rect 122466 9500 122472 9512
rect 121052 9472 121500 9500
rect 122427 9472 122472 9500
rect 121052 9460 121058 9472
rect 120718 9432 120724 9444
rect 115400 9404 120724 9432
rect 120718 9392 120724 9404
rect 120776 9392 120782 9444
rect 121472 9432 121500 9472
rect 122466 9460 122472 9472
rect 122524 9460 122530 9512
rect 124401 9503 124459 9509
rect 124401 9469 124413 9503
rect 124447 9500 124459 9503
rect 124582 9500 124588 9512
rect 124447 9472 124588 9500
rect 124447 9469 124459 9472
rect 124401 9463 124459 9469
rect 124582 9460 124588 9472
rect 124640 9460 124646 9512
rect 125413 9503 125471 9509
rect 125413 9469 125425 9503
rect 125459 9469 125471 9503
rect 125980 9500 126008 9531
rect 127066 9528 127072 9540
rect 127124 9568 127130 9580
rect 129458 9568 129464 9580
rect 127124 9540 129464 9568
rect 127124 9528 127130 9540
rect 129458 9528 129464 9540
rect 129516 9528 129522 9580
rect 131114 9568 131120 9580
rect 131075 9540 131120 9568
rect 131114 9528 131120 9540
rect 131172 9568 131178 9580
rect 131577 9571 131635 9577
rect 131577 9568 131589 9571
rect 131172 9540 131589 9568
rect 131172 9528 131178 9540
rect 131577 9537 131589 9540
rect 131623 9537 131635 9571
rect 131577 9531 131635 9537
rect 132586 9528 132592 9580
rect 132644 9568 132650 9580
rect 136634 9568 136640 9580
rect 132644 9540 136640 9568
rect 132644 9528 132650 9540
rect 136634 9528 136640 9540
rect 136692 9528 136698 9580
rect 136744 9568 136772 9608
rect 137741 9605 137753 9639
rect 137787 9636 137799 9639
rect 138106 9636 138112 9648
rect 137787 9608 138112 9636
rect 137787 9605 137799 9608
rect 137741 9599 137799 9605
rect 138106 9596 138112 9608
rect 138164 9596 138170 9648
rect 139213 9639 139271 9645
rect 139213 9605 139225 9639
rect 139259 9636 139271 9639
rect 140222 9636 140228 9648
rect 139259 9608 140228 9636
rect 139259 9605 139271 9608
rect 139213 9599 139271 9605
rect 140222 9596 140228 9608
rect 140280 9596 140286 9648
rect 141602 9596 141608 9648
rect 141660 9636 141666 9648
rect 142062 9636 142068 9648
rect 141660 9608 142068 9636
rect 141660 9596 141666 9608
rect 142062 9596 142068 9608
rect 142120 9596 142126 9648
rect 142430 9596 142436 9648
rect 142488 9636 142494 9648
rect 147490 9636 147496 9648
rect 142488 9608 147496 9636
rect 142488 9596 142494 9608
rect 147490 9596 147496 9608
rect 147548 9596 147554 9648
rect 147766 9596 147772 9648
rect 147824 9636 147830 9648
rect 151814 9636 151820 9648
rect 147824 9608 150756 9636
rect 151775 9608 151820 9636
rect 147824 9596 147830 9608
rect 138382 9568 138388 9580
rect 136744 9540 138388 9568
rect 138382 9528 138388 9540
rect 138440 9528 138446 9580
rect 138750 9528 138756 9580
rect 138808 9568 138814 9580
rect 142338 9568 142344 9580
rect 138808 9540 142344 9568
rect 138808 9528 138814 9540
rect 142338 9528 142344 9540
rect 142396 9528 142402 9580
rect 143166 9568 143172 9580
rect 143127 9540 143172 9568
rect 143166 9528 143172 9540
rect 143224 9528 143230 9580
rect 147953 9571 148011 9577
rect 147953 9537 147965 9571
rect 147999 9568 148011 9571
rect 148042 9568 148048 9580
rect 147999 9540 148048 9568
rect 147999 9537 148011 9540
rect 147953 9531 148011 9537
rect 148042 9528 148048 9540
rect 148100 9528 148106 9580
rect 148134 9528 148140 9580
rect 148192 9568 148198 9580
rect 148778 9568 148784 9580
rect 148192 9540 148784 9568
rect 148192 9528 148198 9540
rect 148778 9528 148784 9540
rect 148836 9528 148842 9580
rect 150158 9568 150164 9580
rect 150119 9540 150164 9568
rect 150158 9528 150164 9540
rect 150216 9568 150222 9580
rect 150621 9571 150679 9577
rect 150621 9568 150633 9571
rect 150216 9540 150633 9568
rect 150216 9528 150222 9540
rect 150621 9537 150633 9540
rect 150667 9537 150679 9571
rect 150728 9568 150756 9608
rect 151814 9596 151820 9608
rect 151872 9596 151878 9648
rect 157150 9596 157156 9648
rect 157208 9636 157214 9648
rect 158806 9636 158812 9648
rect 157208 9608 158812 9636
rect 157208 9596 157214 9608
rect 158806 9596 158812 9608
rect 158864 9596 158870 9648
rect 160005 9639 160063 9645
rect 160005 9605 160017 9639
rect 160051 9636 160063 9639
rect 160462 9636 160468 9648
rect 160051 9608 160468 9636
rect 160051 9605 160063 9608
rect 160005 9599 160063 9605
rect 160462 9596 160468 9608
rect 160520 9596 160526 9648
rect 162121 9639 162179 9645
rect 162121 9605 162133 9639
rect 162167 9636 162179 9639
rect 162167 9608 165660 9636
rect 162167 9605 162179 9608
rect 162121 9599 162179 9605
rect 154114 9568 154120 9580
rect 150728 9540 154120 9568
rect 150621 9531 150679 9537
rect 154114 9528 154120 9540
rect 154172 9528 154178 9580
rect 154301 9571 154359 9577
rect 154301 9537 154313 9571
rect 154347 9568 154359 9571
rect 154942 9568 154948 9580
rect 154347 9540 154948 9568
rect 154347 9537 154359 9540
rect 154301 9531 154359 9537
rect 154942 9528 154948 9540
rect 155000 9528 155006 9580
rect 155865 9571 155923 9577
rect 155865 9537 155877 9571
rect 155911 9568 155923 9571
rect 156230 9568 156236 9580
rect 155911 9540 156236 9568
rect 155911 9537 155923 9540
rect 155865 9531 155923 9537
rect 156230 9528 156236 9540
rect 156288 9528 156294 9580
rect 159177 9571 159235 9577
rect 159177 9537 159189 9571
rect 159223 9568 159235 9571
rect 159266 9568 159272 9580
rect 159223 9540 159272 9568
rect 159223 9537 159235 9540
rect 159177 9531 159235 9537
rect 159266 9528 159272 9540
rect 159324 9528 159330 9580
rect 163130 9528 163136 9580
rect 163188 9568 163194 9580
rect 164326 9568 164332 9580
rect 163188 9540 163728 9568
rect 164287 9540 164332 9568
rect 163188 9528 163194 9540
rect 127158 9500 127164 9512
rect 125980 9472 127164 9500
rect 125413 9463 125471 9469
rect 123294 9432 123300 9444
rect 121104 9404 121408 9432
rect 121472 9404 123300 9432
rect 108482 9364 108488 9376
rect 104544 9336 108488 9364
rect 99708 9324 99714 9336
rect 108482 9324 108488 9336
rect 108540 9324 108546 9376
rect 112533 9367 112591 9373
rect 112533 9333 112545 9367
rect 112579 9364 112591 9367
rect 121104 9364 121132 9404
rect 121270 9364 121276 9376
rect 112579 9336 121132 9364
rect 121231 9336 121276 9364
rect 112579 9333 112591 9336
rect 112533 9327 112591 9333
rect 121270 9324 121276 9336
rect 121328 9324 121334 9376
rect 121380 9364 121408 9404
rect 123294 9392 123300 9404
rect 123352 9392 123358 9444
rect 125428 9364 125456 9463
rect 127158 9460 127164 9472
rect 127216 9460 127222 9512
rect 129369 9503 129427 9509
rect 129369 9469 129381 9503
rect 129415 9500 129427 9503
rect 129737 9503 129795 9509
rect 129737 9500 129749 9503
rect 129415 9472 129749 9500
rect 129415 9469 129427 9472
rect 129369 9463 129427 9469
rect 129737 9469 129749 9472
rect 129783 9500 129795 9503
rect 129826 9500 129832 9512
rect 129783 9472 129832 9500
rect 129783 9469 129795 9472
rect 129737 9463 129795 9469
rect 129826 9460 129832 9472
rect 129884 9460 129890 9512
rect 130746 9500 130752 9512
rect 130707 9472 130752 9500
rect 130746 9460 130752 9472
rect 130804 9460 130810 9512
rect 131022 9460 131028 9512
rect 131080 9500 131086 9512
rect 134058 9500 134064 9512
rect 131080 9472 134064 9500
rect 131080 9460 131086 9472
rect 134058 9460 134064 9472
rect 134116 9460 134122 9512
rect 138474 9460 138480 9512
rect 138532 9500 138538 9512
rect 138532 9472 141464 9500
rect 138532 9460 138538 9472
rect 132126 9392 132132 9444
rect 132184 9432 132190 9444
rect 134794 9432 134800 9444
rect 132184 9404 134800 9432
rect 132184 9392 132190 9404
rect 134794 9392 134800 9404
rect 134852 9392 134858 9444
rect 139026 9432 139032 9444
rect 135732 9404 139032 9432
rect 127526 9364 127532 9376
rect 121380 9336 125456 9364
rect 127487 9336 127532 9364
rect 127526 9324 127532 9336
rect 127584 9324 127590 9376
rect 133598 9324 133604 9376
rect 133656 9364 133662 9376
rect 135732 9364 135760 9404
rect 139026 9392 139032 9404
rect 139084 9392 139090 9444
rect 141436 9432 141464 9472
rect 141510 9460 141516 9512
rect 141568 9500 141574 9512
rect 141605 9503 141663 9509
rect 141605 9500 141617 9503
rect 141568 9472 141617 9500
rect 141568 9460 141574 9472
rect 141605 9469 141617 9472
rect 141651 9469 141663 9503
rect 142890 9500 142896 9512
rect 141605 9463 141663 9469
rect 141712 9472 142896 9500
rect 141712 9432 141740 9472
rect 142890 9460 142896 9472
rect 142948 9460 142954 9512
rect 143077 9503 143135 9509
rect 143077 9469 143089 9503
rect 143123 9500 143135 9503
rect 144270 9500 144276 9512
rect 143123 9472 144276 9500
rect 143123 9469 143135 9472
rect 143077 9463 143135 9469
rect 144270 9460 144276 9472
rect 144328 9460 144334 9512
rect 145009 9503 145067 9509
rect 145009 9469 145021 9503
rect 145055 9500 145067 9503
rect 145926 9500 145932 9512
rect 145055 9472 145932 9500
rect 145055 9469 145067 9472
rect 145009 9463 145067 9469
rect 145926 9460 145932 9472
rect 145984 9500 145990 9512
rect 146389 9503 146447 9509
rect 146389 9500 146401 9503
rect 145984 9472 146401 9500
rect 145984 9460 145990 9472
rect 146389 9469 146401 9472
rect 146435 9469 146447 9503
rect 146389 9463 146447 9469
rect 147861 9503 147919 9509
rect 147861 9469 147873 9503
rect 147907 9500 147919 9503
rect 148594 9500 148600 9512
rect 147907 9472 148600 9500
rect 147907 9469 147919 9472
rect 147861 9463 147919 9469
rect 148594 9460 148600 9472
rect 148652 9460 148658 9512
rect 148689 9503 148747 9509
rect 148689 9469 148701 9503
rect 148735 9500 148747 9503
rect 149330 9500 149336 9512
rect 148735 9472 149336 9500
rect 148735 9469 148747 9472
rect 148689 9463 148747 9469
rect 149330 9460 149336 9472
rect 149388 9500 149394 9512
rect 152001 9503 152059 9509
rect 152001 9500 152013 9503
rect 149388 9472 152013 9500
rect 149388 9460 149394 9472
rect 152001 9469 152013 9472
rect 152047 9469 152059 9503
rect 155678 9500 155684 9512
rect 155639 9472 155684 9500
rect 152001 9463 152059 9469
rect 155678 9460 155684 9472
rect 155736 9460 155742 9512
rect 157150 9460 157156 9512
rect 157208 9500 157214 9512
rect 157613 9503 157671 9509
rect 157613 9500 157625 9503
rect 157208 9472 157625 9500
rect 157208 9460 157214 9472
rect 157613 9469 157625 9472
rect 157659 9469 157671 9503
rect 157613 9463 157671 9469
rect 157886 9460 157892 9512
rect 157944 9500 157950 9512
rect 158717 9503 158775 9509
rect 158717 9500 158729 9503
rect 157944 9472 158729 9500
rect 157944 9460 157950 9472
rect 158717 9469 158729 9472
rect 158763 9469 158775 9503
rect 158717 9463 158775 9469
rect 160462 9460 160468 9512
rect 160520 9500 160526 9512
rect 160557 9503 160615 9509
rect 160557 9500 160569 9503
rect 160520 9472 160569 9500
rect 160520 9460 160526 9472
rect 160557 9469 160569 9472
rect 160603 9500 160615 9503
rect 161017 9503 161075 9509
rect 161017 9500 161029 9503
rect 160603 9472 161029 9500
rect 160603 9469 160615 9472
rect 160557 9463 160615 9469
rect 161017 9469 161029 9472
rect 161063 9469 161075 9503
rect 163222 9500 163228 9512
rect 163183 9472 163228 9500
rect 161017 9463 161075 9469
rect 163222 9460 163228 9472
rect 163280 9460 163286 9512
rect 163700 9500 163728 9540
rect 164326 9528 164332 9540
rect 164384 9568 164390 9580
rect 165632 9577 165660 9608
rect 165065 9571 165123 9577
rect 165065 9568 165077 9571
rect 164384 9540 165077 9568
rect 164384 9528 164390 9540
rect 165065 9537 165077 9540
rect 165111 9537 165123 9571
rect 165065 9531 165123 9537
rect 165617 9571 165675 9577
rect 165617 9537 165629 9571
rect 165663 9568 165675 9571
rect 165798 9568 165804 9580
rect 165663 9540 165804 9568
rect 165663 9537 165675 9540
rect 165617 9531 165675 9537
rect 165798 9528 165804 9540
rect 165856 9528 165862 9580
rect 166902 9568 166908 9580
rect 166863 9540 166908 9568
rect 166902 9528 166908 9540
rect 166960 9528 166966 9580
rect 164237 9503 164295 9509
rect 164237 9500 164249 9503
rect 163700 9472 164249 9500
rect 164237 9469 164249 9472
rect 164283 9469 164295 9503
rect 164237 9463 164295 9469
rect 166629 9503 166687 9509
rect 166629 9469 166641 9503
rect 166675 9469 166687 9503
rect 166629 9463 166687 9469
rect 141436 9404 141740 9432
rect 141786 9392 141792 9444
rect 141844 9432 141850 9444
rect 145098 9432 145104 9444
rect 141844 9404 145104 9432
rect 141844 9392 141850 9404
rect 145098 9392 145104 9404
rect 145156 9392 145162 9444
rect 149514 9432 149520 9444
rect 145576 9404 149520 9432
rect 133656 9336 135760 9364
rect 133656 9324 133662 9336
rect 135806 9324 135812 9376
rect 135864 9364 135870 9376
rect 138106 9364 138112 9376
rect 135864 9336 138112 9364
rect 135864 9324 135870 9336
rect 138106 9324 138112 9336
rect 138164 9324 138170 9376
rect 138198 9324 138204 9376
rect 138256 9364 138262 9376
rect 142246 9364 142252 9376
rect 138256 9336 142252 9364
rect 138256 9324 138262 9336
rect 142246 9324 142252 9336
rect 142304 9324 142310 9376
rect 143534 9324 143540 9376
rect 143592 9364 143598 9376
rect 145576 9364 145604 9404
rect 149514 9392 149520 9404
rect 149572 9392 149578 9444
rect 150253 9435 150311 9441
rect 150253 9401 150265 9435
rect 150299 9432 150311 9435
rect 150894 9432 150900 9444
rect 150299 9404 150900 9432
rect 150299 9401 150311 9404
rect 150253 9395 150311 9401
rect 150894 9392 150900 9404
rect 150952 9392 150958 9444
rect 163406 9392 163412 9444
rect 163464 9432 163470 9444
rect 166644 9432 166672 9463
rect 163464 9404 166672 9432
rect 163464 9392 163470 9404
rect 143592 9336 145604 9364
rect 143592 9324 143598 9336
rect 145650 9324 145656 9376
rect 145708 9364 145714 9376
rect 151538 9364 151544 9376
rect 145708 9336 151544 9364
rect 145708 9324 145714 9336
rect 151538 9324 151544 9336
rect 151596 9324 151602 9376
rect 151722 9324 151728 9376
rect 151780 9364 151786 9376
rect 153746 9364 153752 9376
rect 151780 9336 153752 9364
rect 151780 9324 151786 9336
rect 153746 9324 153752 9336
rect 153804 9324 153810 9376
rect 156230 9364 156236 9376
rect 156191 9336 156236 9364
rect 156230 9324 156236 9336
rect 156288 9324 156294 9376
rect 157242 9364 157248 9376
rect 157203 9336 157248 9364
rect 157242 9324 157248 9336
rect 157300 9324 157306 9376
rect 159542 9364 159548 9376
rect 159455 9336 159548 9364
rect 159542 9324 159548 9336
rect 159600 9364 159606 9376
rect 160278 9364 160284 9376
rect 159600 9336 160284 9364
rect 159600 9324 159606 9336
rect 160278 9324 160284 9336
rect 160336 9324 160342 9376
rect 160830 9324 160836 9376
rect 160888 9364 160894 9376
rect 164878 9364 164884 9376
rect 160888 9336 164884 9364
rect 160888 9324 160894 9336
rect 164878 9324 164884 9336
rect 164936 9324 164942 9376
rect 368 9274 169556 9296
rect 368 9222 28456 9274
rect 28508 9222 28520 9274
rect 28572 9222 28584 9274
rect 28636 9222 28648 9274
rect 28700 9222 84878 9274
rect 84930 9222 84942 9274
rect 84994 9222 85006 9274
rect 85058 9222 85070 9274
rect 85122 9222 141299 9274
rect 141351 9222 141363 9274
rect 141415 9222 141427 9274
rect 141479 9222 141491 9274
rect 141543 9222 169556 9274
rect 368 9200 169556 9222
rect 3878 9160 3884 9172
rect 3839 9132 3884 9160
rect 3878 9120 3884 9132
rect 3936 9160 3942 9172
rect 3936 9132 4016 9160
rect 3936 9120 3942 9132
rect 3988 9033 4016 9132
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 8846 9160 8852 9172
rect 4672 9132 8852 9160
rect 4672 9120 4678 9132
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 17494 9160 17500 9172
rect 17455 9132 17500 9160
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 19886 9160 19892 9172
rect 19847 9132 19892 9160
rect 19886 9120 19892 9132
rect 19944 9120 19950 9172
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20530 9120 20536 9172
rect 20588 9160 20594 9172
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 20588 9132 21281 9160
rect 20588 9120 20594 9132
rect 21269 9129 21281 9132
rect 21315 9160 21327 9163
rect 21315 9132 21680 9160
rect 21315 9129 21327 9132
rect 21269 9123 21327 9129
rect 5626 9052 5632 9104
rect 5684 9092 5690 9104
rect 5684 9064 16344 9092
rect 5684 9052 5690 9064
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 4062 8984 4068 9036
rect 4120 9024 4126 9036
rect 4985 9027 5043 9033
rect 4985 9024 4997 9027
rect 4120 8996 4997 9024
rect 4120 8984 4126 8996
rect 4985 8993 4997 8996
rect 5031 8993 5043 9027
rect 5442 9024 5448 9036
rect 4985 8987 5043 8993
rect 5092 8996 5448 9024
rect 5092 8965 5120 8996
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 6362 9024 6368 9036
rect 6323 8996 6368 9024
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 7392 8956 7420 8987
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 15194 9024 15200 9036
rect 7800 8996 15200 9024
rect 7800 8984 7806 8996
rect 15194 8984 15200 8996
rect 15252 8984 15258 9036
rect 16316 9033 16344 9064
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 5224 8928 7420 8956
rect 7929 8959 7987 8965
rect 5224 8916 5230 8928
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8956 15347 8959
rect 15378 8956 15384 8968
rect 15335 8928 15384 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 7944 8888 7972 8919
rect 15378 8916 15384 8928
rect 15436 8956 15442 8968
rect 16114 8956 16120 8968
rect 15436 8928 16120 8956
rect 15436 8916 15442 8928
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 17512 8956 17540 9120
rect 18509 9095 18567 9101
rect 18509 9061 18521 9095
rect 18555 9092 18567 9095
rect 18785 9095 18843 9101
rect 18785 9092 18797 9095
rect 18555 9064 18797 9092
rect 18555 9061 18567 9064
rect 18509 9055 18567 9061
rect 18785 9061 18797 9064
rect 18831 9092 18843 9095
rect 21542 9092 21548 9104
rect 18831 9064 21548 9092
rect 18831 9061 18843 9064
rect 18785 9055 18843 9061
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 21652 9024 21680 9132
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 23569 9163 23627 9169
rect 23569 9160 23581 9163
rect 22060 9132 23581 9160
rect 22060 9120 22066 9132
rect 23569 9129 23581 9132
rect 23615 9129 23627 9163
rect 24854 9160 24860 9172
rect 24815 9132 24860 9160
rect 23569 9123 23627 9129
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 25314 9160 25320 9172
rect 25275 9132 25320 9160
rect 25314 9120 25320 9132
rect 25372 9120 25378 9172
rect 25406 9120 25412 9172
rect 25464 9160 25470 9172
rect 25869 9163 25927 9169
rect 25869 9160 25881 9163
rect 25464 9132 25881 9160
rect 25464 9120 25470 9132
rect 25869 9129 25881 9132
rect 25915 9129 25927 9163
rect 25869 9123 25927 9129
rect 25958 9120 25964 9172
rect 26016 9160 26022 9172
rect 28166 9160 28172 9172
rect 26016 9132 28172 9160
rect 26016 9120 26022 9132
rect 28166 9120 28172 9132
rect 28224 9120 28230 9172
rect 28261 9163 28319 9169
rect 28261 9129 28273 9163
rect 28307 9160 28319 9163
rect 28537 9163 28595 9169
rect 28537 9160 28549 9163
rect 28307 9132 28549 9160
rect 28307 9129 28319 9132
rect 28261 9123 28319 9129
rect 28537 9129 28549 9132
rect 28583 9160 28595 9163
rect 28810 9160 28816 9172
rect 28583 9132 28816 9160
rect 28583 9129 28595 9132
rect 28537 9123 28595 9129
rect 28810 9120 28816 9132
rect 28868 9120 28874 9172
rect 30282 9120 30288 9172
rect 30340 9160 30346 9172
rect 30929 9163 30987 9169
rect 30929 9160 30941 9163
rect 30340 9132 30941 9160
rect 30340 9120 30346 9132
rect 30929 9129 30941 9132
rect 30975 9129 30987 9163
rect 30929 9123 30987 9129
rect 31496 9132 34284 9160
rect 22186 9052 22192 9104
rect 22244 9092 22250 9104
rect 31496 9092 31524 9132
rect 31662 9092 31668 9104
rect 22244 9064 31524 9092
rect 31623 9064 31668 9092
rect 22244 9052 22250 9064
rect 31662 9052 31668 9064
rect 31720 9052 31726 9104
rect 22830 9024 22836 9036
rect 17644 8996 21588 9024
rect 21652 8996 22692 9024
rect 22791 8996 22836 9024
rect 17644 8984 17650 8996
rect 17681 8959 17739 8965
rect 17681 8956 17693 8959
rect 16899 8928 17264 8956
rect 17512 8928 17693 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 8294 8888 8300 8900
rect 7944 8860 8300 8888
rect 8294 8848 8300 8860
rect 8352 8848 8358 8900
rect 17236 8832 17264 8928
rect 17681 8925 17693 8928
rect 17727 8925 17739 8959
rect 18046 8956 18052 8968
rect 18007 8928 18052 8956
rect 17681 8919 17739 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8956 18475 8959
rect 18509 8959 18567 8965
rect 18509 8956 18521 8959
rect 18463 8928 18521 8956
rect 18463 8925 18475 8928
rect 18417 8919 18475 8925
rect 18509 8925 18521 8928
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 19518 8916 19524 8968
rect 19576 8956 19582 8968
rect 20165 8959 20223 8965
rect 20165 8956 20177 8959
rect 19576 8928 20177 8956
rect 19576 8916 19582 8928
rect 20165 8925 20177 8928
rect 20211 8925 20223 8959
rect 20165 8919 20223 8925
rect 20901 8959 20959 8965
rect 20901 8925 20913 8959
rect 20947 8956 20959 8959
rect 20993 8959 21051 8965
rect 20993 8956 21005 8959
rect 20947 8928 21005 8956
rect 20947 8925 20959 8928
rect 20901 8919 20959 8925
rect 20993 8925 21005 8928
rect 21039 8925 21051 8959
rect 20993 8919 21051 8925
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 18138 8888 18144 8900
rect 18012 8860 18144 8888
rect 18012 8848 18018 8860
rect 18138 8848 18144 8860
rect 18196 8888 18202 8900
rect 21450 8888 21456 8900
rect 18196 8860 21456 8888
rect 18196 8848 18202 8860
rect 21450 8848 21456 8860
rect 21508 8848 21514 8900
rect 21560 8888 21588 8996
rect 21821 8959 21879 8965
rect 21821 8925 21833 8959
rect 21867 8956 21879 8959
rect 21910 8956 21916 8968
rect 21867 8928 21916 8956
rect 21867 8925 21879 8928
rect 21821 8919 21879 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 22664 8956 22692 8996
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 23569 9027 23627 9033
rect 23308 8996 23520 9024
rect 23308 8956 23336 8996
rect 22664 8928 23336 8956
rect 23385 8959 23443 8965
rect 23385 8925 23397 8959
rect 23431 8925 23443 8959
rect 23492 8956 23520 8996
rect 23569 8993 23581 9027
rect 23615 9024 23627 9027
rect 24213 9027 24271 9033
rect 24213 9024 24225 9027
rect 23615 8996 24225 9024
rect 23615 8993 23627 8996
rect 23569 8987 23627 8993
rect 24213 8993 24225 8996
rect 24259 8993 24271 9027
rect 27522 9024 27528 9036
rect 24213 8987 24271 8993
rect 24320 8996 27528 9024
rect 24320 8956 24348 8996
rect 27522 8984 27528 8996
rect 27580 8984 27586 9036
rect 27614 8984 27620 9036
rect 27672 9024 27678 9036
rect 28997 9027 29055 9033
rect 28997 9024 29009 9027
rect 27672 8996 29009 9024
rect 27672 8984 27678 8996
rect 23492 8928 24348 8956
rect 23385 8919 23443 8925
rect 23290 8888 23296 8900
rect 21560 8860 23296 8888
rect 23290 8848 23296 8860
rect 23348 8848 23354 8900
rect 1486 8780 1492 8832
rect 1544 8820 1550 8832
rect 4614 8820 4620 8832
rect 1544 8792 4620 8820
rect 1544 8780 1550 8792
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5500 8792 5825 8820
rect 5500 8780 5506 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 17034 8820 17040 8832
rect 12584 8792 17040 8820
rect 12584 8780 12590 8792
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17218 8820 17224 8832
rect 17179 8792 17224 8820
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 19518 8820 19524 8832
rect 19479 8792 19524 8820
rect 19518 8780 19524 8792
rect 19576 8780 19582 8832
rect 20993 8823 21051 8829
rect 20993 8789 21005 8823
rect 21039 8820 21051 8823
rect 21637 8823 21695 8829
rect 21637 8820 21649 8823
rect 21039 8792 21649 8820
rect 21039 8789 21051 8792
rect 20993 8783 21051 8789
rect 21637 8789 21649 8792
rect 21683 8820 21695 8823
rect 21726 8820 21732 8832
rect 21683 8792 21732 8820
rect 21683 8789 21695 8792
rect 21637 8783 21695 8789
rect 21726 8780 21732 8792
rect 21784 8780 21790 8832
rect 21818 8780 21824 8832
rect 21876 8820 21882 8832
rect 22186 8820 22192 8832
rect 21876 8792 22192 8820
rect 21876 8780 21882 8792
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 23400 8820 23428 8919
rect 24394 8916 24400 8968
rect 24452 8956 24458 8968
rect 25774 8956 25780 8968
rect 24452 8928 25780 8956
rect 24452 8916 24458 8928
rect 25774 8916 25780 8928
rect 25832 8916 25838 8968
rect 26050 8956 26056 8968
rect 26011 8928 26056 8956
rect 26050 8916 26056 8928
rect 26108 8916 26114 8968
rect 27724 8965 27752 8996
rect 28997 8993 29009 8996
rect 29043 8993 29055 9027
rect 34146 9024 34152 9036
rect 28997 8987 29055 8993
rect 29104 8996 34152 9024
rect 26513 8959 26571 8965
rect 26513 8925 26525 8959
rect 26559 8925 26571 8959
rect 26513 8919 26571 8925
rect 27709 8959 27767 8965
rect 27709 8925 27721 8959
rect 27755 8925 27767 8959
rect 27709 8919 27767 8925
rect 27801 8959 27859 8965
rect 27801 8925 27813 8959
rect 27847 8956 27859 8959
rect 28074 8956 28080 8968
rect 27847 8928 28080 8956
rect 27847 8925 27859 8928
rect 27801 8919 27859 8925
rect 23658 8848 23664 8900
rect 23716 8888 23722 8900
rect 23716 8860 25360 8888
rect 23716 8848 23722 8860
rect 23753 8823 23811 8829
rect 23753 8820 23765 8823
rect 23400 8792 23765 8820
rect 23753 8789 23765 8792
rect 23799 8820 23811 8823
rect 23842 8820 23848 8832
rect 23799 8792 23848 8820
rect 23799 8789 23811 8792
rect 23753 8783 23811 8789
rect 23842 8780 23848 8792
rect 23900 8780 23906 8832
rect 24946 8780 24952 8832
rect 25004 8820 25010 8832
rect 25130 8820 25136 8832
rect 25004 8792 25136 8820
rect 25004 8780 25010 8792
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 25332 8820 25360 8860
rect 25498 8848 25504 8900
rect 25556 8888 25562 8900
rect 26142 8888 26148 8900
rect 25556 8860 26148 8888
rect 25556 8848 25562 8860
rect 26142 8848 26148 8860
rect 26200 8848 26206 8900
rect 26528 8888 26556 8919
rect 28074 8916 28080 8928
rect 28132 8916 28138 8968
rect 28169 8959 28227 8965
rect 28169 8925 28181 8959
rect 28215 8956 28227 8959
rect 28261 8959 28319 8965
rect 28261 8956 28273 8959
rect 28215 8928 28273 8956
rect 28215 8925 28227 8928
rect 28169 8919 28227 8925
rect 28261 8925 28273 8928
rect 28307 8925 28319 8959
rect 28261 8919 28319 8925
rect 28350 8916 28356 8968
rect 28408 8956 28414 8968
rect 29104 8956 29132 8996
rect 34146 8984 34152 8996
rect 34204 8984 34210 9036
rect 34256 9024 34284 9132
rect 34330 9120 34336 9172
rect 34388 9160 34394 9172
rect 34388 9132 38240 9160
rect 34388 9120 34394 9132
rect 34606 9052 34612 9104
rect 34664 9092 34670 9104
rect 38102 9092 38108 9104
rect 34664 9064 38108 9092
rect 34664 9052 34670 9064
rect 38102 9052 38108 9064
rect 38160 9052 38166 9104
rect 38212 9092 38240 9132
rect 38286 9120 38292 9172
rect 38344 9160 38350 9172
rect 38838 9160 38844 9172
rect 38344 9132 38844 9160
rect 38344 9120 38350 9132
rect 38838 9120 38844 9132
rect 38896 9120 38902 9172
rect 39206 9160 39212 9172
rect 39167 9132 39212 9160
rect 39206 9120 39212 9132
rect 39264 9120 39270 9172
rect 39574 9120 39580 9172
rect 39632 9160 39638 9172
rect 40494 9160 40500 9172
rect 39632 9132 40500 9160
rect 39632 9120 39638 9132
rect 40494 9120 40500 9132
rect 40552 9120 40558 9172
rect 40862 9120 40868 9172
rect 40920 9160 40926 9172
rect 41966 9160 41972 9172
rect 40920 9132 41972 9160
rect 40920 9120 40926 9132
rect 41966 9120 41972 9132
rect 42024 9120 42030 9172
rect 42426 9160 42432 9172
rect 42387 9132 42432 9160
rect 42426 9120 42432 9132
rect 42484 9120 42490 9172
rect 42610 9120 42616 9172
rect 42668 9160 42674 9172
rect 42668 9132 43116 9160
rect 42668 9120 42674 9132
rect 39850 9092 39856 9104
rect 38212 9064 39856 9092
rect 39850 9052 39856 9064
rect 39908 9052 39914 9104
rect 39942 9052 39948 9104
rect 40000 9092 40006 9104
rect 42978 9092 42984 9104
rect 40000 9064 42984 9092
rect 40000 9052 40006 9064
rect 42978 9052 42984 9064
rect 43036 9052 43042 9104
rect 43088 9092 43116 9132
rect 43346 9120 43352 9172
rect 43404 9160 43410 9172
rect 43717 9163 43775 9169
rect 43717 9160 43729 9163
rect 43404 9132 43729 9160
rect 43404 9120 43410 9132
rect 43717 9129 43729 9132
rect 43763 9160 43775 9163
rect 51626 9160 51632 9172
rect 43763 9132 51632 9160
rect 43763 9129 43775 9132
rect 43717 9123 43775 9129
rect 51626 9120 51632 9132
rect 51684 9120 51690 9172
rect 51905 9163 51963 9169
rect 51905 9129 51917 9163
rect 51951 9160 51963 9163
rect 52181 9163 52239 9169
rect 52181 9160 52193 9163
rect 51951 9132 52193 9160
rect 51951 9129 51963 9132
rect 51905 9123 51963 9129
rect 52181 9129 52193 9132
rect 52227 9160 52239 9163
rect 53650 9160 53656 9172
rect 52227 9132 53656 9160
rect 52227 9129 52239 9132
rect 52181 9123 52239 9129
rect 53650 9120 53656 9132
rect 53708 9120 53714 9172
rect 55122 9120 55128 9172
rect 55180 9160 55186 9172
rect 55861 9163 55919 9169
rect 55861 9160 55873 9163
rect 55180 9132 55873 9160
rect 55180 9120 55186 9132
rect 55861 9129 55873 9132
rect 55907 9129 55919 9163
rect 55861 9123 55919 9129
rect 55950 9120 55956 9172
rect 56008 9160 56014 9172
rect 57790 9160 57796 9172
rect 56008 9132 57796 9160
rect 56008 9120 56014 9132
rect 57790 9120 57796 9132
rect 57848 9120 57854 9172
rect 57885 9163 57943 9169
rect 57885 9129 57897 9163
rect 57931 9160 57943 9163
rect 57974 9160 57980 9172
rect 57931 9132 57980 9160
rect 57931 9129 57943 9132
rect 57885 9123 57943 9129
rect 57974 9120 57980 9132
rect 58032 9120 58038 9172
rect 58342 9120 58348 9172
rect 58400 9160 58406 9172
rect 58621 9163 58679 9169
rect 58621 9160 58633 9163
rect 58400 9132 58633 9160
rect 58400 9120 58406 9132
rect 58621 9129 58633 9132
rect 58667 9129 58679 9163
rect 58621 9123 58679 9129
rect 59265 9163 59323 9169
rect 59265 9129 59277 9163
rect 59311 9160 59323 9163
rect 59354 9160 59360 9172
rect 59311 9132 59360 9160
rect 59311 9129 59323 9132
rect 59265 9123 59323 9129
rect 59354 9120 59360 9132
rect 59412 9120 59418 9172
rect 59906 9160 59912 9172
rect 59867 9132 59912 9160
rect 59906 9120 59912 9132
rect 59964 9120 59970 9172
rect 60090 9120 60096 9172
rect 60148 9160 60154 9172
rect 61378 9160 61384 9172
rect 60148 9132 61384 9160
rect 60148 9120 60154 9132
rect 61378 9120 61384 9132
rect 61436 9120 61442 9172
rect 74350 9160 74356 9172
rect 74311 9132 74356 9160
rect 74350 9120 74356 9132
rect 74408 9120 74414 9172
rect 74442 9120 74448 9172
rect 74500 9160 74506 9172
rect 75365 9163 75423 9169
rect 75365 9160 75377 9163
rect 74500 9132 75377 9160
rect 74500 9120 74506 9132
rect 75365 9129 75377 9132
rect 75411 9129 75423 9163
rect 75365 9123 75423 9129
rect 76837 9163 76895 9169
rect 76837 9129 76849 9163
rect 76883 9160 76895 9163
rect 76926 9160 76932 9172
rect 76883 9132 76932 9160
rect 76883 9129 76895 9132
rect 76837 9123 76895 9129
rect 76926 9120 76932 9132
rect 76984 9120 76990 9172
rect 80606 9120 80612 9172
rect 80664 9160 80670 9172
rect 80701 9163 80759 9169
rect 80701 9160 80713 9163
rect 80664 9132 80713 9160
rect 80664 9120 80670 9132
rect 80701 9129 80713 9132
rect 80747 9129 80759 9163
rect 83182 9160 83188 9172
rect 83143 9132 83188 9160
rect 80701 9123 80759 9129
rect 83182 9120 83188 9132
rect 83240 9120 83246 9172
rect 85390 9120 85396 9172
rect 85448 9120 85454 9172
rect 86954 9160 86960 9172
rect 86915 9132 86960 9160
rect 86954 9120 86960 9132
rect 87012 9120 87018 9172
rect 92014 9120 92020 9172
rect 92072 9160 92078 9172
rect 92109 9163 92167 9169
rect 92109 9160 92121 9163
rect 92072 9132 92121 9160
rect 92072 9120 92078 9132
rect 92109 9129 92121 9132
rect 92155 9129 92167 9163
rect 92109 9123 92167 9129
rect 93946 9120 93952 9172
rect 94004 9160 94010 9172
rect 96798 9160 96804 9172
rect 94004 9132 96660 9160
rect 96759 9132 96804 9160
rect 94004 9120 94010 9132
rect 46934 9092 46940 9104
rect 43088 9064 46940 9092
rect 46934 9052 46940 9064
rect 46992 9052 46998 9104
rect 47118 9092 47124 9104
rect 47079 9064 47124 9092
rect 47118 9052 47124 9064
rect 47176 9052 47182 9104
rect 47302 9052 47308 9104
rect 47360 9092 47366 9104
rect 54113 9095 54171 9101
rect 54113 9092 54125 9095
rect 47360 9064 54125 9092
rect 47360 9052 47366 9064
rect 54113 9061 54125 9064
rect 54159 9061 54171 9095
rect 54846 9092 54852 9104
rect 54113 9055 54171 9061
rect 54220 9064 54852 9092
rect 34882 9024 34888 9036
rect 34256 8996 34888 9024
rect 34882 8984 34888 8996
rect 34940 8984 34946 9036
rect 34977 9027 35035 9033
rect 34977 8993 34989 9027
rect 35023 9024 35035 9027
rect 35066 9024 35072 9036
rect 35023 8996 35072 9024
rect 35023 8993 35035 8996
rect 34977 8987 35035 8993
rect 35066 8984 35072 8996
rect 35124 8984 35130 9036
rect 36630 9024 36636 9036
rect 35176 8996 36636 9024
rect 28408 8928 29132 8956
rect 28408 8916 28414 8928
rect 29178 8916 29184 8968
rect 29236 8956 29242 8968
rect 31846 8956 31852 8968
rect 29236 8928 31852 8956
rect 29236 8916 29242 8928
rect 31846 8916 31852 8928
rect 31904 8916 31910 8968
rect 31938 8916 31944 8968
rect 31996 8956 32002 8968
rect 35176 8956 35204 8996
rect 36630 8984 36636 8996
rect 36688 8984 36694 9036
rect 36814 9024 36820 9036
rect 36775 8996 36820 9024
rect 36814 8984 36820 8996
rect 36872 8984 36878 9036
rect 36998 9024 37004 9036
rect 36959 8996 37004 9024
rect 36998 8984 37004 8996
rect 37056 8984 37062 9036
rect 37274 8984 37280 9036
rect 37332 9024 37338 9036
rect 37332 8996 39896 9024
rect 37332 8984 37338 8996
rect 31996 8928 35204 8956
rect 31996 8916 32002 8928
rect 36446 8916 36452 8968
rect 36504 8956 36510 8968
rect 38105 8959 38163 8965
rect 38105 8956 38117 8959
rect 36504 8928 38117 8956
rect 36504 8916 36510 8928
rect 38105 8925 38117 8928
rect 38151 8925 38163 8959
rect 38105 8919 38163 8925
rect 38749 8959 38807 8965
rect 38749 8925 38761 8959
rect 38795 8956 38807 8959
rect 39022 8956 39028 8968
rect 38795 8928 39028 8956
rect 38795 8925 38807 8928
rect 38749 8919 38807 8925
rect 39022 8916 39028 8928
rect 39080 8916 39086 8968
rect 26881 8891 26939 8897
rect 26881 8888 26893 8891
rect 26528 8860 26893 8888
rect 26881 8857 26893 8860
rect 26927 8888 26939 8891
rect 39868 8888 39896 8996
rect 40126 8984 40132 9036
rect 40184 9024 40190 9036
rect 40405 9027 40463 9033
rect 40405 9024 40417 9027
rect 40184 8996 40417 9024
rect 40184 8984 40190 8996
rect 40405 8993 40417 8996
rect 40451 8993 40463 9027
rect 40405 8987 40463 8993
rect 40586 8984 40592 9036
rect 40644 9024 40650 9036
rect 41230 9024 41236 9036
rect 40644 8996 41236 9024
rect 40644 8984 40650 8996
rect 41230 8984 41236 8996
rect 41288 8984 41294 9036
rect 41506 8984 41512 9036
rect 41564 9024 41570 9036
rect 41874 9024 41880 9036
rect 41564 8996 41880 9024
rect 41564 8984 41570 8996
rect 41874 8984 41880 8996
rect 41932 8984 41938 9036
rect 41966 8984 41972 9036
rect 42024 9024 42030 9036
rect 46198 9024 46204 9036
rect 42024 8996 46204 9024
rect 42024 8984 42030 8996
rect 46198 8984 46204 8996
rect 46256 8984 46262 9036
rect 46385 9027 46443 9033
rect 46385 8993 46397 9027
rect 46431 9024 46443 9027
rect 46566 9024 46572 9036
rect 46431 8996 46572 9024
rect 46431 8993 46443 8996
rect 46385 8987 46443 8993
rect 46566 8984 46572 8996
rect 46624 9024 46630 9036
rect 47489 9027 47547 9033
rect 47489 9024 47501 9027
rect 46624 8996 47501 9024
rect 46624 8984 46630 8996
rect 47489 8993 47501 8996
rect 47535 8993 47547 9027
rect 47489 8987 47547 8993
rect 47946 8984 47952 9036
rect 48004 9024 48010 9036
rect 49050 9024 49056 9036
rect 48004 8996 49056 9024
rect 48004 8984 48010 8996
rect 49050 8984 49056 8996
rect 49108 8984 49114 9036
rect 50065 9027 50123 9033
rect 50065 8993 50077 9027
rect 50111 9024 50123 9027
rect 50706 9024 50712 9036
rect 50111 8996 50712 9024
rect 50111 8993 50123 8996
rect 50065 8987 50123 8993
rect 50706 8984 50712 8996
rect 50764 8984 50770 9036
rect 52641 9027 52699 9033
rect 52641 9024 52653 9027
rect 51368 8996 52653 9024
rect 39945 8959 40003 8965
rect 39945 8925 39957 8959
rect 39991 8956 40003 8959
rect 40313 8959 40371 8965
rect 40313 8956 40325 8959
rect 39991 8928 40325 8956
rect 39991 8925 40003 8928
rect 39945 8919 40003 8925
rect 40313 8925 40325 8928
rect 40359 8956 40371 8959
rect 40773 8959 40831 8965
rect 40359 8928 40724 8956
rect 40359 8925 40371 8928
rect 40313 8919 40371 8925
rect 40586 8888 40592 8900
rect 26927 8860 39804 8888
rect 39868 8860 40592 8888
rect 26927 8857 26939 8860
rect 26881 8851 26939 8857
rect 26602 8820 26608 8832
rect 25332 8792 26608 8820
rect 26602 8780 26608 8792
rect 26660 8780 26666 8832
rect 26970 8780 26976 8832
rect 27028 8820 27034 8832
rect 27249 8823 27307 8829
rect 27249 8820 27261 8823
rect 27028 8792 27261 8820
rect 27028 8780 27034 8792
rect 27249 8789 27261 8792
rect 27295 8820 27307 8823
rect 27522 8820 27528 8832
rect 27295 8792 27528 8820
rect 27295 8789 27307 8792
rect 27249 8783 27307 8789
rect 27522 8780 27528 8792
rect 27580 8780 27586 8832
rect 27614 8780 27620 8832
rect 27672 8820 27678 8832
rect 33502 8820 33508 8832
rect 27672 8792 33508 8820
rect 27672 8780 27678 8792
rect 33502 8780 33508 8792
rect 33560 8780 33566 8832
rect 33965 8823 34023 8829
rect 33965 8789 33977 8823
rect 34011 8820 34023 8823
rect 34790 8820 34796 8832
rect 34011 8792 34796 8820
rect 34011 8789 34023 8792
rect 33965 8783 34023 8789
rect 34790 8780 34796 8792
rect 34848 8780 34854 8832
rect 34882 8780 34888 8832
rect 34940 8820 34946 8832
rect 38930 8820 38936 8832
rect 34940 8792 38936 8820
rect 34940 8780 34946 8792
rect 38930 8780 38936 8792
rect 38988 8780 38994 8832
rect 39776 8820 39804 8860
rect 40586 8848 40592 8860
rect 40644 8848 40650 8900
rect 40696 8888 40724 8928
rect 40773 8925 40785 8959
rect 40819 8956 40831 8959
rect 41141 8959 41199 8965
rect 41141 8956 41153 8959
rect 40819 8928 41153 8956
rect 40819 8925 40831 8928
rect 40773 8919 40831 8925
rect 41141 8925 41153 8928
rect 41187 8956 41199 8959
rect 41187 8928 41552 8956
rect 41187 8925 41199 8928
rect 41141 8919 41199 8925
rect 41230 8888 41236 8900
rect 40696 8860 41236 8888
rect 41230 8848 41236 8860
rect 41288 8848 41294 8900
rect 41524 8888 41552 8928
rect 41598 8916 41604 8968
rect 41656 8956 41662 8968
rect 42794 8956 42800 8968
rect 41656 8928 42288 8956
rect 41656 8916 41662 8928
rect 42058 8888 42064 8900
rect 41524 8860 42064 8888
rect 42058 8848 42064 8860
rect 42116 8848 42122 8900
rect 40310 8820 40316 8832
rect 39776 8792 40316 8820
rect 40310 8780 40316 8792
rect 40368 8780 40374 8832
rect 41509 8823 41567 8829
rect 41509 8789 41521 8823
rect 41555 8820 41567 8823
rect 42150 8820 42156 8832
rect 41555 8792 42156 8820
rect 41555 8789 41567 8792
rect 41509 8783 41567 8789
rect 42150 8780 42156 8792
rect 42208 8780 42214 8832
rect 42260 8820 42288 8928
rect 42536 8928 42800 8956
rect 42426 8848 42432 8900
rect 42484 8888 42490 8900
rect 42536 8888 42564 8928
rect 42794 8916 42800 8928
rect 42852 8916 42858 8968
rect 42886 8916 42892 8968
rect 42944 8956 42950 8968
rect 42981 8959 43039 8965
rect 42981 8956 42993 8959
rect 42944 8928 42993 8956
rect 42944 8916 42950 8928
rect 42981 8925 42993 8928
rect 43027 8925 43039 8959
rect 43346 8956 43352 8968
rect 43307 8928 43352 8956
rect 42981 8919 43039 8925
rect 43346 8916 43352 8928
rect 43404 8916 43410 8968
rect 46658 8956 46664 8968
rect 43456 8928 46664 8956
rect 42484 8860 42564 8888
rect 42484 8848 42490 8860
rect 43456 8820 43484 8928
rect 46658 8916 46664 8928
rect 46716 8916 46722 8968
rect 47026 8916 47032 8968
rect 47084 8956 47090 8968
rect 51368 8965 51396 8996
rect 52641 8993 52653 8996
rect 52687 8993 52699 9027
rect 52641 8987 52699 8993
rect 53190 8984 53196 9036
rect 53248 9024 53254 9036
rect 53561 9027 53619 9033
rect 53561 9024 53573 9027
rect 53248 8996 53573 9024
rect 53248 8984 53254 8996
rect 53561 8993 53573 8996
rect 53607 9024 53619 9027
rect 54220 9024 54248 9064
rect 54846 9052 54852 9064
rect 54904 9052 54910 9104
rect 55033 9095 55091 9101
rect 55033 9061 55045 9095
rect 55079 9092 55091 9095
rect 60734 9092 60740 9104
rect 55079 9064 60740 9092
rect 55079 9061 55091 9064
rect 55033 9055 55091 9061
rect 54662 9024 54668 9036
rect 53607 8996 54248 9024
rect 54312 8996 54668 9024
rect 53607 8993 53619 8996
rect 53561 8987 53619 8993
rect 50801 8959 50859 8965
rect 50801 8956 50813 8959
rect 47084 8928 50813 8956
rect 47084 8916 47090 8928
rect 50801 8925 50813 8928
rect 50847 8925 50859 8959
rect 50801 8919 50859 8925
rect 50985 8959 51043 8965
rect 50985 8925 50997 8959
rect 51031 8956 51043 8959
rect 51353 8959 51411 8965
rect 51353 8956 51365 8959
rect 51031 8928 51365 8956
rect 51031 8925 51043 8928
rect 50985 8919 51043 8925
rect 51353 8925 51365 8928
rect 51399 8925 51411 8959
rect 51353 8919 51411 8925
rect 51445 8959 51503 8965
rect 51445 8925 51457 8959
rect 51491 8925 51503 8959
rect 51445 8919 51503 8925
rect 51813 8959 51871 8965
rect 51813 8925 51825 8959
rect 51859 8956 51871 8959
rect 51905 8959 51963 8965
rect 51905 8956 51917 8959
rect 51859 8928 51917 8956
rect 51859 8925 51871 8928
rect 51813 8919 51871 8925
rect 51905 8925 51917 8928
rect 51951 8925 51963 8959
rect 51905 8919 51963 8925
rect 43898 8848 43904 8900
rect 43956 8888 43962 8900
rect 48130 8888 48136 8900
rect 43956 8860 48136 8888
rect 43956 8848 43962 8860
rect 48130 8848 48136 8860
rect 48188 8848 48194 8900
rect 48222 8848 48228 8900
rect 48280 8888 48286 8900
rect 48280 8860 48544 8888
rect 48280 8848 48286 8860
rect 42260 8792 43484 8820
rect 43530 8780 43536 8832
rect 43588 8820 43594 8832
rect 48038 8820 48044 8832
rect 43588 8792 48044 8820
rect 43588 8780 43594 8792
rect 48038 8780 48044 8792
rect 48096 8780 48102 8832
rect 48406 8820 48412 8832
rect 48367 8792 48412 8820
rect 48406 8780 48412 8792
rect 48464 8780 48470 8832
rect 48516 8820 48544 8860
rect 48682 8848 48688 8900
rect 48740 8888 48746 8900
rect 51460 8888 51488 8919
rect 52086 8916 52092 8968
rect 52144 8956 52150 8968
rect 52549 8959 52607 8965
rect 52549 8956 52561 8959
rect 52144 8928 52561 8956
rect 52144 8916 52150 8928
rect 52549 8925 52561 8928
rect 52595 8956 52607 8959
rect 54110 8956 54116 8968
rect 52595 8928 54116 8956
rect 52595 8925 52607 8928
rect 52549 8919 52607 8925
rect 54110 8916 54116 8928
rect 54168 8916 54174 8968
rect 54312 8965 54340 8996
rect 54662 8984 54668 8996
rect 54720 8984 54726 9036
rect 54297 8959 54355 8965
rect 54297 8925 54309 8959
rect 54343 8925 54355 8959
rect 54297 8919 54355 8925
rect 54757 8959 54815 8965
rect 54757 8925 54769 8959
rect 54803 8956 54815 8959
rect 55048 8956 55076 9055
rect 60734 9052 60740 9064
rect 60792 9052 60798 9104
rect 62758 9052 62764 9104
rect 62816 9092 62822 9104
rect 63221 9095 63279 9101
rect 63221 9092 63233 9095
rect 62816 9064 63233 9092
rect 62816 9052 62822 9064
rect 63221 9061 63233 9064
rect 63267 9061 63279 9095
rect 63221 9055 63279 9061
rect 82449 9095 82507 9101
rect 82449 9061 82461 9095
rect 82495 9092 82507 9095
rect 83458 9092 83464 9104
rect 82495 9064 83464 9092
rect 82495 9061 82507 9064
rect 82449 9055 82507 9061
rect 83458 9052 83464 9064
rect 83516 9052 83522 9104
rect 85408 9092 85436 9120
rect 85408 9064 88564 9092
rect 55585 9027 55643 9033
rect 55585 8993 55597 9027
rect 55631 9024 55643 9027
rect 55858 9024 55864 9036
rect 55631 8996 55864 9024
rect 55631 8993 55643 8996
rect 55585 8987 55643 8993
rect 55858 8984 55864 8996
rect 55916 8984 55922 9036
rect 56134 8984 56140 9036
rect 56192 9024 56198 9036
rect 57333 9027 57391 9033
rect 57333 9024 57345 9027
rect 56192 8996 56916 9024
rect 56192 8984 56198 8996
rect 54803 8928 55076 8956
rect 54803 8925 54815 8928
rect 54757 8919 54815 8925
rect 55490 8916 55496 8968
rect 55548 8956 55554 8968
rect 56229 8959 56287 8965
rect 56229 8956 56241 8959
rect 55548 8928 56241 8956
rect 55548 8916 55554 8928
rect 56229 8925 56241 8928
rect 56275 8956 56287 8959
rect 56502 8956 56508 8968
rect 56275 8928 56508 8956
rect 56275 8925 56287 8928
rect 56229 8919 56287 8925
rect 56502 8916 56508 8928
rect 56560 8916 56566 8968
rect 56597 8959 56655 8965
rect 56597 8925 56609 8959
rect 56643 8956 56655 8959
rect 56778 8956 56784 8968
rect 56643 8928 56784 8956
rect 56643 8925 56655 8928
rect 56597 8919 56655 8925
rect 56778 8916 56784 8928
rect 56836 8916 56842 8968
rect 48740 8860 51488 8888
rect 48740 8848 48746 8860
rect 51534 8848 51540 8900
rect 51592 8888 51598 8900
rect 51592 8860 52500 8888
rect 51592 8848 51598 8860
rect 50154 8820 50160 8832
rect 48516 8792 50160 8820
rect 50154 8780 50160 8792
rect 50212 8780 50218 8832
rect 50522 8820 50528 8832
rect 50483 8792 50528 8820
rect 50522 8780 50528 8792
rect 50580 8780 50586 8832
rect 50801 8823 50859 8829
rect 50801 8789 50813 8823
rect 50847 8820 50859 8823
rect 52362 8820 52368 8832
rect 50847 8792 52368 8820
rect 50847 8789 50859 8792
rect 50801 8783 50859 8789
rect 52362 8780 52368 8792
rect 52420 8780 52426 8832
rect 52472 8820 52500 8860
rect 53282 8848 53288 8900
rect 53340 8888 53346 8900
rect 55766 8888 55772 8900
rect 53340 8860 55772 8888
rect 53340 8848 53346 8860
rect 55766 8848 55772 8860
rect 55824 8848 55830 8900
rect 55858 8848 55864 8900
rect 55916 8888 55922 8900
rect 56318 8888 56324 8900
rect 55916 8860 56324 8888
rect 55916 8848 55922 8860
rect 56318 8848 56324 8860
rect 56376 8848 56382 8900
rect 56888 8888 56916 8996
rect 56980 8996 57345 9024
rect 56980 8965 57008 8996
rect 57333 8993 57345 8996
rect 57379 9024 57391 9027
rect 58621 9027 58679 9033
rect 57379 8996 58480 9024
rect 57379 8993 57391 8996
rect 57333 8987 57391 8993
rect 56965 8959 57023 8965
rect 56965 8925 56977 8959
rect 57011 8925 57023 8959
rect 57606 8956 57612 8968
rect 56965 8919 57023 8925
rect 57072 8928 57612 8956
rect 57072 8888 57100 8928
rect 57606 8916 57612 8928
rect 57664 8916 57670 8968
rect 58069 8959 58127 8965
rect 58069 8925 58081 8959
rect 58115 8925 58127 8959
rect 58342 8956 58348 8968
rect 58303 8928 58348 8956
rect 58069 8919 58127 8925
rect 56888 8860 57100 8888
rect 57701 8891 57759 8897
rect 57701 8857 57713 8891
rect 57747 8888 57759 8891
rect 58084 8888 58112 8919
rect 58342 8916 58348 8928
rect 58400 8916 58406 8968
rect 58452 8956 58480 8996
rect 58621 8993 58633 9027
rect 58667 9024 58679 9027
rect 58897 9027 58955 9033
rect 58897 9024 58909 9027
rect 58667 8996 58909 9024
rect 58667 8993 58679 8996
rect 58621 8987 58679 8993
rect 58897 8993 58909 8996
rect 58943 9024 58955 9027
rect 61562 9024 61568 9036
rect 58943 8996 61568 9024
rect 58943 8993 58955 8996
rect 58897 8987 58955 8993
rect 61562 8984 61568 8996
rect 61620 8984 61626 9036
rect 63310 8984 63316 9036
rect 63368 9024 63374 9036
rect 64141 9027 64199 9033
rect 64141 9024 64153 9027
rect 63368 8996 64153 9024
rect 63368 8984 63374 8996
rect 60918 8956 60924 8968
rect 58452 8928 60924 8956
rect 60918 8916 60924 8928
rect 60976 8916 60982 8968
rect 61378 8916 61384 8968
rect 61436 8956 61442 8968
rect 63037 8959 63095 8965
rect 61436 8928 61608 8956
rect 61436 8916 61442 8928
rect 61473 8891 61531 8897
rect 61473 8888 61485 8891
rect 57747 8860 61485 8888
rect 57747 8857 57759 8860
rect 57701 8851 57759 8857
rect 61473 8857 61485 8860
rect 61519 8857 61531 8891
rect 61580 8888 61608 8928
rect 63037 8925 63049 8959
rect 63083 8956 63095 8959
rect 63402 8956 63408 8968
rect 63083 8928 63408 8956
rect 63083 8925 63095 8928
rect 63037 8919 63095 8925
rect 63402 8916 63408 8928
rect 63460 8916 63466 8968
rect 63696 8965 63724 8996
rect 64141 8993 64153 8996
rect 64187 8993 64199 9027
rect 64141 8987 64199 8993
rect 71869 9027 71927 9033
rect 71869 8993 71881 9027
rect 71915 9024 71927 9027
rect 72418 9024 72424 9036
rect 71915 8996 72424 9024
rect 71915 8993 71927 8996
rect 71869 8987 71927 8993
rect 72418 8984 72424 8996
rect 72476 8984 72482 9036
rect 72881 9027 72939 9033
rect 72881 8993 72893 9027
rect 72927 9024 72939 9027
rect 73614 9024 73620 9036
rect 72927 8996 73620 9024
rect 72927 8993 72939 8996
rect 72881 8987 72939 8993
rect 73614 8984 73620 8996
rect 73672 8984 73678 9036
rect 73893 9027 73951 9033
rect 73893 8993 73905 9027
rect 73939 9024 73951 9027
rect 74810 9024 74816 9036
rect 73939 8996 74816 9024
rect 73939 8993 73951 8996
rect 73893 8987 73951 8993
rect 74810 8984 74816 8996
rect 74868 8984 74874 9036
rect 74905 9027 74963 9033
rect 74905 8993 74917 9027
rect 74951 9024 74963 9027
rect 76006 9024 76012 9036
rect 74951 8996 76012 9024
rect 74951 8993 74963 8996
rect 74905 8987 74963 8993
rect 76006 8984 76012 8996
rect 76064 8984 76070 9036
rect 76282 9024 76288 9036
rect 76243 8996 76288 9024
rect 76282 8984 76288 8996
rect 76340 8984 76346 9036
rect 80054 8984 80060 9036
rect 80112 9024 80118 9036
rect 82817 9027 82875 9033
rect 82817 9024 82829 9027
rect 80112 8996 80157 9024
rect 81912 8996 82829 9024
rect 80112 8984 80118 8996
rect 81912 8965 81940 8996
rect 82817 8993 82829 8996
rect 82863 9024 82875 9027
rect 84286 9024 84292 9036
rect 82863 8996 84292 9024
rect 82863 8993 82875 8996
rect 82817 8987 82875 8993
rect 84286 8984 84292 8996
rect 84344 8984 84350 9036
rect 85393 9027 85451 9033
rect 85393 8993 85405 9027
rect 85439 9024 85451 9027
rect 87230 9024 87236 9036
rect 85439 8996 87236 9024
rect 85439 8993 85451 8996
rect 85393 8987 85451 8993
rect 87230 8984 87236 8996
rect 87288 8984 87294 9036
rect 88536 9033 88564 9064
rect 89806 9052 89812 9104
rect 89864 9092 89870 9104
rect 96632 9092 96660 9132
rect 96798 9120 96804 9132
rect 96856 9120 96862 9172
rect 98178 9160 98184 9172
rect 98139 9132 98184 9160
rect 98178 9120 98184 9132
rect 98236 9120 98242 9172
rect 99742 9120 99748 9172
rect 99800 9160 99806 9172
rect 99800 9132 99880 9160
rect 99800 9120 99806 9132
rect 89864 9064 95372 9092
rect 96632 9064 99788 9092
rect 89864 9052 89870 9064
rect 88521 9027 88579 9033
rect 88521 8993 88533 9027
rect 88567 8993 88579 9027
rect 90913 9027 90971 9033
rect 90913 9024 90925 9027
rect 88521 8987 88579 8993
rect 88996 8996 90925 9024
rect 63681 8959 63739 8965
rect 63681 8925 63693 8959
rect 63727 8925 63739 8959
rect 63681 8919 63739 8925
rect 81897 8959 81955 8965
rect 81897 8925 81909 8959
rect 81943 8925 81955 8959
rect 87509 8959 87567 8965
rect 87509 8956 87521 8959
rect 81897 8919 81955 8925
rect 87248 8928 87521 8956
rect 67358 8888 67364 8900
rect 61580 8860 67364 8888
rect 61473 8851 61531 8857
rect 67358 8848 67364 8860
rect 67416 8848 67422 8900
rect 81986 8888 81992 8900
rect 81947 8860 81992 8888
rect 81986 8848 81992 8860
rect 82044 8848 82050 8900
rect 87248 8897 87276 8928
rect 87509 8925 87521 8928
rect 87555 8925 87567 8959
rect 87509 8919 87567 8925
rect 86405 8891 86463 8897
rect 86405 8857 86417 8891
rect 86451 8888 86463 8891
rect 87233 8891 87291 8897
rect 87233 8888 87245 8891
rect 86451 8860 87245 8888
rect 86451 8857 86463 8860
rect 86405 8851 86463 8857
rect 87233 8857 87245 8860
rect 87279 8857 87291 8891
rect 87233 8851 87291 8857
rect 59170 8820 59176 8832
rect 52472 8792 59176 8820
rect 59170 8780 59176 8792
rect 59228 8780 59234 8832
rect 59446 8820 59452 8832
rect 59407 8792 59452 8820
rect 59446 8780 59452 8792
rect 59504 8780 59510 8832
rect 60182 8780 60188 8832
rect 60240 8820 60246 8832
rect 60461 8823 60519 8829
rect 60461 8820 60473 8823
rect 60240 8792 60473 8820
rect 60240 8780 60246 8792
rect 60461 8789 60473 8792
rect 60507 8789 60519 8823
rect 60461 8783 60519 8789
rect 60642 8780 60648 8832
rect 60700 8820 60706 8832
rect 64782 8820 64788 8832
rect 60700 8792 64788 8820
rect 60700 8780 60706 8792
rect 64782 8780 64788 8792
rect 64840 8780 64846 8832
rect 86126 8780 86132 8832
rect 86184 8820 86190 8832
rect 88996 8820 89024 8996
rect 90913 8993 90925 8996
rect 90959 8993 90971 9027
rect 93118 9024 93124 9036
rect 93079 8996 93124 9024
rect 90913 8987 90971 8993
rect 93118 8984 93124 8996
rect 93176 8984 93182 9036
rect 95344 9033 95372 9064
rect 95329 9027 95387 9033
rect 95329 8993 95341 9027
rect 95375 8993 95387 9027
rect 95329 8987 95387 8993
rect 97813 9027 97871 9033
rect 97813 8993 97825 9027
rect 97859 9024 97871 9027
rect 97902 9024 97908 9036
rect 97859 8996 97908 9024
rect 97859 8993 97871 8996
rect 97813 8987 97871 8993
rect 97902 8984 97908 8996
rect 97960 9024 97966 9036
rect 99558 9024 99564 9036
rect 97960 8996 99564 9024
rect 97960 8984 97966 8996
rect 99558 8984 99564 8996
rect 99616 8984 99622 9036
rect 99760 9033 99788 9064
rect 99745 9027 99803 9033
rect 99745 8993 99757 9027
rect 99791 8993 99803 9027
rect 99852 9024 99880 9132
rect 99926 9120 99932 9172
rect 99984 9160 99990 9172
rect 108114 9160 108120 9172
rect 99984 9132 108120 9160
rect 99984 9120 99990 9132
rect 108114 9120 108120 9132
rect 108172 9120 108178 9172
rect 108209 9163 108267 9169
rect 108209 9129 108221 9163
rect 108255 9160 108267 9163
rect 108298 9160 108304 9172
rect 108255 9132 108304 9160
rect 108255 9129 108267 9132
rect 108209 9123 108267 9129
rect 108298 9120 108304 9132
rect 108356 9120 108362 9172
rect 120997 9163 121055 9169
rect 120997 9129 121009 9163
rect 121043 9160 121055 9163
rect 121454 9160 121460 9172
rect 121043 9132 121460 9160
rect 121043 9129 121055 9132
rect 120997 9123 121055 9129
rect 121454 9120 121460 9132
rect 121512 9120 121518 9172
rect 124582 9160 124588 9172
rect 124543 9132 124588 9160
rect 124582 9120 124588 9132
rect 124640 9120 124646 9172
rect 127066 9160 127072 9172
rect 127027 9132 127072 9160
rect 127066 9120 127072 9132
rect 127124 9120 127130 9172
rect 133966 9120 133972 9172
rect 134024 9160 134030 9172
rect 143350 9160 143356 9172
rect 134024 9132 143356 9160
rect 134024 9120 134030 9132
rect 143350 9120 143356 9132
rect 143408 9120 143414 9172
rect 143442 9120 143448 9172
rect 143500 9160 143506 9172
rect 145650 9160 145656 9172
rect 143500 9132 145656 9160
rect 143500 9120 143506 9132
rect 145650 9120 145656 9132
rect 145708 9120 145714 9172
rect 145926 9160 145932 9172
rect 145887 9132 145932 9160
rect 145926 9120 145932 9132
rect 145984 9120 145990 9172
rect 146110 9120 146116 9172
rect 146168 9160 146174 9172
rect 154393 9163 154451 9169
rect 146168 9132 152136 9160
rect 146168 9120 146174 9132
rect 100110 9052 100116 9104
rect 100168 9092 100174 9104
rect 100570 9092 100576 9104
rect 100168 9064 100576 9092
rect 100168 9052 100174 9064
rect 100570 9052 100576 9064
rect 100628 9052 100634 9104
rect 101950 9052 101956 9104
rect 102008 9092 102014 9104
rect 109313 9095 109371 9101
rect 102008 9064 106688 9092
rect 102008 9052 102014 9064
rect 104345 9027 104403 9033
rect 104345 9024 104357 9027
rect 99852 8996 104357 9024
rect 99745 8987 99803 8993
rect 104345 8993 104357 8996
rect 104391 8993 104403 9027
rect 104345 8987 104403 8993
rect 105354 8984 105360 9036
rect 105412 9024 105418 9036
rect 106550 9024 106556 9036
rect 105412 8996 106556 9024
rect 105412 8984 105418 8996
rect 106550 8984 106556 8996
rect 106608 8984 106614 9036
rect 89073 8959 89131 8965
rect 89073 8925 89085 8959
rect 89119 8925 89131 8959
rect 89898 8956 89904 8968
rect 89859 8928 89904 8956
rect 89073 8919 89131 8925
rect 86184 8792 89024 8820
rect 89088 8820 89116 8919
rect 89898 8916 89904 8928
rect 89956 8916 89962 8968
rect 91465 8959 91523 8965
rect 91465 8925 91477 8959
rect 91511 8956 91523 8959
rect 94314 8956 94320 8968
rect 91511 8928 91876 8956
rect 94275 8928 94320 8956
rect 91511 8925 91523 8928
rect 91465 8919 91523 8925
rect 89441 8823 89499 8829
rect 89441 8820 89453 8823
rect 89088 8792 89453 8820
rect 86184 8780 86190 8792
rect 89441 8789 89453 8792
rect 89487 8820 89499 8823
rect 89530 8820 89536 8832
rect 89487 8792 89536 8820
rect 89487 8789 89499 8792
rect 89441 8783 89499 8789
rect 89530 8780 89536 8792
rect 89588 8780 89594 8832
rect 91848 8829 91876 8928
rect 94314 8916 94320 8928
rect 94372 8916 94378 8968
rect 95881 8959 95939 8965
rect 95881 8925 95893 8959
rect 95927 8925 95939 8959
rect 95881 8919 95939 8925
rect 96709 8959 96767 8965
rect 96709 8925 96721 8959
rect 96755 8956 96767 8959
rect 98549 8959 98607 8965
rect 96755 8928 97304 8956
rect 96755 8925 96767 8928
rect 96709 8919 96767 8925
rect 91833 8823 91891 8829
rect 91833 8789 91845 8823
rect 91879 8820 91891 8823
rect 92014 8820 92020 8832
rect 91879 8792 92020 8820
rect 91879 8789 91891 8792
rect 91833 8783 91891 8789
rect 92014 8780 92020 8792
rect 92072 8780 92078 8832
rect 92750 8820 92756 8832
rect 92711 8792 92756 8820
rect 92750 8780 92756 8792
rect 92808 8780 92814 8832
rect 95896 8820 95924 8919
rect 97276 8832 97304 8928
rect 98549 8925 98561 8959
rect 98595 8956 98607 8959
rect 98733 8959 98791 8965
rect 98733 8956 98745 8959
rect 98595 8928 98745 8956
rect 98595 8925 98607 8928
rect 98549 8919 98607 8925
rect 98733 8925 98745 8928
rect 98779 8925 98791 8959
rect 98733 8919 98791 8925
rect 98748 8888 98776 8919
rect 99006 8916 99012 8968
rect 99064 8956 99070 8968
rect 99650 8956 99656 8968
rect 99064 8928 99656 8956
rect 99064 8916 99070 8928
rect 99650 8916 99656 8928
rect 99708 8916 99714 8968
rect 100297 8959 100355 8965
rect 100297 8925 100309 8959
rect 100343 8956 100355 8959
rect 100478 8956 100484 8968
rect 100343 8928 100484 8956
rect 100343 8925 100355 8928
rect 100297 8919 100355 8925
rect 100478 8916 100484 8928
rect 100536 8916 100542 8968
rect 100570 8916 100576 8968
rect 100628 8956 100634 8968
rect 103974 8956 103980 8968
rect 100628 8928 103980 8956
rect 100628 8916 100634 8928
rect 103974 8916 103980 8928
rect 104032 8916 104038 8968
rect 106660 8956 106688 9064
rect 109313 9061 109325 9095
rect 109359 9092 109371 9095
rect 109359 9064 115428 9092
rect 109359 9061 109371 9064
rect 109313 9055 109371 9061
rect 107841 9027 107899 9033
rect 107841 8993 107853 9027
rect 107887 9024 107899 9027
rect 108209 9027 108267 9033
rect 108209 9024 108221 9027
rect 107887 8996 108221 9024
rect 107887 8993 107899 8996
rect 107841 8987 107899 8993
rect 108209 8993 108221 8996
rect 108255 8993 108267 9027
rect 112254 9024 112260 9036
rect 112215 8996 112260 9024
rect 108209 8987 108267 8993
rect 112254 8984 112260 8996
rect 112312 8984 112318 9036
rect 113910 9024 113916 9036
rect 113871 8996 113916 9024
rect 113910 8984 113916 8996
rect 113968 9024 113974 9036
rect 114373 9027 114431 9033
rect 114373 9024 114385 9027
rect 113968 8996 114385 9024
rect 113968 8984 113974 8996
rect 114373 8993 114385 8996
rect 114419 8993 114431 9027
rect 114373 8987 114431 8993
rect 115290 8956 115296 8968
rect 106660 8928 115296 8956
rect 115290 8916 115296 8928
rect 115348 8916 115354 8968
rect 115400 8956 115428 9064
rect 116688 9064 118740 9092
rect 115566 9024 115572 9036
rect 115527 8996 115572 9024
rect 115566 8984 115572 8996
rect 115624 8984 115630 9036
rect 115658 8984 115664 9036
rect 115716 9024 115722 9036
rect 116581 9027 116639 9033
rect 116581 9024 116593 9027
rect 115716 8996 116593 9024
rect 115716 8984 115722 8996
rect 116581 8993 116593 8996
rect 116627 8993 116639 9027
rect 116581 8987 116639 8993
rect 116688 8956 116716 9064
rect 118712 9024 118740 9064
rect 120718 9052 120724 9104
rect 120776 9092 120782 9104
rect 122929 9095 122987 9101
rect 122929 9092 122941 9095
rect 120776 9064 122941 9092
rect 120776 9052 120782 9064
rect 122929 9061 122941 9064
rect 122975 9061 122987 9095
rect 122929 9055 122987 9061
rect 123205 9095 123263 9101
rect 123205 9061 123217 9095
rect 123251 9092 123263 9095
rect 123251 9064 124720 9092
rect 123251 9061 123263 9064
rect 123205 9055 123263 9061
rect 119154 9024 119160 9036
rect 118712 8996 119160 9024
rect 119154 8984 119160 8996
rect 119212 8984 119218 9036
rect 119430 8984 119436 9036
rect 119488 9024 119494 9036
rect 122285 9027 122343 9033
rect 122285 9024 122297 9027
rect 119488 8996 122297 9024
rect 119488 8984 119494 8996
rect 122285 8993 122297 8996
rect 122331 8993 122343 9027
rect 123220 9024 123248 9055
rect 122285 8987 122343 8993
rect 122576 8996 123248 9024
rect 124125 9027 124183 9033
rect 115400 8928 116716 8956
rect 117133 8959 117191 8965
rect 117133 8925 117145 8959
rect 117179 8956 117191 8959
rect 117498 8956 117504 8968
rect 117179 8928 117504 8956
rect 117179 8925 117191 8928
rect 117133 8919 117191 8925
rect 117498 8916 117504 8928
rect 117556 8916 117562 8968
rect 118786 8956 118792 8968
rect 118747 8928 118792 8956
rect 118786 8916 118792 8928
rect 118844 8956 118850 8968
rect 119249 8959 119307 8965
rect 119249 8956 119261 8959
rect 118844 8928 119261 8956
rect 118844 8916 118850 8928
rect 119249 8925 119261 8928
rect 119295 8925 119307 8959
rect 121270 8956 121276 8968
rect 121231 8928 121276 8956
rect 119249 8919 119307 8925
rect 121270 8916 121276 8928
rect 121328 8916 121334 8968
rect 122576 8965 122604 8996
rect 124125 8993 124137 9027
rect 124171 9024 124183 9027
rect 124582 9024 124588 9036
rect 124171 8996 124588 9024
rect 124171 8993 124183 8996
rect 124125 8987 124183 8993
rect 124582 8984 124588 8996
rect 124640 8984 124646 9036
rect 124692 9024 124720 9064
rect 124766 9052 124772 9104
rect 124824 9092 124830 9104
rect 130746 9092 130752 9104
rect 124824 9064 130752 9092
rect 124824 9052 124830 9064
rect 130746 9052 130752 9064
rect 130804 9052 130810 9104
rect 136174 9052 136180 9104
rect 136232 9092 136238 9104
rect 147766 9092 147772 9104
rect 136232 9064 147772 9092
rect 136232 9052 136238 9064
rect 147766 9052 147772 9064
rect 147824 9052 147830 9104
rect 147950 9092 147956 9104
rect 147911 9064 147956 9092
rect 147950 9052 147956 9064
rect 148008 9052 148014 9104
rect 150805 9095 150863 9101
rect 148060 9064 149468 9092
rect 125778 9024 125784 9036
rect 124692 8996 125784 9024
rect 125778 8984 125784 8996
rect 125836 8984 125842 9036
rect 127526 9024 127532 9036
rect 127487 8996 127532 9024
rect 127526 8984 127532 8996
rect 127584 8984 127590 9036
rect 128541 9027 128599 9033
rect 128541 8993 128553 9027
rect 128587 8993 128599 9027
rect 129461 9027 129519 9033
rect 129461 9024 129473 9027
rect 128541 8987 128599 8993
rect 129108 8996 129473 9024
rect 122561 8959 122619 8965
rect 122561 8925 122573 8959
rect 122607 8925 122619 8959
rect 122561 8919 122619 8925
rect 122929 8959 122987 8965
rect 122929 8925 122941 8959
rect 122975 8956 122987 8959
rect 128556 8956 128584 8987
rect 129108 8965 129136 8996
rect 129461 8993 129473 8996
rect 129507 9024 129519 9027
rect 130286 9024 130292 9036
rect 129507 8996 130292 9024
rect 129507 8993 129519 8996
rect 129461 8987 129519 8993
rect 130286 8984 130292 8996
rect 130344 8984 130350 9036
rect 131114 9024 131120 9036
rect 131075 8996 131120 9024
rect 131114 8984 131120 8996
rect 131172 8984 131178 9036
rect 138014 8984 138020 9036
rect 138072 9024 138078 9036
rect 139029 9027 139087 9033
rect 138072 8996 138117 9024
rect 138072 8984 138078 8996
rect 139029 8993 139041 9027
rect 139075 9024 139087 9027
rect 140406 9024 140412 9036
rect 139075 8996 140412 9024
rect 139075 8993 139087 8996
rect 139029 8987 139087 8993
rect 140406 8984 140412 8996
rect 140464 8984 140470 9036
rect 142525 9027 142583 9033
rect 140976 8996 142476 9024
rect 122975 8928 128584 8956
rect 129093 8959 129151 8965
rect 122975 8925 122987 8928
rect 122929 8919 122987 8925
rect 129093 8925 129105 8959
rect 129139 8925 129151 8959
rect 129921 8959 129979 8965
rect 129921 8956 129933 8959
rect 129093 8919 129151 8925
rect 129752 8928 129933 8956
rect 101125 8891 101183 8897
rect 101125 8888 101137 8891
rect 98748 8860 101137 8888
rect 101125 8857 101137 8860
rect 101171 8857 101183 8891
rect 103330 8888 103336 8900
rect 103291 8860 103336 8888
rect 101125 8851 101183 8857
rect 103330 8848 103336 8860
rect 103388 8848 103394 8900
rect 104158 8848 104164 8900
rect 104216 8888 104222 8900
rect 104216 8860 106596 8888
rect 104216 8848 104222 8860
rect 96246 8820 96252 8832
rect 95896 8792 96252 8820
rect 96246 8780 96252 8792
rect 96304 8780 96310 8832
rect 96614 8780 96620 8832
rect 96672 8820 96678 8832
rect 97258 8820 97264 8832
rect 96672 8792 96717 8820
rect 97219 8792 97264 8820
rect 96672 8780 96678 8792
rect 97258 8780 97264 8792
rect 97316 8780 97322 8832
rect 100478 8780 100484 8832
rect 100536 8820 100542 8832
rect 100573 8823 100631 8829
rect 100573 8820 100585 8823
rect 100536 8792 100585 8820
rect 100536 8780 100542 8792
rect 100573 8789 100585 8792
rect 100619 8789 100631 8823
rect 101030 8820 101036 8832
rect 100991 8792 101036 8820
rect 100573 8783 100631 8789
rect 101030 8780 101036 8792
rect 101088 8780 101094 8832
rect 102870 8820 102876 8832
rect 102831 8792 102876 8820
rect 102870 8780 102876 8792
rect 102928 8780 102934 8832
rect 104710 8780 104716 8832
rect 104768 8820 104774 8832
rect 104897 8823 104955 8829
rect 104897 8820 104909 8823
rect 104768 8792 104909 8820
rect 104768 8780 104774 8792
rect 104897 8789 104909 8792
rect 104943 8820 104955 8823
rect 106274 8820 106280 8832
rect 104943 8792 106280 8820
rect 104943 8789 104955 8792
rect 104897 8783 104955 8789
rect 106274 8780 106280 8792
rect 106332 8780 106338 8832
rect 106458 8820 106464 8832
rect 106419 8792 106464 8820
rect 106458 8780 106464 8792
rect 106516 8780 106522 8832
rect 106568 8820 106596 8860
rect 106642 8848 106648 8900
rect 106700 8888 106706 8900
rect 118510 8888 118516 8900
rect 106700 8860 118516 8888
rect 106700 8848 106706 8860
rect 118510 8848 118516 8860
rect 118568 8848 118574 8900
rect 121178 8848 121184 8900
rect 121236 8888 121242 8900
rect 126698 8888 126704 8900
rect 121236 8860 126704 8888
rect 121236 8848 121242 8860
rect 126698 8848 126704 8860
rect 126756 8848 126762 8900
rect 129752 8832 129780 8928
rect 129921 8925 129933 8928
rect 129967 8925 129979 8959
rect 131390 8956 131396 8968
rect 131351 8928 131396 8956
rect 129921 8919 129979 8925
rect 131390 8916 131396 8928
rect 131448 8956 131454 8968
rect 131761 8959 131819 8965
rect 131761 8956 131773 8959
rect 131448 8928 131773 8956
rect 131448 8916 131454 8928
rect 131761 8925 131773 8928
rect 131807 8925 131819 8959
rect 131761 8919 131819 8925
rect 140041 8959 140099 8965
rect 140041 8925 140053 8959
rect 140087 8956 140099 8959
rect 140682 8956 140688 8968
rect 140087 8928 140688 8956
rect 140087 8925 140099 8928
rect 140041 8919 140099 8925
rect 140682 8916 140688 8928
rect 140740 8916 140746 8968
rect 139854 8848 139860 8900
rect 139912 8888 139918 8900
rect 140976 8888 141004 8996
rect 141053 8959 141111 8965
rect 141053 8925 141065 8959
rect 141099 8925 141111 8959
rect 141053 8919 141111 8925
rect 142341 8959 142399 8965
rect 142341 8925 142353 8959
rect 142387 8925 142399 8959
rect 142448 8956 142476 8996
rect 142525 8993 142537 9027
rect 142571 9024 142583 9027
rect 142798 9024 142804 9036
rect 142571 8996 142804 9024
rect 142571 8993 142583 8996
rect 142525 8987 142583 8993
rect 142798 8984 142804 8996
rect 142856 8984 142862 9036
rect 143810 9024 143816 9036
rect 143092 8996 143816 9024
rect 143092 8956 143120 8996
rect 143810 8984 143816 8996
rect 143868 8984 143874 9036
rect 144178 8984 144184 9036
rect 144236 9024 144242 9036
rect 144641 9027 144699 9033
rect 144641 9024 144653 9027
rect 144236 8996 144653 9024
rect 144236 8984 144242 8996
rect 144641 8993 144653 8996
rect 144687 8993 144699 9027
rect 148060 9024 148088 9064
rect 148778 9024 148784 9036
rect 144641 8987 144699 8993
rect 147968 8996 148088 9024
rect 148739 8996 148784 9024
rect 142448 8928 143120 8956
rect 142341 8919 142399 8925
rect 139912 8860 141004 8888
rect 139912 8848 139918 8860
rect 109313 8823 109371 8829
rect 109313 8820 109325 8823
rect 106568 8792 109325 8820
rect 109313 8789 109325 8792
rect 109359 8789 109371 8823
rect 109313 8783 109371 8789
rect 109497 8823 109555 8829
rect 109497 8789 109509 8823
rect 109543 8820 109555 8823
rect 109586 8820 109592 8832
rect 109543 8792 109592 8820
rect 109543 8789 109555 8792
rect 109497 8783 109555 8789
rect 109586 8780 109592 8792
rect 109644 8780 109650 8832
rect 115290 8820 115296 8832
rect 115251 8792 115296 8820
rect 115290 8780 115296 8792
rect 115348 8780 115354 8832
rect 117498 8820 117504 8832
rect 117459 8792 117504 8820
rect 117498 8780 117504 8792
rect 117556 8780 117562 8832
rect 120261 8823 120319 8829
rect 120261 8789 120273 8823
rect 120307 8820 120319 8823
rect 120442 8820 120448 8832
rect 120307 8792 120448 8820
rect 120307 8789 120319 8792
rect 120261 8783 120319 8789
rect 120442 8780 120448 8792
rect 120500 8820 120506 8832
rect 120994 8820 121000 8832
rect 120500 8792 121000 8820
rect 120500 8780 120506 8792
rect 120994 8780 121000 8792
rect 121052 8780 121058 8832
rect 123570 8820 123576 8832
rect 123483 8792 123576 8820
rect 123570 8780 123576 8792
rect 123628 8820 123634 8832
rect 125318 8820 125324 8832
rect 123628 8792 125324 8820
rect 123628 8780 123634 8792
rect 125318 8780 125324 8792
rect 125376 8780 125382 8832
rect 125413 8823 125471 8829
rect 125413 8789 125425 8823
rect 125459 8820 125471 8823
rect 125686 8820 125692 8832
rect 125459 8792 125692 8820
rect 125459 8789 125471 8792
rect 125413 8783 125471 8789
rect 125686 8780 125692 8792
rect 125744 8780 125750 8832
rect 125965 8823 126023 8829
rect 125965 8789 125977 8823
rect 126011 8820 126023 8823
rect 127158 8820 127164 8832
rect 126011 8792 127164 8820
rect 126011 8789 126023 8792
rect 125965 8783 126023 8789
rect 127158 8780 127164 8792
rect 127216 8780 127222 8832
rect 129734 8820 129740 8832
rect 129695 8792 129740 8820
rect 129734 8780 129740 8792
rect 129792 8780 129798 8832
rect 140866 8820 140872 8832
rect 140827 8792 140872 8820
rect 140866 8780 140872 8792
rect 140924 8820 140930 8832
rect 141068 8820 141096 8919
rect 142356 8888 142384 8919
rect 143166 8916 143172 8968
rect 143224 8956 143230 8968
rect 143353 8959 143411 8965
rect 143353 8956 143365 8959
rect 143224 8928 143365 8956
rect 143224 8916 143230 8928
rect 143353 8925 143365 8928
rect 143399 8956 143411 8959
rect 146018 8956 146024 8968
rect 143399 8928 146024 8956
rect 143399 8925 143411 8928
rect 143353 8919 143411 8925
rect 146018 8916 146024 8928
rect 146076 8916 146082 8968
rect 146481 8959 146539 8965
rect 146481 8956 146493 8959
rect 146312 8928 146493 8956
rect 142985 8891 143043 8897
rect 142985 8888 142997 8891
rect 142356 8860 142997 8888
rect 142985 8857 142997 8860
rect 143031 8888 143043 8891
rect 145834 8888 145840 8900
rect 143031 8860 145840 8888
rect 143031 8857 143043 8860
rect 142985 8851 143043 8857
rect 145834 8848 145840 8860
rect 145892 8848 145898 8900
rect 146312 8832 146340 8928
rect 146481 8925 146493 8928
rect 146527 8925 146539 8959
rect 146481 8919 146539 8925
rect 146570 8848 146576 8900
rect 146628 8888 146634 8900
rect 147968 8888 147996 8996
rect 148778 8984 148784 8996
rect 148836 8984 148842 9036
rect 149330 9024 149336 9036
rect 149291 8996 149336 9024
rect 149330 8984 149336 8996
rect 149388 8984 149394 9036
rect 149440 9024 149468 9064
rect 150805 9061 150817 9095
rect 150851 9092 150863 9095
rect 151998 9092 152004 9104
rect 150851 9064 152004 9092
rect 150851 9061 150863 9064
rect 150805 9055 150863 9061
rect 151998 9052 152004 9064
rect 152056 9052 152062 9104
rect 152108 9092 152136 9132
rect 154393 9129 154405 9163
rect 154439 9160 154451 9163
rect 154942 9160 154948 9172
rect 154439 9132 154948 9160
rect 154439 9129 154451 9132
rect 154393 9123 154451 9129
rect 154942 9120 154948 9132
rect 155000 9120 155006 9172
rect 157150 9160 157156 9172
rect 157111 9132 157156 9160
rect 157150 9120 157156 9132
rect 157208 9120 157214 9172
rect 165798 9160 165804 9172
rect 165759 9132 165804 9160
rect 165798 9120 165804 9132
rect 165856 9120 165862 9172
rect 156138 9092 156144 9104
rect 152108 9064 156144 9092
rect 156138 9052 156144 9064
rect 156196 9052 156202 9104
rect 158254 9052 158260 9104
rect 158312 9092 158318 9104
rect 160830 9092 160836 9104
rect 158312 9064 160836 9092
rect 158312 9052 158318 9064
rect 160830 9052 160836 9064
rect 160888 9052 160894 9104
rect 162026 9052 162032 9104
rect 162084 9052 162090 9104
rect 163501 9095 163559 9101
rect 163501 9061 163513 9095
rect 163547 9092 163559 9095
rect 166718 9092 166724 9104
rect 163547 9064 166724 9092
rect 163547 9061 163559 9064
rect 163501 9055 163559 9061
rect 151725 9027 151783 9033
rect 149440 8996 151032 9024
rect 148045 8959 148103 8965
rect 148045 8925 148057 8959
rect 148091 8956 148103 8959
rect 150897 8959 150955 8965
rect 148091 8928 148456 8956
rect 148091 8925 148103 8928
rect 148045 8919 148103 8925
rect 146628 8860 147996 8888
rect 146628 8848 146634 8860
rect 140924 8792 141096 8820
rect 140924 8780 140930 8792
rect 141970 8780 141976 8832
rect 142028 8820 142034 8832
rect 143258 8820 143264 8832
rect 142028 8792 143264 8820
rect 142028 8780 142034 8792
rect 143258 8780 143264 8792
rect 143316 8780 143322 8832
rect 143350 8780 143356 8832
rect 143408 8820 143414 8832
rect 143629 8823 143687 8829
rect 143629 8820 143641 8823
rect 143408 8792 143641 8820
rect 143408 8780 143414 8792
rect 143629 8789 143641 8792
rect 143675 8789 143687 8823
rect 146294 8820 146300 8832
rect 146255 8792 146300 8820
rect 143629 8783 143687 8789
rect 146294 8780 146300 8792
rect 146352 8780 146358 8832
rect 148428 8829 148456 8928
rect 150897 8925 150909 8959
rect 150943 8925 150955 8959
rect 150897 8919 150955 8925
rect 148413 8823 148471 8829
rect 148413 8789 148425 8823
rect 148459 8820 148471 8823
rect 149146 8820 149152 8832
rect 148459 8792 149152 8820
rect 148459 8789 148471 8792
rect 148413 8783 148471 8789
rect 149146 8780 149152 8792
rect 149204 8780 149210 8832
rect 150912 8820 150940 8919
rect 151004 8888 151032 8996
rect 151725 8993 151737 9027
rect 151771 9024 151783 9027
rect 151814 9024 151820 9036
rect 151771 8996 151820 9024
rect 151771 8993 151783 8996
rect 151725 8987 151783 8993
rect 151814 8984 151820 8996
rect 151872 8984 151878 9036
rect 153105 9027 153163 9033
rect 153105 8993 153117 9027
rect 153151 9024 153163 9027
rect 153838 9024 153844 9036
rect 153151 8996 153844 9024
rect 153151 8993 153163 8996
rect 153105 8987 153163 8993
rect 153838 8984 153844 8996
rect 153896 8984 153902 9036
rect 156046 9024 156052 9036
rect 156007 8996 156052 9024
rect 156046 8984 156052 8996
rect 156104 8984 156110 9036
rect 158622 9024 158628 9036
rect 158583 8996 158628 9024
rect 158622 8984 158628 8996
rect 158680 8984 158686 9036
rect 160462 9024 160468 9036
rect 160423 8996 160468 9024
rect 160462 8984 160468 8996
rect 160520 8984 160526 9036
rect 161198 8984 161204 9036
rect 161256 9024 161262 9036
rect 161477 9027 161535 9033
rect 161477 9024 161489 9027
rect 161256 8996 161489 9024
rect 161256 8984 161262 8996
rect 161477 8993 161489 8996
rect 161523 8993 161535 9027
rect 162044 9024 162072 9052
rect 163608 9033 163636 9064
rect 166718 9052 166724 9064
rect 166776 9052 166782 9104
rect 163593 9027 163651 9033
rect 162044 8996 163544 9024
rect 161477 8987 161535 8993
rect 153289 8959 153347 8965
rect 153289 8925 153301 8959
rect 153335 8925 153347 8959
rect 154853 8959 154911 8965
rect 154853 8956 154865 8959
rect 153289 8919 153347 8925
rect 153948 8928 154865 8956
rect 151814 8888 151820 8900
rect 151004 8860 151820 8888
rect 151814 8848 151820 8860
rect 151872 8848 151878 8900
rect 151265 8823 151323 8829
rect 151265 8820 151277 8823
rect 150912 8792 151277 8820
rect 151265 8789 151277 8792
rect 151311 8820 151323 8823
rect 151722 8820 151728 8832
rect 151311 8792 151728 8820
rect 151311 8789 151323 8792
rect 151265 8783 151323 8789
rect 151722 8780 151728 8792
rect 151780 8780 151786 8832
rect 153304 8820 153332 8919
rect 153654 8820 153660 8832
rect 153304 8792 153660 8820
rect 153654 8780 153660 8792
rect 153712 8780 153718 8832
rect 153838 8780 153844 8832
rect 153896 8820 153902 8832
rect 153948 8829 153976 8928
rect 154853 8925 154865 8928
rect 154899 8925 154911 8959
rect 155954 8956 155960 8968
rect 155915 8928 155960 8956
rect 154853 8919 154911 8925
rect 155954 8916 155960 8928
rect 156012 8956 156018 8968
rect 156693 8959 156751 8965
rect 156693 8956 156705 8959
rect 156012 8928 156705 8956
rect 156012 8916 156018 8928
rect 156693 8925 156705 8928
rect 156739 8925 156751 8959
rect 157242 8956 157248 8968
rect 157203 8928 157248 8956
rect 156693 8919 156751 8925
rect 157242 8916 157248 8928
rect 157300 8916 157306 8968
rect 158530 8956 158536 8968
rect 158491 8928 158536 8956
rect 158530 8916 158536 8928
rect 158588 8916 158594 8968
rect 162029 8959 162087 8965
rect 162029 8925 162041 8959
rect 162075 8956 162087 8959
rect 163516 8956 163544 8996
rect 163593 8993 163605 9027
rect 163639 9024 163651 9027
rect 164605 9027 164663 9033
rect 164605 9024 164617 9027
rect 163639 8996 163673 9024
rect 163792 8996 164617 9024
rect 163639 8993 163651 8996
rect 163593 8987 163651 8993
rect 163792 8956 163820 8996
rect 164605 8993 164617 8996
rect 164651 8993 164663 9027
rect 164605 8987 164663 8993
rect 162075 8928 162348 8956
rect 163516 8928 163820 8956
rect 162075 8925 162087 8928
rect 162029 8919 162087 8925
rect 162320 8832 162348 8928
rect 164418 8916 164424 8968
rect 164476 8956 164482 8968
rect 164697 8959 164755 8965
rect 164697 8956 164709 8959
rect 164476 8928 164709 8956
rect 164476 8916 164482 8928
rect 164697 8925 164709 8928
rect 164743 8956 164755 8959
rect 165433 8959 165491 8965
rect 165433 8956 165445 8959
rect 164743 8928 165445 8956
rect 164743 8925 164755 8928
rect 164697 8919 164755 8925
rect 165433 8925 165445 8928
rect 165479 8925 165491 8959
rect 165433 8919 165491 8925
rect 163133 8891 163191 8897
rect 163133 8857 163145 8891
rect 163179 8888 163191 8891
rect 163222 8888 163228 8900
rect 163179 8860 163228 8888
rect 163179 8857 163191 8860
rect 163133 8851 163191 8857
rect 163222 8848 163228 8860
rect 163280 8888 163286 8900
rect 166077 8891 166135 8897
rect 166077 8888 166089 8891
rect 163280 8860 166089 8888
rect 163280 8848 163286 8860
rect 166077 8857 166089 8860
rect 166123 8857 166135 8891
rect 166077 8851 166135 8857
rect 153933 8823 153991 8829
rect 153933 8820 153945 8823
rect 153896 8792 153945 8820
rect 153896 8780 153902 8792
rect 153933 8789 153945 8792
rect 153979 8789 153991 8823
rect 153933 8783 153991 8789
rect 159177 8823 159235 8829
rect 159177 8789 159189 8823
rect 159223 8820 159235 8823
rect 159266 8820 159272 8832
rect 159223 8792 159272 8820
rect 159223 8789 159235 8792
rect 159177 8783 159235 8789
rect 159266 8780 159272 8792
rect 159324 8780 159330 8832
rect 162302 8820 162308 8832
rect 162263 8792 162308 8820
rect 162302 8780 162308 8792
rect 162360 8780 162366 8832
rect 166902 8820 166908 8832
rect 166863 8792 166908 8820
rect 166902 8780 166908 8792
rect 166960 8780 166966 8832
rect 368 8730 169556 8752
rect 368 8678 56667 8730
rect 56719 8678 56731 8730
rect 56783 8678 56795 8730
rect 56847 8678 56859 8730
rect 56911 8678 113088 8730
rect 113140 8678 113152 8730
rect 113204 8678 113216 8730
rect 113268 8678 113280 8730
rect 113332 8678 169556 8730
rect 368 8656 169556 8678
rect 1854 8576 1860 8628
rect 1912 8616 1918 8628
rect 5166 8616 5172 8628
rect 1912 8588 5172 8616
rect 1912 8576 1918 8588
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5534 8616 5540 8628
rect 5495 8588 5540 8616
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 6362 8616 6368 8628
rect 6323 8588 6368 8616
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 22278 8616 22284 8628
rect 8772 8588 22284 8616
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 4120 8520 4844 8548
rect 4120 8508 4126 8520
rect 3602 8412 3608 8424
rect 3563 8384 3608 8412
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8381 4675 8415
rect 4816 8412 4844 8520
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 8772 8548 8800 8588
rect 22278 8576 22284 8588
rect 22336 8576 22342 8628
rect 24394 8616 24400 8628
rect 22388 8588 24400 8616
rect 5316 8520 8800 8548
rect 5316 8508 5322 8520
rect 8846 8508 8852 8560
rect 8904 8548 8910 8560
rect 17586 8548 17592 8560
rect 8904 8520 17592 8548
rect 8904 8508 8910 8520
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 17678 8508 17684 8560
rect 17736 8548 17742 8560
rect 17736 8520 18000 8548
rect 17736 8508 17742 8520
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5534 8480 5540 8492
rect 5215 8452 5540 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5644 8452 9076 8480
rect 5644 8412 5672 8452
rect 4816 8384 5672 8412
rect 4617 8375 4675 8381
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 4632 8344 4660 8375
rect 2280 8316 4660 8344
rect 9048 8344 9076 8452
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 14826 8480 14832 8492
rect 10008 8452 14320 8480
rect 14787 8452 14832 8480
rect 10008 8440 10014 8452
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 13354 8412 13360 8424
rect 13311 8384 13360 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 14292 8421 14320 8452
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 15654 8480 15660 8492
rect 15160 8452 15660 8480
rect 15160 8440 15166 8452
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 15838 8480 15844 8492
rect 15799 8452 15844 8480
rect 15838 8440 15844 8452
rect 15896 8440 15902 8492
rect 16393 8483 16451 8489
rect 16393 8449 16405 8483
rect 16439 8480 16451 8483
rect 16666 8480 16672 8492
rect 16439 8452 16672 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 17310 8480 17316 8492
rect 17271 8452 17316 8480
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 17862 8480 17868 8492
rect 17823 8452 17868 8480
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 17972 8480 18000 8520
rect 18598 8508 18604 8560
rect 18656 8548 18662 8560
rect 18693 8551 18751 8557
rect 18693 8548 18705 8551
rect 18656 8520 18705 8548
rect 18656 8508 18662 8520
rect 18693 8517 18705 8520
rect 18739 8517 18751 8551
rect 21634 8548 21640 8560
rect 18693 8511 18751 8517
rect 18800 8520 21640 8548
rect 18800 8480 18828 8520
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 22388 8548 22416 8588
rect 24394 8576 24400 8588
rect 24452 8576 24458 8628
rect 25424 8588 25636 8616
rect 25424 8548 25452 8588
rect 21784 8520 22416 8548
rect 23216 8520 25452 8548
rect 25608 8548 25636 8588
rect 25682 8576 25688 8628
rect 25740 8616 25746 8628
rect 25958 8616 25964 8628
rect 25740 8588 25964 8616
rect 25740 8576 25746 8588
rect 25958 8576 25964 8588
rect 26016 8576 26022 8628
rect 26050 8576 26056 8628
rect 26108 8616 26114 8628
rect 27433 8619 27491 8625
rect 27433 8616 27445 8619
rect 26108 8588 27445 8616
rect 26108 8576 26114 8588
rect 27433 8585 27445 8588
rect 27479 8585 27491 8619
rect 27433 8579 27491 8585
rect 27522 8576 27528 8628
rect 27580 8616 27586 8628
rect 33594 8616 33600 8628
rect 27580 8588 33600 8616
rect 27580 8576 27586 8588
rect 33594 8576 33600 8588
rect 33652 8576 33658 8628
rect 34422 8576 34428 8628
rect 34480 8616 34486 8628
rect 40954 8616 40960 8628
rect 34480 8588 40960 8616
rect 34480 8576 34486 8588
rect 40954 8576 40960 8588
rect 41012 8576 41018 8628
rect 41506 8616 41512 8628
rect 41156 8588 41368 8616
rect 41467 8588 41512 8616
rect 33226 8548 33232 8560
rect 25608 8520 33232 8548
rect 21784 8508 21790 8520
rect 19794 8480 19800 8492
rect 17972 8452 18828 8480
rect 19755 8452 19800 8480
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8480 20315 8483
rect 21085 8483 21143 8489
rect 20303 8452 20668 8480
rect 20303 8449 20315 8452
rect 20257 8443 20315 8449
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 16025 8415 16083 8421
rect 16025 8381 16037 8415
rect 16071 8412 16083 8415
rect 17328 8412 17356 8440
rect 18322 8412 18328 8424
rect 16071 8384 17264 8412
rect 17328 8384 18328 8412
rect 16071 8381 16083 8384
rect 16025 8375 16083 8381
rect 17126 8344 17132 8356
rect 9048 8316 17132 8344
rect 2280 8304 2286 8316
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 15102 8276 15108 8288
rect 9272 8248 15108 8276
rect 9272 8236 9278 8248
rect 15102 8236 15108 8248
rect 15160 8236 15166 8288
rect 17236 8276 17264 8384
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 17402 8344 17408 8356
rect 17363 8316 17408 8344
rect 17402 8304 17408 8316
rect 17460 8304 17466 8356
rect 17954 8344 17960 8356
rect 17512 8316 17960 8344
rect 17512 8276 17540 8316
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 19610 8344 19616 8356
rect 19571 8316 19616 8344
rect 19610 8304 19616 8316
rect 19668 8304 19674 8356
rect 20640 8353 20668 8452
rect 21085 8449 21097 8483
rect 21131 8449 21143 8483
rect 21818 8480 21824 8492
rect 21731 8452 21824 8480
rect 21085 8443 21143 8449
rect 20898 8412 20904 8424
rect 20859 8384 20904 8412
rect 20898 8372 20904 8384
rect 20956 8412 20962 8424
rect 21100 8412 21128 8443
rect 21818 8440 21824 8452
rect 21876 8480 21882 8492
rect 22922 8480 22928 8492
rect 21876 8452 22928 8480
rect 21876 8440 21882 8452
rect 22922 8440 22928 8452
rect 22980 8440 22986 8492
rect 23106 8480 23112 8492
rect 23067 8452 23112 8480
rect 23106 8440 23112 8452
rect 23164 8440 23170 8492
rect 21450 8412 21456 8424
rect 20956 8384 21128 8412
rect 21411 8384 21456 8412
rect 20956 8372 20962 8384
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 23216 8412 23244 8520
rect 33226 8508 33232 8520
rect 33284 8508 33290 8560
rect 34146 8508 34152 8560
rect 34204 8548 34210 8560
rect 36906 8548 36912 8560
rect 34204 8520 36912 8548
rect 34204 8508 34210 8520
rect 36906 8508 36912 8520
rect 36964 8508 36970 8560
rect 37737 8551 37795 8557
rect 37737 8548 37749 8551
rect 37384 8520 37749 8548
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 25041 8483 25099 8489
rect 23716 8452 23761 8480
rect 23716 8440 23722 8452
rect 25041 8449 25053 8483
rect 25087 8449 25099 8483
rect 25222 8480 25228 8492
rect 25183 8452 25228 8480
rect 25041 8443 25099 8449
rect 25056 8412 25084 8443
rect 25222 8440 25228 8452
rect 25280 8440 25286 8492
rect 25590 8480 25596 8492
rect 25551 8452 25596 8480
rect 25590 8440 25596 8452
rect 25648 8440 25654 8492
rect 25774 8440 25780 8492
rect 25832 8480 25838 8492
rect 25832 8452 26556 8480
rect 25832 8440 25838 8452
rect 25130 8412 25136 8424
rect 21928 8384 23244 8412
rect 25043 8384 25136 8412
rect 20625 8347 20683 8353
rect 20625 8313 20637 8347
rect 20671 8344 20683 8347
rect 21928 8344 21956 8384
rect 25130 8372 25136 8384
rect 25188 8412 25194 8424
rect 26421 8415 26479 8421
rect 26421 8412 26433 8415
rect 25188 8384 26433 8412
rect 25188 8372 25194 8384
rect 26421 8381 26433 8384
rect 26467 8381 26479 8415
rect 26421 8375 26479 8381
rect 22094 8344 22100 8356
rect 20671 8316 21956 8344
rect 22055 8316 22100 8344
rect 20671 8313 20683 8316
rect 20625 8307 20683 8313
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 23014 8344 23020 8356
rect 22975 8316 23020 8344
rect 23014 8304 23020 8316
rect 23072 8304 23078 8356
rect 23934 8344 23940 8356
rect 23895 8316 23940 8344
rect 23934 8304 23940 8316
rect 23992 8304 23998 8356
rect 26528 8344 26556 8452
rect 26602 8440 26608 8492
rect 26660 8480 26666 8492
rect 34422 8480 34428 8492
rect 26660 8452 34428 8480
rect 26660 8440 26666 8452
rect 34422 8440 34428 8452
rect 34480 8440 34486 8492
rect 34790 8480 34796 8492
rect 34751 8452 34796 8480
rect 34790 8440 34796 8452
rect 34848 8440 34854 8492
rect 34882 8440 34888 8492
rect 34940 8480 34946 8492
rect 35161 8483 35219 8489
rect 35161 8480 35173 8483
rect 34940 8452 35173 8480
rect 34940 8440 34946 8452
rect 35161 8449 35173 8452
rect 35207 8449 35219 8483
rect 35526 8480 35532 8492
rect 35487 8452 35532 8480
rect 35161 8443 35219 8449
rect 35526 8440 35532 8452
rect 35584 8440 35590 8492
rect 36722 8480 36728 8492
rect 36683 8452 36728 8480
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 37384 8489 37412 8520
rect 37737 8517 37749 8520
rect 37783 8548 37795 8551
rect 41156 8548 41184 8588
rect 37783 8520 41184 8548
rect 41340 8548 41368 8588
rect 41506 8576 41512 8588
rect 41564 8576 41570 8628
rect 45922 8616 45928 8628
rect 41616 8588 45928 8616
rect 41616 8548 41644 8588
rect 45922 8576 45928 8588
rect 45980 8576 45986 8628
rect 46106 8576 46112 8628
rect 46164 8616 46170 8628
rect 47486 8616 47492 8628
rect 46164 8588 47492 8616
rect 46164 8576 46170 8588
rect 47486 8576 47492 8588
rect 47544 8576 47550 8628
rect 47578 8576 47584 8628
rect 47636 8616 47642 8628
rect 48222 8616 48228 8628
rect 47636 8588 48228 8616
rect 47636 8576 47642 8588
rect 48222 8576 48228 8588
rect 48280 8576 48286 8628
rect 48498 8576 48504 8628
rect 48556 8616 48562 8628
rect 49326 8616 49332 8628
rect 48556 8588 49332 8616
rect 48556 8576 48562 8588
rect 49326 8576 49332 8588
rect 49384 8576 49390 8628
rect 49786 8576 49792 8628
rect 49844 8616 49850 8628
rect 50246 8616 50252 8628
rect 49844 8588 50252 8616
rect 49844 8576 49850 8588
rect 50246 8576 50252 8588
rect 50304 8576 50310 8628
rect 50985 8619 51043 8625
rect 50985 8585 50997 8619
rect 51031 8616 51043 8619
rect 51534 8616 51540 8628
rect 51031 8588 51540 8616
rect 51031 8585 51043 8588
rect 50985 8579 51043 8585
rect 51534 8576 51540 8588
rect 51592 8576 51598 8628
rect 51629 8619 51687 8625
rect 51629 8585 51641 8619
rect 51675 8616 51687 8619
rect 51718 8616 51724 8628
rect 51675 8588 51724 8616
rect 51675 8585 51687 8588
rect 51629 8579 51687 8585
rect 51718 8576 51724 8588
rect 51776 8576 51782 8628
rect 52638 8616 52644 8628
rect 51828 8588 52644 8616
rect 41340 8520 41644 8548
rect 37783 8517 37795 8520
rect 37737 8511 37795 8517
rect 42426 8508 42432 8560
rect 42484 8548 42490 8560
rect 42521 8551 42579 8557
rect 42521 8548 42533 8551
rect 42484 8520 42533 8548
rect 42484 8508 42490 8520
rect 42521 8517 42533 8520
rect 42567 8517 42579 8551
rect 42521 8511 42579 8517
rect 42610 8508 42616 8560
rect 42668 8548 42674 8560
rect 43070 8548 43076 8560
rect 42668 8520 43076 8548
rect 42668 8508 42674 8520
rect 43070 8508 43076 8520
rect 43128 8508 43134 8560
rect 48314 8548 48320 8560
rect 43732 8520 48320 8548
rect 37369 8483 37427 8489
rect 36832 8452 37320 8480
rect 26694 8372 26700 8424
rect 26752 8412 26758 8424
rect 29178 8412 29184 8424
rect 26752 8384 29184 8412
rect 26752 8372 26758 8384
rect 29178 8372 29184 8384
rect 29236 8372 29242 8424
rect 29270 8372 29276 8424
rect 29328 8412 29334 8424
rect 29328 8384 34008 8412
rect 29328 8372 29334 8384
rect 33778 8344 33784 8356
rect 24872 8316 26188 8344
rect 26528 8316 33784 8344
rect 17236 8248 17540 8276
rect 17586 8236 17592 8288
rect 17644 8276 17650 8288
rect 24872 8276 24900 8316
rect 17644 8248 24900 8276
rect 17644 8236 17650 8248
rect 25774 8236 25780 8288
rect 25832 8276 25838 8288
rect 25961 8279 26019 8285
rect 25961 8276 25973 8279
rect 25832 8248 25973 8276
rect 25832 8236 25838 8248
rect 25961 8245 25973 8248
rect 26007 8245 26019 8279
rect 26160 8276 26188 8316
rect 33778 8304 33784 8316
rect 33836 8304 33842 8356
rect 33980 8344 34008 8384
rect 34330 8372 34336 8424
rect 34388 8412 34394 8424
rect 36832 8412 36860 8452
rect 34388 8384 36860 8412
rect 37001 8415 37059 8421
rect 34388 8372 34394 8384
rect 37001 8381 37013 8415
rect 37047 8412 37059 8415
rect 37182 8412 37188 8424
rect 37047 8384 37188 8412
rect 37047 8381 37059 8384
rect 37001 8375 37059 8381
rect 37182 8372 37188 8384
rect 37240 8372 37246 8424
rect 37292 8412 37320 8452
rect 37369 8449 37381 8483
rect 37415 8449 37427 8483
rect 37369 8443 37427 8449
rect 37461 8483 37519 8489
rect 37461 8449 37473 8483
rect 37507 8480 37519 8483
rect 38286 8480 38292 8492
rect 37507 8452 38292 8480
rect 37507 8449 37519 8452
rect 37461 8443 37519 8449
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 38657 8483 38715 8489
rect 38657 8449 38669 8483
rect 38703 8480 38715 8483
rect 39390 8480 39396 8492
rect 38703 8452 39396 8480
rect 38703 8449 38715 8452
rect 38657 8443 38715 8449
rect 39390 8440 39396 8452
rect 39448 8480 39454 8492
rect 39761 8483 39819 8489
rect 39761 8480 39773 8483
rect 39448 8452 39773 8480
rect 39448 8440 39454 8452
rect 39761 8449 39773 8452
rect 39807 8449 39819 8483
rect 39761 8443 39819 8449
rect 39850 8440 39856 8492
rect 39908 8480 39914 8492
rect 40129 8483 40187 8489
rect 40129 8480 40141 8483
rect 39908 8452 40141 8480
rect 39908 8440 39914 8452
rect 40129 8449 40141 8452
rect 40175 8449 40187 8483
rect 40129 8443 40187 8449
rect 40497 8483 40555 8489
rect 40497 8449 40509 8483
rect 40543 8480 40555 8483
rect 40954 8480 40960 8492
rect 40543 8452 40960 8480
rect 40543 8449 40555 8452
rect 40497 8443 40555 8449
rect 40954 8440 40960 8452
rect 41012 8480 41018 8492
rect 41598 8480 41604 8492
rect 41012 8452 41604 8480
rect 41012 8440 41018 8452
rect 41598 8440 41604 8452
rect 41656 8440 41662 8492
rect 41690 8440 41696 8492
rect 41748 8480 41754 8492
rect 43530 8480 43536 8492
rect 41748 8452 43536 8480
rect 41748 8440 41754 8452
rect 43530 8440 43536 8452
rect 43588 8440 43594 8492
rect 37292 8384 38700 8412
rect 37461 8347 37519 8353
rect 37461 8344 37473 8347
rect 33980 8316 37473 8344
rect 37461 8313 37473 8316
rect 37507 8313 37519 8347
rect 38672 8344 38700 8384
rect 39206 8372 39212 8424
rect 39264 8412 39270 8424
rect 40678 8412 40684 8424
rect 39264 8384 40684 8412
rect 39264 8372 39270 8384
rect 40678 8372 40684 8384
rect 40736 8372 40742 8424
rect 40770 8372 40776 8424
rect 40828 8412 40834 8424
rect 43732 8412 43760 8520
rect 48314 8508 48320 8520
rect 48372 8508 48378 8560
rect 48406 8508 48412 8560
rect 48464 8548 48470 8560
rect 49605 8551 49663 8557
rect 49605 8548 49617 8551
rect 48464 8520 49617 8548
rect 48464 8508 48470 8520
rect 46474 8480 46480 8492
rect 40828 8384 43760 8412
rect 45480 8452 46480 8480
rect 40828 8372 40834 8384
rect 39758 8344 39764 8356
rect 38672 8316 39764 8344
rect 37461 8307 37519 8313
rect 39758 8304 39764 8316
rect 39816 8304 39822 8356
rect 40034 8304 40040 8356
rect 40092 8344 40098 8356
rect 45480 8344 45508 8452
rect 46474 8440 46480 8452
rect 46532 8440 46538 8492
rect 48774 8480 48780 8492
rect 46584 8452 48780 8480
rect 45554 8372 45560 8424
rect 45612 8412 45618 8424
rect 46584 8412 46612 8452
rect 48774 8440 48780 8452
rect 48832 8440 48838 8492
rect 48884 8489 48912 8520
rect 49605 8517 49617 8520
rect 49651 8517 49663 8551
rect 49605 8511 49663 8517
rect 49970 8508 49976 8560
rect 50028 8548 50034 8560
rect 51828 8548 51856 8588
rect 52638 8576 52644 8588
rect 52696 8576 52702 8628
rect 53190 8576 53196 8628
rect 53248 8616 53254 8628
rect 54018 8616 54024 8628
rect 53248 8588 54024 8616
rect 53248 8576 53254 8588
rect 54018 8576 54024 8588
rect 54076 8576 54082 8628
rect 55766 8576 55772 8628
rect 55824 8616 55830 8628
rect 57790 8616 57796 8628
rect 55824 8588 57796 8616
rect 55824 8576 55830 8588
rect 57790 8576 57796 8588
rect 57848 8576 57854 8628
rect 57882 8576 57888 8628
rect 57940 8616 57946 8628
rect 57977 8619 58035 8625
rect 57977 8616 57989 8619
rect 57940 8588 57989 8616
rect 57940 8576 57946 8588
rect 57977 8585 57989 8588
rect 58023 8585 58035 8619
rect 57977 8579 58035 8585
rect 58526 8576 58532 8628
rect 58584 8616 58590 8628
rect 59262 8616 59268 8628
rect 58584 8588 59268 8616
rect 58584 8576 58590 8588
rect 59262 8576 59268 8588
rect 59320 8576 59326 8628
rect 59446 8616 59452 8628
rect 59407 8588 59452 8616
rect 59446 8576 59452 8588
rect 59504 8576 59510 8628
rect 63034 8616 63040 8628
rect 59556 8588 63040 8616
rect 50028 8520 51856 8548
rect 50028 8508 50034 8520
rect 52362 8508 52368 8560
rect 52420 8548 52426 8560
rect 56778 8548 56784 8560
rect 52420 8520 56784 8548
rect 52420 8508 52426 8520
rect 56778 8508 56784 8520
rect 56836 8508 56842 8560
rect 57701 8551 57759 8557
rect 57701 8548 57713 8551
rect 57348 8520 57713 8548
rect 48869 8483 48927 8489
rect 48869 8449 48881 8483
rect 48915 8449 48927 8483
rect 48869 8443 48927 8449
rect 49329 8483 49387 8489
rect 49329 8449 49341 8483
rect 49375 8480 49387 8483
rect 49988 8480 50016 8508
rect 51994 8480 52000 8492
rect 49375 8452 50016 8480
rect 50080 8452 52000 8480
rect 49375 8449 49387 8452
rect 49329 8443 49387 8449
rect 45612 8384 46612 8412
rect 46661 8415 46719 8421
rect 45612 8372 45618 8384
rect 46661 8381 46673 8415
rect 46707 8412 46719 8415
rect 46750 8412 46756 8424
rect 46707 8384 46756 8412
rect 46707 8381 46719 8384
rect 46661 8375 46719 8381
rect 46750 8372 46756 8384
rect 46808 8372 46814 8424
rect 46842 8372 46848 8424
rect 46900 8412 46906 8424
rect 49878 8412 49884 8424
rect 46900 8384 49884 8412
rect 46900 8372 46906 8384
rect 49878 8372 49884 8384
rect 49936 8372 49942 8424
rect 40092 8316 45508 8344
rect 45572 8316 45876 8344
rect 40092 8304 40098 8316
rect 45572 8276 45600 8316
rect 45738 8276 45744 8288
rect 26160 8248 45600 8276
rect 45699 8248 45744 8276
rect 25961 8239 26019 8245
rect 45738 8236 45744 8248
rect 45796 8236 45802 8288
rect 45848 8276 45876 8316
rect 45922 8304 45928 8356
rect 45980 8344 45986 8356
rect 47854 8344 47860 8356
rect 45980 8316 47860 8344
rect 45980 8304 45986 8316
rect 47854 8304 47860 8316
rect 47912 8304 47918 8356
rect 48406 8304 48412 8356
rect 48464 8344 48470 8356
rect 48685 8347 48743 8353
rect 48685 8344 48697 8347
rect 48464 8316 48697 8344
rect 48464 8304 48470 8316
rect 48685 8313 48697 8316
rect 48731 8313 48743 8347
rect 48685 8307 48743 8313
rect 50080 8276 50108 8452
rect 51994 8440 52000 8452
rect 52052 8440 52058 8492
rect 52273 8483 52331 8489
rect 52273 8449 52285 8483
rect 52319 8480 52331 8483
rect 52730 8480 52736 8492
rect 52319 8452 52592 8480
rect 52643 8452 52736 8480
rect 52319 8449 52331 8452
rect 52273 8443 52331 8449
rect 50154 8372 50160 8424
rect 50212 8412 50218 8424
rect 52362 8412 52368 8424
rect 50212 8384 52368 8412
rect 50212 8372 50218 8384
rect 52362 8372 52368 8384
rect 52420 8372 52426 8424
rect 52564 8412 52592 8452
rect 52730 8440 52736 8452
rect 52788 8480 52794 8492
rect 54754 8480 54760 8492
rect 52788 8452 54760 8480
rect 52788 8440 52794 8452
rect 54754 8440 54760 8452
rect 54812 8440 54818 8492
rect 55125 8483 55183 8489
rect 55125 8449 55137 8483
rect 55171 8449 55183 8483
rect 55125 8443 55183 8449
rect 55585 8483 55643 8489
rect 55585 8449 55597 8483
rect 55631 8480 55643 8483
rect 55674 8480 55680 8492
rect 55631 8452 55680 8480
rect 55631 8449 55643 8452
rect 55585 8443 55643 8449
rect 53006 8412 53012 8424
rect 52564 8384 53012 8412
rect 53006 8372 53012 8384
rect 53064 8412 53070 8424
rect 53561 8415 53619 8421
rect 53561 8412 53573 8415
rect 53064 8384 53573 8412
rect 53064 8372 53070 8384
rect 53561 8381 53573 8384
rect 53607 8381 53619 8415
rect 53561 8375 53619 8381
rect 54846 8372 54852 8424
rect 54904 8412 54910 8424
rect 55140 8412 55168 8443
rect 55674 8440 55680 8452
rect 55732 8480 55738 8492
rect 55950 8480 55956 8492
rect 55732 8452 55956 8480
rect 55732 8440 55738 8452
rect 55950 8440 55956 8452
rect 56008 8440 56014 8492
rect 56042 8440 56048 8492
rect 56100 8440 56106 8492
rect 56226 8440 56232 8492
rect 56284 8480 56290 8492
rect 57348 8489 57376 8520
rect 57701 8517 57713 8520
rect 57747 8548 57759 8551
rect 58250 8548 58256 8560
rect 57747 8520 58256 8548
rect 57747 8517 57759 8520
rect 57701 8511 57759 8517
rect 58250 8508 58256 8520
rect 58308 8508 58314 8560
rect 59464 8548 59492 8576
rect 58636 8520 59492 8548
rect 56597 8483 56655 8489
rect 56597 8480 56609 8483
rect 56284 8452 56609 8480
rect 56284 8440 56290 8452
rect 56597 8449 56609 8452
rect 56643 8449 56655 8483
rect 56597 8443 56655 8449
rect 57333 8483 57391 8489
rect 57333 8449 57345 8483
rect 57379 8449 57391 8483
rect 57333 8443 57391 8449
rect 57422 8440 57428 8492
rect 57480 8480 57486 8492
rect 57606 8480 57612 8492
rect 57480 8452 57612 8480
rect 57480 8440 57486 8452
rect 57606 8440 57612 8452
rect 57664 8440 57670 8492
rect 58636 8489 58664 8520
rect 58621 8483 58679 8489
rect 58621 8449 58633 8483
rect 58667 8449 58679 8483
rect 58986 8480 58992 8492
rect 58947 8452 58992 8480
rect 58621 8443 58679 8449
rect 58986 8440 58992 8452
rect 59044 8440 59050 8492
rect 59078 8440 59084 8492
rect 59136 8480 59142 8492
rect 59556 8480 59584 8588
rect 63034 8576 63040 8588
rect 63092 8576 63098 8628
rect 63402 8576 63408 8628
rect 63460 8616 63466 8628
rect 65245 8619 65303 8625
rect 65245 8616 65257 8619
rect 63460 8588 65257 8616
rect 63460 8576 63466 8588
rect 65245 8585 65257 8588
rect 65291 8585 65303 8619
rect 65245 8579 65303 8585
rect 73433 8619 73491 8625
rect 73433 8585 73445 8619
rect 73479 8616 73491 8619
rect 74074 8616 74080 8628
rect 73479 8588 74080 8616
rect 73479 8585 73491 8588
rect 73433 8579 73491 8585
rect 74074 8576 74080 8588
rect 74132 8576 74138 8628
rect 74350 8576 74356 8628
rect 74408 8616 74414 8628
rect 74445 8619 74503 8625
rect 74445 8616 74457 8619
rect 74408 8588 74457 8616
rect 74408 8576 74414 8588
rect 74445 8585 74457 8588
rect 74491 8585 74503 8619
rect 80146 8616 80152 8628
rect 80107 8588 80152 8616
rect 74445 8579 74503 8585
rect 80146 8576 80152 8588
rect 80204 8576 80210 8628
rect 85850 8576 85856 8628
rect 85908 8616 85914 8628
rect 88334 8616 88340 8628
rect 85908 8588 88340 8616
rect 85908 8576 85914 8588
rect 88334 8576 88340 8588
rect 88392 8576 88398 8628
rect 89993 8619 90051 8625
rect 89993 8585 90005 8619
rect 90039 8616 90051 8619
rect 90266 8616 90272 8628
rect 90039 8588 90272 8616
rect 90039 8585 90051 8588
rect 89993 8579 90051 8585
rect 90266 8576 90272 8588
rect 90324 8576 90330 8628
rect 94777 8619 94835 8625
rect 94777 8616 94789 8619
rect 94424 8588 94789 8616
rect 59998 8508 60004 8560
rect 60056 8548 60062 8560
rect 65058 8548 65064 8560
rect 60056 8520 60504 8548
rect 60056 8508 60062 8520
rect 60182 8480 60188 8492
rect 59136 8452 59584 8480
rect 60143 8452 60188 8480
rect 59136 8440 59142 8452
rect 60182 8440 60188 8452
rect 60240 8440 60246 8492
rect 60277 8483 60335 8489
rect 60277 8449 60289 8483
rect 60323 8480 60335 8483
rect 60366 8480 60372 8492
rect 60323 8452 60372 8480
rect 60323 8449 60335 8452
rect 60277 8443 60335 8449
rect 60366 8440 60372 8452
rect 60424 8440 60430 8492
rect 60476 8489 60504 8520
rect 60660 8520 65064 8548
rect 60461 8483 60519 8489
rect 60461 8449 60473 8483
rect 60507 8480 60519 8483
rect 60550 8480 60556 8492
rect 60507 8452 60556 8480
rect 60507 8449 60519 8452
rect 60461 8443 60519 8449
rect 60550 8440 60556 8452
rect 60608 8440 60614 8492
rect 55861 8415 55919 8421
rect 55861 8412 55873 8415
rect 54904 8384 55873 8412
rect 54904 8372 54910 8384
rect 55861 8381 55873 8384
rect 55907 8381 55919 8415
rect 56060 8412 56088 8440
rect 58342 8412 58348 8424
rect 56060 8384 58348 8412
rect 55861 8375 55919 8381
rect 58342 8372 58348 8384
rect 58400 8372 58406 8424
rect 58713 8415 58771 8421
rect 58713 8381 58725 8415
rect 58759 8412 58771 8415
rect 59170 8412 59176 8424
rect 58759 8384 59176 8412
rect 58759 8381 58771 8384
rect 58713 8375 58771 8381
rect 59170 8372 59176 8384
rect 59228 8372 59234 8424
rect 59814 8372 59820 8424
rect 59872 8412 59878 8424
rect 60660 8412 60688 8520
rect 65058 8508 65064 8520
rect 65116 8508 65122 8560
rect 66254 8508 66260 8560
rect 66312 8548 66318 8560
rect 76558 8548 76564 8560
rect 66312 8520 76564 8548
rect 66312 8508 66318 8520
rect 76558 8508 76564 8520
rect 76616 8508 76622 8560
rect 85669 8551 85727 8557
rect 85669 8517 85681 8551
rect 85715 8548 85727 8551
rect 90450 8548 90456 8560
rect 85715 8520 90456 8548
rect 85715 8517 85727 8520
rect 85669 8511 85727 8517
rect 90450 8508 90456 8520
rect 90508 8508 90514 8560
rect 60826 8440 60832 8492
rect 60884 8480 60890 8492
rect 64414 8480 64420 8492
rect 60884 8452 64000 8480
rect 64375 8452 64420 8480
rect 60884 8440 60890 8452
rect 62850 8412 62856 8424
rect 59872 8384 60688 8412
rect 62811 8384 62856 8412
rect 59872 8372 59878 8384
rect 62850 8372 62856 8384
rect 62908 8372 62914 8424
rect 63862 8412 63868 8424
rect 63823 8384 63868 8412
rect 63862 8372 63868 8384
rect 63920 8372 63926 8424
rect 63972 8412 64000 8452
rect 64414 8440 64420 8452
rect 64472 8440 64478 8492
rect 83458 8480 83464 8492
rect 83419 8452 83464 8480
rect 83458 8440 83464 8452
rect 83516 8440 83522 8492
rect 87598 8440 87604 8492
rect 87656 8480 87662 8492
rect 87656 8452 89208 8480
rect 87656 8440 87662 8452
rect 68094 8412 68100 8424
rect 63972 8384 68100 8412
rect 68094 8372 68100 8384
rect 68152 8372 68158 8424
rect 71774 8412 71780 8424
rect 71735 8384 71780 8412
rect 71774 8372 71780 8384
rect 71832 8372 71838 8424
rect 79045 8415 79103 8421
rect 79045 8381 79057 8415
rect 79091 8412 79103 8415
rect 81986 8412 81992 8424
rect 79091 8384 79456 8412
rect 81947 8384 81992 8412
rect 79091 8381 79103 8384
rect 79045 8375 79103 8381
rect 50706 8304 50712 8356
rect 50764 8344 50770 8356
rect 50764 8316 51580 8344
rect 50764 8304 50770 8316
rect 45848 8248 50108 8276
rect 50522 8236 50528 8288
rect 50580 8276 50586 8288
rect 51074 8276 51080 8288
rect 50580 8248 51080 8276
rect 50580 8236 50586 8248
rect 51074 8236 51080 8248
rect 51132 8236 51138 8288
rect 51552 8276 51580 8316
rect 51626 8304 51632 8356
rect 51684 8344 51690 8356
rect 52089 8347 52147 8353
rect 52089 8344 52101 8347
rect 51684 8316 52101 8344
rect 51684 8304 51690 8316
rect 52089 8313 52101 8316
rect 52135 8313 52147 8347
rect 52089 8307 52147 8313
rect 52178 8304 52184 8356
rect 52236 8344 52242 8356
rect 53282 8344 53288 8356
rect 52236 8316 53288 8344
rect 52236 8304 52242 8316
rect 53282 8304 53288 8316
rect 53340 8304 53346 8356
rect 54938 8344 54944 8356
rect 54036 8316 54524 8344
rect 54899 8316 54944 8344
rect 51810 8276 51816 8288
rect 51552 8248 51816 8276
rect 51810 8236 51816 8248
rect 51868 8236 51874 8288
rect 51902 8236 51908 8288
rect 51960 8276 51966 8288
rect 54036 8276 54064 8316
rect 54386 8276 54392 8288
rect 51960 8248 54064 8276
rect 54347 8248 54392 8276
rect 51960 8236 51966 8248
rect 54386 8236 54392 8248
rect 54444 8236 54450 8288
rect 54496 8276 54524 8316
rect 54938 8304 54944 8316
rect 54996 8304 55002 8356
rect 55306 8304 55312 8356
rect 55364 8344 55370 8356
rect 56689 8347 56747 8353
rect 56689 8344 56701 8347
rect 55364 8316 56701 8344
rect 55364 8304 55370 8316
rect 56689 8313 56701 8316
rect 56735 8313 56747 8347
rect 56689 8307 56747 8313
rect 56778 8304 56784 8356
rect 56836 8344 56842 8356
rect 64322 8344 64328 8356
rect 56836 8316 64328 8344
rect 56836 8304 56842 8316
rect 64322 8304 64328 8316
rect 64380 8304 64386 8356
rect 79428 8288 79456 8384
rect 81986 8372 81992 8384
rect 82044 8372 82050 8424
rect 82998 8412 83004 8424
rect 82959 8384 83004 8412
rect 82998 8372 83004 8384
rect 83056 8372 83062 8424
rect 86681 8415 86739 8421
rect 86681 8381 86693 8415
rect 86727 8412 86739 8415
rect 87230 8412 87236 8424
rect 86727 8384 87236 8412
rect 86727 8381 86739 8384
rect 86681 8375 86739 8381
rect 87230 8372 87236 8384
rect 87288 8412 87294 8424
rect 87693 8415 87751 8421
rect 87693 8412 87705 8415
rect 87288 8384 87705 8412
rect 87288 8372 87294 8384
rect 87693 8381 87705 8384
rect 87739 8381 87751 8415
rect 87693 8375 87751 8381
rect 87966 8372 87972 8424
rect 88024 8412 88030 8424
rect 89180 8412 89208 8452
rect 89254 8440 89260 8492
rect 89312 8480 89318 8492
rect 91646 8480 91652 8492
rect 89312 8452 89357 8480
rect 90192 8452 91324 8480
rect 91607 8452 91652 8480
rect 89312 8440 89318 8452
rect 90192 8412 90220 8452
rect 88024 8384 89116 8412
rect 89180 8384 90220 8412
rect 90269 8415 90327 8421
rect 88024 8372 88030 8384
rect 86862 8304 86868 8356
rect 86920 8344 86926 8356
rect 88981 8347 89039 8353
rect 88981 8344 88993 8347
rect 86920 8316 88993 8344
rect 86920 8304 86926 8316
rect 88981 8313 88993 8316
rect 89027 8313 89039 8347
rect 89088 8344 89116 8384
rect 90269 8381 90281 8415
rect 90315 8412 90327 8415
rect 90450 8412 90456 8424
rect 90315 8384 90456 8412
rect 90315 8381 90327 8384
rect 90269 8375 90327 8381
rect 90450 8372 90456 8384
rect 90508 8372 90514 8424
rect 91296 8421 91324 8452
rect 91646 8440 91652 8452
rect 91704 8440 91710 8492
rect 92842 8480 92848 8492
rect 92803 8452 92848 8480
rect 92842 8440 92848 8452
rect 92900 8440 92906 8492
rect 94424 8489 94452 8588
rect 94777 8585 94789 8588
rect 94823 8616 94835 8619
rect 98270 8616 98276 8628
rect 94823 8588 98276 8616
rect 94823 8585 94835 8588
rect 94777 8579 94835 8585
rect 98270 8576 98276 8588
rect 98328 8576 98334 8628
rect 98365 8619 98423 8625
rect 98365 8585 98377 8619
rect 98411 8616 98423 8619
rect 103330 8616 103336 8628
rect 98411 8588 103336 8616
rect 98411 8585 98423 8588
rect 98365 8579 98423 8585
rect 94958 8508 94964 8560
rect 95016 8548 95022 8560
rect 98089 8551 98147 8557
rect 98089 8548 98101 8551
rect 95016 8520 98101 8548
rect 95016 8508 95022 8520
rect 98089 8517 98101 8520
rect 98135 8517 98147 8551
rect 98089 8511 98147 8517
rect 94409 8483 94467 8489
rect 94409 8449 94421 8483
rect 94455 8449 94467 8483
rect 94409 8443 94467 8449
rect 94590 8440 94596 8492
rect 94648 8480 94654 8492
rect 97629 8483 97687 8489
rect 94648 8452 96200 8480
rect 94648 8440 94654 8452
rect 91281 8415 91339 8421
rect 91281 8381 91293 8415
rect 91327 8381 91339 8415
rect 91281 8375 91339 8381
rect 92106 8372 92112 8424
rect 92164 8412 92170 8424
rect 93857 8415 93915 8421
rect 93857 8412 93869 8415
rect 92164 8384 93869 8412
rect 92164 8372 92170 8384
rect 93857 8381 93869 8384
rect 93903 8381 93915 8415
rect 96065 8415 96123 8421
rect 96065 8412 96077 8415
rect 93857 8375 93915 8381
rect 95620 8384 96077 8412
rect 95620 8356 95648 8384
rect 96065 8381 96077 8384
rect 96111 8381 96123 8415
rect 96065 8375 96123 8381
rect 91094 8344 91100 8356
rect 89088 8316 91100 8344
rect 88981 8307 89039 8313
rect 91094 8304 91100 8316
rect 91152 8304 91158 8356
rect 95602 8344 95608 8356
rect 95563 8316 95608 8344
rect 95602 8304 95608 8316
rect 95660 8304 95666 8356
rect 96172 8344 96200 8452
rect 97629 8449 97641 8483
rect 97675 8480 97687 8483
rect 97994 8480 98000 8492
rect 97675 8452 98000 8480
rect 97675 8449 97687 8452
rect 97629 8443 97687 8449
rect 97994 8440 98000 8452
rect 98052 8440 98058 8492
rect 98472 8489 98500 8588
rect 103330 8576 103336 8588
rect 103388 8576 103394 8628
rect 108390 8576 108396 8628
rect 108448 8616 108454 8628
rect 113269 8619 113327 8625
rect 113269 8616 113281 8619
rect 108448 8588 113281 8616
rect 108448 8576 108454 8588
rect 113269 8585 113281 8588
rect 113315 8585 113327 8619
rect 119890 8616 119896 8628
rect 113269 8579 113327 8585
rect 113836 8588 119896 8616
rect 101493 8551 101551 8557
rect 101493 8548 101505 8551
rect 99576 8520 101505 8548
rect 98457 8483 98515 8489
rect 98457 8449 98469 8483
rect 98503 8449 98515 8483
rect 99576 8480 99604 8520
rect 101493 8517 101505 8520
rect 101539 8517 101551 8551
rect 101493 8511 101551 8517
rect 102686 8508 102692 8560
rect 102744 8548 102750 8560
rect 113836 8548 113864 8588
rect 119890 8576 119896 8588
rect 119948 8576 119954 8628
rect 121270 8576 121276 8628
rect 121328 8616 121334 8628
rect 122285 8619 122343 8625
rect 122285 8616 122297 8619
rect 121328 8588 122297 8616
rect 121328 8576 121334 8588
rect 122285 8585 122297 8588
rect 122331 8585 122343 8619
rect 124674 8616 124680 8628
rect 124635 8588 124680 8616
rect 122285 8579 122343 8585
rect 124674 8576 124680 8588
rect 124732 8576 124738 8628
rect 128078 8616 128084 8628
rect 128039 8588 128084 8616
rect 128078 8576 128084 8588
rect 128136 8576 128142 8628
rect 139673 8619 139731 8625
rect 139673 8585 139685 8619
rect 139719 8616 139731 8619
rect 141602 8616 141608 8628
rect 139719 8588 141608 8616
rect 139719 8585 139731 8588
rect 139673 8579 139731 8585
rect 141602 8576 141608 8588
rect 141660 8616 141666 8628
rect 142157 8619 142215 8625
rect 142157 8616 142169 8619
rect 141660 8588 142169 8616
rect 141660 8576 141666 8588
rect 142157 8585 142169 8588
rect 142203 8585 142215 8619
rect 142157 8579 142215 8585
rect 142246 8576 142252 8628
rect 142304 8616 142310 8628
rect 145098 8616 145104 8628
rect 142304 8588 145104 8616
rect 142304 8576 142310 8588
rect 145098 8576 145104 8588
rect 145156 8576 145162 8628
rect 145285 8619 145343 8625
rect 145285 8585 145297 8619
rect 145331 8616 145343 8619
rect 146294 8616 146300 8628
rect 145331 8588 146300 8616
rect 145331 8585 145343 8588
rect 145285 8579 145343 8585
rect 146294 8576 146300 8588
rect 146352 8576 146358 8628
rect 152734 8576 152740 8628
rect 152792 8616 152798 8628
rect 153930 8616 153936 8628
rect 152792 8588 153936 8616
rect 152792 8576 152798 8588
rect 153930 8576 153936 8588
rect 153988 8576 153994 8628
rect 157150 8576 157156 8628
rect 157208 8616 157214 8628
rect 157613 8619 157671 8625
rect 157613 8616 157625 8619
rect 157208 8588 157625 8616
rect 157208 8576 157214 8588
rect 157613 8585 157625 8588
rect 157659 8585 157671 8619
rect 157613 8579 157671 8585
rect 161658 8576 161664 8628
rect 161716 8616 161722 8628
rect 164786 8616 164792 8628
rect 161716 8588 164792 8616
rect 161716 8576 161722 8588
rect 164786 8576 164792 8588
rect 164844 8576 164850 8628
rect 120902 8548 120908 8560
rect 102744 8520 113864 8548
rect 113928 8520 120908 8548
rect 102744 8508 102750 8520
rect 98457 8443 98515 8449
rect 98564 8452 99604 8480
rect 100021 8483 100079 8489
rect 96614 8372 96620 8424
rect 96672 8412 96678 8424
rect 98564 8412 98592 8452
rect 100021 8449 100033 8483
rect 100067 8480 100079 8483
rect 100294 8480 100300 8492
rect 100067 8452 100300 8480
rect 100067 8449 100079 8452
rect 100021 8443 100079 8449
rect 100294 8440 100300 8452
rect 100352 8440 100358 8492
rect 102870 8440 102876 8492
rect 102928 8480 102934 8492
rect 103057 8483 103115 8489
rect 103057 8480 103069 8483
rect 102928 8452 103069 8480
rect 102928 8440 102934 8452
rect 103057 8449 103069 8452
rect 103103 8449 103115 8483
rect 103057 8443 103115 8449
rect 103974 8440 103980 8492
rect 104032 8480 104038 8492
rect 104618 8480 104624 8492
rect 104032 8452 104480 8480
rect 104579 8452 104624 8480
rect 104032 8440 104038 8452
rect 96672 8384 98592 8412
rect 99469 8415 99527 8421
rect 96672 8372 96678 8384
rect 99469 8381 99481 8415
rect 99515 8381 99527 8415
rect 104069 8415 104127 8421
rect 104069 8412 104081 8415
rect 99469 8375 99527 8381
rect 99576 8384 104081 8412
rect 97353 8347 97411 8353
rect 97353 8344 97365 8347
rect 96172 8316 97365 8344
rect 97353 8313 97365 8316
rect 97399 8313 97411 8347
rect 97353 8307 97411 8313
rect 98089 8347 98147 8353
rect 98089 8313 98101 8347
rect 98135 8344 98147 8347
rect 99484 8344 99512 8375
rect 98135 8316 99512 8344
rect 98135 8313 98147 8316
rect 98089 8307 98147 8313
rect 55858 8276 55864 8288
rect 54496 8248 55864 8276
rect 55858 8236 55864 8248
rect 55916 8236 55922 8288
rect 56134 8236 56140 8288
rect 56192 8276 56198 8288
rect 57238 8276 57244 8288
rect 56192 8248 57244 8276
rect 56192 8236 56198 8248
rect 57238 8236 57244 8248
rect 57296 8236 57302 8288
rect 57422 8236 57428 8288
rect 57480 8276 57486 8288
rect 60826 8276 60832 8288
rect 57480 8248 60832 8276
rect 57480 8236 57486 8248
rect 60826 8236 60832 8248
rect 60884 8236 60890 8288
rect 61010 8276 61016 8288
rect 60971 8248 61016 8276
rect 61010 8236 61016 8248
rect 61068 8236 61074 8288
rect 79410 8236 79416 8288
rect 79468 8276 79474 8288
rect 79505 8279 79563 8285
rect 79505 8276 79517 8279
rect 79468 8248 79517 8276
rect 79468 8236 79474 8248
rect 79505 8245 79517 8248
rect 79551 8245 79563 8279
rect 83826 8276 83832 8288
rect 83787 8248 83832 8276
rect 79505 8239 79563 8245
rect 83826 8236 83832 8248
rect 83884 8236 83890 8288
rect 87506 8276 87512 8288
rect 87467 8248 87512 8276
rect 87506 8236 87512 8248
rect 87564 8236 87570 8288
rect 97994 8276 98000 8288
rect 97955 8248 98000 8276
rect 97994 8236 98000 8248
rect 98052 8236 98058 8288
rect 99374 8236 99380 8288
rect 99432 8276 99438 8288
rect 99576 8276 99604 8384
rect 104069 8381 104081 8384
rect 104115 8381 104127 8415
rect 104452 8412 104480 8452
rect 104618 8440 104624 8452
rect 104676 8440 104682 8492
rect 106458 8440 106464 8492
rect 106516 8480 106522 8492
rect 107102 8480 107108 8492
rect 106516 8452 107108 8480
rect 106516 8440 106522 8452
rect 107102 8440 107108 8452
rect 107160 8440 107166 8492
rect 108482 8480 108488 8492
rect 108040 8452 108252 8480
rect 108443 8452 108488 8480
rect 108040 8412 108068 8452
rect 104452 8384 108068 8412
rect 108117 8415 108175 8421
rect 104069 8375 104127 8381
rect 108117 8381 108129 8415
rect 108163 8381 108175 8415
rect 108224 8412 108252 8452
rect 108482 8440 108488 8452
rect 108540 8440 108546 8492
rect 113928 8480 113956 8520
rect 120902 8508 120908 8520
rect 120960 8508 120966 8560
rect 127066 8548 127072 8560
rect 126808 8520 127072 8548
rect 111076 8452 113956 8480
rect 114373 8483 114431 8489
rect 111076 8412 111104 8452
rect 114373 8449 114385 8483
rect 114419 8480 114431 8483
rect 115842 8480 115848 8492
rect 114419 8452 115848 8480
rect 114419 8449 114431 8452
rect 114373 8443 114431 8449
rect 115842 8440 115848 8452
rect 115900 8440 115906 8492
rect 118510 8440 118516 8492
rect 118568 8480 118574 8492
rect 121178 8480 121184 8492
rect 118568 8452 121184 8480
rect 118568 8440 118574 8452
rect 121178 8440 121184 8452
rect 121236 8440 121242 8492
rect 121362 8480 121368 8492
rect 121323 8452 121368 8480
rect 121362 8440 121368 8452
rect 121420 8440 121426 8492
rect 125686 8480 125692 8492
rect 125647 8452 125692 8480
rect 125686 8440 125692 8452
rect 125744 8440 125750 8492
rect 126808 8489 126836 8520
rect 127066 8508 127072 8520
rect 127124 8508 127130 8560
rect 138106 8508 138112 8560
rect 138164 8548 138170 8560
rect 138164 8520 144040 8548
rect 138164 8508 138170 8520
rect 126793 8483 126851 8489
rect 126793 8449 126805 8483
rect 126839 8449 126851 8483
rect 131022 8480 131028 8492
rect 126793 8443 126851 8449
rect 126900 8452 130608 8480
rect 130983 8452 131028 8480
rect 108224 8384 111104 8412
rect 113361 8415 113419 8421
rect 108117 8375 108175 8381
rect 113361 8381 113373 8415
rect 113407 8412 113419 8415
rect 113450 8412 113456 8424
rect 113407 8384 113456 8412
rect 113407 8381 113419 8384
rect 113361 8375 113419 8381
rect 100294 8344 100300 8356
rect 100255 8316 100300 8344
rect 100294 8304 100300 8316
rect 100352 8304 100358 8356
rect 101214 8304 101220 8356
rect 101272 8344 101278 8356
rect 108132 8344 108160 8375
rect 113450 8372 113456 8384
rect 113508 8372 113514 8424
rect 115937 8415 115995 8421
rect 115937 8381 115949 8415
rect 115983 8412 115995 8415
rect 116397 8415 116455 8421
rect 116397 8412 116409 8415
rect 115983 8384 116409 8412
rect 115983 8381 115995 8384
rect 115937 8375 115995 8381
rect 116397 8381 116409 8384
rect 116443 8412 116455 8415
rect 116578 8412 116584 8424
rect 116443 8384 116584 8412
rect 116443 8381 116455 8384
rect 116397 8375 116455 8381
rect 116578 8372 116584 8384
rect 116636 8372 116642 8424
rect 119890 8412 119896 8424
rect 119851 8384 119896 8412
rect 119890 8372 119896 8384
rect 119948 8372 119954 8424
rect 120902 8412 120908 8424
rect 120863 8384 120908 8412
rect 120902 8372 120908 8384
rect 120960 8372 120966 8424
rect 120994 8372 121000 8424
rect 121052 8412 121058 8424
rect 125962 8412 125968 8424
rect 121052 8384 125968 8412
rect 121052 8372 121058 8384
rect 125962 8372 125968 8384
rect 126020 8372 126026 8424
rect 126698 8412 126704 8424
rect 126659 8384 126704 8412
rect 126698 8372 126704 8384
rect 126756 8372 126762 8424
rect 113269 8347 113327 8353
rect 101272 8316 108160 8344
rect 112088 8316 112392 8344
rect 101272 8304 101278 8316
rect 99432 8248 99604 8276
rect 99432 8236 99438 8248
rect 102318 8236 102324 8288
rect 102376 8276 102382 8288
rect 108574 8276 108580 8288
rect 102376 8248 108580 8276
rect 102376 8236 102382 8248
rect 108574 8236 108580 8248
rect 108632 8236 108638 8288
rect 109770 8236 109776 8288
rect 109828 8276 109834 8288
rect 112088 8276 112116 8316
rect 112254 8276 112260 8288
rect 109828 8248 112116 8276
rect 112215 8248 112260 8276
rect 109828 8236 109834 8248
rect 112254 8236 112260 8248
rect 112312 8236 112318 8288
rect 112364 8276 112392 8316
rect 113269 8313 113281 8347
rect 113315 8344 113327 8347
rect 126900 8344 126928 8452
rect 129550 8412 129556 8424
rect 129511 8384 129556 8412
rect 129550 8372 129556 8384
rect 129608 8372 129614 8424
rect 130580 8421 130608 8452
rect 131022 8440 131028 8452
rect 131080 8440 131086 8492
rect 139210 8440 139216 8492
rect 139268 8480 139274 8492
rect 142341 8483 142399 8489
rect 139268 8452 141924 8480
rect 139268 8440 139274 8452
rect 130565 8415 130623 8421
rect 130565 8381 130577 8415
rect 130611 8381 130623 8415
rect 130565 8375 130623 8381
rect 132681 8415 132739 8421
rect 132681 8381 132693 8415
rect 132727 8381 132739 8415
rect 132681 8375 132739 8381
rect 141329 8415 141387 8421
rect 141329 8381 141341 8415
rect 141375 8412 141387 8415
rect 141786 8412 141792 8424
rect 141375 8384 141792 8412
rect 141375 8381 141387 8384
rect 141329 8375 141387 8381
rect 113315 8316 126928 8344
rect 113315 8313 113327 8316
rect 113269 8307 113327 8313
rect 115842 8276 115848 8288
rect 112364 8248 115848 8276
rect 115842 8236 115848 8248
rect 115900 8236 115906 8288
rect 116486 8236 116492 8288
rect 116544 8276 116550 8288
rect 131206 8276 131212 8288
rect 116544 8248 131212 8276
rect 116544 8236 116550 8248
rect 131206 8236 131212 8248
rect 131264 8236 131270 8288
rect 132696 8276 132724 8375
rect 141786 8372 141792 8384
rect 141844 8372 141850 8424
rect 141896 8412 141924 8452
rect 142341 8449 142353 8483
rect 142387 8480 142399 8483
rect 142430 8480 142436 8492
rect 142387 8452 142436 8480
rect 142387 8449 142399 8452
rect 142341 8443 142399 8449
rect 142430 8440 142436 8452
rect 142488 8480 142494 8492
rect 143350 8480 143356 8492
rect 142488 8452 143356 8480
rect 142488 8440 142494 8452
rect 143350 8440 143356 8452
rect 143408 8440 143414 8492
rect 143902 8480 143908 8492
rect 143863 8452 143908 8480
rect 143902 8440 143908 8452
rect 143960 8440 143966 8492
rect 144012 8480 144040 8520
rect 146846 8508 146852 8560
rect 146904 8548 146910 8560
rect 153010 8548 153016 8560
rect 146904 8520 153016 8548
rect 146904 8508 146910 8520
rect 153010 8508 153016 8520
rect 153068 8508 153074 8560
rect 154206 8508 154212 8560
rect 154264 8548 154270 8560
rect 155310 8548 155316 8560
rect 154264 8520 155316 8548
rect 154264 8508 154270 8520
rect 155310 8508 155316 8520
rect 155368 8508 155374 8560
rect 157518 8508 157524 8560
rect 157576 8548 157582 8560
rect 159358 8548 159364 8560
rect 157576 8520 159364 8548
rect 157576 8508 157582 8520
rect 159358 8508 159364 8520
rect 159416 8508 159422 8560
rect 160094 8508 160100 8560
rect 160152 8548 160158 8560
rect 162394 8548 162400 8560
rect 160152 8520 162400 8548
rect 160152 8508 160158 8520
rect 162394 8508 162400 8520
rect 162452 8508 162458 8560
rect 162762 8508 162768 8560
rect 162820 8548 162826 8560
rect 165154 8548 165160 8560
rect 162820 8520 165160 8548
rect 162820 8508 162826 8520
rect 165154 8508 165160 8520
rect 165212 8508 165218 8560
rect 146202 8480 146208 8492
rect 144012 8452 146208 8480
rect 146202 8440 146208 8452
rect 146260 8440 146266 8492
rect 146386 8489 146392 8492
rect 146384 8443 146392 8489
rect 146444 8480 146450 8492
rect 147766 8480 147772 8492
rect 146444 8452 146484 8480
rect 147727 8452 147772 8480
rect 146386 8440 146392 8443
rect 146444 8440 146450 8452
rect 147766 8440 147772 8452
rect 147824 8480 147830 8492
rect 148229 8483 148287 8489
rect 148229 8480 148241 8483
rect 147824 8452 148241 8480
rect 147824 8440 147830 8452
rect 148229 8449 148241 8452
rect 148275 8449 148287 8483
rect 148229 8443 148287 8449
rect 150805 8483 150863 8489
rect 150805 8449 150817 8483
rect 150851 8480 150863 8483
rect 151170 8480 151176 8492
rect 150851 8452 151176 8480
rect 150851 8449 150863 8452
rect 150805 8443 150863 8449
rect 151170 8440 151176 8452
rect 151228 8440 151234 8492
rect 152369 8483 152427 8489
rect 152369 8449 152381 8483
rect 152415 8480 152427 8483
rect 152458 8480 152464 8492
rect 152415 8452 152464 8480
rect 152415 8449 152427 8452
rect 152369 8443 152427 8449
rect 152458 8440 152464 8452
rect 152516 8480 152522 8492
rect 153194 8480 153200 8492
rect 152516 8452 153200 8480
rect 152516 8440 152522 8452
rect 153194 8440 153200 8452
rect 153252 8440 153258 8492
rect 153933 8483 153991 8489
rect 153933 8449 153945 8483
rect 153979 8480 153991 8483
rect 154761 8483 154819 8489
rect 153979 8452 154344 8480
rect 153979 8449 153991 8452
rect 153933 8443 153991 8449
rect 143537 8415 143595 8421
rect 143537 8412 143549 8415
rect 141896 8384 143549 8412
rect 143537 8381 143549 8384
rect 143583 8381 143595 8415
rect 147401 8415 147459 8421
rect 147401 8412 147413 8415
rect 143537 8375 143595 8381
rect 144840 8384 147413 8412
rect 140590 8304 140596 8356
rect 140648 8344 140654 8356
rect 142798 8344 142804 8356
rect 140648 8316 142804 8344
rect 140648 8304 140654 8316
rect 142798 8304 142804 8316
rect 142856 8304 142862 8356
rect 143258 8304 143264 8356
rect 143316 8344 143322 8356
rect 144840 8344 144868 8384
rect 147401 8381 147413 8384
rect 147447 8381 147459 8415
rect 149238 8412 149244 8424
rect 149199 8384 149244 8412
rect 147401 8375 147459 8381
rect 149238 8372 149244 8384
rect 149296 8372 149302 8424
rect 150526 8412 150532 8424
rect 150487 8384 150532 8412
rect 150526 8372 150532 8384
rect 150584 8372 150590 8424
rect 153102 8372 153108 8424
rect 153160 8412 153166 8424
rect 153381 8415 153439 8421
rect 153381 8412 153393 8415
rect 153160 8384 153393 8412
rect 153160 8372 153166 8384
rect 153381 8381 153393 8384
rect 153427 8381 153439 8415
rect 153381 8375 153439 8381
rect 154316 8356 154344 8452
rect 154761 8449 154773 8483
rect 154807 8480 154819 8483
rect 154850 8480 154856 8492
rect 154807 8452 154856 8480
rect 154807 8449 154819 8452
rect 154761 8443 154819 8449
rect 154850 8440 154856 8452
rect 154908 8440 154914 8492
rect 156046 8480 156052 8492
rect 156007 8452 156052 8480
rect 156046 8440 156052 8452
rect 156104 8480 156110 8492
rect 156601 8483 156659 8489
rect 156601 8480 156613 8483
rect 156104 8452 156613 8480
rect 156104 8440 156110 8452
rect 156601 8449 156613 8452
rect 156647 8449 156659 8483
rect 156601 8443 156659 8449
rect 158990 8440 158996 8492
rect 159048 8480 159054 8492
rect 160738 8480 160744 8492
rect 159048 8452 160508 8480
rect 160699 8452 160744 8480
rect 159048 8440 159054 8452
rect 155402 8372 155408 8424
rect 155460 8412 155466 8424
rect 155957 8415 156015 8421
rect 155957 8412 155969 8415
rect 155460 8384 155969 8412
rect 155460 8372 155466 8384
rect 155957 8381 155969 8384
rect 156003 8381 156015 8415
rect 159450 8412 159456 8424
rect 159411 8384 159456 8412
rect 155957 8375 156015 8381
rect 159450 8372 159456 8384
rect 159508 8372 159514 8424
rect 160480 8421 160508 8452
rect 160738 8440 160744 8452
rect 160796 8440 160802 8492
rect 163774 8440 163780 8492
rect 163832 8480 163838 8492
rect 164694 8480 164700 8492
rect 163832 8452 164700 8480
rect 163832 8440 163838 8452
rect 164694 8440 164700 8452
rect 164752 8440 164758 8492
rect 165614 8480 165620 8492
rect 165575 8452 165620 8480
rect 165614 8440 165620 8452
rect 165672 8440 165678 8492
rect 160465 8415 160523 8421
rect 160465 8381 160477 8415
rect 160511 8381 160523 8415
rect 160465 8375 160523 8381
rect 161106 8372 161112 8424
rect 161164 8412 161170 8424
rect 161385 8415 161443 8421
rect 161385 8412 161397 8415
rect 161164 8384 161397 8412
rect 161164 8372 161170 8384
rect 161385 8381 161397 8384
rect 161431 8412 161443 8415
rect 161845 8415 161903 8421
rect 161845 8412 161857 8415
rect 161431 8384 161857 8412
rect 161431 8381 161443 8384
rect 161385 8375 161443 8381
rect 161845 8381 161857 8384
rect 161891 8381 161903 8415
rect 161845 8375 161903 8381
rect 163501 8415 163559 8421
rect 163501 8381 163513 8415
rect 163547 8412 163559 8415
rect 164513 8415 164571 8421
rect 164513 8412 164525 8415
rect 163547 8384 164525 8412
rect 163547 8381 163559 8384
rect 163501 8375 163559 8381
rect 164513 8381 164525 8384
rect 164559 8412 164571 8415
rect 166166 8412 166172 8424
rect 164559 8384 166172 8412
rect 164559 8381 164571 8384
rect 164513 8375 164571 8381
rect 166166 8372 166172 8384
rect 166224 8372 166230 8424
rect 143316 8316 144868 8344
rect 143316 8304 143322 8316
rect 145190 8304 145196 8356
rect 145248 8344 145254 8356
rect 150894 8344 150900 8356
rect 145248 8316 150900 8344
rect 145248 8304 145254 8316
rect 150894 8304 150900 8316
rect 150952 8304 150958 8356
rect 154298 8344 154304 8356
rect 154259 8316 154304 8344
rect 154298 8304 154304 8316
rect 154356 8304 154362 8356
rect 155034 8304 155040 8356
rect 155092 8344 155098 8356
rect 156506 8344 156512 8356
rect 155092 8316 156512 8344
rect 155092 8304 155098 8316
rect 156506 8304 156512 8316
rect 156564 8304 156570 8356
rect 158530 8344 158536 8356
rect 158491 8316 158536 8344
rect 158530 8304 158536 8316
rect 158588 8304 158594 8356
rect 159726 8304 159732 8356
rect 159784 8344 159790 8356
rect 162118 8344 162124 8356
rect 159784 8316 162124 8344
rect 159784 8304 159790 8316
rect 162118 8304 162124 8316
rect 162176 8304 162182 8356
rect 164602 8304 164608 8356
rect 164660 8344 164666 8356
rect 165801 8347 165859 8353
rect 165801 8344 165813 8347
rect 164660 8316 165813 8344
rect 164660 8304 164666 8316
rect 165801 8313 165813 8316
rect 165847 8313 165859 8347
rect 165801 8307 165859 8313
rect 133046 8276 133052 8288
rect 132696 8248 133052 8276
rect 133046 8236 133052 8248
rect 133104 8276 133110 8288
rect 133141 8279 133199 8285
rect 133141 8276 133153 8279
rect 133104 8248 133153 8276
rect 133104 8236 133110 8248
rect 133141 8245 133153 8248
rect 133187 8245 133199 8279
rect 145006 8276 145012 8288
rect 144967 8248 145012 8276
rect 133141 8239 133199 8245
rect 145006 8236 145012 8248
rect 145064 8236 145070 8288
rect 151170 8276 151176 8288
rect 151131 8248 151176 8276
rect 151170 8236 151176 8248
rect 151228 8236 151234 8288
rect 368 8186 169556 8208
rect 368 8134 28456 8186
rect 28508 8134 28520 8186
rect 28572 8134 28584 8186
rect 28636 8134 28648 8186
rect 28700 8134 84878 8186
rect 84930 8134 84942 8186
rect 84994 8134 85006 8186
rect 85058 8134 85070 8186
rect 85122 8134 141299 8186
rect 141351 8134 141363 8186
rect 141415 8134 141427 8186
rect 141479 8134 141491 8186
rect 141543 8134 169556 8186
rect 368 8112 169556 8134
rect 750 8032 756 8084
rect 808 8072 814 8084
rect 8018 8072 8024 8084
rect 808 8044 8024 8072
rect 808 8032 814 8044
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 15838 8072 15844 8084
rect 15799 8044 15844 8072
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 16666 8072 16672 8084
rect 16579 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8072 16730 8084
rect 17678 8072 17684 8084
rect 16724 8044 17684 8072
rect 16724 8032 16730 8044
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 18049 8075 18107 8081
rect 18049 8041 18061 8075
rect 18095 8072 18107 8075
rect 18138 8072 18144 8084
rect 18095 8044 18144 8072
rect 18095 8041 18107 8044
rect 18049 8035 18107 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 18322 8072 18328 8084
rect 18283 8044 18328 8072
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 20346 8032 20352 8084
rect 20404 8072 20410 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 20404 8044 20545 8072
rect 20404 8032 20410 8044
rect 20533 8041 20545 8044
rect 20579 8041 20591 8075
rect 21818 8072 21824 8084
rect 21779 8044 21824 8072
rect 20533 8035 20591 8041
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 23658 8032 23664 8084
rect 23716 8072 23722 8084
rect 23937 8075 23995 8081
rect 23937 8072 23949 8075
rect 23716 8044 23949 8072
rect 23716 8032 23722 8044
rect 23937 8041 23949 8044
rect 23983 8041 23995 8075
rect 25130 8072 25136 8084
rect 25091 8044 25136 8072
rect 23937 8035 23995 8041
rect 25130 8032 25136 8044
rect 25188 8032 25194 8084
rect 25590 8072 25596 8084
rect 25551 8044 25596 8072
rect 25590 8032 25596 8044
rect 25648 8032 25654 8084
rect 26050 8032 26056 8084
rect 26108 8072 26114 8084
rect 26510 8072 26516 8084
rect 26108 8044 26516 8072
rect 26108 8032 26114 8044
rect 26510 8032 26516 8044
rect 26568 8032 26574 8084
rect 26605 8075 26663 8081
rect 26605 8041 26617 8075
rect 26651 8072 26663 8075
rect 26881 8075 26939 8081
rect 26881 8072 26893 8075
rect 26651 8044 26893 8072
rect 26651 8041 26663 8044
rect 26605 8035 26663 8041
rect 26881 8041 26893 8044
rect 26927 8072 26939 8075
rect 34606 8072 34612 8084
rect 26927 8044 34612 8072
rect 26927 8041 26939 8044
rect 26881 8035 26939 8041
rect 34606 8032 34612 8044
rect 34664 8032 34670 8084
rect 34790 8072 34796 8084
rect 34751 8044 34796 8072
rect 34790 8032 34796 8044
rect 34848 8032 34854 8084
rect 35526 8072 35532 8084
rect 35487 8044 35532 8072
rect 35526 8032 35532 8044
rect 35584 8032 35590 8084
rect 35894 8032 35900 8084
rect 35952 8072 35958 8084
rect 39206 8072 39212 8084
rect 35952 8044 39212 8072
rect 35952 8032 35958 8044
rect 39206 8032 39212 8044
rect 39264 8032 39270 8084
rect 39390 8072 39396 8084
rect 39351 8044 39396 8072
rect 39390 8032 39396 8044
rect 39448 8032 39454 8084
rect 39485 8075 39543 8081
rect 39485 8041 39497 8075
rect 39531 8072 39543 8075
rect 39945 8075 40003 8081
rect 39945 8072 39957 8075
rect 39531 8044 39957 8072
rect 39531 8041 39543 8044
rect 39485 8035 39543 8041
rect 39945 8041 39957 8044
rect 39991 8041 40003 8075
rect 39945 8035 40003 8041
rect 40034 8032 40040 8084
rect 40092 8072 40098 8084
rect 40770 8072 40776 8084
rect 40092 8044 40776 8072
rect 40092 8032 40098 8044
rect 40770 8032 40776 8044
rect 40828 8032 40834 8084
rect 40880 8044 41552 8072
rect 2777 8007 2835 8013
rect 2777 7973 2789 8007
rect 2823 8004 2835 8007
rect 3602 8004 3608 8016
rect 2823 7976 3608 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 3602 7964 3608 7976
rect 3660 8004 3666 8016
rect 3660 7976 6040 8004
rect 3660 7964 3666 7976
rect 4614 7936 4620 7948
rect 4575 7908 4620 7936
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 6012 7945 6040 7976
rect 6086 7964 6092 8016
rect 6144 8004 6150 8016
rect 12250 8004 12256 8016
rect 6144 7976 12256 8004
rect 6144 7964 6150 7976
rect 12250 7964 12256 7976
rect 12308 7964 12314 8016
rect 14090 7964 14096 8016
rect 14148 8004 14154 8016
rect 25498 8004 25504 8016
rect 14148 7976 25504 8004
rect 14148 7964 14154 7976
rect 25498 7964 25504 7976
rect 25556 7964 25562 8016
rect 25866 8004 25872 8016
rect 25827 7976 25872 8004
rect 25866 7964 25872 7976
rect 25924 7964 25930 8016
rect 26142 7964 26148 8016
rect 26200 8004 26206 8016
rect 40880 8004 40908 8044
rect 41230 8004 41236 8016
rect 26200 7976 40908 8004
rect 41191 7976 41236 8004
rect 26200 7964 26206 7976
rect 41230 7964 41236 7976
rect 41288 7964 41294 8016
rect 41524 8004 41552 8044
rect 41598 8032 41604 8084
rect 41656 8072 41662 8084
rect 44726 8072 44732 8084
rect 41656 8044 44732 8072
rect 41656 8032 41662 8044
rect 44726 8032 44732 8044
rect 44784 8032 44790 8084
rect 44818 8032 44824 8084
rect 44876 8072 44882 8084
rect 49786 8072 49792 8084
rect 44876 8044 49792 8072
rect 44876 8032 44882 8044
rect 49786 8032 49792 8044
rect 49844 8032 49850 8084
rect 49970 8072 49976 8084
rect 49931 8044 49976 8072
rect 49970 8032 49976 8044
rect 50028 8032 50034 8084
rect 50154 8032 50160 8084
rect 50212 8072 50218 8084
rect 51902 8072 51908 8084
rect 50212 8044 51908 8072
rect 50212 8032 50218 8044
rect 51902 8032 51908 8044
rect 51960 8032 51966 8084
rect 52730 8032 52736 8084
rect 52788 8072 52794 8084
rect 53006 8072 53012 8084
rect 52788 8044 52833 8072
rect 52967 8044 53012 8072
rect 52788 8032 52794 8044
rect 53006 8032 53012 8044
rect 53064 8032 53070 8084
rect 55674 8072 55680 8084
rect 55635 8044 55680 8072
rect 55674 8032 55680 8044
rect 55732 8032 55738 8084
rect 56870 8072 56876 8084
rect 55784 8044 56876 8072
rect 41524 7976 46796 8004
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7936 15163 7939
rect 15838 7936 15844 7948
rect 15151 7908 15844 7936
rect 15151 7905 15163 7908
rect 15105 7899 15163 7905
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 16114 7936 16120 7948
rect 16075 7908 16120 7936
rect 16114 7896 16120 7908
rect 16172 7896 16178 7948
rect 19613 7939 19671 7945
rect 19613 7936 19625 7939
rect 19260 7908 19625 7936
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 5169 7871 5227 7877
rect 3660 7840 3705 7868
rect 3660 7828 3666 7840
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 14826 7868 14832 7880
rect 14739 7840 14832 7868
rect 5169 7831 5227 7837
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7732 2283 7735
rect 3053 7735 3111 7741
rect 3053 7732 3065 7735
rect 2271 7704 3065 7732
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 3053 7701 3065 7704
rect 3099 7732 3111 7735
rect 3602 7732 3608 7744
rect 3099 7704 3608 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 5184 7732 5212 7831
rect 14826 7828 14832 7840
rect 14884 7868 14890 7880
rect 17586 7868 17592 7880
rect 14884 7840 17592 7868
rect 14884 7828 14890 7840
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 18598 7868 18604 7880
rect 18559 7840 18604 7868
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 18874 7868 18880 7880
rect 18835 7840 18880 7868
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19260 7877 19288 7908
rect 19613 7905 19625 7908
rect 19659 7936 19671 7939
rect 21634 7936 21640 7948
rect 19659 7908 21640 7936
rect 19659 7905 19671 7908
rect 19613 7899 19671 7905
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 22278 7896 22284 7948
rect 22336 7936 22342 7948
rect 23109 7939 23167 7945
rect 23109 7936 23121 7939
rect 22336 7908 23121 7936
rect 22336 7896 22342 7908
rect 23109 7905 23121 7908
rect 23155 7905 23167 7939
rect 23109 7899 23167 7905
rect 23382 7896 23388 7948
rect 23440 7896 23446 7948
rect 27341 7939 27399 7945
rect 27341 7936 27353 7939
rect 25884 7908 27353 7936
rect 19245 7871 19303 7877
rect 19245 7837 19257 7871
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 21726 7868 21732 7880
rect 21223 7840 21732 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 17497 7803 17555 7809
rect 17497 7769 17509 7803
rect 17543 7800 17555 7803
rect 20456 7800 20484 7831
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 22094 7868 22100 7880
rect 22007 7840 22100 7868
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 23400 7868 23428 7896
rect 23661 7871 23719 7877
rect 23661 7868 23673 7871
rect 23400 7840 23673 7868
rect 23661 7837 23673 7840
rect 23707 7868 23719 7871
rect 23934 7868 23940 7880
rect 23707 7840 23940 7868
rect 23707 7837 23719 7840
rect 23661 7831 23719 7837
rect 23934 7828 23940 7840
rect 23992 7828 23998 7880
rect 25590 7868 25596 7880
rect 24596 7840 25596 7868
rect 17543 7772 20484 7800
rect 17543 7769 17555 7772
rect 17497 7763 17555 7769
rect 5534 7732 5540 7744
rect 5184 7704 5540 7732
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 8938 7732 8944 7744
rect 8899 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 13354 7732 13360 7744
rect 13315 7704 13360 7732
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 13449 7735 13507 7741
rect 13449 7701 13461 7735
rect 13495 7732 13507 7735
rect 14090 7732 14096 7744
rect 13495 7704 14096 7732
rect 13495 7701 13507 7704
rect 13449 7695 13507 7701
rect 14090 7692 14096 7704
rect 14148 7692 14154 7744
rect 14458 7692 14464 7744
rect 14516 7732 14522 7744
rect 19150 7732 19156 7744
rect 14516 7704 19156 7732
rect 14516 7692 14522 7704
rect 19150 7692 19156 7704
rect 19208 7692 19214 7744
rect 19794 7692 19800 7744
rect 19852 7732 19858 7744
rect 19889 7735 19947 7741
rect 19889 7732 19901 7735
rect 19852 7704 19901 7732
rect 19852 7692 19858 7704
rect 19889 7701 19901 7704
rect 19935 7701 19947 7735
rect 20456 7732 20484 7772
rect 20806 7760 20812 7812
rect 20864 7800 20870 7812
rect 22112 7800 22140 7828
rect 24489 7803 24547 7809
rect 24489 7800 24501 7803
rect 20864 7772 21128 7800
rect 22112 7772 24501 7800
rect 20864 7760 20870 7772
rect 20990 7732 20996 7744
rect 20456 7704 20996 7732
rect 19889 7695 19947 7701
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 21100 7732 21128 7772
rect 24489 7769 24501 7772
rect 24535 7769 24547 7803
rect 24489 7763 24547 7769
rect 24596 7732 24624 7840
rect 25590 7828 25596 7840
rect 25648 7828 25654 7880
rect 25774 7868 25780 7880
rect 25735 7840 25780 7868
rect 25774 7828 25780 7840
rect 25832 7868 25838 7880
rect 25884 7868 25912 7908
rect 27341 7905 27353 7908
rect 27387 7905 27399 7939
rect 38105 7939 38163 7945
rect 38105 7936 38117 7939
rect 27341 7899 27399 7905
rect 27448 7908 38117 7936
rect 25832 7840 25912 7868
rect 26513 7871 26571 7877
rect 25832 7828 25838 7840
rect 26513 7837 26525 7871
rect 26559 7868 26571 7871
rect 26605 7871 26663 7877
rect 26605 7868 26617 7871
rect 26559 7840 26617 7868
rect 26559 7837 26571 7840
rect 26513 7831 26571 7837
rect 26605 7837 26617 7840
rect 26651 7837 26663 7871
rect 26605 7831 26663 7837
rect 24854 7760 24860 7812
rect 24912 7800 24918 7812
rect 27448 7800 27476 7908
rect 38105 7905 38117 7908
rect 38151 7905 38163 7939
rect 38105 7899 38163 7905
rect 38212 7908 38884 7936
rect 27522 7828 27528 7880
rect 27580 7868 27586 7880
rect 35526 7868 35532 7880
rect 27580 7840 35532 7868
rect 27580 7828 27586 7840
rect 35526 7828 35532 7840
rect 35584 7828 35590 7880
rect 35897 7871 35955 7877
rect 35897 7837 35909 7871
rect 35943 7868 35955 7871
rect 36722 7868 36728 7880
rect 35943 7840 36728 7868
rect 35943 7837 35955 7840
rect 35897 7831 35955 7837
rect 36722 7828 36728 7840
rect 36780 7828 36786 7880
rect 37093 7871 37151 7877
rect 37093 7837 37105 7871
rect 37139 7837 37151 7871
rect 37093 7831 37151 7837
rect 33778 7800 33784 7812
rect 24912 7772 27476 7800
rect 27540 7772 33784 7800
rect 24912 7760 24918 7772
rect 21100 7704 24624 7732
rect 24762 7692 24768 7744
rect 24820 7732 24826 7744
rect 27540 7732 27568 7772
rect 33778 7760 33784 7772
rect 33836 7760 33842 7812
rect 33870 7760 33876 7812
rect 33928 7800 33934 7812
rect 34422 7800 34428 7812
rect 33928 7772 34428 7800
rect 33928 7760 33934 7772
rect 34422 7760 34428 7772
rect 34480 7760 34486 7812
rect 34885 7803 34943 7809
rect 34885 7769 34897 7803
rect 34931 7800 34943 7803
rect 36357 7803 36415 7809
rect 36357 7800 36369 7803
rect 34931 7772 36369 7800
rect 34931 7769 34943 7772
rect 34885 7763 34943 7769
rect 36357 7769 36369 7772
rect 36403 7800 36415 7803
rect 37108 7800 37136 7831
rect 37182 7828 37188 7880
rect 37240 7868 37246 7880
rect 38212 7868 38240 7908
rect 37240 7840 38240 7868
rect 38657 7871 38715 7877
rect 37240 7828 37246 7840
rect 38657 7837 38669 7871
rect 38703 7868 38715 7871
rect 38746 7868 38752 7880
rect 38703 7840 38752 7868
rect 38703 7837 38715 7840
rect 38657 7831 38715 7837
rect 38746 7828 38752 7840
rect 38804 7828 38810 7880
rect 38856 7868 38884 7908
rect 38930 7896 38936 7948
rect 38988 7936 38994 7948
rect 39025 7939 39083 7945
rect 39025 7936 39037 7939
rect 38988 7908 39037 7936
rect 38988 7896 38994 7908
rect 39025 7905 39037 7908
rect 39071 7936 39083 7939
rect 39666 7936 39672 7948
rect 39071 7908 39672 7936
rect 39071 7905 39083 7908
rect 39025 7899 39083 7905
rect 39666 7896 39672 7908
rect 39724 7896 39730 7948
rect 39758 7896 39764 7948
rect 39816 7936 39822 7948
rect 39816 7908 41276 7936
rect 39816 7896 39822 7908
rect 39485 7871 39543 7877
rect 39485 7868 39497 7871
rect 38856 7840 39497 7868
rect 39485 7837 39497 7840
rect 39531 7837 39543 7871
rect 39485 7831 39543 7837
rect 40129 7871 40187 7877
rect 40129 7837 40141 7871
rect 40175 7837 40187 7871
rect 40129 7831 40187 7837
rect 40589 7871 40647 7877
rect 40589 7837 40601 7871
rect 40635 7868 40647 7871
rect 40957 7871 41015 7877
rect 40957 7868 40969 7871
rect 40635 7840 40969 7868
rect 40635 7837 40647 7840
rect 40589 7831 40647 7837
rect 40957 7837 40969 7840
rect 41003 7868 41015 7871
rect 41138 7868 41144 7880
rect 41003 7840 41144 7868
rect 41003 7837 41015 7840
rect 40957 7831 41015 7837
rect 39761 7803 39819 7809
rect 36403 7772 37136 7800
rect 37200 7772 39712 7800
rect 36403 7769 36415 7772
rect 36357 7763 36415 7769
rect 24820 7704 27568 7732
rect 24820 7692 24826 7704
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 35158 7732 35164 7744
rect 27672 7704 35164 7732
rect 27672 7692 27678 7704
rect 35158 7692 35164 7704
rect 35216 7692 35222 7744
rect 36262 7692 36268 7744
rect 36320 7732 36326 7744
rect 37200 7732 37228 7772
rect 36320 7704 37228 7732
rect 36320 7692 36326 7704
rect 37458 7692 37464 7744
rect 37516 7732 37522 7744
rect 39574 7732 39580 7744
rect 37516 7704 39580 7732
rect 37516 7692 37522 7704
rect 39574 7692 39580 7704
rect 39632 7692 39638 7744
rect 39684 7732 39712 7772
rect 39761 7769 39773 7803
rect 39807 7800 39819 7803
rect 40144 7800 40172 7831
rect 41138 7828 41144 7840
rect 41196 7828 41202 7880
rect 41248 7868 41276 7908
rect 41322 7896 41328 7948
rect 41380 7936 41386 7948
rect 42613 7939 42671 7945
rect 42613 7936 42625 7939
rect 41380 7908 42625 7936
rect 41380 7896 41386 7908
rect 42613 7905 42625 7908
rect 42659 7905 42671 7939
rect 42613 7899 42671 7905
rect 42702 7896 42708 7948
rect 42760 7936 42766 7948
rect 44818 7936 44824 7948
rect 42760 7908 44824 7936
rect 42760 7896 42766 7908
rect 44818 7896 44824 7908
rect 44876 7896 44882 7948
rect 45738 7936 45744 7948
rect 45699 7908 45744 7936
rect 45738 7896 45744 7908
rect 45796 7896 45802 7948
rect 45830 7896 45836 7948
rect 45888 7936 45894 7948
rect 46768 7945 46796 7976
rect 47486 7964 47492 8016
rect 47544 8004 47550 8016
rect 48866 8004 48872 8016
rect 47544 7976 48872 8004
rect 47544 7964 47550 7976
rect 48866 7964 48872 7976
rect 48924 7964 48930 8016
rect 49329 8007 49387 8013
rect 49329 8004 49341 8007
rect 48976 7976 49341 8004
rect 46753 7939 46811 7945
rect 45888 7908 46520 7936
rect 45888 7896 45894 7908
rect 41248 7840 41368 7868
rect 41340 7800 41368 7840
rect 41414 7828 41420 7880
rect 41472 7868 41478 7880
rect 42058 7868 42064 7880
rect 41472 7840 42064 7868
rect 41472 7828 41478 7840
rect 42058 7828 42064 7840
rect 42116 7828 42122 7880
rect 46382 7868 46388 7880
rect 42168 7840 46388 7868
rect 42168 7800 42196 7840
rect 46382 7828 46388 7840
rect 46440 7828 46446 7880
rect 46492 7868 46520 7908
rect 46753 7905 46765 7939
rect 46799 7905 46811 7939
rect 46753 7899 46811 7905
rect 46934 7896 46940 7948
rect 46992 7936 46998 7948
rect 48976 7936 49004 7976
rect 49329 7973 49341 7976
rect 49375 7973 49387 8007
rect 49605 8007 49663 8013
rect 49605 8004 49617 8007
rect 49329 7967 49387 7973
rect 49436 7976 49617 8004
rect 46992 7908 49004 7936
rect 46992 7896 46998 7908
rect 49050 7896 49056 7948
rect 49108 7896 49114 7948
rect 49436 7936 49464 7976
rect 49605 7973 49617 7976
rect 49651 8004 49663 8007
rect 50062 8004 50068 8016
rect 49651 7976 50068 8004
rect 49651 7973 49663 7976
rect 49605 7967 49663 7973
rect 50062 7964 50068 7976
rect 50120 7964 50126 8016
rect 50246 7964 50252 8016
rect 50304 8004 50310 8016
rect 55784 8004 55812 8044
rect 56870 8032 56876 8044
rect 56928 8032 56934 8084
rect 57054 8032 57060 8084
rect 57112 8072 57118 8084
rect 58986 8072 58992 8084
rect 57112 8044 58664 8072
rect 58947 8044 58992 8072
rect 57112 8032 57118 8044
rect 50304 7976 55812 8004
rect 55876 7976 58572 8004
rect 50304 7964 50310 7976
rect 49252 7908 49464 7936
rect 47305 7871 47363 7877
rect 46492 7840 47072 7868
rect 46934 7800 46940 7812
rect 39807 7772 41276 7800
rect 41340 7772 42196 7800
rect 42260 7772 46940 7800
rect 39807 7769 39819 7772
rect 39761 7763 39819 7769
rect 40862 7732 40868 7744
rect 39684 7704 40868 7732
rect 40862 7692 40868 7704
rect 40920 7692 40926 7744
rect 40954 7692 40960 7744
rect 41012 7732 41018 7744
rect 41138 7732 41144 7744
rect 41012 7704 41144 7732
rect 41012 7692 41018 7704
rect 41138 7692 41144 7704
rect 41196 7692 41202 7744
rect 41248 7732 41276 7772
rect 41417 7735 41475 7741
rect 41417 7732 41429 7735
rect 41248 7704 41429 7732
rect 41417 7701 41429 7704
rect 41463 7701 41475 7735
rect 41417 7695 41475 7701
rect 41598 7692 41604 7744
rect 41656 7732 41662 7744
rect 42260 7732 42288 7772
rect 46934 7760 46940 7772
rect 46992 7760 46998 7812
rect 47044 7800 47072 7840
rect 47305 7837 47317 7871
rect 47351 7868 47363 7871
rect 47578 7868 47584 7880
rect 47351 7840 47584 7868
rect 47351 7837 47363 7840
rect 47305 7831 47363 7837
rect 47578 7828 47584 7840
rect 47636 7828 47642 7880
rect 48774 7868 48780 7880
rect 47688 7840 48636 7868
rect 48735 7840 48780 7868
rect 47688 7800 47716 7840
rect 47044 7772 47716 7800
rect 47762 7760 47768 7812
rect 47820 7800 47826 7812
rect 48498 7800 48504 7812
rect 47820 7772 48504 7800
rect 47820 7760 47826 7772
rect 48498 7760 48504 7772
rect 48556 7760 48562 7812
rect 48608 7800 48636 7840
rect 48774 7828 48780 7840
rect 48832 7828 48838 7880
rect 48869 7871 48927 7877
rect 48869 7837 48881 7871
rect 48915 7868 48927 7871
rect 49068 7868 49096 7896
rect 49252 7877 49280 7908
rect 49510 7896 49516 7948
rect 49568 7936 49574 7948
rect 55876 7936 55904 7976
rect 49568 7908 55904 7936
rect 49568 7896 49574 7908
rect 56042 7896 56048 7948
rect 56100 7936 56106 7948
rect 56100 7908 57100 7936
rect 56100 7896 56106 7908
rect 48915 7840 49096 7868
rect 49237 7871 49295 7877
rect 48915 7837 48927 7840
rect 48869 7831 48927 7837
rect 49237 7837 49249 7871
rect 49283 7837 49295 7871
rect 49970 7868 49976 7880
rect 49237 7831 49295 7837
rect 49344 7840 49976 7868
rect 49344 7800 49372 7840
rect 49970 7828 49976 7840
rect 50028 7828 50034 7880
rect 50065 7871 50123 7877
rect 50065 7837 50077 7871
rect 50111 7868 50123 7871
rect 50522 7868 50528 7880
rect 50111 7840 50528 7868
rect 50111 7837 50123 7840
rect 50065 7831 50123 7837
rect 50522 7828 50528 7840
rect 50580 7828 50586 7880
rect 51350 7868 51356 7880
rect 50632 7840 51356 7868
rect 48608 7772 49372 7800
rect 49421 7803 49479 7809
rect 49421 7769 49433 7803
rect 49467 7800 49479 7803
rect 49510 7800 49516 7812
rect 49467 7772 49516 7800
rect 49467 7769 49479 7772
rect 49421 7763 49479 7769
rect 49510 7760 49516 7772
rect 49568 7760 49574 7812
rect 49602 7760 49608 7812
rect 49660 7800 49666 7812
rect 50632 7800 50660 7840
rect 51350 7828 51356 7840
rect 51408 7828 51414 7880
rect 51534 7868 51540 7880
rect 51495 7840 51540 7868
rect 51534 7828 51540 7840
rect 51592 7828 51598 7880
rect 51718 7868 51724 7880
rect 51679 7840 51724 7868
rect 51718 7828 51724 7840
rect 51776 7828 51782 7880
rect 52086 7868 52092 7880
rect 52047 7840 52092 7868
rect 52086 7828 52092 7840
rect 52144 7828 52150 7880
rect 52270 7828 52276 7880
rect 52328 7868 52334 7880
rect 54018 7868 54024 7880
rect 52328 7840 54024 7868
rect 52328 7828 52334 7840
rect 54018 7828 54024 7840
rect 54076 7828 54082 7880
rect 54386 7868 54392 7880
rect 54347 7840 54392 7868
rect 54386 7828 54392 7840
rect 54444 7828 54450 7880
rect 54570 7868 54576 7880
rect 54531 7840 54576 7868
rect 54570 7828 54576 7840
rect 54628 7828 54634 7880
rect 54941 7871 54999 7877
rect 54941 7837 54953 7871
rect 54987 7868 54999 7871
rect 55309 7871 55367 7877
rect 55309 7868 55321 7871
rect 54987 7840 55321 7868
rect 54987 7837 54999 7840
rect 54941 7831 54999 7837
rect 55309 7837 55321 7840
rect 55355 7868 55367 7871
rect 56781 7871 56839 7877
rect 56781 7868 56793 7871
rect 55355 7840 55812 7868
rect 55355 7837 55367 7840
rect 55309 7831 55367 7837
rect 55582 7800 55588 7812
rect 49660 7772 50660 7800
rect 50724 7772 55588 7800
rect 49660 7760 49666 7772
rect 41656 7704 42288 7732
rect 41656 7692 41662 7704
rect 42334 7692 42340 7744
rect 42392 7732 42398 7744
rect 47302 7732 47308 7744
rect 42392 7704 47308 7732
rect 42392 7692 42398 7704
rect 47302 7692 47308 7704
rect 47360 7692 47366 7744
rect 47578 7732 47584 7744
rect 47539 7704 47584 7732
rect 47578 7692 47584 7704
rect 47636 7692 47642 7744
rect 47670 7692 47676 7744
rect 47728 7732 47734 7744
rect 50154 7732 50160 7744
rect 47728 7704 50160 7732
rect 47728 7692 47734 7704
rect 50154 7692 50160 7704
rect 50212 7692 50218 7744
rect 50246 7692 50252 7744
rect 50304 7732 50310 7744
rect 50724 7732 50752 7772
rect 55582 7760 55588 7772
rect 55640 7760 55646 7812
rect 55784 7800 55812 7840
rect 55968 7840 56793 7868
rect 55858 7800 55864 7812
rect 55784 7772 55864 7800
rect 55858 7760 55864 7772
rect 55916 7760 55922 7812
rect 55968 7809 55996 7840
rect 56781 7837 56793 7840
rect 56827 7868 56839 7871
rect 56965 7871 57023 7877
rect 56965 7868 56977 7871
rect 56827 7840 56977 7868
rect 56827 7837 56839 7840
rect 56781 7831 56839 7837
rect 56965 7837 56977 7840
rect 57011 7837 57023 7871
rect 57072 7868 57100 7908
rect 57330 7896 57336 7948
rect 57388 7936 57394 7948
rect 57514 7936 57520 7948
rect 57388 7908 57520 7936
rect 57388 7896 57394 7908
rect 57514 7896 57520 7908
rect 57572 7896 57578 7948
rect 57974 7936 57980 7948
rect 57935 7908 57980 7936
rect 57974 7896 57980 7908
rect 58032 7896 58038 7948
rect 58434 7936 58440 7948
rect 58084 7908 58440 7936
rect 58084 7868 58112 7908
rect 58434 7896 58440 7908
rect 58492 7896 58498 7948
rect 58342 7868 58348 7880
rect 57072 7840 58112 7868
rect 58303 7840 58348 7868
rect 56965 7831 57023 7837
rect 58342 7828 58348 7840
rect 58400 7828 58406 7880
rect 58544 7868 58572 7976
rect 58636 7936 58664 8044
rect 58986 8032 58992 8044
rect 59044 8032 59050 8084
rect 60182 8072 60188 8084
rect 60143 8044 60188 8072
rect 60182 8032 60188 8044
rect 60240 8032 60246 8084
rect 60550 8072 60556 8084
rect 60511 8044 60556 8072
rect 60550 8032 60556 8044
rect 60608 8032 60614 8084
rect 62850 8032 62856 8084
rect 62908 8072 62914 8084
rect 63129 8075 63187 8081
rect 63129 8072 63141 8075
rect 62908 8044 63141 8072
rect 62908 8032 62914 8044
rect 63129 8041 63141 8044
rect 63175 8072 63187 8075
rect 63221 8075 63279 8081
rect 63221 8072 63233 8075
rect 63175 8044 63233 8072
rect 63175 8041 63187 8044
rect 63129 8035 63187 8041
rect 63221 8041 63233 8044
rect 63267 8041 63279 8075
rect 63221 8035 63279 8041
rect 71685 8075 71743 8081
rect 71685 8041 71697 8075
rect 71731 8072 71743 8075
rect 71774 8072 71780 8084
rect 71731 8044 71780 8072
rect 71731 8041 71743 8044
rect 71685 8035 71743 8041
rect 71774 8032 71780 8044
rect 71832 8032 71838 8084
rect 87230 8072 87236 8084
rect 87191 8044 87236 8072
rect 87230 8032 87236 8044
rect 87288 8032 87294 8084
rect 92661 8075 92719 8081
rect 92661 8041 92673 8075
rect 92707 8072 92719 8075
rect 92842 8072 92848 8084
rect 92707 8044 92848 8072
rect 92707 8041 92719 8044
rect 92661 8035 92719 8041
rect 92842 8032 92848 8044
rect 92900 8032 92906 8084
rect 102870 8032 102876 8084
rect 102928 8072 102934 8084
rect 103057 8075 103115 8081
rect 103057 8072 103069 8075
rect 102928 8044 103069 8072
rect 102928 8032 102934 8044
rect 103057 8041 103069 8044
rect 103103 8041 103115 8075
rect 107102 8072 107108 8084
rect 107063 8044 107108 8072
rect 103057 8035 103115 8041
rect 107102 8032 107108 8044
rect 107160 8032 107166 8084
rect 108482 8072 108488 8084
rect 108443 8044 108488 8072
rect 108482 8032 108488 8044
rect 108540 8072 108546 8084
rect 124950 8072 124956 8084
rect 108540 8044 124956 8072
rect 108540 8032 108546 8044
rect 124950 8032 124956 8044
rect 125008 8032 125014 8084
rect 125686 8032 125692 8084
rect 125744 8072 125750 8084
rect 125965 8075 126023 8081
rect 125965 8072 125977 8075
rect 125744 8044 125977 8072
rect 125744 8032 125750 8044
rect 125965 8041 125977 8044
rect 126011 8041 126023 8075
rect 129550 8072 129556 8084
rect 125965 8035 126023 8041
rect 128740 8044 129556 8072
rect 59265 8007 59323 8013
rect 59265 7973 59277 8007
rect 59311 8004 59323 8007
rect 59311 7976 84516 8004
rect 59311 7973 59323 7976
rect 59265 7967 59323 7973
rect 61010 7936 61016 7948
rect 58636 7908 60872 7936
rect 60971 7908 61016 7936
rect 59265 7871 59323 7877
rect 59265 7868 59277 7871
rect 58544 7840 59277 7868
rect 59265 7837 59277 7840
rect 59311 7837 59323 7871
rect 59265 7831 59323 7837
rect 59354 7828 59360 7880
rect 59412 7868 59418 7880
rect 60642 7868 60648 7880
rect 59412 7840 60648 7868
rect 59412 7828 59418 7840
rect 60642 7828 60648 7840
rect 60700 7828 60706 7880
rect 55953 7803 56011 7809
rect 55953 7769 55965 7803
rect 55999 7769 56011 7803
rect 55953 7763 56011 7769
rect 57054 7760 57060 7812
rect 57112 7800 57118 7812
rect 60844 7800 60872 7908
rect 61010 7896 61016 7908
rect 61068 7896 61074 7948
rect 62114 7936 62120 7948
rect 62075 7908 62120 7936
rect 62114 7896 62120 7908
rect 62172 7896 62178 7948
rect 63129 7939 63187 7945
rect 63129 7905 63141 7939
rect 63175 7936 63187 7939
rect 63405 7939 63463 7945
rect 63405 7936 63417 7939
rect 63175 7908 63417 7936
rect 63175 7905 63187 7908
rect 63129 7899 63187 7905
rect 63405 7905 63417 7908
rect 63451 7905 63463 7939
rect 63405 7899 63463 7905
rect 64049 7939 64107 7945
rect 64049 7905 64061 7939
rect 64095 7936 64107 7939
rect 68002 7936 68008 7948
rect 64095 7908 68008 7936
rect 64095 7905 64107 7908
rect 64049 7899 64107 7905
rect 68002 7896 68008 7908
rect 68060 7896 68066 7948
rect 71774 7936 71780 7948
rect 71735 7908 71780 7936
rect 71774 7896 71780 7908
rect 71832 7896 71838 7948
rect 72786 7936 72792 7948
rect 72747 7908 72792 7936
rect 72786 7896 72792 7908
rect 72844 7896 72850 7948
rect 79410 7936 79416 7948
rect 79371 7908 79416 7936
rect 79410 7896 79416 7908
rect 79468 7896 79474 7948
rect 80422 7936 80428 7948
rect 80383 7908 80428 7936
rect 80422 7896 80428 7908
rect 80480 7896 80486 7948
rect 81897 7939 81955 7945
rect 81897 7905 81909 7939
rect 81943 7936 81955 7939
rect 81986 7936 81992 7948
rect 81943 7908 81992 7936
rect 81943 7905 81955 7908
rect 81897 7899 81955 7905
rect 81986 7896 81992 7908
rect 82044 7936 82050 7948
rect 82357 7939 82415 7945
rect 82357 7936 82369 7939
rect 82044 7908 82369 7936
rect 82044 7896 82050 7908
rect 82357 7905 82369 7908
rect 82403 7905 82415 7939
rect 82357 7899 82415 7905
rect 83366 7896 83372 7948
rect 83424 7936 83430 7948
rect 83461 7939 83519 7945
rect 83461 7936 83473 7939
rect 83424 7908 83473 7936
rect 83424 7896 83430 7908
rect 83461 7905 83473 7908
rect 83507 7936 83519 7939
rect 83826 7936 83832 7948
rect 83507 7908 83832 7936
rect 83507 7905 83519 7908
rect 83461 7899 83519 7905
rect 83826 7896 83832 7908
rect 83884 7896 83890 7948
rect 84488 7945 84516 7976
rect 89254 7964 89260 8016
rect 89312 8004 89318 8016
rect 89809 8007 89867 8013
rect 89809 8004 89821 8007
rect 89312 7976 89821 8004
rect 89312 7964 89318 7976
rect 89809 7973 89821 7976
rect 89855 8004 89867 8007
rect 101769 8007 101827 8013
rect 101769 8004 101781 8007
rect 89855 7976 101781 8004
rect 89855 7973 89867 7976
rect 89809 7967 89867 7973
rect 101769 7973 101781 7976
rect 101815 7973 101827 8007
rect 101769 7967 101827 7973
rect 101861 8007 101919 8013
rect 101861 7973 101873 8007
rect 101907 8004 101919 8007
rect 101907 7976 117360 8004
rect 101907 7973 101919 7976
rect 101861 7967 101919 7973
rect 84473 7939 84531 7945
rect 84473 7905 84485 7939
rect 84519 7905 84531 7939
rect 84473 7899 84531 7905
rect 86405 7939 86463 7945
rect 86405 7905 86417 7939
rect 86451 7936 86463 7939
rect 87506 7936 87512 7948
rect 86451 7908 87512 7936
rect 86451 7905 86463 7908
rect 86405 7899 86463 7905
rect 87506 7896 87512 7908
rect 87564 7896 87570 7948
rect 88334 7896 88340 7948
rect 88392 7936 88398 7948
rect 88521 7939 88579 7945
rect 88521 7936 88533 7939
rect 88392 7908 88533 7936
rect 88392 7896 88398 7908
rect 88521 7905 88533 7908
rect 88567 7905 88579 7939
rect 88521 7899 88579 7905
rect 89901 7939 89959 7945
rect 89901 7905 89913 7939
rect 89947 7936 89959 7939
rect 90266 7936 90272 7948
rect 89947 7908 90272 7936
rect 89947 7905 89959 7908
rect 89901 7899 89959 7905
rect 90266 7896 90272 7908
rect 90324 7896 90330 7948
rect 91094 7936 91100 7948
rect 91055 7908 91100 7936
rect 91094 7896 91100 7908
rect 91152 7896 91158 7948
rect 98454 7896 98460 7948
rect 98512 7936 98518 7948
rect 98512 7908 100340 7936
rect 98512 7896 98518 7908
rect 62577 7871 62635 7877
rect 62577 7837 62589 7871
rect 62623 7868 62635 7871
rect 62945 7871 63003 7877
rect 62945 7868 62957 7871
rect 62623 7840 62957 7868
rect 62623 7837 62635 7840
rect 62577 7831 62635 7837
rect 62945 7837 62957 7840
rect 62991 7868 63003 7871
rect 72878 7868 72884 7880
rect 62991 7840 72884 7868
rect 62991 7837 63003 7840
rect 62945 7831 63003 7837
rect 72878 7828 72884 7840
rect 72936 7828 72942 7880
rect 73341 7871 73399 7877
rect 73341 7837 73353 7871
rect 73387 7868 73399 7871
rect 80882 7868 80888 7880
rect 73387 7840 73752 7868
rect 80843 7840 80888 7868
rect 73387 7837 73399 7840
rect 73341 7831 73399 7837
rect 64049 7803 64107 7809
rect 64049 7800 64061 7803
rect 57112 7772 59584 7800
rect 60844 7772 64061 7800
rect 57112 7760 57118 7772
rect 50304 7704 50752 7732
rect 50304 7692 50310 7704
rect 50798 7692 50804 7744
rect 50856 7732 50862 7744
rect 52270 7732 52276 7744
rect 50856 7704 52276 7732
rect 50856 7692 50862 7704
rect 52270 7692 52276 7704
rect 52328 7692 52334 7744
rect 52362 7692 52368 7744
rect 52420 7732 52426 7744
rect 55766 7732 55772 7744
rect 52420 7704 55772 7732
rect 52420 7692 52426 7704
rect 55766 7692 55772 7704
rect 55824 7692 55830 7744
rect 56226 7692 56232 7744
rect 56284 7732 56290 7744
rect 56413 7735 56471 7741
rect 56413 7732 56425 7735
rect 56284 7704 56425 7732
rect 56284 7692 56290 7704
rect 56413 7701 56425 7704
rect 56459 7701 56471 7735
rect 56413 7695 56471 7701
rect 56502 7692 56508 7744
rect 56560 7732 56566 7744
rect 57238 7732 57244 7744
rect 56560 7704 57244 7732
rect 56560 7692 56566 7704
rect 57238 7692 57244 7704
rect 57296 7692 57302 7744
rect 59078 7692 59084 7744
rect 59136 7732 59142 7744
rect 59449 7735 59507 7741
rect 59449 7732 59461 7735
rect 59136 7704 59461 7732
rect 59136 7692 59142 7704
rect 59449 7701 59461 7704
rect 59495 7701 59507 7735
rect 59556 7732 59584 7772
rect 64049 7769 64061 7772
rect 64095 7769 64107 7803
rect 64049 7763 64107 7769
rect 64233 7803 64291 7809
rect 64233 7769 64245 7803
rect 64279 7800 64291 7803
rect 64414 7800 64420 7812
rect 64279 7772 64420 7800
rect 64279 7769 64291 7772
rect 64233 7763 64291 7769
rect 64414 7760 64420 7772
rect 64472 7800 64478 7812
rect 71130 7800 71136 7812
rect 64472 7772 71136 7800
rect 64472 7760 64478 7772
rect 71130 7760 71136 7772
rect 71188 7760 71194 7812
rect 67726 7732 67732 7744
rect 59556 7704 67732 7732
rect 59449 7695 59507 7701
rect 67726 7692 67732 7704
rect 67784 7692 67790 7744
rect 68830 7732 68836 7744
rect 68791 7704 68836 7732
rect 68830 7692 68836 7704
rect 68888 7692 68894 7744
rect 73724 7741 73752 7840
rect 80882 7828 80888 7840
rect 80940 7868 80946 7880
rect 81253 7871 81311 7877
rect 81253 7868 81265 7871
rect 80940 7840 81265 7868
rect 80940 7828 80946 7840
rect 81253 7837 81265 7840
rect 81299 7837 81311 7871
rect 84746 7868 84752 7880
rect 84707 7840 84752 7868
rect 81253 7831 81311 7837
rect 84746 7828 84752 7840
rect 84804 7868 84810 7880
rect 85301 7871 85359 7877
rect 85301 7868 85313 7871
rect 84804 7840 85313 7868
rect 84804 7828 84810 7840
rect 85301 7837 85313 7840
rect 85347 7837 85359 7871
rect 85301 7831 85359 7837
rect 89073 7871 89131 7877
rect 89073 7837 89085 7871
rect 89119 7837 89131 7871
rect 89073 7831 89131 7837
rect 73709 7735 73767 7741
rect 73709 7701 73721 7735
rect 73755 7732 73767 7735
rect 80146 7732 80152 7744
rect 73755 7704 80152 7732
rect 73755 7701 73767 7704
rect 73709 7695 73767 7701
rect 80146 7692 80152 7704
rect 80204 7692 80210 7744
rect 83369 7735 83427 7741
rect 83369 7701 83381 7735
rect 83415 7732 83427 7735
rect 83458 7732 83464 7744
rect 83415 7704 83464 7732
rect 83415 7701 83427 7704
rect 83369 7695 83427 7701
rect 83458 7692 83464 7704
rect 83516 7692 83522 7744
rect 89088 7732 89116 7831
rect 91278 7828 91284 7880
rect 91336 7868 91342 7880
rect 91465 7871 91523 7877
rect 91465 7868 91477 7871
rect 91336 7840 91477 7868
rect 91336 7828 91342 7840
rect 91465 7837 91477 7840
rect 91511 7868 91523 7871
rect 100205 7871 100263 7877
rect 100205 7868 100217 7871
rect 91511 7840 100217 7868
rect 91511 7837 91523 7840
rect 91465 7831 91523 7837
rect 100205 7837 100217 7840
rect 100251 7837 100263 7871
rect 100312 7868 100340 7908
rect 100386 7896 100392 7948
rect 100444 7936 100450 7948
rect 102965 7939 103023 7945
rect 102965 7936 102977 7939
rect 100444 7908 102977 7936
rect 100444 7896 100450 7908
rect 102965 7905 102977 7908
rect 103011 7905 103023 7939
rect 103330 7936 103336 7948
rect 103291 7908 103336 7936
rect 102965 7899 103023 7905
rect 103330 7896 103336 7908
rect 103388 7896 103394 7948
rect 103790 7896 103796 7948
rect 103848 7936 103854 7948
rect 110417 7939 110475 7945
rect 110417 7936 110429 7939
rect 103848 7908 110429 7936
rect 103848 7896 103854 7908
rect 110417 7905 110429 7908
rect 110463 7905 110475 7939
rect 112254 7936 112260 7948
rect 112215 7908 112260 7936
rect 110417 7899 110475 7905
rect 112254 7896 112260 7908
rect 112312 7896 112318 7948
rect 113269 7939 113327 7945
rect 113269 7905 113281 7939
rect 113315 7905 113327 7939
rect 113269 7899 113327 7905
rect 113376 7908 114048 7936
rect 113284 7868 113312 7899
rect 100312 7840 113312 7868
rect 100205 7831 100263 7837
rect 91646 7760 91652 7812
rect 91704 7800 91710 7812
rect 91833 7803 91891 7809
rect 91833 7800 91845 7803
rect 91704 7772 91845 7800
rect 91704 7760 91710 7772
rect 91833 7769 91845 7772
rect 91879 7800 91891 7803
rect 99745 7803 99803 7809
rect 99745 7800 99757 7803
rect 91879 7772 99757 7800
rect 91879 7769 91891 7772
rect 91833 7763 91891 7769
rect 99745 7769 99757 7772
rect 99791 7769 99803 7803
rect 99745 7763 99803 7769
rect 101769 7803 101827 7809
rect 101769 7769 101781 7803
rect 101815 7800 101827 7803
rect 106550 7800 106556 7812
rect 101815 7772 106556 7800
rect 101815 7769 101827 7772
rect 101769 7763 101827 7769
rect 106550 7760 106556 7772
rect 106608 7760 106614 7812
rect 110417 7803 110475 7809
rect 110417 7769 110429 7803
rect 110463 7800 110475 7803
rect 113376 7800 113404 7908
rect 113821 7871 113879 7877
rect 113821 7837 113833 7871
rect 113867 7868 113879 7871
rect 113913 7871 113971 7877
rect 113913 7868 113925 7871
rect 113867 7840 113925 7868
rect 113867 7837 113879 7840
rect 113821 7831 113879 7837
rect 113913 7837 113925 7840
rect 113959 7837 113971 7871
rect 114020 7868 114048 7908
rect 114094 7896 114100 7948
rect 114152 7936 114158 7948
rect 117332 7945 117360 7976
rect 117317 7939 117375 7945
rect 114152 7908 117268 7936
rect 114152 7896 114158 7908
rect 116118 7868 116124 7880
rect 114020 7840 116124 7868
rect 113913 7831 113971 7837
rect 116118 7828 116124 7840
rect 116176 7828 116182 7880
rect 116305 7871 116363 7877
rect 116305 7837 116317 7871
rect 116351 7837 116363 7871
rect 117240 7868 117268 7908
rect 117317 7905 117329 7939
rect 117363 7905 117375 7939
rect 117317 7899 117375 7905
rect 117424 7908 119844 7936
rect 117424 7868 117452 7908
rect 117240 7840 117452 7868
rect 117869 7871 117927 7877
rect 116305 7831 116363 7837
rect 117869 7837 117881 7871
rect 117915 7868 117927 7871
rect 118145 7871 118203 7877
rect 118145 7868 118157 7871
rect 117915 7840 118157 7868
rect 117915 7837 117927 7840
rect 117869 7831 117927 7837
rect 118145 7837 118157 7840
rect 118191 7837 118203 7871
rect 119816 7868 119844 7908
rect 119890 7896 119896 7948
rect 119948 7936 119954 7948
rect 119985 7939 120043 7945
rect 119985 7936 119997 7939
rect 119948 7908 119997 7936
rect 119948 7896 119954 7908
rect 119985 7905 119997 7908
rect 120031 7936 120043 7939
rect 120445 7939 120503 7945
rect 120445 7936 120457 7939
rect 120031 7908 120457 7936
rect 120031 7905 120043 7908
rect 119985 7899 120043 7905
rect 120445 7905 120457 7908
rect 120491 7905 120503 7939
rect 120445 7899 120503 7905
rect 125505 7939 125563 7945
rect 125505 7905 125517 7939
rect 125551 7936 125563 7939
rect 126238 7936 126244 7948
rect 125551 7908 126244 7936
rect 125551 7905 125563 7908
rect 125505 7899 125563 7905
rect 126238 7896 126244 7908
rect 126296 7896 126302 7948
rect 127437 7939 127495 7945
rect 127437 7905 127449 7939
rect 127483 7936 127495 7939
rect 127526 7936 127532 7948
rect 127483 7908 127532 7936
rect 127483 7905 127495 7908
rect 127437 7899 127495 7905
rect 127526 7896 127532 7908
rect 127584 7896 127590 7948
rect 128740 7945 128768 8044
rect 129550 8032 129556 8044
rect 129608 8032 129614 8084
rect 146386 8032 146392 8084
rect 146444 8072 146450 8084
rect 147030 8072 147036 8084
rect 146444 8044 147036 8072
rect 146444 8032 146450 8044
rect 147030 8032 147036 8044
rect 147088 8072 147094 8084
rect 147217 8075 147275 8081
rect 147217 8072 147229 8075
rect 147088 8044 147229 8072
rect 147088 8032 147094 8044
rect 147217 8041 147229 8044
rect 147263 8041 147275 8075
rect 152458 8072 152464 8084
rect 152419 8044 152464 8072
rect 147217 8035 147275 8041
rect 152458 8032 152464 8044
rect 152516 8032 152522 8084
rect 154850 8032 154856 8084
rect 154908 8072 154914 8084
rect 155221 8075 155279 8081
rect 155221 8072 155233 8075
rect 154908 8044 155233 8072
rect 154908 8032 154914 8044
rect 155221 8041 155233 8044
rect 155267 8041 155279 8075
rect 166166 8072 166172 8084
rect 166127 8044 166172 8072
rect 155221 8035 155279 8041
rect 166166 8032 166172 8044
rect 166224 8032 166230 8084
rect 131206 7964 131212 8016
rect 131264 8004 131270 8016
rect 148873 8007 148931 8013
rect 131264 7976 134104 8004
rect 131264 7964 131270 7976
rect 128725 7939 128783 7945
rect 128725 7905 128737 7939
rect 128771 7905 128783 7939
rect 129734 7936 129740 7948
rect 129695 7908 129740 7936
rect 128725 7899 128783 7905
rect 129734 7896 129740 7908
rect 129792 7896 129798 7948
rect 129826 7896 129832 7948
rect 129884 7936 129890 7948
rect 130749 7939 130807 7945
rect 130749 7936 130761 7939
rect 129884 7908 130761 7936
rect 129884 7896 129890 7908
rect 130749 7905 130761 7908
rect 130795 7905 130807 7939
rect 133046 7936 133052 7948
rect 133007 7908 133052 7936
rect 130749 7899 130807 7905
rect 133046 7896 133052 7908
rect 133104 7896 133110 7948
rect 134076 7945 134104 7976
rect 148873 7973 148885 8007
rect 148919 8004 148931 8007
rect 149422 8004 149428 8016
rect 148919 7976 149428 8004
rect 148919 7973 148931 7976
rect 148873 7967 148931 7973
rect 149422 7964 149428 7976
rect 149480 7964 149486 8016
rect 156782 8004 156788 8016
rect 156743 7976 156788 8004
rect 156782 7964 156788 7976
rect 156840 7964 156846 8016
rect 164786 8004 164792 8016
rect 164747 7976 164792 8004
rect 164786 7964 164792 7976
rect 164844 7964 164850 8016
rect 134061 7939 134119 7945
rect 134061 7905 134073 7939
rect 134107 7905 134119 7939
rect 134061 7899 134119 7905
rect 140685 7939 140743 7945
rect 140685 7905 140697 7939
rect 140731 7936 140743 7939
rect 140866 7936 140872 7948
rect 140731 7908 140872 7936
rect 140731 7905 140743 7908
rect 140685 7899 140743 7905
rect 140866 7896 140872 7908
rect 140924 7896 140930 7948
rect 141786 7936 141792 7948
rect 141747 7908 141792 7936
rect 141786 7896 141792 7908
rect 141844 7896 141850 7948
rect 142798 7936 142804 7948
rect 142759 7908 142804 7936
rect 142798 7896 142804 7908
rect 142856 7896 142862 7948
rect 145006 7936 145012 7948
rect 144967 7908 145012 7936
rect 145006 7896 145012 7908
rect 145064 7896 145070 7948
rect 145098 7896 145104 7948
rect 145156 7936 145162 7948
rect 146021 7939 146079 7945
rect 146021 7936 146033 7939
rect 145156 7908 146033 7936
rect 145156 7896 145162 7908
rect 146021 7905 146033 7908
rect 146067 7905 146079 7939
rect 146021 7899 146079 7905
rect 147122 7896 147128 7948
rect 147180 7936 147186 7948
rect 147401 7939 147459 7945
rect 147401 7936 147413 7939
rect 147180 7908 147413 7936
rect 147180 7896 147186 7908
rect 147401 7905 147413 7908
rect 147447 7905 147459 7939
rect 150894 7936 150900 7948
rect 150855 7908 150900 7936
rect 147401 7899 147459 7905
rect 150894 7896 150900 7908
rect 150952 7896 150958 7948
rect 153470 7896 153476 7948
rect 153528 7936 153534 7948
rect 154025 7939 154083 7945
rect 154025 7936 154037 7939
rect 153528 7908 154037 7936
rect 153528 7896 153534 7908
rect 154025 7905 154037 7908
rect 154071 7905 154083 7939
rect 159358 7936 159364 7948
rect 154025 7899 154083 7905
rect 156984 7908 157472 7936
rect 159319 7908 159364 7936
rect 133414 7868 133420 7880
rect 119816 7840 133420 7868
rect 118145 7831 118203 7837
rect 116210 7800 116216 7812
rect 110463 7772 113404 7800
rect 113468 7772 116216 7800
rect 110463 7769 110475 7772
rect 110417 7763 110475 7769
rect 89441 7735 89499 7741
rect 89441 7732 89453 7735
rect 89088 7704 89453 7732
rect 89441 7701 89453 7704
rect 89487 7732 89499 7735
rect 89487 7704 93072 7732
rect 89487 7701 89499 7704
rect 89441 7695 89499 7701
rect 368 7642 93012 7664
rect 368 7590 56667 7642
rect 56719 7590 56731 7642
rect 56783 7590 56795 7642
rect 56847 7590 56859 7642
rect 56911 7590 93012 7642
rect 368 7568 93012 7590
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 14458 7528 14464 7540
rect 5592 7500 14464 7528
rect 5592 7488 5598 7500
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 19150 7488 19156 7540
rect 19208 7528 19214 7540
rect 27522 7528 27528 7540
rect 19208 7500 27528 7528
rect 19208 7488 19214 7500
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 27614 7488 27620 7540
rect 27672 7528 27678 7540
rect 33962 7528 33968 7540
rect 27672 7500 33968 7528
rect 27672 7488 27678 7500
rect 33962 7488 33968 7500
rect 34020 7488 34026 7540
rect 34606 7488 34612 7540
rect 34664 7528 34670 7540
rect 40586 7528 40592 7540
rect 34664 7500 40592 7528
rect 34664 7488 34670 7500
rect 40586 7488 40592 7500
rect 40644 7488 40650 7540
rect 40678 7488 40684 7540
rect 40736 7528 40742 7540
rect 42242 7528 42248 7540
rect 40736 7500 42248 7528
rect 40736 7488 40742 7500
rect 42242 7488 42248 7500
rect 42300 7488 42306 7540
rect 42352 7500 42564 7528
rect 4062 7420 4068 7472
rect 4120 7460 4126 7472
rect 18690 7460 18696 7472
rect 4120 7432 16160 7460
rect 18651 7432 18696 7460
rect 4120 7420 4126 7432
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7392 9551 7395
rect 9582 7392 9588 7404
rect 9539 7364 9588 7392
rect 9539 7361 9551 7364
rect 9493 7355 9551 7361
rect 3602 7324 3608 7336
rect 3563 7296 3608 7324
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 4580 7296 4629 7324
rect 4580 7284 4586 7296
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 5092 7324 5120 7355
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7392 9735 7395
rect 13906 7392 13912 7404
rect 9723 7364 13912 7392
rect 9723 7361 9735 7364
rect 9677 7355 9735 7361
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 14090 7392 14096 7404
rect 14051 7364 14096 7392
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 5534 7324 5540 7336
rect 5092 7296 5540 7324
rect 4617 7287 4675 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 7926 7324 7932 7336
rect 7887 7296 7932 7324
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8018 7284 8024 7336
rect 8076 7324 8082 7336
rect 8941 7327 8999 7333
rect 8941 7324 8953 7327
rect 8076 7296 8953 7324
rect 8076 7284 8082 7296
rect 8941 7293 8953 7296
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 14274 7324 14280 7336
rect 13127 7296 14280 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 15194 7324 15200 7336
rect 15155 7296 15200 7324
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 15672 7324 15700 7355
rect 16022 7324 16028 7336
rect 15672 7296 16028 7324
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 16132 7324 16160 7432
rect 18690 7420 18696 7432
rect 18748 7420 18754 7472
rect 19242 7420 19248 7472
rect 19300 7460 19306 7472
rect 19794 7460 19800 7472
rect 19300 7432 19800 7460
rect 19300 7420 19306 7432
rect 19794 7420 19800 7432
rect 19852 7420 19858 7472
rect 20809 7463 20867 7469
rect 19996 7432 20760 7460
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 17727 7364 19717 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 19705 7361 19717 7364
rect 19751 7392 19763 7395
rect 19886 7392 19892 7404
rect 19751 7364 19892 7392
rect 19751 7361 19763 7364
rect 19705 7355 19763 7361
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 19150 7324 19156 7336
rect 16132 7296 19156 7324
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 19996 7324 20024 7432
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20487 7364 20545 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 19300 7296 20024 7324
rect 20073 7327 20131 7333
rect 19300 7284 19306 7296
rect 20073 7293 20085 7327
rect 20119 7324 20131 7327
rect 20622 7324 20628 7336
rect 20119 7296 20628 7324
rect 20119 7293 20131 7296
rect 20073 7287 20131 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 20732 7324 20760 7432
rect 20809 7429 20821 7463
rect 20855 7460 20867 7463
rect 20990 7460 20996 7472
rect 20855 7432 20996 7460
rect 20855 7429 20867 7432
rect 20809 7423 20867 7429
rect 20990 7420 20996 7432
rect 21048 7420 21054 7472
rect 21358 7420 21364 7472
rect 21416 7460 21422 7472
rect 34146 7460 34152 7472
rect 21416 7432 29592 7460
rect 34107 7432 34152 7460
rect 21416 7420 21422 7432
rect 21545 7395 21603 7401
rect 21545 7361 21557 7395
rect 21591 7392 21603 7395
rect 21910 7392 21916 7404
rect 21591 7364 21916 7392
rect 21591 7361 21603 7364
rect 21545 7355 21603 7361
rect 21910 7352 21916 7364
rect 21968 7352 21974 7404
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7392 22063 7395
rect 22373 7395 22431 7401
rect 22373 7392 22385 7395
rect 22051 7364 22385 7392
rect 22051 7361 22063 7364
rect 22005 7355 22063 7361
rect 22373 7361 22385 7364
rect 22419 7392 22431 7395
rect 25038 7392 25044 7404
rect 22419 7364 24808 7392
rect 24999 7364 25044 7392
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 23566 7324 23572 7336
rect 20732 7296 23572 7324
rect 23566 7284 23572 7296
rect 23624 7284 23630 7336
rect 23658 7284 23664 7336
rect 23716 7324 23722 7336
rect 24670 7324 24676 7336
rect 23716 7296 23761 7324
rect 24631 7296 24676 7324
rect 23716 7284 23722 7296
rect 24670 7284 24676 7296
rect 24728 7284 24734 7336
rect 24780 7324 24808 7364
rect 25038 7352 25044 7364
rect 25096 7352 25102 7404
rect 28902 7392 28908 7404
rect 25148 7364 28908 7392
rect 25148 7324 25176 7364
rect 28902 7352 28908 7364
rect 28960 7352 28966 7404
rect 29564 7392 29592 7432
rect 34146 7420 34152 7432
rect 34204 7420 34210 7472
rect 34238 7420 34244 7472
rect 34296 7460 34302 7472
rect 37369 7463 37427 7469
rect 37369 7460 37381 7463
rect 34296 7432 37381 7460
rect 34296 7420 34302 7432
rect 37369 7429 37381 7432
rect 37415 7429 37427 7463
rect 37369 7423 37427 7429
rect 37476 7432 39620 7460
rect 35894 7392 35900 7404
rect 29564 7364 35900 7392
rect 35894 7352 35900 7364
rect 35952 7352 35958 7404
rect 36262 7392 36268 7404
rect 36223 7364 36268 7392
rect 36262 7352 36268 7364
rect 36320 7352 36326 7404
rect 36633 7395 36691 7401
rect 36633 7361 36645 7395
rect 36679 7361 36691 7395
rect 36633 7355 36691 7361
rect 26418 7324 26424 7336
rect 24780 7296 25176 7324
rect 25240 7296 26424 7324
rect 8202 7216 8208 7268
rect 8260 7256 8266 7268
rect 9677 7259 9735 7265
rect 9677 7256 9689 7259
rect 8260 7228 9689 7256
rect 8260 7216 8266 7228
rect 9677 7225 9689 7228
rect 9723 7225 9735 7259
rect 9677 7219 9735 7225
rect 18690 7216 18696 7268
rect 18748 7256 18754 7268
rect 18966 7256 18972 7268
rect 18748 7228 18972 7256
rect 18748 7216 18754 7228
rect 18966 7216 18972 7228
rect 19024 7216 19030 7268
rect 20806 7256 20812 7268
rect 20456 7228 20812 7256
rect 9582 7148 9588 7200
rect 9640 7188 9646 7200
rect 9769 7191 9827 7197
rect 9769 7188 9781 7191
rect 9640 7160 9781 7188
rect 9640 7148 9646 7160
rect 9769 7157 9781 7160
rect 9815 7157 9827 7191
rect 9769 7151 9827 7157
rect 13906 7148 13912 7200
rect 13964 7188 13970 7200
rect 20456 7188 20484 7228
rect 20806 7216 20812 7228
rect 20864 7216 20870 7268
rect 21177 7259 21235 7265
rect 21177 7225 21189 7259
rect 21223 7256 21235 7259
rect 21726 7256 21732 7268
rect 21223 7228 21732 7256
rect 21223 7225 21235 7228
rect 21177 7219 21235 7225
rect 21726 7216 21732 7228
rect 21784 7256 21790 7268
rect 25240 7256 25268 7296
rect 26418 7284 26424 7296
rect 26476 7284 26482 7336
rect 26510 7284 26516 7336
rect 26568 7324 26574 7336
rect 26568 7296 26613 7324
rect 26568 7284 26574 7296
rect 26694 7284 26700 7336
rect 26752 7324 26758 7336
rect 27614 7324 27620 7336
rect 26752 7296 27620 7324
rect 26752 7284 26758 7296
rect 27614 7284 27620 7296
rect 27672 7284 27678 7336
rect 34422 7284 34428 7336
rect 34480 7324 34486 7336
rect 34790 7324 34796 7336
rect 34480 7296 34796 7324
rect 34480 7284 34486 7296
rect 34790 7284 34796 7296
rect 34848 7284 34854 7336
rect 35250 7284 35256 7336
rect 35308 7324 35314 7336
rect 35308 7296 36492 7324
rect 35308 7284 35314 7296
rect 21784 7228 25268 7256
rect 21784 7216 21790 7228
rect 32490 7216 32496 7268
rect 32548 7256 32554 7268
rect 36081 7259 36139 7265
rect 36081 7256 36093 7259
rect 32548 7228 36093 7256
rect 32548 7216 32554 7228
rect 36081 7225 36093 7228
rect 36127 7225 36139 7259
rect 36081 7219 36139 7225
rect 13964 7160 20484 7188
rect 20533 7191 20591 7197
rect 13964 7148 13970 7160
rect 20533 7157 20545 7191
rect 20579 7188 20591 7191
rect 21266 7188 21272 7200
rect 20579 7160 21272 7188
rect 20579 7157 20591 7160
rect 20533 7151 20591 7157
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 21361 7191 21419 7197
rect 21361 7157 21373 7191
rect 21407 7188 21419 7191
rect 21542 7188 21548 7200
rect 21407 7160 21548 7188
rect 21407 7157 21419 7160
rect 21361 7151 21419 7157
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 23106 7188 23112 7200
rect 23067 7160 23112 7188
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 23198 7148 23204 7200
rect 23256 7188 23262 7200
rect 28810 7188 28816 7200
rect 23256 7160 28816 7188
rect 23256 7148 23262 7160
rect 28810 7148 28816 7160
rect 28868 7148 28874 7200
rect 28902 7148 28908 7200
rect 28960 7188 28966 7200
rect 33686 7188 33692 7200
rect 28960 7160 33692 7188
rect 28960 7148 28966 7160
rect 33686 7148 33692 7160
rect 33744 7148 33750 7200
rect 33962 7188 33968 7200
rect 33923 7160 33968 7188
rect 33962 7148 33968 7160
rect 34020 7148 34026 7200
rect 34606 7148 34612 7200
rect 34664 7188 34670 7200
rect 36354 7188 36360 7200
rect 34664 7160 36360 7188
rect 34664 7148 34670 7160
rect 36354 7148 36360 7160
rect 36412 7148 36418 7200
rect 36464 7188 36492 7296
rect 36648 7256 36676 7355
rect 37182 7352 37188 7404
rect 37240 7392 37246 7404
rect 37476 7392 37504 7432
rect 37240 7364 37504 7392
rect 37829 7395 37887 7401
rect 37240 7352 37246 7364
rect 37829 7361 37841 7395
rect 37875 7361 37887 7395
rect 37829 7355 37887 7361
rect 38289 7395 38347 7401
rect 38289 7361 38301 7395
rect 38335 7392 38347 7395
rect 38470 7392 38476 7404
rect 38335 7364 38476 7392
rect 38335 7361 38347 7364
rect 38289 7355 38347 7361
rect 37274 7284 37280 7336
rect 37332 7324 37338 7336
rect 37332 7296 37377 7324
rect 37332 7284 37338 7296
rect 37458 7284 37464 7336
rect 37516 7324 37522 7336
rect 37844 7324 37872 7355
rect 38470 7352 38476 7364
rect 38528 7392 38534 7404
rect 39482 7392 39488 7404
rect 38528 7364 39488 7392
rect 38528 7352 38534 7364
rect 39482 7352 39488 7364
rect 39540 7352 39546 7404
rect 39592 7392 39620 7432
rect 39666 7420 39672 7472
rect 39724 7460 39730 7472
rect 42352 7460 42380 7500
rect 39724 7432 42380 7460
rect 42429 7463 42487 7469
rect 39724 7420 39730 7432
rect 42429 7429 42441 7463
rect 42475 7429 42487 7463
rect 42536 7460 42564 7500
rect 42610 7488 42616 7540
rect 42668 7528 42674 7540
rect 45554 7528 45560 7540
rect 42668 7500 45560 7528
rect 42668 7488 42674 7500
rect 45554 7488 45560 7500
rect 45612 7488 45618 7540
rect 45738 7488 45744 7540
rect 45796 7528 45802 7540
rect 45833 7531 45891 7537
rect 45833 7528 45845 7531
rect 45796 7500 45845 7528
rect 45796 7488 45802 7500
rect 45833 7497 45845 7500
rect 45879 7497 45891 7531
rect 71682 7528 71688 7540
rect 45833 7491 45891 7497
rect 45940 7500 71688 7528
rect 45940 7460 45968 7500
rect 71682 7488 71688 7500
rect 71740 7488 71746 7540
rect 83366 7528 83372 7540
rect 83327 7500 83372 7528
rect 83366 7488 83372 7500
rect 83424 7488 83430 7540
rect 93044 7528 93072 7704
rect 97166 7692 97172 7744
rect 97224 7732 97230 7744
rect 101861 7735 101919 7741
rect 101861 7732 101873 7735
rect 97224 7704 101873 7732
rect 97224 7692 97230 7704
rect 101861 7701 101873 7704
rect 101907 7701 101919 7735
rect 102318 7732 102324 7744
rect 102279 7704 102324 7732
rect 101861 7695 101919 7701
rect 102318 7692 102324 7704
rect 102376 7692 102382 7744
rect 102965 7735 103023 7741
rect 102965 7701 102977 7735
rect 103011 7732 103023 7735
rect 104342 7732 104348 7744
rect 103011 7704 104348 7732
rect 103011 7701 103023 7704
rect 102965 7695 103023 7701
rect 104342 7692 104348 7704
rect 104400 7692 104406 7744
rect 104437 7735 104495 7741
rect 104437 7701 104449 7735
rect 104483 7732 104495 7735
rect 104618 7732 104624 7744
rect 104483 7704 104624 7732
rect 104483 7701 104495 7704
rect 104437 7695 104495 7701
rect 104618 7692 104624 7704
rect 104676 7732 104682 7744
rect 113468 7732 113496 7772
rect 116210 7760 116216 7772
rect 116268 7760 116274 7812
rect 116320 7800 116348 7831
rect 116578 7800 116584 7812
rect 116320 7772 116584 7800
rect 116578 7760 116584 7772
rect 116636 7760 116642 7812
rect 118160 7800 118188 7831
rect 133414 7828 133420 7840
rect 133472 7828 133478 7880
rect 134242 7868 134248 7880
rect 134203 7840 134248 7868
rect 134242 7828 134248 7840
rect 134300 7868 134306 7880
rect 134889 7871 134947 7877
rect 134889 7868 134901 7871
rect 134300 7840 134901 7868
rect 134300 7828 134306 7840
rect 134889 7837 134901 7840
rect 134935 7837 134947 7871
rect 134889 7831 134947 7837
rect 143353 7871 143411 7877
rect 143353 7837 143365 7871
rect 143399 7837 143411 7871
rect 146386 7868 146392 7880
rect 146347 7840 146392 7868
rect 143353 7831 143411 7837
rect 120810 7800 120816 7812
rect 118160 7772 120816 7800
rect 120810 7760 120816 7772
rect 120868 7760 120874 7812
rect 121273 7803 121331 7809
rect 121273 7769 121285 7803
rect 121319 7800 121331 7803
rect 121362 7800 121368 7812
rect 121319 7772 121368 7800
rect 121319 7769 121331 7772
rect 121273 7763 121331 7769
rect 121362 7760 121368 7772
rect 121420 7800 121426 7812
rect 122466 7800 122472 7812
rect 121420 7772 122472 7800
rect 121420 7760 121426 7772
rect 122466 7760 122472 7772
rect 122524 7760 122530 7812
rect 104676 7704 113496 7732
rect 113913 7735 113971 7741
rect 104676 7692 104682 7704
rect 113913 7701 113925 7735
rect 113959 7732 113971 7735
rect 114189 7735 114247 7741
rect 114189 7732 114201 7735
rect 113959 7704 114201 7732
rect 113959 7701 113971 7704
rect 113913 7695 113971 7701
rect 114189 7701 114201 7704
rect 114235 7732 114247 7735
rect 118786 7732 118792 7744
rect 114235 7704 118792 7732
rect 114235 7701 114247 7704
rect 114189 7695 114247 7701
rect 118786 7692 118792 7704
rect 118844 7692 118850 7744
rect 118970 7732 118976 7744
rect 118931 7704 118976 7732
rect 118970 7692 118976 7704
rect 119028 7692 119034 7744
rect 121454 7692 121460 7744
rect 121512 7732 121518 7744
rect 121825 7735 121883 7741
rect 121825 7732 121837 7735
rect 121512 7704 121837 7732
rect 121512 7692 121518 7704
rect 121825 7701 121837 7704
rect 121871 7701 121883 7735
rect 127066 7732 127072 7744
rect 126979 7704 127072 7732
rect 121825 7695 121883 7701
rect 127066 7692 127072 7704
rect 127124 7732 127130 7744
rect 127986 7732 127992 7744
rect 127124 7704 127992 7732
rect 127124 7692 127130 7704
rect 127986 7692 127992 7704
rect 128044 7692 128050 7744
rect 131022 7692 131028 7744
rect 131080 7732 131086 7744
rect 131209 7735 131267 7741
rect 131209 7732 131221 7735
rect 131080 7704 131221 7732
rect 131080 7692 131086 7704
rect 131209 7701 131221 7704
rect 131255 7701 131267 7735
rect 143368 7732 143396 7831
rect 146386 7828 146392 7840
rect 146444 7868 146450 7880
rect 146849 7871 146907 7877
rect 146849 7868 146861 7871
rect 146444 7840 146861 7868
rect 146444 7828 146450 7840
rect 146849 7837 146861 7840
rect 146895 7837 146907 7871
rect 146849 7831 146907 7837
rect 148965 7871 149023 7877
rect 148965 7837 148977 7871
rect 149011 7868 149023 7871
rect 149701 7871 149759 7877
rect 149011 7840 149376 7868
rect 149011 7837 149023 7840
rect 148965 7831 149023 7837
rect 143721 7803 143779 7809
rect 143721 7769 143733 7803
rect 143767 7800 143779 7803
rect 143902 7800 143908 7812
rect 143767 7772 143908 7800
rect 143767 7769 143779 7772
rect 143721 7763 143779 7769
rect 143902 7760 143908 7772
rect 143960 7800 143966 7812
rect 145374 7800 145380 7812
rect 143960 7772 145380 7800
rect 143960 7760 143966 7772
rect 145374 7760 145380 7772
rect 145432 7760 145438 7812
rect 144089 7735 144147 7741
rect 144089 7732 144101 7735
rect 143368 7704 144101 7732
rect 131209 7695 131267 7701
rect 144089 7701 144101 7704
rect 144135 7732 144147 7735
rect 146478 7732 146484 7744
rect 144135 7704 146484 7732
rect 144135 7701 144147 7704
rect 144089 7695 144147 7701
rect 146478 7692 146484 7704
rect 146536 7692 146542 7744
rect 149348 7741 149376 7840
rect 149701 7837 149713 7871
rect 149747 7868 149759 7871
rect 149885 7871 149943 7877
rect 149885 7868 149897 7871
rect 149747 7840 149897 7868
rect 149747 7837 149759 7840
rect 149701 7831 149759 7837
rect 149885 7837 149897 7840
rect 149931 7868 149943 7871
rect 150434 7868 150440 7880
rect 149931 7840 150440 7868
rect 149931 7837 149943 7840
rect 149885 7831 149943 7837
rect 150434 7828 150440 7840
rect 150492 7828 150498 7880
rect 150986 7868 150992 7880
rect 150947 7840 150992 7868
rect 150986 7828 150992 7840
rect 151044 7868 151050 7880
rect 151725 7871 151783 7877
rect 151725 7868 151737 7871
rect 151044 7840 151737 7868
rect 151044 7828 151050 7840
rect 151725 7837 151737 7840
rect 151771 7837 151783 7871
rect 151725 7831 151783 7837
rect 153013 7871 153071 7877
rect 153013 7837 153025 7871
rect 153059 7837 153071 7871
rect 153013 7831 153071 7837
rect 154577 7871 154635 7877
rect 154577 7837 154589 7871
rect 154623 7837 154635 7871
rect 154577 7831 154635 7837
rect 155497 7871 155555 7877
rect 155497 7837 155509 7871
rect 155543 7868 155555 7871
rect 156138 7868 156144 7880
rect 155543 7840 156144 7868
rect 155543 7837 155555 7840
rect 155497 7831 155555 7837
rect 149333 7735 149391 7741
rect 149333 7701 149345 7735
rect 149379 7732 149391 7735
rect 149422 7732 149428 7744
rect 149379 7704 149428 7732
rect 149379 7701 149391 7704
rect 149333 7695 149391 7701
rect 149422 7692 149428 7704
rect 149480 7692 149486 7744
rect 152918 7732 152924 7744
rect 152879 7704 152924 7732
rect 152918 7692 152924 7704
rect 152976 7732 152982 7744
rect 153028 7732 153056 7831
rect 152976 7704 153056 7732
rect 154592 7732 154620 7831
rect 156138 7828 156144 7840
rect 156196 7828 156202 7880
rect 156984 7877 157012 7908
rect 156969 7871 157027 7877
rect 156969 7837 156981 7871
rect 157015 7837 157027 7871
rect 156969 7831 157027 7837
rect 157444 7809 157472 7908
rect 159358 7896 159364 7908
rect 159416 7896 159422 7948
rect 161106 7936 161112 7948
rect 161067 7908 161112 7936
rect 161106 7896 161112 7908
rect 161164 7896 161170 7948
rect 162118 7936 162124 7948
rect 162079 7908 162124 7936
rect 162118 7896 162124 7908
rect 162176 7896 162182 7948
rect 166718 7936 166724 7948
rect 166679 7908 166724 7936
rect 166718 7896 166724 7908
rect 166776 7896 166782 7948
rect 158257 7871 158315 7877
rect 158257 7837 158269 7871
rect 158303 7868 158315 7871
rect 158349 7871 158407 7877
rect 158349 7868 158361 7871
rect 158303 7840 158361 7868
rect 158303 7837 158315 7840
rect 158257 7831 158315 7837
rect 158349 7837 158361 7840
rect 158395 7868 158407 7871
rect 158714 7868 158720 7880
rect 158395 7840 158720 7868
rect 158395 7837 158407 7840
rect 158349 7831 158407 7837
rect 158714 7828 158720 7840
rect 158772 7828 158778 7880
rect 159726 7868 159732 7880
rect 159687 7840 159732 7868
rect 159726 7828 159732 7840
rect 159784 7868 159790 7880
rect 160189 7871 160247 7877
rect 160189 7868 160201 7871
rect 159784 7840 160201 7868
rect 159784 7828 159790 7840
rect 160189 7837 160201 7840
rect 160235 7837 160247 7871
rect 160189 7831 160247 7837
rect 161934 7828 161940 7880
rect 161992 7868 161998 7880
rect 162213 7871 162271 7877
rect 162213 7868 162225 7871
rect 161992 7840 162225 7868
rect 161992 7828 161998 7840
rect 162213 7837 162225 7840
rect 162259 7868 162271 7871
rect 162949 7871 163007 7877
rect 162949 7868 162961 7871
rect 162259 7840 162961 7868
rect 162259 7837 162271 7840
rect 162213 7831 162271 7837
rect 162949 7837 162961 7840
rect 162995 7837 163007 7871
rect 162949 7831 163007 7837
rect 163501 7871 163559 7877
rect 163501 7837 163513 7871
rect 163547 7837 163559 7871
rect 164602 7868 164608 7880
rect 164563 7840 164608 7868
rect 163501 7831 163559 7837
rect 157429 7803 157487 7809
rect 157429 7769 157441 7803
rect 157475 7800 157487 7803
rect 157518 7800 157524 7812
rect 157475 7772 157524 7800
rect 157475 7769 157487 7772
rect 157429 7763 157487 7769
rect 157518 7760 157524 7772
rect 157576 7760 157582 7812
rect 154942 7732 154948 7744
rect 154592 7704 154948 7732
rect 152976 7692 152982 7704
rect 154942 7692 154948 7704
rect 155000 7692 155006 7744
rect 160738 7732 160744 7744
rect 160699 7704 160744 7732
rect 160738 7692 160744 7704
rect 160796 7692 160802 7744
rect 163406 7732 163412 7744
rect 163367 7704 163412 7732
rect 163406 7692 163412 7704
rect 163464 7732 163470 7744
rect 163516 7732 163544 7831
rect 164602 7828 164608 7840
rect 164660 7868 164666 7880
rect 165341 7871 165399 7877
rect 165341 7868 165353 7871
rect 164660 7840 165353 7868
rect 164660 7828 164666 7840
rect 165341 7837 165353 7840
rect 165387 7837 165399 7871
rect 165341 7831 165399 7837
rect 163464 7704 163544 7732
rect 163464 7692 163470 7704
rect 165614 7692 165620 7744
rect 165672 7732 165678 7744
rect 165801 7735 165859 7741
rect 165801 7732 165813 7735
rect 165672 7704 165813 7732
rect 165672 7692 165678 7704
rect 165801 7701 165813 7704
rect 165847 7701 165859 7735
rect 165801 7695 165859 7701
rect 96430 7624 96436 7676
rect 96488 7664 96494 7676
rect 101401 7667 101459 7673
rect 101401 7664 101413 7667
rect 96488 7636 101413 7664
rect 96488 7624 96494 7636
rect 101401 7633 101413 7636
rect 101447 7633 101459 7667
rect 101401 7627 101459 7633
rect 102028 7642 169556 7664
rect 99745 7599 99803 7605
rect 99745 7565 99757 7599
rect 99791 7596 99803 7599
rect 99791 7568 100524 7596
rect 102028 7590 113088 7642
rect 113140 7590 113152 7642
rect 113204 7590 113216 7642
rect 113268 7590 113280 7642
rect 113332 7590 169556 7642
rect 102028 7568 169556 7590
rect 99791 7565 99803 7568
rect 99745 7559 99803 7565
rect 100386 7528 100392 7540
rect 93044 7500 100392 7528
rect 100386 7488 100392 7500
rect 100444 7488 100450 7540
rect 100496 7528 100524 7568
rect 108482 7528 108488 7540
rect 100496 7500 108488 7528
rect 108482 7488 108488 7500
rect 108540 7488 108546 7540
rect 108574 7488 108580 7540
rect 108632 7528 108638 7540
rect 142430 7528 142436 7540
rect 108632 7500 116808 7528
rect 142391 7500 142436 7528
rect 108632 7488 108638 7500
rect 47854 7460 47860 7472
rect 42536 7432 45968 7460
rect 46032 7432 47860 7460
rect 42429 7423 42487 7429
rect 40586 7392 40592 7404
rect 39592 7364 40592 7392
rect 40586 7352 40592 7364
rect 40644 7352 40650 7404
rect 41325 7395 41383 7401
rect 41325 7361 41337 7395
rect 41371 7361 41383 7395
rect 41325 7355 41383 7361
rect 38565 7327 38623 7333
rect 38565 7324 38577 7327
rect 37516 7296 38577 7324
rect 37516 7284 37522 7296
rect 38565 7293 38577 7296
rect 38611 7293 38623 7327
rect 38565 7287 38623 7293
rect 38654 7284 38660 7336
rect 38712 7324 38718 7336
rect 39298 7324 39304 7336
rect 38712 7296 39304 7324
rect 38712 7284 38718 7296
rect 39298 7284 39304 7296
rect 39356 7284 39362 7336
rect 39390 7284 39396 7336
rect 39448 7324 39454 7336
rect 39761 7327 39819 7333
rect 39761 7324 39773 7327
rect 39448 7296 39773 7324
rect 39448 7284 39454 7296
rect 39761 7293 39773 7296
rect 39807 7293 39819 7327
rect 40678 7324 40684 7336
rect 39761 7287 39819 7293
rect 39868 7296 40684 7324
rect 36998 7256 37004 7268
rect 36648 7228 37004 7256
rect 36998 7216 37004 7228
rect 37056 7256 37062 7268
rect 39868 7256 39896 7296
rect 40678 7284 40684 7296
rect 40736 7284 40742 7336
rect 40773 7327 40831 7333
rect 40773 7293 40785 7327
rect 40819 7293 40831 7327
rect 41340 7324 41368 7355
rect 41782 7352 41788 7404
rect 41840 7392 41846 7404
rect 42242 7392 42248 7404
rect 41840 7364 42248 7392
rect 41840 7352 41846 7364
rect 42242 7352 42248 7364
rect 42300 7352 42306 7404
rect 41414 7324 41420 7336
rect 41340 7296 41420 7324
rect 40773 7287 40831 7293
rect 37056 7228 39896 7256
rect 37056 7216 37062 7228
rect 39942 7216 39948 7268
rect 40000 7256 40006 7268
rect 40788 7256 40816 7287
rect 41414 7284 41420 7296
rect 41472 7284 41478 7336
rect 41598 7324 41604 7336
rect 41559 7296 41604 7324
rect 41598 7284 41604 7296
rect 41656 7284 41662 7336
rect 41690 7284 41696 7336
rect 41748 7324 41754 7336
rect 42150 7324 42156 7336
rect 41748 7296 42156 7324
rect 41748 7284 41754 7296
rect 42150 7284 42156 7296
rect 42208 7284 42214 7336
rect 42444 7324 42472 7423
rect 42705 7395 42763 7401
rect 42705 7361 42717 7395
rect 42751 7392 42763 7395
rect 42751 7364 44404 7392
rect 42751 7361 42763 7364
rect 42705 7355 42763 7361
rect 42610 7324 42616 7336
rect 42444 7296 42616 7324
rect 42610 7284 42616 7296
rect 42668 7324 42674 7336
rect 42889 7327 42947 7333
rect 42889 7324 42901 7327
rect 42668 7296 42901 7324
rect 42668 7284 42674 7296
rect 42889 7293 42901 7296
rect 42935 7293 42947 7327
rect 44266 7324 44272 7336
rect 44227 7296 44272 7324
rect 42889 7287 42947 7293
rect 44266 7284 44272 7296
rect 44324 7284 44330 7336
rect 44376 7324 44404 7364
rect 44542 7352 44548 7404
rect 44600 7392 44606 7404
rect 46032 7392 46060 7432
rect 47854 7420 47860 7432
rect 47912 7420 47918 7472
rect 48498 7460 48504 7472
rect 47964 7432 48504 7460
rect 44600 7364 46060 7392
rect 44600 7352 44606 7364
rect 46750 7352 46756 7404
rect 46808 7392 46814 7404
rect 46845 7395 46903 7401
rect 46845 7392 46857 7395
rect 46808 7364 46857 7392
rect 46808 7352 46814 7364
rect 46845 7361 46857 7364
rect 46891 7361 46903 7395
rect 46845 7355 46903 7361
rect 46934 7352 46940 7404
rect 46992 7392 46998 7404
rect 47762 7392 47768 7404
rect 46992 7364 47768 7392
rect 46992 7352 46998 7364
rect 47762 7352 47768 7364
rect 47820 7352 47826 7404
rect 47964 7401 47992 7432
rect 48498 7420 48504 7432
rect 48556 7420 48562 7472
rect 48777 7463 48835 7469
rect 48777 7429 48789 7463
rect 48823 7460 48835 7463
rect 48866 7460 48872 7472
rect 48823 7432 48872 7460
rect 48823 7429 48835 7432
rect 48777 7423 48835 7429
rect 48866 7420 48872 7432
rect 48924 7460 48930 7472
rect 49237 7463 49295 7469
rect 49237 7460 49249 7463
rect 48924 7432 49249 7460
rect 48924 7420 48930 7432
rect 49237 7429 49249 7432
rect 49283 7429 49295 7463
rect 49237 7423 49295 7429
rect 49786 7420 49792 7472
rect 49844 7460 49850 7472
rect 50798 7460 50804 7472
rect 49844 7432 50804 7460
rect 49844 7420 49850 7432
rect 50798 7420 50804 7432
rect 50856 7420 50862 7472
rect 50985 7463 51043 7469
rect 50985 7429 50997 7463
rect 51031 7460 51043 7463
rect 51442 7460 51448 7472
rect 51031 7432 51448 7460
rect 51031 7429 51043 7432
rect 50985 7423 51043 7429
rect 51442 7420 51448 7432
rect 51500 7420 51506 7472
rect 51537 7463 51595 7469
rect 51537 7429 51549 7463
rect 51583 7460 51595 7463
rect 51626 7460 51632 7472
rect 51583 7432 51632 7460
rect 51583 7429 51595 7432
rect 51537 7423 51595 7429
rect 51626 7420 51632 7432
rect 51684 7420 51690 7472
rect 51994 7420 52000 7472
rect 52052 7460 52058 7472
rect 52730 7460 52736 7472
rect 52052 7432 52736 7460
rect 52052 7420 52058 7432
rect 52730 7420 52736 7432
rect 52788 7420 52794 7472
rect 52825 7463 52883 7469
rect 52825 7429 52837 7463
rect 52871 7460 52883 7463
rect 53558 7460 53564 7472
rect 52871 7432 53564 7460
rect 52871 7429 52883 7432
rect 52825 7423 52883 7429
rect 53558 7420 53564 7432
rect 53616 7420 53622 7472
rect 53837 7463 53895 7469
rect 53837 7429 53849 7463
rect 53883 7460 53895 7463
rect 54386 7460 54392 7472
rect 53883 7432 54392 7460
rect 53883 7429 53895 7432
rect 53837 7423 53895 7429
rect 54386 7420 54392 7432
rect 54444 7420 54450 7472
rect 54846 7460 54852 7472
rect 54807 7432 54852 7460
rect 54846 7420 54852 7432
rect 54904 7420 54910 7472
rect 60921 7463 60979 7469
rect 55324 7432 59952 7460
rect 47949 7395 48007 7401
rect 47949 7361 47961 7395
rect 47995 7361 48007 7395
rect 55324 7392 55352 7432
rect 47949 7355 48007 7361
rect 48056 7364 55352 7392
rect 48056 7324 48084 7364
rect 55582 7352 55588 7404
rect 55640 7392 55646 7404
rect 55640 7364 55904 7392
rect 55640 7352 55646 7364
rect 44376 7296 48084 7324
rect 48130 7284 48136 7336
rect 48188 7324 48194 7336
rect 48188 7296 48233 7324
rect 48188 7284 48194 7296
rect 48866 7284 48872 7336
rect 48924 7324 48930 7336
rect 54846 7324 54852 7336
rect 48924 7296 54852 7324
rect 48924 7284 48930 7296
rect 54846 7284 54852 7296
rect 54904 7284 54910 7336
rect 55876 7324 55904 7364
rect 56134 7352 56140 7404
rect 56192 7392 56198 7404
rect 56597 7395 56655 7401
rect 56597 7392 56609 7395
rect 56192 7364 56609 7392
rect 56192 7352 56198 7364
rect 56597 7361 56609 7364
rect 56643 7361 56655 7395
rect 56597 7355 56655 7361
rect 56778 7352 56784 7404
rect 56836 7352 56842 7404
rect 56962 7352 56968 7404
rect 57020 7352 57026 7404
rect 57333 7395 57391 7401
rect 57333 7361 57345 7395
rect 57379 7392 57391 7395
rect 57422 7392 57428 7404
rect 57379 7364 57428 7392
rect 57379 7361 57391 7364
rect 57333 7355 57391 7361
rect 57422 7352 57428 7364
rect 57480 7352 57486 7404
rect 59814 7392 59820 7404
rect 59775 7364 59820 7392
rect 59814 7352 59820 7364
rect 59872 7352 59878 7404
rect 59924 7392 59952 7432
rect 60921 7429 60933 7463
rect 60967 7460 60979 7463
rect 61010 7460 61016 7472
rect 60967 7432 61016 7460
rect 60967 7429 60979 7432
rect 60921 7423 60979 7429
rect 61010 7420 61016 7432
rect 61068 7420 61074 7472
rect 90450 7460 90456 7472
rect 90411 7432 90456 7460
rect 90450 7420 90456 7432
rect 90508 7420 90514 7472
rect 91278 7460 91284 7472
rect 91239 7432 91284 7460
rect 91278 7420 91284 7432
rect 91336 7420 91342 7472
rect 91741 7463 91799 7469
rect 91741 7429 91753 7463
rect 91787 7460 91799 7463
rect 94314 7460 94320 7472
rect 91787 7432 94320 7460
rect 91787 7429 91799 7432
rect 91741 7423 91799 7429
rect 94314 7420 94320 7432
rect 94372 7420 94378 7472
rect 98638 7420 98644 7472
rect 98696 7460 98702 7472
rect 98696 7432 116072 7460
rect 98696 7420 98702 7432
rect 63862 7392 63868 7404
rect 59924 7364 63868 7392
rect 63862 7352 63868 7364
rect 63920 7352 63926 7404
rect 68830 7392 68836 7404
rect 68791 7364 68836 7392
rect 68830 7352 68836 7364
rect 68888 7352 68894 7404
rect 70118 7392 70124 7404
rect 70079 7364 70124 7392
rect 70118 7352 70124 7364
rect 70176 7352 70182 7404
rect 81342 7392 81348 7404
rect 81303 7364 81348 7392
rect 81342 7352 81348 7364
rect 81400 7352 81406 7404
rect 89349 7395 89407 7401
rect 89349 7361 89361 7395
rect 89395 7361 89407 7395
rect 89349 7355 89407 7361
rect 56796 7324 56824 7352
rect 55876 7296 56824 7324
rect 56980 7324 57008 7352
rect 57974 7324 57980 7336
rect 56980 7296 57980 7324
rect 57974 7284 57980 7296
rect 58032 7284 58038 7336
rect 58437 7327 58495 7333
rect 58437 7293 58449 7327
rect 58483 7324 58495 7327
rect 59078 7324 59084 7336
rect 58483 7296 59084 7324
rect 58483 7293 58495 7296
rect 58437 7287 58495 7293
rect 59078 7284 59084 7296
rect 59136 7284 59142 7336
rect 59449 7327 59507 7333
rect 59449 7293 59461 7327
rect 59495 7293 59507 7327
rect 69842 7324 69848 7336
rect 69803 7296 69848 7324
rect 59449 7287 59507 7293
rect 40000 7228 40816 7256
rect 40000 7216 40006 7228
rect 40862 7216 40868 7268
rect 40920 7256 40926 7268
rect 42426 7256 42432 7268
rect 40920 7228 42432 7256
rect 40920 7216 40926 7228
rect 42426 7216 42432 7228
rect 42484 7216 42490 7268
rect 42794 7216 42800 7268
rect 42852 7256 42858 7268
rect 42852 7228 45048 7256
rect 42852 7216 42858 7228
rect 37182 7188 37188 7200
rect 36464 7160 37188 7188
rect 37182 7148 37188 7160
rect 37240 7148 37246 7200
rect 37369 7191 37427 7197
rect 37369 7157 37381 7191
rect 37415 7188 37427 7191
rect 37645 7191 37703 7197
rect 37645 7188 37657 7191
rect 37415 7160 37657 7188
rect 37415 7157 37427 7160
rect 37369 7151 37427 7157
rect 37645 7157 37657 7160
rect 37691 7157 37703 7191
rect 37645 7151 37703 7157
rect 38562 7148 38568 7200
rect 38620 7188 38626 7200
rect 42705 7191 42763 7197
rect 42705 7188 42717 7191
rect 38620 7160 42717 7188
rect 38620 7148 38626 7160
rect 42705 7157 42717 7160
rect 42751 7157 42763 7191
rect 42705 7151 42763 7157
rect 43530 7148 43536 7200
rect 43588 7188 43594 7200
rect 44174 7188 44180 7200
rect 43588 7160 44180 7188
rect 43588 7148 43594 7160
rect 44174 7148 44180 7160
rect 44232 7148 44238 7200
rect 44266 7148 44272 7200
rect 44324 7188 44330 7200
rect 44910 7188 44916 7200
rect 44324 7160 44916 7188
rect 44324 7148 44330 7160
rect 44910 7148 44916 7160
rect 44968 7148 44974 7200
rect 45020 7188 45048 7228
rect 45094 7216 45100 7268
rect 45152 7256 45158 7268
rect 45152 7228 55996 7256
rect 45152 7216 45158 7228
rect 46934 7188 46940 7200
rect 45020 7160 46940 7188
rect 46934 7148 46940 7160
rect 46992 7148 46998 7200
rect 47026 7148 47032 7200
rect 47084 7188 47090 7200
rect 51902 7188 51908 7200
rect 47084 7160 51908 7188
rect 47084 7148 47090 7160
rect 51902 7148 51908 7160
rect 51960 7148 51966 7200
rect 52086 7188 52092 7200
rect 51999 7160 52092 7188
rect 52086 7148 52092 7160
rect 52144 7188 52150 7200
rect 55490 7188 55496 7200
rect 52144 7160 55496 7188
rect 52144 7148 52150 7160
rect 55490 7148 55496 7160
rect 55548 7148 55554 7200
rect 55968 7188 55996 7228
rect 56042 7216 56048 7268
rect 56100 7256 56106 7268
rect 56689 7259 56747 7265
rect 56689 7256 56701 7259
rect 56100 7228 56701 7256
rect 56100 7216 56106 7228
rect 56689 7225 56701 7228
rect 56735 7225 56747 7259
rect 56689 7219 56747 7225
rect 56962 7216 56968 7268
rect 57020 7256 57026 7268
rect 59464 7256 59492 7287
rect 69842 7284 69848 7296
rect 69900 7284 69906 7336
rect 79778 7324 79784 7336
rect 79739 7296 79784 7324
rect 79778 7284 79784 7296
rect 79836 7284 79842 7336
rect 80790 7324 80796 7336
rect 80751 7296 80796 7324
rect 80790 7284 80796 7296
rect 80848 7284 80854 7336
rect 86773 7327 86831 7333
rect 86773 7293 86785 7327
rect 86819 7324 86831 7327
rect 87598 7324 87604 7336
rect 86819 7296 87604 7324
rect 86819 7293 86831 7296
rect 86773 7287 86831 7293
rect 87598 7284 87604 7296
rect 87656 7284 87662 7336
rect 87782 7324 87788 7336
rect 87743 7296 87788 7324
rect 87782 7284 87788 7296
rect 87840 7284 87846 7336
rect 89070 7324 89076 7336
rect 89031 7296 89076 7324
rect 89070 7284 89076 7296
rect 89128 7284 89134 7336
rect 89364 7324 89392 7355
rect 102318 7352 102324 7404
rect 102376 7392 102382 7404
rect 102597 7395 102655 7401
rect 102597 7392 102609 7395
rect 102376 7364 102609 7392
rect 102376 7352 102382 7364
rect 102597 7361 102609 7364
rect 102643 7361 102655 7395
rect 103974 7392 103980 7404
rect 103935 7364 103980 7392
rect 102597 7355 102655 7361
rect 103974 7352 103980 7364
rect 104032 7352 104038 7404
rect 109310 7352 109316 7404
rect 109368 7392 109374 7404
rect 114094 7392 114100 7404
rect 109368 7364 114100 7392
rect 109368 7352 109374 7364
rect 114094 7352 114100 7364
rect 114152 7352 114158 7404
rect 114925 7395 114983 7401
rect 114925 7361 114937 7395
rect 114971 7392 114983 7395
rect 115293 7395 115351 7401
rect 115293 7392 115305 7395
rect 114971 7364 115305 7392
rect 114971 7361 114983 7364
rect 114925 7355 114983 7361
rect 115293 7361 115305 7364
rect 115339 7392 115351 7395
rect 115934 7392 115940 7404
rect 115339 7364 115940 7392
rect 115339 7361 115351 7364
rect 115293 7355 115351 7361
rect 115934 7352 115940 7364
rect 115992 7352 115998 7404
rect 89717 7327 89775 7333
rect 89717 7324 89729 7327
rect 89364 7296 89729 7324
rect 89717 7293 89729 7296
rect 89763 7324 89775 7327
rect 96522 7324 96528 7336
rect 89763 7296 96528 7324
rect 89763 7293 89775 7296
rect 89717 7287 89775 7293
rect 96522 7284 96528 7296
rect 96580 7284 96586 7336
rect 96890 7284 96896 7336
rect 96948 7324 96954 7336
rect 96948 7296 104112 7324
rect 96948 7284 96954 7296
rect 57020 7228 59492 7256
rect 101401 7259 101459 7265
rect 57020 7216 57026 7228
rect 101401 7225 101413 7259
rect 101447 7256 101459 7259
rect 103885 7259 103943 7265
rect 103885 7256 103897 7259
rect 101447 7228 103897 7256
rect 101447 7225 101459 7228
rect 101401 7219 101459 7225
rect 103885 7225 103897 7228
rect 103931 7225 103943 7259
rect 104084 7256 104112 7296
rect 104526 7284 104532 7336
rect 104584 7324 104590 7336
rect 113266 7324 113272 7336
rect 104584 7296 113272 7324
rect 104584 7284 104590 7296
rect 113266 7284 113272 7296
rect 113324 7284 113330 7336
rect 113361 7327 113419 7333
rect 113361 7293 113373 7327
rect 113407 7324 113419 7327
rect 113450 7324 113456 7336
rect 113407 7296 113456 7324
rect 113407 7293 113419 7296
rect 113361 7287 113419 7293
rect 113450 7284 113456 7296
rect 113508 7284 113514 7336
rect 114373 7327 114431 7333
rect 114373 7293 114385 7327
rect 114419 7293 114431 7327
rect 115750 7324 115756 7336
rect 115711 7296 115756 7324
rect 114373 7287 114431 7293
rect 114388 7256 114416 7287
rect 115750 7284 115756 7296
rect 115808 7284 115814 7336
rect 116044 7256 116072 7432
rect 116780 7333 116808 7500
rect 142430 7488 142436 7500
rect 142488 7488 142494 7540
rect 145006 7488 145012 7540
rect 145064 7528 145070 7540
rect 145193 7531 145251 7537
rect 145193 7528 145205 7531
rect 145064 7500 145205 7528
rect 145064 7488 145070 7500
rect 145193 7497 145205 7500
rect 145239 7497 145251 7531
rect 147030 7528 147036 7540
rect 146991 7500 147036 7528
rect 145193 7491 145251 7497
rect 147030 7488 147036 7500
rect 147088 7488 147094 7540
rect 147122 7488 147128 7540
rect 147180 7528 147186 7540
rect 147493 7531 147551 7537
rect 147493 7528 147505 7531
rect 147180 7500 147505 7528
rect 147180 7488 147186 7500
rect 147493 7497 147505 7500
rect 147539 7497 147551 7531
rect 147493 7491 147551 7497
rect 149238 7488 149244 7540
rect 149296 7528 149302 7540
rect 149885 7531 149943 7537
rect 149885 7528 149897 7531
rect 149296 7500 149897 7528
rect 149296 7488 149302 7500
rect 149885 7497 149897 7500
rect 149931 7497 149943 7531
rect 150434 7528 150440 7540
rect 150395 7500 150440 7528
rect 149885 7491 149943 7497
rect 116946 7420 116952 7472
rect 117004 7460 117010 7472
rect 149900 7460 149928 7491
rect 150434 7488 150440 7500
rect 150492 7488 150498 7540
rect 156138 7528 156144 7540
rect 156099 7500 156144 7528
rect 156138 7488 156144 7500
rect 156196 7488 156202 7540
rect 158714 7528 158720 7540
rect 158675 7500 158720 7528
rect 158714 7488 158720 7500
rect 158772 7488 158778 7540
rect 159450 7528 159456 7540
rect 159411 7500 159456 7528
rect 159450 7488 159456 7500
rect 159508 7488 159514 7540
rect 163406 7488 163412 7540
rect 163464 7528 163470 7540
rect 166261 7531 166319 7537
rect 166261 7528 166273 7531
rect 163464 7500 166273 7528
rect 163464 7488 163470 7500
rect 166261 7497 166273 7500
rect 166307 7497 166319 7531
rect 166261 7491 166319 7497
rect 151449 7463 151507 7469
rect 151449 7460 151461 7463
rect 117004 7432 126468 7460
rect 149900 7432 151461 7460
rect 117004 7420 117010 7432
rect 117130 7392 117136 7404
rect 117091 7364 117136 7392
rect 117130 7352 117136 7364
rect 117188 7352 117194 7404
rect 118970 7392 118976 7404
rect 118931 7364 118976 7392
rect 118970 7352 118976 7364
rect 119028 7352 119034 7404
rect 120537 7395 120595 7401
rect 120537 7361 120549 7395
rect 120583 7392 120595 7395
rect 120626 7392 120632 7404
rect 120583 7364 120632 7392
rect 120583 7361 120595 7364
rect 120537 7355 120595 7361
rect 120626 7352 120632 7364
rect 120684 7352 120690 7404
rect 122926 7392 122932 7404
rect 122887 7364 122932 7392
rect 122926 7352 122932 7364
rect 122984 7392 122990 7404
rect 123205 7395 123263 7401
rect 123205 7392 123217 7395
rect 122984 7364 123217 7392
rect 122984 7352 122990 7364
rect 123205 7361 123217 7364
rect 123251 7361 123263 7395
rect 123205 7355 123263 7361
rect 116765 7327 116823 7333
rect 116765 7293 116777 7327
rect 116811 7293 116823 7327
rect 116765 7287 116823 7293
rect 119985 7327 120043 7333
rect 119985 7293 119997 7327
rect 120031 7293 120043 7327
rect 121362 7324 121368 7336
rect 121323 7296 121368 7324
rect 119985 7287 120043 7293
rect 120000 7256 120028 7287
rect 121362 7284 121368 7296
rect 121420 7284 121426 7336
rect 122377 7327 122435 7333
rect 122377 7293 122389 7327
rect 122423 7293 122435 7327
rect 125410 7324 125416 7336
rect 125371 7296 125416 7324
rect 122377 7287 122435 7293
rect 104084 7228 114416 7256
rect 114480 7228 115336 7256
rect 116044 7228 120028 7256
rect 103885 7219 103943 7225
rect 56594 7188 56600 7200
rect 55968 7160 56600 7188
rect 56594 7148 56600 7160
rect 56652 7148 56658 7200
rect 57606 7188 57612 7200
rect 57567 7160 57612 7188
rect 57606 7148 57612 7160
rect 57664 7148 57670 7200
rect 58342 7188 58348 7200
rect 58303 7160 58348 7188
rect 58342 7148 58348 7160
rect 58400 7148 58406 7200
rect 60274 7188 60280 7200
rect 60235 7160 60280 7188
rect 60274 7148 60280 7160
rect 60332 7148 60338 7200
rect 81894 7188 81900 7200
rect 81855 7160 81900 7188
rect 81894 7148 81900 7160
rect 81952 7148 81958 7200
rect 104342 7148 104348 7200
rect 104400 7188 104406 7200
rect 114480 7188 114508 7228
rect 104400 7160 114508 7188
rect 115308 7188 115336 7228
rect 122392 7188 122420 7287
rect 125410 7284 125416 7296
rect 125468 7284 125474 7336
rect 126440 7333 126468 7432
rect 151449 7429 151461 7432
rect 151495 7429 151507 7463
rect 151449 7423 151507 7429
rect 152918 7420 152924 7472
rect 152976 7460 152982 7472
rect 156693 7463 156751 7469
rect 156693 7460 156705 7463
rect 152976 7432 156705 7460
rect 152976 7420 152982 7432
rect 156693 7429 156705 7432
rect 156739 7429 156751 7463
rect 156693 7423 156751 7429
rect 126882 7392 126888 7404
rect 126843 7364 126888 7392
rect 126882 7352 126888 7364
rect 126940 7352 126946 7404
rect 133230 7352 133236 7404
rect 133288 7392 133294 7404
rect 133325 7395 133383 7401
rect 133325 7392 133337 7395
rect 133288 7364 133337 7392
rect 133288 7352 133294 7364
rect 133325 7361 133337 7364
rect 133371 7361 133383 7395
rect 144362 7392 144368 7404
rect 144323 7364 144368 7392
rect 133325 7355 133383 7361
rect 144362 7352 144368 7364
rect 144420 7352 144426 7404
rect 149330 7392 149336 7404
rect 149291 7364 149336 7392
rect 149330 7352 149336 7364
rect 149388 7352 149394 7404
rect 155862 7392 155868 7404
rect 155823 7364 155868 7392
rect 155862 7352 155868 7364
rect 155920 7352 155926 7404
rect 160922 7352 160928 7404
rect 160980 7392 160986 7404
rect 161017 7395 161075 7401
rect 161017 7392 161029 7395
rect 160980 7364 161029 7392
rect 160980 7352 160986 7364
rect 161017 7361 161029 7364
rect 161063 7392 161075 7395
rect 161753 7395 161811 7401
rect 161753 7392 161765 7395
rect 161063 7364 161765 7392
rect 161063 7361 161075 7364
rect 161017 7355 161075 7361
rect 161753 7361 161765 7364
rect 161799 7361 161811 7395
rect 164970 7392 164976 7404
rect 164931 7364 164976 7392
rect 161753 7355 161811 7361
rect 164970 7352 164976 7364
rect 165028 7352 165034 7404
rect 126425 7327 126483 7333
rect 126425 7293 126437 7327
rect 126471 7293 126483 7327
rect 126425 7287 126483 7293
rect 127434 7284 127440 7336
rect 127492 7324 127498 7336
rect 127529 7327 127587 7333
rect 127529 7324 127541 7327
rect 127492 7296 127541 7324
rect 127492 7284 127498 7296
rect 127529 7293 127541 7296
rect 127575 7324 127587 7327
rect 127805 7327 127863 7333
rect 127805 7324 127817 7327
rect 127575 7296 127817 7324
rect 127575 7293 127587 7296
rect 127529 7287 127587 7293
rect 127805 7293 127817 7296
rect 127851 7293 127863 7327
rect 127805 7287 127863 7293
rect 129826 7284 129832 7336
rect 129884 7324 129890 7336
rect 129921 7327 129979 7333
rect 129921 7324 129933 7327
rect 129884 7296 129933 7324
rect 129884 7284 129890 7296
rect 129921 7293 129933 7296
rect 129967 7324 129979 7327
rect 130197 7327 130255 7333
rect 130197 7324 130209 7327
rect 129967 7296 130209 7324
rect 129967 7293 129979 7296
rect 129921 7287 129979 7293
rect 130197 7293 130209 7296
rect 130243 7293 130255 7327
rect 132218 7324 132224 7336
rect 132179 7296 132224 7324
rect 130197 7287 130255 7293
rect 132218 7284 132224 7296
rect 132276 7284 132282 7336
rect 133414 7324 133420 7336
rect 133375 7296 133420 7324
rect 133414 7284 133420 7296
rect 133472 7284 133478 7336
rect 142798 7324 142804 7336
rect 142759 7296 142804 7324
rect 142798 7284 142804 7296
rect 142856 7284 142862 7336
rect 143810 7324 143816 7336
rect 143771 7296 143816 7324
rect 143810 7284 143816 7296
rect 143868 7284 143874 7336
rect 148042 7324 148048 7336
rect 148003 7296 148048 7324
rect 148042 7284 148048 7296
rect 148100 7284 148106 7336
rect 149514 7324 149520 7336
rect 149475 7296 149520 7324
rect 149514 7284 149520 7296
rect 149572 7284 149578 7336
rect 153289 7327 153347 7333
rect 153289 7293 153301 7327
rect 153335 7324 153347 7327
rect 154301 7327 154359 7333
rect 154301 7324 154313 7327
rect 153335 7296 154313 7324
rect 153335 7293 153347 7296
rect 153289 7287 153347 7293
rect 154301 7293 154313 7296
rect 154347 7324 154359 7327
rect 155218 7324 155224 7336
rect 154347 7296 155224 7324
rect 154347 7293 154359 7296
rect 154301 7287 154359 7293
rect 155218 7284 155224 7296
rect 155276 7284 155282 7336
rect 155310 7284 155316 7336
rect 155368 7324 155374 7336
rect 159910 7324 159916 7336
rect 155368 7296 155413 7324
rect 159871 7296 159916 7324
rect 155368 7284 155374 7296
rect 159910 7284 159916 7296
rect 159968 7284 159974 7336
rect 160830 7284 160836 7336
rect 160888 7324 160894 7336
rect 161109 7327 161167 7333
rect 161109 7324 161121 7327
rect 160888 7296 161121 7324
rect 160888 7284 160894 7296
rect 161109 7293 161121 7296
rect 161155 7293 161167 7327
rect 161109 7287 161167 7293
rect 162765 7327 162823 7333
rect 162765 7293 162777 7327
rect 162811 7324 162823 7327
rect 163314 7324 163320 7336
rect 162811 7296 163320 7324
rect 162811 7293 162823 7296
rect 162765 7287 162823 7293
rect 163314 7284 163320 7296
rect 163372 7324 163378 7336
rect 163869 7327 163927 7333
rect 163869 7324 163881 7327
rect 163372 7296 163881 7324
rect 163372 7284 163378 7296
rect 163869 7293 163881 7296
rect 163915 7293 163927 7327
rect 163869 7287 163927 7293
rect 164234 7284 164240 7336
rect 164292 7324 164298 7336
rect 164881 7327 164939 7333
rect 164881 7324 164893 7327
rect 164292 7296 164893 7324
rect 164292 7284 164298 7296
rect 164881 7293 164893 7296
rect 164927 7293 164939 7327
rect 164881 7287 164939 7293
rect 134886 7188 134892 7200
rect 115308 7160 122420 7188
rect 134847 7160 134892 7188
rect 104400 7148 104406 7160
rect 134886 7148 134892 7160
rect 134944 7148 134950 7200
rect 141786 7188 141792 7200
rect 141747 7160 141792 7188
rect 141786 7148 141792 7160
rect 141844 7148 141850 7200
rect 153010 7188 153016 7200
rect 152971 7160 153016 7188
rect 153010 7148 153016 7160
rect 153068 7148 153074 7200
rect 163498 7188 163504 7200
rect 163459 7160 163504 7188
rect 163498 7148 163504 7160
rect 163556 7148 163562 7200
rect 368 7098 93012 7120
rect 368 7046 28456 7098
rect 28508 7046 28520 7098
rect 28572 7046 28584 7098
rect 28636 7046 28648 7098
rect 28700 7046 84878 7098
rect 84930 7046 84942 7098
rect 84994 7046 85006 7098
rect 85058 7046 85070 7098
rect 85122 7046 93012 7098
rect 368 7024 93012 7046
rect 102028 7098 169556 7120
rect 102028 7046 141299 7098
rect 141351 7046 141363 7098
rect 141415 7046 141427 7098
rect 141479 7046 141491 7098
rect 141543 7046 169556 7098
rect 102028 7024 169556 7046
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 14001 6987 14059 6993
rect 4856 6956 11008 6984
rect 4856 6944 4862 6956
rect 5718 6916 5724 6928
rect 5679 6888 5724 6916
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 10229 6919 10287 6925
rect 10229 6916 10241 6919
rect 9824 6888 10241 6916
rect 9824 6876 9830 6888
rect 10229 6885 10241 6888
rect 10275 6885 10287 6919
rect 10980 6916 11008 6956
rect 14001 6953 14013 6987
rect 14047 6984 14059 6987
rect 14090 6984 14096 6996
rect 14047 6956 14096 6984
rect 14047 6953 14059 6956
rect 14001 6947 14059 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 23658 6984 23664 6996
rect 15528 6956 23520 6984
rect 23619 6956 23664 6984
rect 15528 6944 15534 6956
rect 22741 6919 22799 6925
rect 22741 6916 22753 6919
rect 10980 6888 22753 6916
rect 10229 6879 10287 6885
rect 22741 6885 22753 6888
rect 22787 6885 22799 6919
rect 23492 6916 23520 6956
rect 23658 6944 23664 6956
rect 23716 6944 23722 6996
rect 23842 6944 23848 6996
rect 23900 6984 23906 6996
rect 26234 6984 26240 6996
rect 23900 6956 26240 6984
rect 23900 6944 23906 6956
rect 26234 6944 26240 6956
rect 26292 6944 26298 6996
rect 26421 6987 26479 6993
rect 26421 6953 26433 6987
rect 26467 6984 26479 6987
rect 26510 6984 26516 6996
rect 26467 6956 26516 6984
rect 26467 6953 26479 6956
rect 26421 6947 26479 6953
rect 26510 6944 26516 6956
rect 26568 6944 26574 6996
rect 26602 6944 26608 6996
rect 26660 6984 26666 6996
rect 28810 6984 28816 6996
rect 26660 6956 28816 6984
rect 26660 6944 26666 6956
rect 28810 6944 28816 6956
rect 28868 6944 28874 6996
rect 33778 6944 33784 6996
rect 33836 6984 33842 6996
rect 36446 6984 36452 6996
rect 33836 6956 36452 6984
rect 33836 6944 33842 6956
rect 36446 6944 36452 6956
rect 36504 6944 36510 6996
rect 36906 6944 36912 6996
rect 36964 6984 36970 6996
rect 38286 6984 38292 6996
rect 36964 6956 38292 6984
rect 36964 6944 36970 6956
rect 38286 6944 38292 6956
rect 38344 6944 38350 6996
rect 38470 6984 38476 6996
rect 38431 6956 38476 6984
rect 38470 6944 38476 6956
rect 38528 6944 38534 6996
rect 38838 6944 38844 6996
rect 38896 6984 38902 6996
rect 39390 6984 39396 6996
rect 38896 6956 39396 6984
rect 38896 6944 38902 6956
rect 39390 6944 39396 6956
rect 39448 6944 39454 6996
rect 39482 6944 39488 6996
rect 39540 6984 39546 6996
rect 41414 6984 41420 6996
rect 39540 6956 41420 6984
rect 39540 6944 39546 6956
rect 41414 6944 41420 6956
rect 41472 6944 41478 6996
rect 41782 6984 41788 6996
rect 41616 6956 41788 6984
rect 37093 6919 37151 6925
rect 37093 6916 37105 6919
rect 23492 6888 36676 6916
rect 22741 6879 22799 6885
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 3602 6848 3608 6860
rect 3467 6820 3608 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 3602 6808 3608 6820
rect 3660 6848 3666 6860
rect 3881 6851 3939 6857
rect 3881 6848 3893 6851
rect 3660 6820 3893 6848
rect 3660 6808 3666 6820
rect 3881 6817 3893 6820
rect 3927 6817 3939 6851
rect 6362 6848 6368 6860
rect 3881 6811 3939 6817
rect 6012 6820 6368 6848
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 6012 6789 6040 6820
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 7837 6851 7895 6857
rect 7837 6817 7849 6851
rect 7883 6848 7895 6851
rect 7926 6848 7932 6860
rect 7883 6820 7932 6848
rect 7883 6817 7895 6820
rect 7837 6811 7895 6817
rect 7926 6808 7932 6820
rect 7984 6848 7990 6860
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 7984 6820 8309 6848
rect 7984 6808 7990 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 8938 6848 8944 6860
rect 8803 6820 8944 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13412 6820 13461 6848
rect 13412 6808 13418 6820
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 14274 6848 14280 6860
rect 14235 6820 14280 6848
rect 13449 6811 13507 6817
rect 14274 6808 14280 6820
rect 14332 6848 14338 6860
rect 14553 6851 14611 6857
rect 14553 6848 14565 6851
rect 14332 6820 14565 6848
rect 14332 6808 14338 6820
rect 14553 6817 14565 6820
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 15286 6808 15292 6860
rect 15344 6848 15350 6860
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15344 6820 15577 6848
rect 15344 6808 15350 6820
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 19061 6851 19119 6857
rect 19061 6817 19073 6851
rect 19107 6848 19119 6851
rect 19518 6848 19524 6860
rect 19107 6820 19524 6848
rect 19107 6817 19119 6820
rect 19061 6811 19119 6817
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 19886 6848 19892 6860
rect 19847 6820 19892 6848
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 20441 6851 20499 6857
rect 20441 6817 20453 6851
rect 20487 6848 20499 6851
rect 20898 6848 20904 6860
rect 20487 6820 20904 6848
rect 20487 6817 20499 6820
rect 20441 6811 20499 6817
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 20993 6851 21051 6857
rect 20993 6817 21005 6851
rect 21039 6848 21051 6851
rect 21358 6848 21364 6860
rect 21039 6820 21364 6848
rect 21039 6817 21051 6820
rect 20993 6811 21051 6817
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 23658 6808 23664 6860
rect 23716 6848 23722 6860
rect 23845 6851 23903 6857
rect 23845 6848 23857 6851
rect 23716 6820 23857 6848
rect 23716 6808 23722 6820
rect 23845 6817 23857 6820
rect 23891 6817 23903 6851
rect 26510 6848 26516 6860
rect 26471 6820 26516 6848
rect 23845 6811 23903 6817
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 26786 6808 26792 6860
rect 26844 6848 26850 6860
rect 27525 6851 27583 6857
rect 27525 6848 27537 6851
rect 26844 6820 27537 6848
rect 26844 6808 26850 6820
rect 27525 6817 27537 6820
rect 27571 6817 27583 6851
rect 29270 6848 29276 6860
rect 27525 6811 27583 6817
rect 27632 6820 29276 6848
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4304 6752 4353 6780
rect 4304 6740 4310 6752
rect 4341 6749 4353 6752
rect 4387 6780 4399 6783
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 4387 6752 4445 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4433 6749 4445 6752
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 21082 6780 21088 6792
rect 18095 6752 21088 6780
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 10520 6644 10548 6743
rect 16132 6712 16160 6743
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 16482 6712 16488 6724
rect 16132 6684 16488 6712
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 10870 6644 10876 6656
rect 10520 6616 10876 6644
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 21266 6644 21272 6656
rect 21227 6616 21272 6644
rect 21266 6604 21272 6616
rect 21324 6644 21330 6656
rect 21468 6644 21496 6743
rect 22462 6740 22468 6792
rect 22520 6780 22526 6792
rect 22557 6783 22615 6789
rect 22557 6780 22569 6783
rect 22520 6752 22569 6780
rect 22520 6740 22526 6752
rect 22557 6749 22569 6752
rect 22603 6780 22615 6783
rect 23293 6783 23351 6789
rect 23293 6780 23305 6783
rect 22603 6752 23305 6780
rect 22603 6749 22615 6752
rect 22557 6743 22615 6749
rect 23293 6749 23305 6752
rect 23339 6749 23351 6783
rect 23293 6743 23351 6749
rect 26234 6740 26240 6792
rect 26292 6780 26298 6792
rect 27632 6780 27660 6820
rect 29270 6808 29276 6820
rect 29328 6808 29334 6860
rect 33597 6851 33655 6857
rect 29380 6820 30236 6848
rect 27982 6780 27988 6792
rect 26292 6752 27660 6780
rect 27943 6752 27988 6780
rect 26292 6740 26298 6752
rect 27982 6740 27988 6752
rect 28040 6740 28046 6792
rect 28166 6740 28172 6792
rect 28224 6780 28230 6792
rect 29380 6780 29408 6820
rect 28224 6752 29408 6780
rect 30208 6780 30236 6820
rect 33597 6817 33609 6851
rect 33643 6848 33655 6851
rect 34057 6851 34115 6857
rect 34057 6848 34069 6851
rect 33643 6820 34069 6848
rect 33643 6817 33655 6820
rect 33597 6811 33655 6817
rect 34057 6817 34069 6820
rect 34103 6817 34115 6851
rect 34793 6851 34851 6857
rect 34793 6848 34805 6851
rect 34057 6811 34115 6817
rect 34440 6820 34805 6848
rect 33778 6780 33784 6792
rect 30208 6752 33784 6780
rect 28224 6740 28230 6752
rect 33778 6740 33784 6752
rect 33836 6740 33842 6792
rect 33962 6780 33968 6792
rect 33875 6752 33968 6780
rect 33962 6740 33968 6752
rect 34020 6740 34026 6792
rect 34440 6789 34468 6820
rect 34793 6817 34805 6820
rect 34839 6848 34851 6851
rect 35434 6848 35440 6860
rect 34839 6820 35440 6848
rect 34839 6817 34851 6820
rect 34793 6811 34851 6817
rect 35434 6808 35440 6820
rect 35492 6808 35498 6860
rect 35526 6808 35532 6860
rect 35584 6848 35590 6860
rect 36354 6848 36360 6860
rect 35584 6820 36360 6848
rect 35584 6808 35590 6820
rect 36354 6808 36360 6820
rect 36412 6808 36418 6860
rect 34425 6783 34483 6789
rect 34425 6749 34437 6783
rect 34471 6749 34483 6783
rect 34425 6743 34483 6749
rect 34698 6740 34704 6792
rect 34756 6780 34762 6792
rect 36078 6780 36084 6792
rect 34756 6752 36084 6780
rect 34756 6740 34762 6752
rect 36078 6740 36084 6752
rect 36136 6740 36142 6792
rect 36262 6780 36268 6792
rect 36223 6752 36268 6780
rect 36262 6740 36268 6752
rect 36320 6740 36326 6792
rect 36648 6780 36676 6888
rect 36740 6888 37105 6916
rect 36740 6860 36768 6888
rect 37093 6885 37105 6888
rect 37139 6885 37151 6919
rect 41141 6919 41199 6925
rect 41141 6916 41153 6919
rect 37093 6879 37151 6885
rect 37200 6888 41153 6916
rect 36722 6808 36728 6860
rect 36780 6808 36786 6860
rect 37200 6848 37228 6888
rect 41141 6885 41153 6888
rect 41187 6885 41199 6919
rect 41616 6916 41644 6956
rect 41782 6944 41788 6956
rect 41840 6944 41846 6996
rect 45094 6984 45100 6996
rect 41892 6956 45100 6984
rect 41141 6879 41199 6885
rect 41248 6888 41644 6916
rect 36832 6820 37228 6848
rect 37829 6851 37887 6857
rect 36832 6780 36860 6820
rect 37829 6817 37841 6851
rect 37875 6848 37887 6851
rect 40310 6848 40316 6860
rect 37875 6820 40316 6848
rect 37875 6817 37887 6820
rect 37829 6811 37887 6817
rect 40310 6808 40316 6820
rect 40368 6808 40374 6860
rect 40586 6808 40592 6860
rect 40644 6848 40650 6860
rect 41248 6848 41276 6888
rect 41690 6876 41696 6928
rect 41748 6916 41754 6928
rect 41892 6916 41920 6956
rect 45094 6944 45100 6956
rect 45152 6944 45158 6996
rect 45462 6944 45468 6996
rect 45520 6984 45526 6996
rect 46658 6984 46664 6996
rect 45520 6956 46664 6984
rect 45520 6944 45526 6956
rect 46658 6944 46664 6956
rect 46716 6944 46722 6996
rect 46750 6944 46756 6996
rect 46808 6984 46814 6996
rect 46845 6987 46903 6993
rect 46845 6984 46857 6987
rect 46808 6956 46857 6984
rect 46808 6944 46814 6956
rect 46845 6953 46857 6956
rect 46891 6953 46903 6987
rect 46845 6947 46903 6953
rect 47118 6944 47124 6996
rect 47176 6984 47182 6996
rect 48866 6984 48872 6996
rect 47176 6956 48872 6984
rect 47176 6944 47182 6956
rect 48866 6944 48872 6956
rect 48924 6944 48930 6996
rect 48958 6944 48964 6996
rect 49016 6984 49022 6996
rect 50246 6984 50252 6996
rect 49016 6956 50252 6984
rect 49016 6944 49022 6956
rect 50246 6944 50252 6956
rect 50304 6944 50310 6996
rect 50338 6944 50344 6996
rect 50396 6984 50402 6996
rect 51077 6987 51135 6993
rect 51077 6984 51089 6987
rect 50396 6956 51089 6984
rect 50396 6944 50402 6956
rect 51077 6953 51089 6956
rect 51123 6953 51135 6987
rect 51077 6947 51135 6953
rect 51442 6944 51448 6996
rect 51500 6984 51506 6996
rect 52454 6984 52460 6996
rect 51500 6956 52460 6984
rect 51500 6944 51506 6956
rect 52454 6944 52460 6956
rect 52512 6944 52518 6996
rect 52730 6944 52736 6996
rect 52788 6984 52794 6996
rect 54110 6984 54116 6996
rect 52788 6956 54116 6984
rect 52788 6944 52794 6956
rect 54110 6944 54116 6956
rect 54168 6944 54174 6996
rect 55122 6944 55128 6996
rect 55180 6984 55186 6996
rect 57057 6987 57115 6993
rect 57057 6984 57069 6987
rect 55180 6956 57069 6984
rect 55180 6944 55186 6956
rect 57057 6953 57069 6956
rect 57103 6953 57115 6987
rect 57330 6984 57336 6996
rect 57291 6956 57336 6984
rect 57057 6947 57115 6953
rect 57330 6944 57336 6956
rect 57388 6944 57394 6996
rect 57514 6944 57520 6996
rect 57572 6984 57578 6996
rect 57698 6984 57704 6996
rect 57572 6956 57704 6984
rect 57572 6944 57578 6956
rect 57698 6944 57704 6956
rect 57756 6944 57762 6996
rect 58897 6987 58955 6993
rect 58897 6953 58909 6987
rect 58943 6984 58955 6987
rect 59078 6984 59084 6996
rect 58943 6956 59084 6984
rect 58943 6953 58955 6956
rect 58897 6947 58955 6953
rect 59078 6944 59084 6956
rect 59136 6944 59142 6996
rect 68830 6984 68836 6996
rect 68791 6956 68836 6984
rect 68830 6944 68836 6956
rect 68888 6944 68894 6996
rect 70118 6984 70124 6996
rect 70079 6956 70124 6984
rect 70118 6944 70124 6956
rect 70176 6944 70182 6996
rect 80977 6987 81035 6993
rect 80977 6953 80989 6987
rect 81023 6984 81035 6987
rect 88150 6984 88156 6996
rect 81023 6956 88156 6984
rect 81023 6953 81035 6956
rect 80977 6947 81035 6953
rect 88150 6944 88156 6956
rect 88208 6944 88214 6996
rect 95326 6944 95332 6996
rect 95384 6984 95390 6996
rect 113361 6987 113419 6993
rect 95384 6956 111840 6984
rect 95384 6944 95390 6956
rect 41748 6888 41920 6916
rect 41748 6876 41754 6888
rect 42150 6876 42156 6928
rect 42208 6916 42214 6928
rect 42705 6919 42763 6925
rect 42705 6916 42717 6919
rect 42208 6888 42717 6916
rect 42208 6876 42214 6888
rect 42705 6885 42717 6888
rect 42751 6885 42763 6919
rect 50706 6916 50712 6928
rect 42705 6879 42763 6885
rect 42812 6888 50712 6916
rect 40644 6820 41276 6848
rect 40644 6808 40650 6820
rect 41414 6808 41420 6860
rect 41472 6848 41478 6860
rect 42518 6848 42524 6860
rect 41472 6820 42524 6848
rect 41472 6808 41478 6820
rect 42518 6808 42524 6820
rect 42576 6808 42582 6860
rect 42610 6808 42616 6860
rect 42668 6848 42674 6860
rect 42668 6820 42748 6848
rect 42668 6808 42674 6820
rect 37274 6780 37280 6792
rect 36648 6752 36860 6780
rect 37235 6752 37280 6780
rect 37274 6740 37280 6752
rect 37332 6740 37338 6792
rect 37737 6783 37795 6789
rect 37737 6749 37749 6783
rect 37783 6780 37795 6783
rect 38010 6780 38016 6792
rect 37783 6752 38016 6780
rect 37783 6749 37795 6752
rect 37737 6743 37795 6749
rect 38010 6740 38016 6752
rect 38068 6740 38074 6792
rect 39758 6780 39764 6792
rect 39671 6752 39764 6780
rect 39758 6740 39764 6752
rect 39816 6780 39822 6792
rect 39853 6783 39911 6789
rect 39853 6780 39865 6783
rect 39816 6752 39865 6780
rect 39816 6740 39822 6752
rect 39853 6749 39865 6752
rect 39899 6749 39911 6783
rect 39853 6743 39911 6749
rect 39942 6740 39948 6792
rect 40000 6780 40006 6792
rect 41230 6780 41236 6792
rect 40000 6752 41236 6780
rect 40000 6740 40006 6752
rect 41230 6740 41236 6752
rect 41288 6740 41294 6792
rect 41325 6783 41383 6789
rect 41325 6749 41337 6783
rect 41371 6780 41383 6783
rect 41598 6780 41604 6792
rect 41371 6752 41604 6780
rect 41371 6749 41383 6752
rect 41325 6743 41383 6749
rect 41598 6740 41604 6752
rect 41656 6780 41662 6792
rect 41966 6780 41972 6792
rect 41656 6752 41972 6780
rect 41656 6740 41662 6752
rect 41966 6740 41972 6752
rect 42024 6740 42030 6792
rect 42242 6740 42248 6792
rect 42300 6780 42306 6792
rect 42720 6789 42748 6820
rect 42705 6783 42763 6789
rect 42300 6752 42656 6780
rect 42300 6740 42306 6752
rect 21634 6672 21640 6724
rect 21692 6712 21698 6724
rect 24762 6712 24768 6724
rect 21692 6684 24768 6712
rect 21692 6672 21698 6684
rect 24762 6672 24768 6684
rect 24820 6672 24826 6724
rect 25130 6672 25136 6724
rect 25188 6712 25194 6724
rect 33597 6715 33655 6721
rect 33597 6712 33609 6715
rect 25188 6684 33609 6712
rect 25188 6672 25194 6684
rect 33597 6681 33609 6684
rect 33643 6681 33655 6715
rect 33980 6712 34008 6740
rect 35253 6715 35311 6721
rect 35253 6712 35265 6715
rect 33980 6684 35265 6712
rect 33597 6675 33655 6681
rect 35253 6681 35265 6684
rect 35299 6681 35311 6715
rect 36630 6712 36636 6724
rect 35253 6675 35311 6681
rect 35360 6684 36636 6712
rect 25038 6644 25044 6656
rect 21324 6616 21496 6644
rect 24951 6616 25044 6644
rect 21324 6604 21330 6616
rect 25038 6604 25044 6616
rect 25096 6644 25102 6656
rect 27798 6644 27804 6656
rect 25096 6616 27804 6644
rect 25096 6604 25102 6616
rect 27798 6604 27804 6616
rect 27856 6604 27862 6656
rect 27982 6604 27988 6656
rect 28040 6644 28046 6656
rect 28258 6644 28264 6656
rect 28040 6616 28264 6644
rect 28040 6604 28046 6616
rect 28258 6604 28264 6616
rect 28316 6604 28322 6656
rect 28350 6604 28356 6656
rect 28408 6644 28414 6656
rect 28445 6647 28503 6653
rect 28445 6644 28457 6647
rect 28408 6616 28457 6644
rect 28408 6604 28414 6616
rect 28445 6613 28457 6616
rect 28491 6644 28503 6647
rect 35360 6644 35388 6684
rect 36630 6672 36636 6684
rect 36688 6672 36694 6724
rect 36725 6715 36783 6721
rect 36725 6681 36737 6715
rect 36771 6712 36783 6715
rect 36906 6712 36912 6724
rect 36771 6684 36912 6712
rect 36771 6681 36783 6684
rect 36725 6675 36783 6681
rect 36906 6672 36912 6684
rect 36964 6672 36970 6724
rect 36998 6672 37004 6724
rect 37056 6712 37062 6724
rect 42518 6712 42524 6724
rect 37056 6684 42524 6712
rect 37056 6672 37062 6684
rect 42518 6672 42524 6684
rect 42576 6672 42582 6724
rect 42628 6712 42656 6752
rect 42705 6749 42717 6783
rect 42751 6749 42763 6783
rect 42705 6743 42763 6749
rect 42812 6712 42840 6888
rect 50706 6876 50712 6888
rect 50764 6876 50770 6928
rect 50890 6876 50896 6928
rect 50948 6916 50954 6928
rect 55674 6916 55680 6928
rect 50948 6888 55680 6916
rect 50948 6876 50954 6888
rect 55674 6876 55680 6888
rect 55732 6876 55738 6928
rect 56502 6876 56508 6928
rect 56560 6916 56566 6928
rect 57422 6916 57428 6928
rect 56560 6888 57428 6916
rect 56560 6876 56566 6888
rect 57422 6876 57428 6888
rect 57480 6876 57486 6928
rect 57974 6876 57980 6928
rect 58032 6916 58038 6928
rect 79965 6919 80023 6925
rect 79965 6916 79977 6919
rect 58032 6888 79977 6916
rect 58032 6876 58038 6888
rect 79965 6885 79977 6888
rect 80011 6885 80023 6919
rect 83182 6916 83188 6928
rect 83143 6888 83188 6916
rect 79965 6879 80023 6885
rect 83182 6876 83188 6888
rect 83240 6876 83246 6928
rect 87782 6916 87788 6928
rect 87743 6888 87788 6916
rect 87782 6876 87788 6888
rect 87840 6876 87846 6928
rect 101692 6888 101904 6916
rect 43622 6808 43628 6860
rect 43680 6848 43686 6860
rect 45554 6848 45560 6860
rect 43680 6820 45560 6848
rect 43680 6808 43686 6820
rect 45554 6808 45560 6820
rect 45612 6808 45618 6860
rect 45649 6851 45707 6857
rect 45649 6817 45661 6851
rect 45695 6848 45707 6851
rect 51813 6851 51871 6857
rect 45695 6820 51672 6848
rect 45695 6817 45707 6820
rect 45649 6811 45707 6817
rect 43349 6783 43407 6789
rect 43349 6749 43361 6783
rect 43395 6780 43407 6783
rect 43714 6780 43720 6792
rect 43395 6752 43720 6780
rect 43395 6749 43407 6752
rect 43349 6743 43407 6749
rect 43714 6740 43720 6752
rect 43772 6740 43778 6792
rect 44910 6780 44916 6792
rect 44871 6752 44916 6780
rect 44910 6740 44916 6752
rect 44968 6740 44974 6792
rect 45097 6783 45155 6789
rect 45097 6749 45109 6783
rect 45143 6780 45155 6783
rect 45370 6780 45376 6792
rect 45143 6752 45376 6780
rect 45143 6749 45155 6752
rect 45097 6743 45155 6749
rect 45370 6740 45376 6752
rect 45428 6740 45434 6792
rect 45465 6783 45523 6789
rect 45465 6749 45477 6783
rect 45511 6780 45523 6783
rect 45833 6783 45891 6789
rect 45833 6780 45845 6783
rect 45511 6752 45845 6780
rect 45511 6749 45523 6752
rect 45465 6743 45523 6749
rect 45833 6749 45845 6752
rect 45879 6780 45891 6783
rect 46934 6780 46940 6792
rect 45879 6752 46940 6780
rect 45879 6749 45891 6752
rect 45833 6743 45891 6749
rect 46934 6740 46940 6752
rect 46992 6740 46998 6792
rect 47394 6740 47400 6792
rect 47452 6780 47458 6792
rect 48130 6780 48136 6792
rect 47452 6752 48136 6780
rect 47452 6740 47458 6752
rect 48130 6740 48136 6752
rect 48188 6740 48194 6792
rect 48317 6783 48375 6789
rect 48317 6749 48329 6783
rect 48363 6780 48375 6783
rect 49786 6780 49792 6792
rect 48363 6752 49792 6780
rect 48363 6749 48375 6752
rect 48317 6743 48375 6749
rect 49786 6740 49792 6752
rect 49844 6740 49850 6792
rect 49973 6783 50031 6789
rect 49973 6749 49985 6783
rect 50019 6780 50031 6783
rect 51258 6780 51264 6792
rect 50019 6752 51264 6780
rect 50019 6749 50031 6752
rect 49973 6743 50031 6749
rect 51258 6740 51264 6752
rect 51316 6740 51322 6792
rect 51537 6783 51595 6789
rect 51537 6749 51549 6783
rect 51583 6749 51595 6783
rect 51644 6780 51672 6820
rect 51813 6817 51825 6851
rect 51859 6848 51871 6851
rect 52089 6851 52147 6857
rect 52089 6848 52101 6851
rect 51859 6820 52101 6848
rect 51859 6817 51871 6820
rect 51813 6811 51871 6817
rect 52089 6817 52101 6820
rect 52135 6848 52147 6851
rect 52178 6848 52184 6860
rect 52135 6820 52184 6848
rect 52135 6817 52147 6820
rect 52089 6811 52147 6817
rect 52178 6808 52184 6820
rect 52236 6808 52242 6860
rect 52270 6808 52276 6860
rect 52328 6848 52334 6860
rect 53190 6848 53196 6860
rect 52328 6820 53196 6848
rect 52328 6808 52334 6820
rect 53190 6808 53196 6820
rect 53248 6808 53254 6860
rect 54389 6851 54447 6857
rect 54389 6817 54401 6851
rect 54435 6848 54447 6851
rect 56134 6848 56140 6860
rect 54435 6820 56140 6848
rect 54435 6817 54447 6820
rect 54389 6811 54447 6817
rect 56134 6808 56140 6820
rect 56192 6848 56198 6860
rect 56873 6851 56931 6857
rect 56873 6848 56885 6851
rect 56192 6820 56885 6848
rect 56192 6808 56198 6820
rect 56873 6817 56885 6820
rect 56919 6817 56931 6851
rect 56873 6811 56931 6817
rect 57057 6851 57115 6857
rect 57057 6817 57069 6851
rect 57103 6848 57115 6851
rect 57330 6848 57336 6860
rect 57103 6820 57336 6848
rect 57103 6817 57115 6820
rect 57057 6811 57115 6817
rect 57330 6808 57336 6820
rect 57388 6808 57394 6860
rect 58250 6848 58256 6860
rect 57440 6820 58256 6848
rect 54754 6780 54760 6792
rect 51644 6752 54760 6780
rect 51537 6743 51595 6749
rect 42628 6684 42840 6712
rect 42886 6672 42892 6724
rect 42944 6712 42950 6724
rect 45649 6715 45707 6721
rect 45649 6712 45661 6715
rect 42944 6684 45661 6712
rect 42944 6672 42950 6684
rect 45649 6681 45661 6684
rect 45695 6681 45707 6715
rect 50522 6712 50528 6724
rect 45649 6675 45707 6681
rect 45756 6684 50528 6712
rect 28491 6616 35388 6644
rect 28491 6613 28503 6616
rect 28445 6607 28503 6613
rect 35434 6604 35440 6656
rect 35492 6644 35498 6656
rect 37829 6647 37887 6653
rect 37829 6644 37841 6647
rect 35492 6616 37841 6644
rect 35492 6604 35498 6616
rect 37829 6613 37841 6616
rect 37875 6613 37887 6647
rect 38010 6644 38016 6656
rect 37971 6616 38016 6644
rect 37829 6607 37887 6613
rect 38010 6604 38016 6616
rect 38068 6604 38074 6656
rect 38838 6644 38844 6656
rect 38799 6616 38844 6644
rect 38838 6604 38844 6616
rect 38896 6604 38902 6656
rect 38930 6604 38936 6656
rect 38988 6644 38994 6656
rect 41414 6644 41420 6656
rect 38988 6616 41420 6644
rect 38988 6604 38994 6616
rect 41414 6604 41420 6616
rect 41472 6604 41478 6656
rect 41506 6604 41512 6656
rect 41564 6644 41570 6656
rect 41693 6647 41751 6653
rect 41693 6644 41705 6647
rect 41564 6616 41705 6644
rect 41564 6604 41570 6616
rect 41693 6613 41705 6616
rect 41739 6644 41751 6647
rect 45756 6644 45784 6684
rect 50522 6672 50528 6684
rect 50580 6672 50586 6724
rect 50614 6672 50620 6724
rect 50672 6712 50678 6724
rect 51442 6712 51448 6724
rect 50672 6684 51448 6712
rect 50672 6672 50678 6684
rect 51442 6672 51448 6684
rect 51500 6672 51506 6724
rect 51552 6712 51580 6743
rect 54754 6740 54760 6752
rect 54812 6740 54818 6792
rect 55401 6783 55459 6789
rect 55401 6749 55413 6783
rect 55447 6780 55459 6783
rect 56226 6780 56232 6792
rect 55447 6752 56232 6780
rect 55447 6749 55459 6752
rect 55401 6743 55459 6749
rect 56226 6740 56232 6752
rect 56284 6740 56290 6792
rect 56318 6740 56324 6792
rect 56376 6780 56382 6792
rect 57440 6780 57468 6820
rect 58250 6808 58256 6820
rect 58308 6808 58314 6860
rect 59909 6851 59967 6857
rect 59909 6817 59921 6851
rect 59955 6848 59967 6851
rect 60274 6848 60280 6860
rect 59955 6820 60280 6848
rect 59955 6817 59967 6820
rect 59909 6811 59967 6817
rect 60274 6808 60280 6820
rect 60332 6808 60338 6860
rect 60458 6808 60464 6860
rect 60516 6848 60522 6860
rect 60921 6851 60979 6857
rect 60921 6848 60933 6851
rect 60516 6820 60933 6848
rect 60516 6808 60522 6820
rect 60921 6817 60933 6820
rect 60967 6817 60979 6851
rect 63402 6848 63408 6860
rect 60921 6811 60979 6817
rect 61396 6820 63408 6848
rect 57606 6780 57612 6792
rect 56376 6752 57468 6780
rect 57567 6752 57612 6780
rect 56376 6740 56382 6752
rect 57606 6740 57612 6752
rect 57664 6740 57670 6792
rect 57793 6783 57851 6789
rect 57793 6749 57805 6783
rect 57839 6780 57851 6783
rect 57882 6780 57888 6792
rect 57839 6752 57888 6780
rect 57839 6749 57851 6752
rect 57793 6743 57851 6749
rect 57882 6740 57888 6752
rect 57940 6740 57946 6792
rect 58158 6780 58164 6792
rect 58119 6752 58164 6780
rect 58158 6740 58164 6752
rect 58216 6780 58222 6792
rect 58437 6783 58495 6789
rect 58437 6780 58449 6783
rect 58216 6752 58449 6780
rect 58216 6740 58222 6752
rect 58437 6749 58449 6752
rect 58483 6749 58495 6783
rect 58437 6743 58495 6749
rect 58526 6740 58532 6792
rect 58584 6780 58590 6792
rect 61396 6780 61424 6820
rect 63402 6808 63408 6820
rect 63460 6808 63466 6860
rect 65426 6808 65432 6860
rect 65484 6848 65490 6860
rect 73246 6848 73252 6860
rect 65484 6820 73252 6848
rect 65484 6808 65490 6820
rect 73246 6808 73252 6820
rect 73304 6808 73310 6860
rect 79597 6851 79655 6857
rect 79597 6817 79609 6851
rect 79643 6848 79655 6851
rect 79778 6848 79784 6860
rect 79643 6820 79784 6848
rect 79643 6817 79655 6820
rect 79597 6811 79655 6817
rect 79778 6808 79784 6820
rect 79836 6848 79842 6860
rect 80057 6851 80115 6857
rect 80057 6848 80069 6851
rect 79836 6820 80069 6848
rect 79836 6808 79842 6820
rect 80057 6817 80069 6820
rect 80103 6817 80115 6851
rect 81894 6848 81900 6860
rect 81855 6820 81900 6848
rect 80057 6811 80115 6817
rect 81894 6808 81900 6820
rect 81952 6808 81958 6860
rect 87598 6808 87604 6860
rect 87656 6848 87662 6860
rect 88153 6851 88211 6857
rect 88153 6848 88165 6851
rect 87656 6820 88165 6848
rect 87656 6808 87662 6820
rect 88153 6817 88165 6820
rect 88199 6848 88211 6851
rect 88337 6851 88395 6857
rect 88337 6848 88349 6851
rect 88199 6820 88349 6848
rect 88199 6817 88211 6820
rect 88153 6811 88211 6817
rect 88337 6817 88349 6820
rect 88383 6817 88395 6851
rect 88337 6811 88395 6817
rect 88426 6808 88432 6860
rect 88484 6848 88490 6860
rect 89349 6851 89407 6857
rect 89349 6848 89361 6851
rect 88484 6820 89361 6848
rect 88484 6808 88490 6820
rect 89349 6817 89361 6820
rect 89395 6817 89407 6851
rect 89349 6811 89407 6817
rect 91741 6851 91799 6857
rect 91741 6817 91753 6851
rect 91787 6848 91799 6851
rect 95602 6848 95608 6860
rect 91787 6820 95608 6848
rect 91787 6817 91799 6820
rect 91741 6811 91799 6817
rect 95602 6808 95608 6820
rect 95660 6808 95666 6860
rect 101493 6851 101551 6857
rect 101493 6848 101505 6851
rect 95712 6820 101505 6848
rect 58584 6752 61424 6780
rect 61473 6783 61531 6789
rect 58584 6740 58590 6752
rect 61473 6749 61485 6783
rect 61519 6780 61531 6783
rect 61841 6783 61899 6789
rect 61841 6780 61853 6783
rect 61519 6752 61853 6780
rect 61519 6749 61531 6752
rect 61473 6743 61531 6749
rect 61841 6749 61853 6752
rect 61887 6780 61899 6783
rect 74718 6780 74724 6792
rect 61887 6752 74724 6780
rect 61887 6749 61899 6752
rect 61841 6743 61899 6749
rect 74718 6740 74724 6752
rect 74776 6740 74782 6792
rect 82814 6740 82820 6792
rect 82872 6780 82878 6792
rect 83001 6783 83059 6789
rect 83001 6780 83013 6783
rect 82872 6752 83013 6780
rect 82872 6740 82878 6752
rect 83001 6749 83013 6752
rect 83047 6780 83059 6783
rect 83737 6783 83795 6789
rect 83737 6780 83749 6783
rect 83047 6752 83749 6780
rect 83047 6749 83059 6752
rect 83001 6743 83059 6749
rect 83737 6749 83749 6752
rect 83783 6749 83795 6783
rect 83737 6743 83795 6749
rect 89901 6783 89959 6789
rect 89901 6749 89913 6783
rect 89947 6749 89959 6783
rect 89901 6743 89959 6749
rect 51813 6715 51871 6721
rect 51813 6712 51825 6715
rect 51552 6684 51825 6712
rect 51813 6681 51825 6684
rect 51859 6681 51871 6715
rect 72050 6712 72056 6724
rect 51813 6675 51871 6681
rect 52196 6684 72056 6712
rect 41739 6616 45784 6644
rect 41739 6613 41751 6616
rect 41693 6607 41751 6613
rect 45830 6604 45836 6656
rect 45888 6644 45894 6656
rect 46293 6647 46351 6653
rect 46293 6644 46305 6647
rect 45888 6616 46305 6644
rect 45888 6604 45894 6616
rect 46293 6613 46305 6616
rect 46339 6613 46351 6647
rect 46293 6607 46351 6613
rect 46474 6604 46480 6656
rect 46532 6644 46538 6656
rect 48317 6647 48375 6653
rect 48317 6644 48329 6647
rect 46532 6616 48329 6644
rect 46532 6604 46538 6616
rect 48317 6613 48329 6616
rect 48363 6613 48375 6647
rect 48498 6644 48504 6656
rect 48411 6616 48504 6644
rect 48317 6607 48375 6613
rect 48498 6604 48504 6616
rect 48556 6644 48562 6656
rect 52196 6644 52224 6684
rect 72050 6672 72056 6684
rect 72108 6672 72114 6724
rect 79965 6715 80023 6721
rect 79965 6681 79977 6715
rect 80011 6712 80023 6715
rect 80977 6715 81035 6721
rect 80977 6712 80989 6715
rect 80011 6684 80989 6712
rect 80011 6681 80023 6684
rect 79965 6675 80023 6681
rect 80977 6681 80989 6684
rect 81023 6681 81035 6715
rect 89916 6712 89944 6743
rect 91370 6740 91376 6792
rect 91428 6780 91434 6792
rect 95712 6780 95740 6820
rect 101493 6817 101505 6820
rect 101539 6817 101551 6851
rect 101493 6811 101551 6817
rect 101692 6780 101720 6888
rect 101876 6848 101904 6888
rect 102318 6876 102324 6928
rect 102376 6916 102382 6928
rect 102781 6919 102839 6925
rect 102781 6916 102793 6919
rect 102376 6888 102793 6916
rect 102376 6876 102382 6888
rect 102781 6885 102793 6888
rect 102827 6885 102839 6919
rect 103974 6916 103980 6928
rect 103935 6888 103980 6916
rect 102781 6879 102839 6885
rect 103974 6876 103980 6888
rect 104032 6876 104038 6928
rect 104066 6876 104072 6928
rect 104124 6916 104130 6928
rect 110874 6916 110880 6928
rect 104124 6888 110880 6916
rect 104124 6876 104130 6888
rect 110874 6876 110880 6888
rect 110932 6876 110938 6928
rect 111812 6916 111840 6956
rect 113361 6953 113373 6987
rect 113407 6984 113419 6987
rect 113450 6984 113456 6996
rect 113407 6956 113456 6984
rect 113407 6953 113419 6956
rect 113361 6947 113419 6953
rect 113450 6944 113456 6956
rect 113508 6944 113514 6996
rect 113542 6944 113548 6996
rect 113600 6984 113606 6996
rect 118970 6984 118976 6996
rect 113600 6956 118280 6984
rect 118931 6956 118976 6984
rect 113600 6944 113606 6956
rect 114741 6919 114799 6925
rect 114741 6916 114753 6919
rect 111812 6888 114753 6916
rect 114741 6885 114753 6888
rect 114787 6885 114799 6919
rect 118252 6916 118280 6956
rect 118970 6944 118976 6956
rect 119028 6944 119034 6996
rect 120445 6987 120503 6993
rect 120445 6953 120457 6987
rect 120491 6984 120503 6987
rect 121362 6984 121368 6996
rect 120491 6956 121368 6984
rect 120491 6953 120503 6956
rect 120445 6947 120503 6953
rect 121362 6944 121368 6956
rect 121420 6944 121426 6996
rect 132218 6984 132224 6996
rect 132179 6956 132224 6984
rect 132218 6944 132224 6956
rect 132276 6944 132282 6996
rect 155218 6984 155224 6996
rect 155179 6956 155224 6984
rect 155218 6944 155224 6956
rect 155276 6944 155282 6996
rect 163314 6984 163320 6996
rect 163275 6956 163320 6984
rect 163314 6944 163320 6956
rect 163372 6944 163378 6996
rect 128725 6919 128783 6925
rect 128725 6916 128737 6919
rect 118252 6888 128737 6916
rect 114741 6879 114799 6885
rect 128725 6885 128737 6888
rect 128771 6885 128783 6919
rect 128725 6879 128783 6885
rect 109494 6848 109500 6860
rect 101876 6820 109500 6848
rect 109494 6808 109500 6820
rect 109552 6808 109558 6860
rect 112165 6851 112223 6857
rect 112165 6817 112177 6851
rect 112211 6848 112223 6851
rect 112254 6848 112260 6860
rect 112211 6820 112260 6848
rect 112211 6817 112223 6820
rect 112165 6811 112223 6817
rect 112254 6808 112260 6820
rect 112312 6808 112318 6860
rect 113284 6820 114784 6848
rect 91428 6752 95740 6780
rect 95896 6752 101720 6780
rect 91428 6740 91434 6752
rect 90269 6715 90327 6721
rect 90269 6712 90281 6715
rect 89916 6684 90281 6712
rect 80977 6675 81035 6681
rect 90269 6681 90281 6684
rect 90315 6712 90327 6715
rect 95896 6712 95924 6752
rect 102134 6740 102140 6792
rect 102192 6780 102198 6792
rect 102321 6783 102379 6789
rect 102321 6780 102333 6783
rect 102192 6752 102333 6780
rect 102192 6740 102198 6752
rect 102321 6749 102333 6752
rect 102367 6749 102379 6783
rect 108666 6780 108672 6792
rect 102321 6743 102379 6749
rect 102428 6752 108672 6780
rect 90315 6684 95924 6712
rect 90315 6681 90327 6684
rect 90269 6675 90327 6681
rect 96246 6672 96252 6724
rect 96304 6712 96310 6724
rect 102428 6712 102456 6752
rect 108666 6740 108672 6752
rect 108724 6740 108730 6792
rect 113284 6780 113312 6820
rect 108776 6752 113312 6780
rect 113453 6783 113511 6789
rect 96304 6684 102456 6712
rect 96304 6672 96310 6684
rect 106366 6672 106372 6724
rect 106424 6712 106430 6724
rect 108776 6712 108804 6752
rect 113453 6749 113465 6783
rect 113499 6749 113511 6783
rect 114646 6780 114652 6792
rect 114607 6752 114652 6780
rect 113453 6743 113511 6749
rect 106424 6684 108804 6712
rect 106424 6672 106430 6684
rect 113468 6656 113496 6743
rect 114646 6740 114652 6752
rect 114704 6740 114710 6792
rect 114756 6780 114784 6820
rect 114830 6808 114836 6860
rect 114888 6848 114894 6860
rect 115385 6851 115443 6857
rect 115385 6848 115397 6851
rect 114888 6820 115397 6848
rect 114888 6808 114894 6820
rect 115385 6817 115397 6820
rect 115431 6848 115443 6851
rect 117774 6848 117780 6860
rect 115431 6820 117780 6848
rect 115431 6817 115443 6820
rect 115385 6811 115443 6817
rect 117774 6808 117780 6820
rect 117832 6808 117838 6860
rect 122837 6851 122895 6857
rect 122837 6817 122849 6851
rect 122883 6817 122895 6851
rect 125410 6848 125416 6860
rect 125371 6820 125416 6848
rect 122837 6811 122895 6817
rect 118602 6780 118608 6792
rect 114756 6752 118608 6780
rect 118602 6740 118608 6752
rect 118660 6740 118666 6792
rect 120077 6783 120135 6789
rect 120077 6749 120089 6783
rect 120123 6780 120135 6783
rect 120445 6783 120503 6789
rect 120445 6780 120457 6783
rect 120123 6752 120457 6780
rect 120123 6749 120135 6752
rect 120077 6743 120135 6749
rect 120445 6749 120457 6752
rect 120491 6749 120503 6783
rect 120445 6743 120503 6749
rect 121089 6783 121147 6789
rect 121089 6749 121101 6783
rect 121135 6780 121147 6783
rect 121822 6780 121828 6792
rect 121135 6752 121828 6780
rect 121135 6749 121147 6752
rect 121089 6743 121147 6749
rect 121822 6740 121828 6752
rect 121880 6740 121886 6792
rect 113634 6672 113640 6724
rect 113692 6712 113698 6724
rect 122852 6712 122880 6811
rect 125410 6808 125416 6820
rect 125468 6848 125474 6860
rect 125873 6851 125931 6857
rect 125873 6848 125885 6851
rect 125468 6820 125885 6848
rect 125468 6808 125474 6820
rect 125873 6817 125885 6820
rect 125919 6817 125931 6851
rect 127434 6848 127440 6860
rect 127395 6820 127440 6848
rect 125873 6811 125931 6817
rect 127434 6808 127440 6820
rect 127492 6808 127498 6860
rect 129826 6848 129832 6860
rect 129787 6820 129832 6848
rect 129826 6808 129832 6820
rect 129884 6808 129890 6860
rect 130841 6851 130899 6857
rect 130841 6817 130853 6851
rect 130887 6817 130899 6851
rect 132236 6848 132264 6944
rect 136174 6916 136180 6928
rect 136135 6888 136180 6916
rect 136174 6876 136180 6888
rect 136232 6876 136238 6928
rect 142890 6876 142896 6928
rect 142948 6916 142954 6928
rect 143077 6919 143135 6925
rect 143077 6916 143089 6919
rect 142948 6888 143089 6916
rect 142948 6876 142954 6888
rect 143077 6885 143089 6888
rect 143123 6885 143135 6919
rect 143077 6879 143135 6885
rect 153746 6876 153752 6928
rect 153804 6916 153810 6928
rect 154301 6919 154359 6925
rect 154301 6916 154313 6919
rect 153804 6888 154313 6916
rect 153804 6876 153810 6888
rect 154301 6885 154313 6888
rect 154347 6885 154359 6919
rect 162394 6916 162400 6928
rect 162355 6888 162400 6916
rect 154301 6879 154359 6885
rect 162394 6876 162400 6888
rect 162452 6876 162458 6928
rect 164789 6919 164847 6925
rect 164789 6885 164801 6919
rect 164835 6916 164847 6919
rect 164878 6916 164884 6928
rect 164835 6888 164884 6916
rect 164835 6885 164847 6888
rect 164789 6879 164847 6885
rect 164878 6876 164884 6888
rect 164936 6876 164942 6928
rect 133049 6851 133107 6857
rect 133049 6848 133061 6851
rect 132236 6820 133061 6848
rect 130841 6811 130899 6817
rect 133049 6817 133061 6820
rect 133095 6817 133107 6851
rect 141786 6848 141792 6860
rect 141747 6820 141792 6848
rect 133049 6811 133107 6817
rect 123389 6783 123447 6789
rect 123389 6749 123401 6783
rect 123435 6780 123447 6783
rect 123481 6783 123539 6789
rect 123481 6780 123493 6783
rect 123435 6752 123493 6780
rect 123435 6749 123447 6752
rect 123389 6743 123447 6749
rect 123481 6749 123493 6752
rect 123527 6749 123539 6783
rect 128538 6780 128544 6792
rect 128499 6752 128544 6780
rect 123481 6743 123539 6749
rect 128538 6740 128544 6752
rect 128596 6780 128602 6792
rect 129277 6783 129335 6789
rect 129277 6780 129289 6783
rect 128596 6752 129289 6780
rect 128596 6740 128602 6752
rect 129277 6749 129289 6752
rect 129323 6749 129335 6783
rect 129277 6743 129335 6749
rect 113692 6684 122880 6712
rect 113692 6672 113698 6684
rect 123018 6672 123024 6724
rect 123076 6712 123082 6724
rect 130856 6712 130884 6811
rect 141786 6808 141792 6820
rect 141844 6808 141850 6860
rect 146021 6851 146079 6857
rect 146021 6817 146033 6851
rect 146067 6848 146079 6851
rect 146938 6848 146944 6860
rect 146067 6820 146944 6848
rect 146067 6817 146079 6820
rect 146021 6811 146079 6817
rect 146938 6808 146944 6820
rect 146996 6808 147002 6860
rect 148042 6808 148048 6860
rect 148100 6848 148106 6860
rect 148137 6851 148195 6857
rect 148137 6848 148149 6851
rect 148100 6820 148149 6848
rect 148100 6808 148106 6820
rect 148137 6817 148149 6820
rect 148183 6848 148195 6851
rect 148597 6851 148655 6857
rect 148597 6848 148609 6851
rect 148183 6820 148609 6848
rect 148183 6817 148195 6820
rect 148137 6811 148195 6817
rect 148597 6817 148609 6820
rect 148643 6817 148655 6851
rect 151814 6848 151820 6860
rect 151775 6820 151820 6848
rect 148597 6811 148655 6817
rect 151814 6808 151820 6820
rect 151872 6808 151878 6860
rect 156138 6808 156144 6860
rect 156196 6848 156202 6860
rect 156509 6851 156567 6857
rect 156509 6848 156521 6851
rect 156196 6820 156521 6848
rect 156196 6808 156202 6820
rect 156509 6817 156521 6820
rect 156555 6817 156567 6851
rect 156509 6811 156567 6817
rect 159910 6808 159916 6860
rect 159968 6848 159974 6860
rect 160005 6851 160063 6857
rect 160005 6848 160017 6851
rect 159968 6820 160017 6848
rect 159968 6808 159974 6820
rect 160005 6817 160017 6820
rect 160051 6848 160063 6851
rect 160465 6851 160523 6857
rect 160465 6848 160477 6851
rect 160051 6820 160477 6848
rect 160051 6817 160063 6820
rect 160005 6811 160063 6817
rect 160465 6817 160477 6820
rect 160511 6817 160523 6851
rect 163498 6848 163504 6860
rect 163459 6820 163504 6848
rect 160465 6811 160523 6817
rect 163498 6808 163504 6820
rect 163556 6808 163562 6860
rect 131114 6780 131120 6792
rect 131075 6752 131120 6780
rect 131114 6740 131120 6752
rect 131172 6780 131178 6792
rect 131669 6783 131727 6789
rect 131669 6780 131681 6783
rect 131172 6752 131681 6780
rect 131172 6740 131178 6752
rect 131669 6749 131681 6752
rect 131715 6749 131727 6783
rect 134886 6780 134892 6792
rect 134847 6752 134892 6780
rect 131669 6743 131727 6749
rect 134886 6740 134892 6752
rect 134944 6740 134950 6792
rect 135990 6780 135996 6792
rect 135951 6752 135996 6780
rect 135990 6740 135996 6752
rect 136048 6780 136054 6792
rect 136729 6783 136787 6789
rect 136729 6780 136741 6783
rect 136048 6752 136741 6780
rect 136048 6740 136054 6752
rect 136729 6749 136741 6752
rect 136775 6749 136787 6783
rect 142890 6780 142896 6792
rect 142851 6752 142896 6780
rect 136729 6743 136787 6749
rect 142890 6740 142896 6752
rect 142948 6780 142954 6792
rect 143629 6783 143687 6789
rect 143629 6780 143641 6783
rect 142948 6752 143641 6780
rect 142948 6740 142954 6752
rect 143629 6749 143641 6752
rect 143675 6749 143687 6783
rect 143629 6743 143687 6749
rect 150529 6783 150587 6789
rect 150529 6749 150541 6783
rect 150575 6780 150587 6783
rect 150621 6783 150679 6789
rect 150621 6780 150633 6783
rect 150575 6752 150633 6780
rect 150575 6749 150587 6752
rect 150529 6743 150587 6749
rect 150621 6749 150633 6752
rect 150667 6780 150679 6783
rect 150802 6780 150808 6792
rect 150667 6752 150808 6780
rect 150667 6749 150679 6752
rect 150621 6743 150679 6749
rect 150802 6740 150808 6752
rect 150860 6740 150866 6792
rect 152090 6780 152096 6792
rect 152051 6752 152096 6780
rect 152090 6740 152096 6752
rect 152148 6780 152154 6792
rect 152461 6783 152519 6789
rect 152461 6780 152473 6783
rect 152148 6752 152473 6780
rect 152148 6740 152154 6752
rect 152461 6749 152473 6752
rect 152507 6749 152519 6783
rect 153010 6780 153016 6792
rect 152971 6752 153016 6780
rect 152461 6743 152519 6749
rect 153010 6740 153016 6752
rect 153068 6740 153074 6792
rect 153746 6740 153752 6792
rect 153804 6780 153810 6792
rect 154117 6783 154175 6789
rect 154117 6780 154129 6783
rect 153804 6752 154129 6780
rect 153804 6740 153810 6752
rect 154117 6749 154129 6752
rect 154163 6780 154175 6783
rect 154853 6783 154911 6789
rect 154853 6780 154865 6783
rect 154163 6752 154865 6780
rect 154163 6749 154175 6752
rect 154117 6743 154175 6749
rect 154853 6749 154865 6752
rect 154899 6749 154911 6783
rect 154853 6743 154911 6749
rect 160925 6783 160983 6789
rect 160925 6749 160937 6783
rect 160971 6780 160983 6783
rect 161109 6783 161167 6789
rect 161109 6780 161121 6783
rect 160971 6752 161121 6780
rect 160971 6749 160983 6752
rect 160925 6743 160983 6749
rect 161109 6749 161121 6752
rect 161155 6780 161167 6783
rect 161474 6780 161480 6792
rect 161155 6752 161480 6780
rect 161155 6749 161167 6752
rect 161109 6743 161167 6749
rect 161474 6740 161480 6752
rect 161532 6740 161538 6792
rect 162489 6783 162547 6789
rect 162489 6749 162501 6783
rect 162535 6749 162547 6783
rect 162489 6743 162547 6749
rect 123076 6684 130884 6712
rect 123076 6672 123082 6684
rect 162394 6672 162400 6724
rect 162452 6712 162458 6724
rect 162504 6712 162532 6743
rect 164234 6740 164240 6792
rect 164292 6780 164298 6792
rect 164605 6783 164663 6789
rect 164605 6780 164617 6783
rect 164292 6752 164617 6780
rect 164292 6740 164298 6752
rect 164605 6749 164617 6752
rect 164651 6780 164663 6783
rect 165709 6783 165767 6789
rect 165709 6780 165721 6783
rect 164651 6752 165721 6780
rect 164651 6749 164663 6752
rect 164605 6743 164663 6749
rect 165709 6749 165721 6752
rect 165755 6749 165767 6783
rect 165709 6743 165767 6749
rect 162949 6715 163007 6721
rect 162949 6712 162961 6715
rect 162452 6684 162961 6712
rect 162452 6672 162458 6684
rect 162949 6681 162961 6684
rect 162995 6681 163007 6715
rect 162949 6675 163007 6681
rect 48556 6616 52224 6644
rect 48556 6604 48562 6616
rect 52362 6604 52368 6656
rect 52420 6644 52426 6656
rect 56318 6644 56324 6656
rect 52420 6616 56324 6644
rect 52420 6604 52426 6616
rect 56318 6604 56324 6616
rect 56376 6604 56382 6656
rect 56410 6604 56416 6656
rect 56468 6644 56474 6656
rect 56468 6616 56513 6644
rect 56468 6604 56474 6616
rect 56962 6604 56968 6656
rect 57020 6644 57026 6656
rect 59446 6644 59452 6656
rect 57020 6616 59452 6644
rect 57020 6604 57026 6616
rect 59446 6604 59452 6616
rect 59504 6604 59510 6656
rect 59814 6644 59820 6656
rect 59775 6616 59820 6644
rect 59814 6604 59820 6616
rect 59872 6604 59878 6656
rect 64506 6604 64512 6656
rect 64564 6644 64570 6656
rect 65061 6647 65119 6653
rect 65061 6644 65073 6647
rect 64564 6616 65073 6644
rect 64564 6604 64570 6616
rect 65061 6613 65073 6616
rect 65107 6613 65119 6647
rect 65061 6607 65119 6613
rect 69569 6647 69627 6653
rect 69569 6613 69581 6647
rect 69615 6644 69627 6647
rect 69934 6644 69940 6656
rect 69615 6616 69940 6644
rect 69615 6613 69627 6616
rect 69569 6607 69627 6613
rect 69934 6604 69940 6616
rect 69992 6604 69998 6656
rect 70118 6604 70124 6656
rect 70176 6644 70182 6656
rect 79134 6644 79140 6656
rect 70176 6616 79140 6644
rect 70176 6604 70182 6616
rect 79134 6604 79140 6616
rect 79192 6604 79198 6656
rect 81161 6647 81219 6653
rect 81161 6613 81173 6647
rect 81207 6644 81219 6647
rect 81342 6644 81348 6656
rect 81207 6616 81348 6644
rect 81207 6613 81219 6616
rect 81161 6607 81219 6613
rect 81342 6604 81348 6616
rect 81400 6644 81406 6656
rect 81986 6644 81992 6656
rect 81400 6616 81992 6644
rect 81400 6604 81406 6616
rect 81986 6604 81992 6616
rect 82044 6604 82050 6656
rect 88518 6604 88524 6656
rect 88576 6644 88582 6656
rect 100570 6644 100576 6656
rect 88576 6616 100576 6644
rect 88576 6604 88582 6616
rect 100570 6604 100576 6616
rect 100628 6604 100634 6656
rect 103054 6604 103060 6656
rect 103112 6644 103118 6656
rect 108942 6644 108948 6656
rect 103112 6616 108948 6644
rect 103112 6604 103118 6616
rect 108942 6604 108948 6616
rect 109000 6604 109006 6656
rect 112993 6647 113051 6653
rect 112993 6613 113005 6647
rect 113039 6644 113051 6647
rect 113450 6644 113456 6656
rect 113039 6616 113456 6644
rect 113039 6613 113051 6616
rect 112993 6607 113051 6613
rect 113450 6604 113456 6616
rect 113508 6604 113514 6656
rect 115750 6644 115756 6656
rect 115711 6616 115756 6644
rect 115750 6604 115756 6616
rect 115808 6604 115814 6656
rect 117130 6644 117136 6656
rect 117091 6616 117136 6644
rect 117130 6604 117136 6616
rect 117188 6604 117194 6656
rect 120626 6644 120632 6656
rect 120587 6616 120632 6644
rect 120626 6604 120632 6616
rect 120684 6604 120690 6656
rect 123481 6647 123539 6653
rect 123481 6613 123493 6647
rect 123527 6644 123539 6647
rect 123757 6647 123815 6653
rect 123757 6644 123769 6647
rect 123527 6616 123769 6644
rect 123527 6613 123539 6616
rect 123481 6607 123539 6613
rect 123757 6613 123769 6616
rect 123803 6644 123815 6647
rect 124214 6644 124220 6656
rect 123803 6616 124220 6644
rect 123803 6613 123815 6616
rect 123757 6607 123815 6613
rect 124214 6604 124220 6616
rect 124272 6604 124278 6656
rect 126793 6647 126851 6653
rect 126793 6613 126805 6647
rect 126839 6644 126851 6647
rect 126974 6644 126980 6656
rect 126839 6616 126980 6644
rect 126839 6613 126851 6616
rect 126793 6607 126851 6613
rect 126974 6604 126980 6616
rect 127032 6604 127038 6656
rect 133230 6604 133236 6656
rect 133288 6644 133294 6656
rect 133509 6647 133567 6653
rect 133509 6644 133521 6647
rect 133288 6616 133521 6644
rect 133288 6604 133294 6616
rect 133509 6613 133521 6616
rect 133555 6613 133567 6647
rect 133509 6607 133567 6613
rect 144362 6604 144368 6656
rect 144420 6644 144426 6656
rect 144549 6647 144607 6653
rect 144549 6644 144561 6647
rect 144420 6616 144561 6644
rect 144420 6604 144426 6616
rect 144549 6613 144561 6616
rect 144595 6644 144607 6647
rect 145190 6644 145196 6656
rect 144595 6616 145196 6644
rect 144595 6613 144607 6616
rect 144549 6607 144607 6613
rect 145190 6604 145196 6616
rect 145248 6604 145254 6656
rect 149330 6644 149336 6656
rect 149291 6616 149336 6644
rect 149330 6604 149336 6616
rect 149388 6604 149394 6656
rect 155494 6644 155500 6656
rect 155455 6616 155500 6644
rect 155494 6604 155500 6616
rect 155552 6604 155558 6656
rect 155862 6604 155868 6656
rect 155920 6644 155926 6656
rect 155957 6647 156015 6653
rect 155957 6644 155969 6647
rect 155920 6616 155969 6644
rect 155920 6604 155926 6616
rect 155957 6613 155969 6616
rect 156003 6613 156015 6647
rect 155957 6607 156015 6613
rect 164510 6604 164516 6656
rect 164568 6644 164574 6656
rect 164970 6644 164976 6656
rect 164568 6616 164976 6644
rect 164568 6604 164574 6616
rect 164970 6604 164976 6616
rect 165028 6644 165034 6656
rect 165341 6647 165399 6653
rect 165341 6644 165353 6647
rect 165028 6616 165353 6644
rect 165028 6604 165034 6616
rect 165341 6613 165353 6616
rect 165387 6613 165399 6647
rect 165341 6607 165399 6613
rect 368 6554 93012 6576
rect 368 6502 56667 6554
rect 56719 6502 56731 6554
rect 56783 6502 56795 6554
rect 56847 6502 56859 6554
rect 56911 6502 93012 6554
rect 368 6480 93012 6502
rect 102028 6554 169556 6576
rect 102028 6502 113088 6554
rect 113140 6502 113152 6554
rect 113204 6502 113216 6554
rect 113268 6502 113280 6554
rect 113332 6502 169556 6554
rect 102028 6480 169556 6502
rect 4246 6440 4252 6452
rect 4207 6412 4252 6440
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 21821 6443 21879 6449
rect 21821 6409 21833 6443
rect 21867 6440 21879 6443
rect 21910 6440 21916 6452
rect 21867 6412 21916 6440
rect 21867 6409 21879 6412
rect 21821 6403 21879 6409
rect 21910 6400 21916 6412
rect 21968 6400 21974 6452
rect 23676 6412 31064 6440
rect 3694 6332 3700 6384
rect 3752 6372 3758 6384
rect 8202 6372 8208 6384
rect 3752 6344 8208 6372
rect 3752 6332 3758 6344
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 10686 6332 10692 6384
rect 10744 6372 10750 6384
rect 23676 6372 23704 6412
rect 10744 6344 23704 6372
rect 23768 6344 27752 6372
rect 10744 6332 10750 6344
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6304 9091 6307
rect 9214 6304 9220 6316
rect 9079 6276 9220 6304
rect 9079 6273 9091 6276
rect 9033 6267 9091 6273
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 21082 6304 21088 6316
rect 15160 6276 20576 6304
rect 21043 6276 21088 6304
rect 15160 6264 15166 6276
rect 3234 6236 3240 6248
rect 3195 6208 3240 6236
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 5905 6239 5963 6245
rect 5905 6236 5917 6239
rect 5868 6208 5917 6236
rect 5868 6196 5874 6208
rect 5905 6205 5917 6208
rect 5951 6236 5963 6239
rect 6089 6239 6147 6245
rect 6089 6236 6101 6239
rect 5951 6208 6101 6236
rect 5951 6205 5963 6208
rect 5905 6199 5963 6205
rect 6089 6205 6101 6208
rect 6135 6205 6147 6239
rect 6089 6199 6147 6205
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6236 7527 6239
rect 8018 6236 8024 6248
rect 7515 6208 8024 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8570 6236 8576 6248
rect 8531 6208 8576 6236
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6236 9919 6239
rect 10410 6236 10416 6248
rect 9907 6208 10416 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 15930 6196 15936 6248
rect 15988 6236 15994 6248
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15988 6208 16037 6236
rect 15988 6196 15994 6208
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 19518 6236 19524 6248
rect 19479 6208 19524 6236
rect 16025 6199 16083 6205
rect 19518 6196 19524 6208
rect 19576 6196 19582 6248
rect 20548 6245 20576 6276
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 22002 6264 22008 6316
rect 22060 6304 22066 6316
rect 23768 6304 23796 6344
rect 22060 6276 23796 6304
rect 24029 6307 24087 6313
rect 22060 6264 22066 6276
rect 24029 6273 24041 6307
rect 24075 6304 24087 6307
rect 24946 6304 24952 6316
rect 24075 6276 24952 6304
rect 24075 6273 24087 6276
rect 24029 6267 24087 6273
rect 24946 6264 24952 6276
rect 25004 6264 25010 6316
rect 26053 6307 26111 6313
rect 26053 6273 26065 6307
rect 26099 6273 26111 6307
rect 26053 6267 26111 6273
rect 26145 6307 26203 6313
rect 26145 6273 26157 6307
rect 26191 6304 26203 6307
rect 26234 6304 26240 6316
rect 26191 6276 26240 6304
rect 26191 6273 26203 6276
rect 26145 6267 26203 6273
rect 20533 6239 20591 6245
rect 20533 6205 20545 6239
rect 20579 6205 20591 6239
rect 20533 6199 20591 6205
rect 22646 6196 22652 6248
rect 22704 6236 22710 6248
rect 23385 6239 23443 6245
rect 23385 6236 23397 6239
rect 22704 6208 23397 6236
rect 22704 6196 22710 6208
rect 23385 6205 23397 6208
rect 23431 6205 23443 6239
rect 23385 6199 23443 6205
rect 25590 6196 25596 6248
rect 25648 6236 25654 6248
rect 26068 6236 26096 6267
rect 26234 6264 26240 6276
rect 26292 6264 26298 6316
rect 26510 6304 26516 6316
rect 26471 6276 26516 6304
rect 26510 6264 26516 6276
rect 26568 6264 26574 6316
rect 27341 6239 27399 6245
rect 27341 6236 27353 6239
rect 25648 6208 27353 6236
rect 25648 6196 25654 6208
rect 27341 6205 27353 6208
rect 27387 6205 27399 6239
rect 27724 6236 27752 6344
rect 27798 6332 27804 6384
rect 27856 6372 27862 6384
rect 31036 6372 31064 6412
rect 31110 6400 31116 6452
rect 31168 6440 31174 6452
rect 36170 6440 36176 6452
rect 31168 6412 36176 6440
rect 31168 6400 31174 6412
rect 36170 6400 36176 6412
rect 36228 6400 36234 6452
rect 36262 6400 36268 6452
rect 36320 6440 36326 6452
rect 36541 6443 36599 6449
rect 36541 6440 36553 6443
rect 36320 6412 36553 6440
rect 36320 6400 36326 6412
rect 36541 6409 36553 6412
rect 36587 6409 36599 6443
rect 36541 6403 36599 6409
rect 36630 6400 36636 6452
rect 36688 6440 36694 6452
rect 39574 6440 39580 6452
rect 36688 6412 39580 6440
rect 36688 6400 36694 6412
rect 39574 6400 39580 6412
rect 39632 6400 39638 6452
rect 39758 6440 39764 6452
rect 39719 6412 39764 6440
rect 39758 6400 39764 6412
rect 39816 6400 39822 6452
rect 39850 6400 39856 6452
rect 39908 6440 39914 6452
rect 40862 6440 40868 6452
rect 39908 6412 40868 6440
rect 39908 6400 39914 6412
rect 40862 6400 40868 6412
rect 40920 6400 40926 6452
rect 41138 6400 41144 6452
rect 41196 6440 41202 6452
rect 43530 6440 43536 6452
rect 41196 6412 43536 6440
rect 41196 6400 41202 6412
rect 43530 6400 43536 6412
rect 43588 6400 43594 6452
rect 43714 6400 43720 6452
rect 43772 6440 43778 6452
rect 47670 6440 47676 6452
rect 43772 6412 47676 6440
rect 43772 6400 43778 6412
rect 47670 6400 47676 6412
rect 47728 6400 47734 6452
rect 47762 6400 47768 6452
rect 47820 6440 47826 6452
rect 50706 6440 50712 6452
rect 47820 6412 50712 6440
rect 47820 6400 47826 6412
rect 50706 6400 50712 6412
rect 50764 6400 50770 6452
rect 50798 6400 50804 6452
rect 50856 6440 50862 6452
rect 51258 6440 51264 6452
rect 50856 6412 51264 6440
rect 50856 6400 50862 6412
rect 51258 6400 51264 6412
rect 51316 6400 51322 6452
rect 51442 6400 51448 6452
rect 51500 6440 51506 6452
rect 52362 6440 52368 6452
rect 51500 6412 52368 6440
rect 51500 6400 51506 6412
rect 52362 6400 52368 6412
rect 52420 6400 52426 6452
rect 52730 6400 52736 6452
rect 52788 6440 52794 6452
rect 53929 6443 53987 6449
rect 53929 6440 53941 6443
rect 52788 6412 53941 6440
rect 52788 6400 52794 6412
rect 53929 6409 53941 6412
rect 53975 6409 53987 6443
rect 53929 6403 53987 6409
rect 54018 6400 54024 6452
rect 54076 6440 54082 6452
rect 56597 6443 56655 6449
rect 56597 6440 56609 6443
rect 54076 6412 56609 6440
rect 54076 6400 54082 6412
rect 56597 6409 56609 6412
rect 56643 6409 56655 6443
rect 56597 6403 56655 6409
rect 56689 6443 56747 6449
rect 56689 6409 56701 6443
rect 56735 6440 56747 6443
rect 57606 6440 57612 6452
rect 56735 6412 57612 6440
rect 56735 6409 56747 6412
rect 56689 6403 56747 6409
rect 57606 6400 57612 6412
rect 57664 6400 57670 6452
rect 60093 6443 60151 6449
rect 60093 6409 60105 6443
rect 60139 6440 60151 6443
rect 60274 6440 60280 6452
rect 60139 6412 60280 6440
rect 60139 6409 60151 6412
rect 60093 6403 60151 6409
rect 60274 6400 60280 6412
rect 60332 6400 60338 6452
rect 81345 6443 81403 6449
rect 81345 6409 81357 6443
rect 81391 6440 81403 6443
rect 81894 6440 81900 6452
rect 81391 6412 81900 6440
rect 81391 6409 81403 6412
rect 81345 6403 81403 6409
rect 81894 6400 81900 6412
rect 81952 6400 81958 6452
rect 87782 6400 87788 6452
rect 87840 6440 87846 6452
rect 87969 6443 88027 6449
rect 87969 6440 87981 6443
rect 87840 6412 87981 6440
rect 87840 6400 87846 6412
rect 87969 6409 87981 6412
rect 88015 6409 88027 6443
rect 87969 6403 88027 6409
rect 89530 6400 89536 6452
rect 89588 6440 89594 6452
rect 95053 6443 95111 6449
rect 95053 6440 95065 6443
rect 89588 6412 95065 6440
rect 89588 6400 89594 6412
rect 95053 6409 95065 6412
rect 95099 6409 95111 6443
rect 95053 6403 95111 6409
rect 97994 6400 98000 6452
rect 98052 6440 98058 6452
rect 104434 6440 104440 6452
rect 98052 6412 104440 6440
rect 98052 6400 98058 6412
rect 104434 6400 104440 6412
rect 104492 6400 104498 6452
rect 104710 6400 104716 6452
rect 104768 6440 104774 6452
rect 104768 6412 159404 6440
rect 104768 6400 104774 6412
rect 27856 6344 30972 6372
rect 31036 6344 37412 6372
rect 27856 6332 27862 6344
rect 29822 6304 29828 6316
rect 29783 6276 29828 6304
rect 29822 6264 29828 6276
rect 29880 6264 29886 6316
rect 30285 6307 30343 6313
rect 30285 6273 30297 6307
rect 30331 6304 30343 6307
rect 30374 6304 30380 6316
rect 30331 6276 30380 6304
rect 30331 6273 30343 6276
rect 30285 6267 30343 6273
rect 30374 6264 30380 6276
rect 30432 6304 30438 6316
rect 30834 6304 30840 6316
rect 30432 6276 30840 6304
rect 30432 6264 30438 6276
rect 30834 6264 30840 6276
rect 30892 6264 30898 6316
rect 30944 6304 30972 6344
rect 34698 6304 34704 6316
rect 30944 6276 34704 6304
rect 34698 6264 34704 6276
rect 34756 6264 34762 6316
rect 35066 6264 35072 6316
rect 35124 6304 35130 6316
rect 35713 6307 35771 6313
rect 35124 6276 35296 6304
rect 35124 6264 35130 6276
rect 31110 6236 31116 6248
rect 27724 6208 31116 6236
rect 27341 6199 27399 6205
rect 31110 6196 31116 6208
rect 31168 6196 31174 6248
rect 33686 6196 33692 6248
rect 33744 6236 33750 6248
rect 34149 6239 34207 6245
rect 34149 6236 34161 6239
rect 33744 6208 34161 6236
rect 33744 6196 33750 6208
rect 34149 6205 34161 6208
rect 34195 6205 34207 6239
rect 34149 6199 34207 6205
rect 35161 6239 35219 6245
rect 35161 6205 35173 6239
rect 35207 6205 35219 6239
rect 35268 6236 35296 6276
rect 35713 6273 35725 6307
rect 35759 6304 35771 6307
rect 35986 6304 35992 6316
rect 35759 6276 35992 6304
rect 35759 6273 35771 6276
rect 35713 6267 35771 6273
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 36078 6264 36084 6316
rect 36136 6304 36142 6316
rect 37274 6304 37280 6316
rect 36136 6276 37280 6304
rect 36136 6264 36142 6276
rect 37274 6264 37280 6276
rect 37332 6264 37338 6316
rect 37384 6304 37412 6344
rect 37458 6332 37464 6384
rect 37516 6372 37522 6384
rect 37553 6375 37611 6381
rect 37553 6372 37565 6375
rect 37516 6344 37565 6372
rect 37516 6332 37522 6344
rect 37553 6341 37565 6344
rect 37599 6341 37611 6375
rect 41322 6372 41328 6384
rect 37553 6335 37611 6341
rect 37660 6344 41328 6372
rect 37660 6304 37688 6344
rect 41322 6332 41328 6344
rect 41380 6332 41386 6384
rect 41414 6332 41420 6384
rect 41472 6372 41478 6384
rect 42978 6372 42984 6384
rect 41472 6344 42984 6372
rect 41472 6332 41478 6344
rect 42978 6332 42984 6344
rect 43036 6332 43042 6384
rect 43162 6332 43168 6384
rect 43220 6332 43226 6384
rect 43438 6372 43444 6384
rect 43272 6344 43444 6372
rect 37384 6276 37688 6304
rect 37826 6264 37832 6316
rect 37884 6304 37890 6316
rect 38930 6304 38936 6316
rect 37884 6276 38936 6304
rect 37884 6264 37890 6276
rect 38930 6264 38936 6276
rect 38988 6264 38994 6316
rect 41138 6304 41144 6316
rect 39408 6276 41144 6304
rect 39408 6236 39436 6276
rect 41138 6264 41144 6276
rect 41196 6264 41202 6316
rect 41598 6304 41604 6316
rect 41248 6276 41604 6304
rect 35268 6208 39436 6236
rect 35161 6199 35219 6205
rect 4890 6128 4896 6180
rect 4948 6168 4954 6180
rect 4948 6140 29224 6168
rect 4948 6128 4954 6140
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 3697 6103 3755 6109
rect 3697 6100 3709 6103
rect 3476 6072 3709 6100
rect 3476 6060 3482 6072
rect 3697 6069 3709 6072
rect 3743 6069 3755 6103
rect 21358 6100 21364 6112
rect 21319 6072 21364 6100
rect 3697 6063 3755 6069
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 24302 6060 24308 6112
rect 24360 6100 24366 6112
rect 29086 6100 29092 6112
rect 24360 6072 29092 6100
rect 24360 6060 24366 6072
rect 29086 6060 29092 6072
rect 29144 6060 29150 6112
rect 29196 6100 29224 6140
rect 29270 6128 29276 6180
rect 29328 6168 29334 6180
rect 35176 6168 35204 6199
rect 39482 6196 39488 6248
rect 39540 6236 39546 6248
rect 41248 6236 41276 6276
rect 41598 6264 41604 6276
rect 41656 6264 41662 6316
rect 41690 6264 41696 6316
rect 41748 6304 41754 6316
rect 41748 6276 41793 6304
rect 41748 6264 41754 6276
rect 41874 6264 41880 6316
rect 41932 6304 41938 6316
rect 42150 6304 42156 6316
rect 41932 6276 42156 6304
rect 41932 6264 41938 6276
rect 42150 6264 42156 6276
rect 42208 6264 42214 6316
rect 42794 6264 42800 6316
rect 42852 6304 42858 6316
rect 43180 6304 43208 6332
rect 43272 6313 43300 6344
rect 43438 6332 43444 6344
rect 43496 6372 43502 6384
rect 52270 6372 52276 6384
rect 43496 6344 52276 6372
rect 43496 6332 43502 6344
rect 52270 6332 52276 6344
rect 52328 6332 52334 6384
rect 54662 6372 54668 6384
rect 52656 6344 54668 6372
rect 52656 6316 52684 6344
rect 54662 6332 54668 6344
rect 54720 6332 54726 6384
rect 55490 6372 55496 6384
rect 55451 6344 55496 6372
rect 55490 6332 55496 6344
rect 55548 6332 55554 6384
rect 58526 6372 58532 6384
rect 55600 6344 58532 6372
rect 42852 6276 43208 6304
rect 43257 6307 43315 6313
rect 42852 6264 42858 6276
rect 43257 6273 43269 6307
rect 43303 6273 43315 6307
rect 47210 6304 47216 6316
rect 43257 6267 43315 6273
rect 43364 6276 46704 6304
rect 47171 6276 47216 6304
rect 39540 6208 41276 6236
rect 39540 6196 39546 6208
rect 41322 6196 41328 6248
rect 41380 6236 41386 6248
rect 42705 6239 42763 6245
rect 42705 6236 42717 6239
rect 41380 6208 42717 6236
rect 41380 6196 41386 6208
rect 42705 6205 42717 6208
rect 42751 6205 42763 6239
rect 43364 6236 43392 6276
rect 42705 6199 42763 6205
rect 43272 6208 43392 6236
rect 43272 6168 43300 6208
rect 43530 6196 43536 6248
rect 43588 6236 43594 6248
rect 45462 6236 45468 6248
rect 43588 6208 45468 6236
rect 43588 6196 43594 6208
rect 45462 6196 45468 6208
rect 45520 6196 45526 6248
rect 45646 6236 45652 6248
rect 45559 6208 45652 6236
rect 45646 6196 45652 6208
rect 45704 6236 45710 6248
rect 45830 6236 45836 6248
rect 45704 6208 45836 6236
rect 45704 6196 45710 6208
rect 45830 6196 45836 6208
rect 45888 6196 45894 6248
rect 45922 6196 45928 6248
rect 45980 6236 45986 6248
rect 46474 6236 46480 6248
rect 45980 6208 46480 6236
rect 45980 6196 45986 6208
rect 46474 6196 46480 6208
rect 46532 6196 46538 6248
rect 46676 6245 46704 6276
rect 47210 6264 47216 6276
rect 47268 6264 47274 6316
rect 47302 6264 47308 6316
rect 47360 6304 47366 6316
rect 50154 6304 50160 6316
rect 47360 6276 50160 6304
rect 47360 6264 47366 6276
rect 50154 6264 50160 6276
rect 50212 6264 50218 6316
rect 50706 6264 50712 6316
rect 50764 6304 50770 6316
rect 50764 6276 50936 6304
rect 50764 6264 50770 6276
rect 46661 6239 46719 6245
rect 46661 6205 46673 6239
rect 46707 6205 46719 6239
rect 46661 6199 46719 6205
rect 46842 6196 46848 6248
rect 46900 6236 46906 6248
rect 50908 6236 50936 6276
rect 51166 6264 51172 6316
rect 51224 6304 51230 6316
rect 51261 6307 51319 6313
rect 51261 6304 51273 6307
rect 51224 6276 51273 6304
rect 51224 6264 51230 6276
rect 51261 6273 51273 6276
rect 51307 6273 51319 6307
rect 51261 6267 51319 6273
rect 51626 6264 51632 6316
rect 51684 6304 51690 6316
rect 52454 6304 52460 6316
rect 51684 6276 52460 6304
rect 51684 6264 51690 6276
rect 52454 6264 52460 6276
rect 52512 6264 52518 6316
rect 52638 6304 52644 6316
rect 52551 6276 52644 6304
rect 52638 6264 52644 6276
rect 52696 6264 52702 6316
rect 55600 6304 55628 6344
rect 58526 6332 58532 6344
rect 58584 6332 58590 6384
rect 58636 6344 59400 6372
rect 53116 6276 55628 6304
rect 46900 6208 50844 6236
rect 50908 6208 51580 6236
rect 46900 6196 46906 6208
rect 29328 6140 35204 6168
rect 35912 6140 43300 6168
rect 29328 6128 29334 6140
rect 35912 6100 35940 6140
rect 43346 6128 43352 6180
rect 43404 6168 43410 6180
rect 48038 6168 48044 6180
rect 43404 6140 48044 6168
rect 43404 6128 43410 6140
rect 48038 6128 48044 6140
rect 48096 6128 48102 6180
rect 48130 6128 48136 6180
rect 48188 6168 48194 6180
rect 50706 6168 50712 6180
rect 48188 6140 50712 6168
rect 48188 6128 48194 6140
rect 50706 6128 50712 6140
rect 50764 6128 50770 6180
rect 50816 6168 50844 6208
rect 51442 6168 51448 6180
rect 50816 6140 51448 6168
rect 51442 6128 51448 6140
rect 51500 6128 51506 6180
rect 51552 6168 51580 6208
rect 51902 6196 51908 6248
rect 51960 6236 51966 6248
rect 52273 6239 52331 6245
rect 52273 6236 52285 6239
rect 51960 6208 52285 6236
rect 51960 6196 51966 6208
rect 52273 6205 52285 6208
rect 52319 6205 52331 6239
rect 52273 6199 52331 6205
rect 52362 6196 52368 6248
rect 52420 6236 52426 6248
rect 53116 6236 53144 6276
rect 56410 6264 56416 6316
rect 56468 6304 56474 6316
rect 57422 6304 57428 6316
rect 56468 6276 57428 6304
rect 56468 6264 56474 6276
rect 57422 6264 57428 6276
rect 57480 6304 57486 6316
rect 57701 6307 57759 6313
rect 57701 6304 57713 6307
rect 57480 6276 57713 6304
rect 57480 6264 57486 6276
rect 57701 6273 57713 6276
rect 57747 6273 57759 6307
rect 57701 6267 57759 6273
rect 52420 6208 53144 6236
rect 52420 6196 52426 6208
rect 55030 6196 55036 6248
rect 55088 6236 55094 6248
rect 58636 6236 58664 6344
rect 59262 6304 59268 6316
rect 59223 6276 59268 6304
rect 59262 6264 59268 6276
rect 59320 6264 59326 6316
rect 59372 6304 59400 6344
rect 59446 6332 59452 6384
rect 59504 6372 59510 6384
rect 89990 6372 89996 6384
rect 59504 6344 89996 6372
rect 59504 6332 59510 6344
rect 89990 6332 89996 6344
rect 90048 6332 90054 6384
rect 92014 6332 92020 6384
rect 92072 6372 92078 6384
rect 104342 6372 104348 6384
rect 92072 6344 104348 6372
rect 92072 6332 92078 6344
rect 104342 6332 104348 6344
rect 104400 6332 104406 6384
rect 104618 6332 104624 6384
rect 104676 6372 104682 6384
rect 106274 6372 106280 6384
rect 104676 6344 106280 6372
rect 104676 6332 104682 6344
rect 106274 6332 106280 6344
rect 106332 6332 106338 6384
rect 130010 6372 130016 6384
rect 108224 6344 130016 6372
rect 63862 6304 63868 6316
rect 59372 6276 63868 6304
rect 63862 6264 63868 6276
rect 63920 6264 63926 6316
rect 64506 6304 64512 6316
rect 64467 6276 64512 6304
rect 64506 6264 64512 6276
rect 64564 6264 64570 6316
rect 66070 6304 66076 6316
rect 66031 6276 66076 6304
rect 66070 6264 66076 6276
rect 66128 6264 66134 6316
rect 69934 6304 69940 6316
rect 69895 6276 69940 6304
rect 69934 6264 69940 6276
rect 69992 6264 69998 6316
rect 71501 6307 71559 6313
rect 71501 6273 71513 6307
rect 71547 6304 71559 6307
rect 71774 6304 71780 6316
rect 71547 6276 71780 6304
rect 71547 6273 71559 6276
rect 71501 6267 71559 6273
rect 71774 6264 71780 6276
rect 71832 6264 71838 6316
rect 91830 6304 91836 6316
rect 86420 6276 91508 6304
rect 91791 6276 91836 6304
rect 65518 6236 65524 6248
rect 55088 6208 58664 6236
rect 58912 6208 59400 6236
rect 65479 6208 65524 6236
rect 55088 6196 55094 6208
rect 55858 6168 55864 6180
rect 51552 6140 55864 6168
rect 55858 6128 55864 6140
rect 55916 6128 55922 6180
rect 56597 6171 56655 6177
rect 56597 6137 56609 6171
rect 56643 6168 56655 6171
rect 57606 6168 57612 6180
rect 56643 6140 57612 6168
rect 56643 6137 56655 6140
rect 56597 6131 56655 6137
rect 57606 6128 57612 6140
rect 57664 6128 57670 6180
rect 57790 6128 57796 6180
rect 57848 6168 57854 6180
rect 58912 6168 58940 6208
rect 57848 6140 58940 6168
rect 58989 6171 59047 6177
rect 57848 6128 57854 6140
rect 58989 6137 59001 6171
rect 59035 6137 59047 6171
rect 59372 6168 59400 6208
rect 65518 6196 65524 6208
rect 65576 6196 65582 6248
rect 70946 6236 70952 6248
rect 70907 6208 70952 6236
rect 70946 6196 70952 6208
rect 71004 6196 71010 6248
rect 81253 6239 81311 6245
rect 81253 6205 81265 6239
rect 81299 6236 81311 6239
rect 86420 6236 86448 6276
rect 81299 6208 86448 6236
rect 86497 6239 86555 6245
rect 81299 6205 81311 6208
rect 81253 6199 81311 6205
rect 86497 6205 86509 6239
rect 86543 6236 86555 6239
rect 87506 6236 87512 6248
rect 86543 6208 87512 6236
rect 86543 6205 86555 6208
rect 86497 6199 86555 6205
rect 87506 6196 87512 6208
rect 87564 6196 87570 6248
rect 88981 6239 89039 6245
rect 88981 6205 88993 6239
rect 89027 6236 89039 6239
rect 90266 6236 90272 6248
rect 89027 6208 90272 6236
rect 89027 6205 89039 6208
rect 88981 6199 89039 6205
rect 90266 6196 90272 6208
rect 90324 6196 90330 6248
rect 91186 6196 91192 6248
rect 91244 6236 91250 6248
rect 91281 6239 91339 6245
rect 91281 6236 91293 6239
rect 91244 6208 91293 6236
rect 91244 6196 91250 6208
rect 91281 6205 91293 6208
rect 91327 6205 91339 6239
rect 91480 6236 91508 6276
rect 91830 6264 91836 6276
rect 91888 6264 91894 6316
rect 97258 6264 97264 6316
rect 97316 6304 97322 6316
rect 97316 6276 107424 6304
rect 97316 6264 97322 6276
rect 91480 6208 95188 6236
rect 91281 6199 91339 6205
rect 75730 6168 75736 6180
rect 59372 6140 75736 6168
rect 58989 6131 59047 6137
rect 36078 6100 36084 6112
rect 29196 6072 35940 6100
rect 36039 6072 36084 6100
rect 36078 6060 36084 6072
rect 36136 6060 36142 6112
rect 36170 6060 36176 6112
rect 36228 6100 36234 6112
rect 51258 6100 51264 6112
rect 36228 6072 51264 6100
rect 36228 6060 36234 6072
rect 51258 6060 51264 6072
rect 51316 6060 51322 6112
rect 51350 6060 51356 6112
rect 51408 6100 51414 6112
rect 59004 6100 59032 6131
rect 75730 6128 75736 6140
rect 75788 6128 75794 6180
rect 95160 6168 95188 6208
rect 101674 6196 101680 6248
rect 101732 6236 101738 6248
rect 103330 6236 103336 6248
rect 101732 6208 103336 6236
rect 101732 6196 101738 6208
rect 103330 6196 103336 6208
rect 103388 6196 103394 6248
rect 104802 6196 104808 6248
rect 104860 6236 104866 6248
rect 106274 6236 106280 6248
rect 104860 6208 106280 6236
rect 104860 6196 104866 6208
rect 106274 6196 106280 6208
rect 106332 6196 106338 6248
rect 103514 6168 103520 6180
rect 95160 6140 103520 6168
rect 103514 6128 103520 6140
rect 103572 6128 103578 6180
rect 107396 6168 107424 6276
rect 107470 6196 107476 6248
rect 107528 6236 107534 6248
rect 108224 6236 108252 6344
rect 130010 6332 130016 6344
rect 130068 6332 130074 6384
rect 134886 6332 134892 6384
rect 134944 6372 134950 6384
rect 135809 6375 135867 6381
rect 135809 6372 135821 6375
rect 134944 6344 135821 6372
rect 134944 6332 134950 6344
rect 135809 6341 135821 6344
rect 135855 6341 135867 6375
rect 135809 6335 135867 6341
rect 141786 6332 141792 6384
rect 141844 6372 141850 6384
rect 142157 6375 142215 6381
rect 142157 6372 142169 6375
rect 141844 6344 142169 6372
rect 141844 6332 141850 6344
rect 142157 6341 142169 6344
rect 142203 6341 142215 6375
rect 142798 6372 142804 6384
rect 142759 6344 142804 6372
rect 142157 6335 142215 6341
rect 142798 6332 142804 6344
rect 142856 6372 142862 6384
rect 143169 6375 143227 6381
rect 143169 6372 143181 6375
rect 142856 6344 143181 6372
rect 142856 6332 142862 6344
rect 143169 6341 143181 6344
rect 143215 6341 143227 6375
rect 150802 6372 150808 6384
rect 150763 6344 150808 6372
rect 143169 6335 143227 6341
rect 150802 6332 150808 6344
rect 150860 6332 150866 6384
rect 153010 6332 153016 6384
rect 153068 6372 153074 6384
rect 155773 6375 155831 6381
rect 155773 6372 155785 6375
rect 153068 6344 155785 6372
rect 153068 6332 153074 6344
rect 155773 6341 155785 6344
rect 155819 6341 155831 6375
rect 155773 6335 155831 6341
rect 156785 6375 156843 6381
rect 156785 6341 156797 6375
rect 156831 6372 156843 6375
rect 157242 6372 157248 6384
rect 156831 6344 157248 6372
rect 156831 6341 156843 6344
rect 156785 6335 156843 6341
rect 157242 6332 157248 6344
rect 157300 6332 157306 6384
rect 159376 6372 159404 6412
rect 159450 6400 159456 6452
rect 159508 6440 159514 6452
rect 159729 6443 159787 6449
rect 159729 6440 159741 6443
rect 159508 6412 159741 6440
rect 159508 6400 159514 6412
rect 159729 6409 159741 6412
rect 159775 6409 159787 6443
rect 161474 6440 161480 6452
rect 161435 6412 161480 6440
rect 159729 6403 159787 6409
rect 161474 6400 161480 6412
rect 161532 6400 161538 6452
rect 162489 6443 162547 6449
rect 162489 6409 162501 6443
rect 162535 6440 162547 6443
rect 163498 6440 163504 6452
rect 162535 6412 163504 6440
rect 162535 6409 162547 6412
rect 162489 6403 162547 6409
rect 163498 6400 163504 6412
rect 163556 6400 163562 6452
rect 164786 6372 164792 6384
rect 159376 6344 164792 6372
rect 164786 6332 164792 6344
rect 164844 6332 164850 6384
rect 122469 6307 122527 6313
rect 113284 6276 121960 6304
rect 107528 6208 108252 6236
rect 107528 6196 107534 6208
rect 108298 6196 108304 6248
rect 108356 6236 108362 6248
rect 113284 6236 113312 6276
rect 108356 6208 113312 6236
rect 113361 6239 113419 6245
rect 108356 6196 108362 6208
rect 113361 6205 113373 6239
rect 113407 6236 113419 6239
rect 113450 6236 113456 6248
rect 113407 6208 113456 6236
rect 113407 6205 113419 6208
rect 113361 6199 113419 6205
rect 113450 6196 113456 6208
rect 113508 6196 113514 6248
rect 115201 6239 115259 6245
rect 115201 6205 115213 6239
rect 115247 6236 115259 6239
rect 115750 6236 115756 6248
rect 115247 6208 115756 6236
rect 115247 6205 115259 6208
rect 115201 6199 115259 6205
rect 115750 6196 115756 6208
rect 115808 6196 115814 6248
rect 120905 6239 120963 6245
rect 120905 6205 120917 6239
rect 120951 6236 120963 6239
rect 121454 6236 121460 6248
rect 120951 6208 121460 6236
rect 120951 6205 120963 6208
rect 120905 6199 120963 6205
rect 121454 6196 121460 6208
rect 121512 6196 121518 6248
rect 121932 6245 121960 6276
rect 122469 6273 122481 6307
rect 122515 6304 122527 6307
rect 123018 6304 123024 6316
rect 122515 6276 123024 6304
rect 122515 6273 122527 6276
rect 122469 6267 122527 6273
rect 123018 6264 123024 6276
rect 123076 6264 123082 6316
rect 145742 6264 145748 6316
rect 145800 6304 145806 6316
rect 149977 6307 150035 6313
rect 145800 6276 149468 6304
rect 145800 6264 145806 6276
rect 121917 6239 121975 6245
rect 121917 6205 121929 6239
rect 121963 6205 121975 6239
rect 121917 6199 121975 6205
rect 122834 6196 122840 6248
rect 122892 6236 122898 6248
rect 122929 6239 122987 6245
rect 122929 6236 122941 6239
rect 122892 6208 122941 6236
rect 122892 6196 122898 6208
rect 122929 6205 122941 6208
rect 122975 6236 122987 6239
rect 123297 6239 123355 6245
rect 123297 6236 123309 6239
rect 122975 6208 123309 6236
rect 122975 6205 122987 6208
rect 122929 6199 122987 6205
rect 123297 6205 123309 6208
rect 123343 6205 123355 6239
rect 123297 6199 123355 6205
rect 128906 6196 128912 6248
rect 128964 6236 128970 6248
rect 129093 6239 129151 6245
rect 129093 6236 129105 6239
rect 128964 6208 129105 6236
rect 128964 6196 128970 6208
rect 129093 6205 129105 6208
rect 129139 6205 129151 6239
rect 148410 6236 148416 6248
rect 148371 6208 148416 6236
rect 129093 6199 129151 6205
rect 148410 6196 148416 6208
rect 148468 6196 148474 6248
rect 149440 6245 149468 6276
rect 149977 6273 149989 6307
rect 150023 6304 150035 6307
rect 150066 6304 150072 6316
rect 150023 6276 150072 6304
rect 150023 6273 150035 6276
rect 149977 6267 150035 6273
rect 150066 6264 150072 6276
rect 150124 6264 150130 6316
rect 153105 6307 153163 6313
rect 153105 6273 153117 6307
rect 153151 6304 153163 6307
rect 153470 6304 153476 6316
rect 153151 6276 153476 6304
rect 153151 6273 153163 6276
rect 153105 6267 153163 6273
rect 153470 6264 153476 6276
rect 153528 6264 153534 6316
rect 154850 6304 154856 6316
rect 154811 6276 154856 6304
rect 154850 6264 154856 6276
rect 154908 6264 154914 6316
rect 164970 6304 164976 6316
rect 164931 6276 164976 6304
rect 164970 6264 164976 6276
rect 165028 6264 165034 6316
rect 149425 6239 149483 6245
rect 149425 6205 149437 6239
rect 149471 6205 149483 6239
rect 153378 6236 153384 6248
rect 153291 6208 153384 6236
rect 149425 6199 149483 6205
rect 153378 6196 153384 6208
rect 153436 6236 153442 6248
rect 154574 6236 154580 6248
rect 153436 6208 154580 6236
rect 153436 6196 153442 6208
rect 154574 6196 154580 6208
rect 154632 6196 154638 6248
rect 158254 6236 158260 6248
rect 158215 6208 158260 6236
rect 158254 6196 158260 6208
rect 158312 6196 158318 6248
rect 163498 6196 163504 6248
rect 163556 6236 163562 6248
rect 163869 6239 163927 6245
rect 163869 6236 163881 6239
rect 163556 6208 163881 6236
rect 163556 6196 163562 6208
rect 163869 6205 163881 6208
rect 163915 6236 163927 6239
rect 166261 6239 166319 6245
rect 166261 6236 166273 6239
rect 163915 6208 166273 6236
rect 163915 6205 163927 6208
rect 163869 6199 163927 6205
rect 166261 6205 166273 6208
rect 166307 6205 166319 6239
rect 166261 6199 166319 6205
rect 114830 6168 114836 6180
rect 107396 6140 114836 6168
rect 114830 6128 114836 6140
rect 114888 6128 114894 6180
rect 148870 6168 148876 6180
rect 124140 6140 143488 6168
rect 124140 6112 124168 6140
rect 51408 6072 59032 6100
rect 51408 6060 51414 6072
rect 75822 6060 75828 6112
rect 75880 6100 75886 6112
rect 81253 6103 81311 6109
rect 81253 6100 81265 6103
rect 75880 6072 81265 6100
rect 75880 6060 75886 6072
rect 81253 6069 81265 6072
rect 81299 6069 81311 6103
rect 100938 6100 100944 6112
rect 81253 6063 81311 6069
rect 93044 6072 100944 6100
rect 368 6010 93012 6032
rect 368 5958 28456 6010
rect 28508 5958 28520 6010
rect 28572 5958 28584 6010
rect 28636 5958 28648 6010
rect 28700 5958 84878 6010
rect 84930 5958 84942 6010
rect 84994 5958 85006 6010
rect 85058 5958 85070 6010
rect 85122 5958 93012 6010
rect 368 5936 93012 5958
rect 9214 5896 9220 5908
rect 9175 5868 9220 5896
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 12342 5896 12348 5908
rect 12303 5868 12348 5896
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 15930 5896 15936 5908
rect 15891 5868 15936 5896
rect 15930 5856 15936 5868
rect 15988 5856 15994 5908
rect 19518 5896 19524 5908
rect 19076 5868 19524 5896
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 11885 5831 11943 5837
rect 3844 5800 8064 5828
rect 3844 5788 3850 5800
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 3418 5760 3424 5772
rect 2271 5732 3424 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4212 5732 4445 5760
rect 4212 5720 4218 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 5810 5760 5816 5772
rect 5771 5732 5816 5760
rect 4433 5723 4491 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 6914 5760 6920 5772
rect 6875 5732 6920 5760
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7742 5760 7748 5772
rect 7392 5732 7748 5760
rect 7392 5701 7420 5732
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 5000 5624 5028 5655
rect 5350 5624 5356 5636
rect 5000 5596 5356 5624
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 8036 5624 8064 5800
rect 11885 5797 11897 5831
rect 11931 5828 11943 5831
rect 14734 5828 14740 5840
rect 11931 5800 14740 5828
rect 11931 5797 11943 5800
rect 11885 5791 11943 5797
rect 14734 5788 14740 5800
rect 14792 5788 14798 5840
rect 10410 5760 10416 5772
rect 10371 5732 10416 5760
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 15948 5760 15976 5856
rect 19076 5769 19104 5868
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20901 5899 20959 5905
rect 20901 5865 20913 5899
rect 20947 5896 20959 5899
rect 21082 5896 21088 5908
rect 20947 5868 21088 5896
rect 20947 5865 20959 5868
rect 20901 5859 20959 5865
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 23385 5899 23443 5905
rect 23385 5865 23397 5899
rect 23431 5896 23443 5899
rect 24946 5896 24952 5908
rect 23431 5868 24952 5896
rect 23431 5865 23443 5868
rect 23385 5859 23443 5865
rect 24946 5856 24952 5868
rect 25004 5856 25010 5908
rect 25590 5896 25596 5908
rect 25551 5868 25596 5896
rect 25590 5856 25596 5868
rect 25648 5856 25654 5908
rect 26786 5856 26792 5908
rect 26844 5896 26850 5908
rect 28810 5896 28816 5908
rect 26844 5868 28816 5896
rect 26844 5856 26850 5868
rect 28810 5856 28816 5868
rect 28868 5856 28874 5908
rect 30285 5899 30343 5905
rect 30285 5865 30297 5899
rect 30331 5896 30343 5899
rect 30374 5896 30380 5908
rect 30331 5868 30380 5896
rect 30331 5865 30343 5868
rect 30285 5859 30343 5865
rect 30374 5856 30380 5868
rect 30432 5856 30438 5908
rect 31113 5899 31171 5905
rect 31113 5865 31125 5899
rect 31159 5896 31171 5899
rect 33413 5899 33471 5905
rect 31159 5868 32076 5896
rect 31159 5865 31171 5868
rect 31113 5859 31171 5865
rect 21174 5788 21180 5840
rect 21232 5828 21238 5840
rect 21232 5800 26096 5828
rect 21232 5788 21238 5800
rect 16025 5763 16083 5769
rect 16025 5760 16037 5763
rect 15948 5732 16037 5760
rect 16025 5729 16037 5732
rect 16071 5729 16083 5763
rect 16025 5723 16083 5729
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 19061 5763 19119 5769
rect 19061 5729 19073 5763
rect 19107 5729 19119 5763
rect 19061 5723 19119 5729
rect 21085 5763 21143 5769
rect 21085 5729 21097 5763
rect 21131 5760 21143 5763
rect 21358 5760 21364 5772
rect 21131 5732 21364 5760
rect 21131 5729 21143 5732
rect 21085 5723 21143 5729
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5692 12035 5695
rect 12342 5692 12348 5704
rect 12023 5664 12348 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 17052 5624 17080 5723
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 22097 5763 22155 5769
rect 22097 5729 22109 5763
rect 22143 5729 22155 5763
rect 22097 5723 22155 5729
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5692 17647 5695
rect 17957 5695 18015 5701
rect 17957 5692 17969 5695
rect 17635 5664 17969 5692
rect 17635 5661 17647 5664
rect 17589 5655 17647 5661
rect 17957 5661 17969 5664
rect 18003 5692 18015 5695
rect 22002 5692 22008 5704
rect 18003 5664 22008 5692
rect 18003 5661 18015 5664
rect 17957 5655 18015 5661
rect 22002 5652 22008 5664
rect 22060 5652 22066 5704
rect 8036 5596 17080 5624
rect 17126 5584 17132 5636
rect 17184 5624 17190 5636
rect 22112 5624 22140 5723
rect 22649 5695 22707 5701
rect 22649 5661 22661 5695
rect 22695 5692 22707 5695
rect 22741 5695 22799 5701
rect 22741 5692 22753 5695
rect 22695 5664 22753 5692
rect 22695 5661 22707 5664
rect 22649 5655 22707 5661
rect 22741 5661 22753 5664
rect 22787 5661 22799 5695
rect 24026 5692 24032 5704
rect 23987 5664 24032 5692
rect 22741 5655 22799 5661
rect 24026 5652 24032 5664
rect 24084 5692 24090 5704
rect 24489 5695 24547 5701
rect 24489 5692 24501 5695
rect 24084 5664 24501 5692
rect 24084 5652 24090 5664
rect 24489 5661 24501 5664
rect 24535 5661 24547 5695
rect 24489 5655 24547 5661
rect 23477 5627 23535 5633
rect 23477 5624 23489 5627
rect 17184 5596 22140 5624
rect 22664 5596 23489 5624
rect 17184 5584 17190 5596
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 5718 5556 5724 5568
rect 3752 5528 5724 5556
rect 3752 5516 3758 5528
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 8018 5556 8024 5568
rect 7979 5528 8024 5556
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 21174 5516 21180 5568
rect 21232 5556 21238 5568
rect 22664 5556 22692 5596
rect 23477 5593 23489 5596
rect 23523 5593 23535 5627
rect 23477 5587 23535 5593
rect 24854 5584 24860 5636
rect 24912 5624 24918 5636
rect 25777 5627 25835 5633
rect 25777 5624 25789 5627
rect 24912 5596 25789 5624
rect 24912 5584 24918 5596
rect 25777 5593 25789 5596
rect 25823 5593 25835 5627
rect 26068 5624 26096 5800
rect 26510 5788 26516 5840
rect 26568 5828 26574 5840
rect 26881 5831 26939 5837
rect 26881 5828 26893 5831
rect 26568 5800 26893 5828
rect 26568 5788 26574 5800
rect 26881 5797 26893 5800
rect 26927 5828 26939 5831
rect 32048 5828 32076 5868
rect 33413 5865 33425 5899
rect 33459 5896 33471 5899
rect 33686 5896 33692 5908
rect 33459 5868 33692 5896
rect 33459 5865 33471 5868
rect 33413 5859 33471 5865
rect 33686 5856 33692 5868
rect 33744 5856 33750 5908
rect 35342 5896 35348 5908
rect 34164 5868 35348 5896
rect 34164 5828 34192 5868
rect 35342 5856 35348 5868
rect 35400 5856 35406 5908
rect 36078 5856 36084 5908
rect 36136 5896 36142 5908
rect 37918 5896 37924 5908
rect 36136 5868 37924 5896
rect 36136 5856 36142 5868
rect 37918 5856 37924 5868
rect 37976 5856 37982 5908
rect 38010 5856 38016 5908
rect 38068 5896 38074 5908
rect 42702 5896 42708 5908
rect 38068 5868 42708 5896
rect 38068 5856 38074 5868
rect 42702 5856 42708 5868
rect 42760 5856 42766 5908
rect 42812 5868 43116 5896
rect 35066 5828 35072 5840
rect 26927 5800 31984 5828
rect 32048 5800 34192 5828
rect 34256 5800 35072 5828
rect 26927 5797 26939 5800
rect 26881 5791 26939 5797
rect 28074 5760 28080 5772
rect 26436 5732 28080 5760
rect 26436 5704 26464 5732
rect 28074 5720 28080 5732
rect 28132 5720 28138 5772
rect 26418 5692 26424 5704
rect 26331 5664 26424 5692
rect 26418 5652 26424 5664
rect 26476 5652 26482 5704
rect 27982 5652 27988 5704
rect 28040 5692 28046 5704
rect 31956 5692 31984 5800
rect 33137 5763 33195 5769
rect 33137 5729 33149 5763
rect 33183 5760 33195 5763
rect 33413 5763 33471 5769
rect 33413 5760 33425 5763
rect 33183 5732 33425 5760
rect 33183 5729 33195 5732
rect 33137 5723 33195 5729
rect 33413 5729 33425 5732
rect 33459 5729 33471 5763
rect 34256 5760 34284 5800
rect 35066 5788 35072 5800
rect 35124 5788 35130 5840
rect 35250 5788 35256 5840
rect 35308 5828 35314 5840
rect 42812 5828 42840 5868
rect 42978 5828 42984 5840
rect 35308 5800 42840 5828
rect 42939 5800 42984 5828
rect 35308 5788 35314 5800
rect 42978 5788 42984 5800
rect 43036 5788 43042 5840
rect 43088 5828 43116 5868
rect 44358 5856 44364 5908
rect 44416 5896 44422 5908
rect 45922 5896 45928 5908
rect 44416 5868 45928 5896
rect 44416 5856 44422 5868
rect 45922 5856 45928 5868
rect 45980 5856 45986 5908
rect 46201 5899 46259 5905
rect 46201 5865 46213 5899
rect 46247 5896 46259 5899
rect 46385 5899 46443 5905
rect 46385 5896 46397 5899
rect 46247 5868 46397 5896
rect 46247 5865 46259 5868
rect 46201 5859 46259 5865
rect 46385 5865 46397 5868
rect 46431 5896 46443 5899
rect 48590 5896 48596 5908
rect 46431 5868 48596 5896
rect 46431 5865 46443 5868
rect 46385 5859 46443 5865
rect 48590 5856 48596 5868
rect 48648 5856 48654 5908
rect 49786 5856 49792 5908
rect 49844 5896 49850 5908
rect 50433 5899 50491 5905
rect 49844 5868 50016 5896
rect 49844 5856 49850 5868
rect 49881 5831 49939 5837
rect 49881 5828 49893 5831
rect 43088 5800 49893 5828
rect 49881 5797 49893 5800
rect 49927 5797 49939 5831
rect 49988 5828 50016 5868
rect 50433 5865 50445 5899
rect 50479 5896 50491 5899
rect 50709 5899 50767 5905
rect 50709 5896 50721 5899
rect 50479 5868 50721 5896
rect 50479 5865 50491 5868
rect 50433 5859 50491 5865
rect 50709 5865 50721 5868
rect 50755 5896 50767 5899
rect 51074 5896 51080 5908
rect 50755 5868 51080 5896
rect 50755 5865 50767 5868
rect 50709 5859 50767 5865
rect 51074 5856 51080 5868
rect 51132 5856 51138 5908
rect 51258 5856 51264 5908
rect 51316 5896 51322 5908
rect 56873 5899 56931 5905
rect 56873 5896 56885 5899
rect 51316 5868 56885 5896
rect 51316 5856 51322 5868
rect 56873 5865 56885 5868
rect 56919 5865 56931 5899
rect 56873 5859 56931 5865
rect 56962 5856 56968 5908
rect 57020 5896 57026 5908
rect 57238 5896 57244 5908
rect 57020 5868 57244 5896
rect 57020 5856 57026 5868
rect 57238 5856 57244 5868
rect 57296 5856 57302 5908
rect 57422 5896 57428 5908
rect 57383 5868 57428 5896
rect 57422 5856 57428 5868
rect 57480 5856 57486 5908
rect 57885 5899 57943 5905
rect 57885 5896 57897 5899
rect 57532 5868 57897 5896
rect 57532 5828 57560 5868
rect 57885 5865 57897 5868
rect 57931 5865 57943 5899
rect 57885 5859 57943 5865
rect 58437 5899 58495 5905
rect 58437 5865 58449 5899
rect 58483 5896 58495 5899
rect 58713 5899 58771 5905
rect 58713 5896 58725 5899
rect 58483 5868 58725 5896
rect 58483 5865 58495 5868
rect 58437 5859 58495 5865
rect 58713 5865 58725 5868
rect 58759 5896 58771 5899
rect 59722 5896 59728 5908
rect 58759 5868 59728 5896
rect 58759 5865 58771 5868
rect 58713 5859 58771 5865
rect 59722 5856 59728 5868
rect 59780 5856 59786 5908
rect 64506 5896 64512 5908
rect 64467 5868 64512 5896
rect 64506 5856 64512 5868
rect 64564 5856 64570 5908
rect 69934 5896 69940 5908
rect 69895 5868 69940 5896
rect 69934 5856 69940 5868
rect 69992 5856 69998 5908
rect 90266 5896 90272 5908
rect 90227 5868 90272 5896
rect 90266 5856 90272 5868
rect 90324 5856 90330 5908
rect 65426 5828 65432 5840
rect 49988 5800 57560 5828
rect 57624 5800 65432 5828
rect 49881 5791 49939 5797
rect 33413 5723 33471 5729
rect 33520 5732 34284 5760
rect 33520 5692 33548 5732
rect 34974 5720 34980 5772
rect 35032 5760 35038 5772
rect 35161 5763 35219 5769
rect 35161 5760 35173 5763
rect 35032 5732 35173 5760
rect 35032 5720 35038 5732
rect 35161 5729 35173 5732
rect 35207 5729 35219 5763
rect 35161 5723 35219 5729
rect 35342 5720 35348 5772
rect 35400 5760 35406 5772
rect 36630 5760 36636 5772
rect 35400 5732 36636 5760
rect 35400 5720 35406 5732
rect 36630 5720 36636 5732
rect 36688 5720 36694 5772
rect 37001 5763 37059 5769
rect 37001 5729 37013 5763
rect 37047 5760 37059 5763
rect 37090 5760 37096 5772
rect 37047 5732 37096 5760
rect 37047 5729 37059 5732
rect 37001 5723 37059 5729
rect 37090 5720 37096 5732
rect 37148 5720 37154 5772
rect 37274 5720 37280 5772
rect 37332 5760 37338 5772
rect 37826 5760 37832 5772
rect 37332 5732 37832 5760
rect 37332 5720 37338 5732
rect 37826 5720 37832 5732
rect 37884 5720 37890 5772
rect 37918 5720 37924 5772
rect 37976 5760 37982 5772
rect 40494 5760 40500 5772
rect 37976 5732 40500 5760
rect 37976 5720 37982 5732
rect 40494 5720 40500 5732
rect 40552 5720 40558 5772
rect 41509 5763 41567 5769
rect 41509 5729 41521 5763
rect 41555 5760 41567 5763
rect 41690 5760 41696 5772
rect 41555 5732 41696 5760
rect 41555 5729 41567 5732
rect 41509 5723 41567 5729
rect 41690 5720 41696 5732
rect 41748 5760 41754 5772
rect 41969 5763 42027 5769
rect 41969 5760 41981 5763
rect 41748 5732 41981 5760
rect 41748 5720 41754 5732
rect 41969 5729 41981 5732
rect 42015 5729 42027 5763
rect 47486 5760 47492 5772
rect 41969 5723 42027 5729
rect 42076 5732 47492 5760
rect 28040 5664 31248 5692
rect 31956 5664 33548 5692
rect 34057 5695 34115 5701
rect 28040 5652 28046 5664
rect 31113 5627 31171 5633
rect 31113 5624 31125 5627
rect 26068 5596 31125 5624
rect 25777 5587 25835 5593
rect 31113 5593 31125 5596
rect 31159 5593 31171 5627
rect 31220 5624 31248 5664
rect 34057 5661 34069 5695
rect 34103 5692 34115 5695
rect 34146 5692 34152 5704
rect 34103 5664 34152 5692
rect 34103 5661 34115 5664
rect 34057 5655 34115 5661
rect 34146 5652 34152 5664
rect 34204 5652 34210 5704
rect 35621 5695 35679 5701
rect 35621 5661 35633 5695
rect 35667 5692 35679 5695
rect 35667 5664 36124 5692
rect 35667 5661 35679 5664
rect 35621 5655 35679 5661
rect 34238 5624 34244 5636
rect 31220 5596 34244 5624
rect 31113 5587 31171 5593
rect 34238 5584 34244 5596
rect 34296 5584 34302 5636
rect 34790 5584 34796 5636
rect 34848 5624 34854 5636
rect 35894 5624 35900 5636
rect 34848 5596 35900 5624
rect 34848 5584 34854 5596
rect 35894 5584 35900 5596
rect 35952 5584 35958 5636
rect 36096 5633 36124 5664
rect 36262 5652 36268 5704
rect 36320 5692 36326 5704
rect 39850 5692 39856 5704
rect 36320 5664 39856 5692
rect 36320 5652 36326 5664
rect 39850 5652 39856 5664
rect 39908 5652 39914 5704
rect 40310 5652 40316 5704
rect 40368 5692 40374 5704
rect 42076 5692 42104 5732
rect 47486 5720 47492 5732
rect 47544 5720 47550 5772
rect 47854 5720 47860 5772
rect 47912 5760 47918 5772
rect 51166 5760 51172 5772
rect 47912 5732 50568 5760
rect 51127 5732 51172 5760
rect 47912 5720 47918 5732
rect 40368 5664 42104 5692
rect 40368 5652 40374 5664
rect 42150 5652 42156 5704
rect 42208 5692 42214 5704
rect 44542 5692 44548 5704
rect 42208 5664 44548 5692
rect 42208 5652 42214 5664
rect 44542 5652 44548 5664
rect 44600 5652 44606 5704
rect 45925 5695 45983 5701
rect 45112 5664 45416 5692
rect 36081 5627 36139 5633
rect 36081 5593 36093 5627
rect 36127 5624 36139 5627
rect 45112 5624 45140 5664
rect 45278 5624 45284 5636
rect 36127 5596 45140 5624
rect 45239 5596 45284 5624
rect 36127 5593 36139 5596
rect 36081 5587 36139 5593
rect 45278 5584 45284 5596
rect 45336 5584 45342 5636
rect 45388 5624 45416 5664
rect 45925 5661 45937 5695
rect 45971 5692 45983 5695
rect 46201 5695 46259 5701
rect 46201 5692 46213 5695
rect 45971 5664 46213 5692
rect 45971 5661 45983 5664
rect 45925 5655 45983 5661
rect 46201 5661 46213 5664
rect 46247 5661 46259 5695
rect 46201 5655 46259 5661
rect 46290 5652 46296 5704
rect 46348 5692 46354 5704
rect 50062 5692 50068 5704
rect 46348 5664 50068 5692
rect 46348 5652 46354 5664
rect 50062 5652 50068 5664
rect 50120 5652 50126 5704
rect 50249 5695 50307 5701
rect 50249 5661 50261 5695
rect 50295 5692 50307 5695
rect 50433 5695 50491 5701
rect 50433 5692 50445 5695
rect 50295 5664 50445 5692
rect 50295 5661 50307 5664
rect 50249 5655 50307 5661
rect 50433 5661 50445 5664
rect 50479 5661 50491 5695
rect 50540 5692 50568 5732
rect 51166 5720 51172 5732
rect 51224 5760 51230 5772
rect 51629 5763 51687 5769
rect 51629 5760 51641 5763
rect 51224 5732 51641 5760
rect 51224 5720 51230 5732
rect 51629 5729 51641 5732
rect 51675 5729 51687 5763
rect 52638 5760 52644 5772
rect 52599 5732 52644 5760
rect 51629 5723 51687 5729
rect 52638 5720 52644 5732
rect 52696 5720 52702 5772
rect 52730 5720 52736 5772
rect 52788 5760 52794 5772
rect 54481 5763 54539 5769
rect 54481 5760 54493 5763
rect 52788 5732 54493 5760
rect 52788 5720 52794 5732
rect 54481 5729 54493 5732
rect 54527 5729 54539 5763
rect 54481 5723 54539 5729
rect 54662 5720 54668 5772
rect 54720 5760 54726 5772
rect 55309 5763 55367 5769
rect 54720 5732 55260 5760
rect 54720 5720 54726 5732
rect 55122 5692 55128 5704
rect 50540 5664 54984 5692
rect 55083 5664 55128 5692
rect 50433 5655 50491 5661
rect 47394 5624 47400 5636
rect 45388 5596 47400 5624
rect 47394 5584 47400 5596
rect 47452 5584 47458 5636
rect 47486 5584 47492 5636
rect 47544 5624 47550 5636
rect 54846 5624 54852 5636
rect 47544 5596 54852 5624
rect 47544 5584 47550 5596
rect 54846 5584 54852 5596
rect 54904 5584 54910 5636
rect 54956 5624 54984 5664
rect 55122 5652 55128 5664
rect 55180 5652 55186 5704
rect 55232 5692 55260 5732
rect 55309 5729 55321 5763
rect 55355 5760 55367 5763
rect 56045 5763 56103 5769
rect 56045 5760 56057 5763
rect 55355 5732 56057 5760
rect 55355 5729 55367 5732
rect 55309 5723 55367 5729
rect 56045 5729 56057 5732
rect 56091 5729 56103 5763
rect 57624 5760 57652 5800
rect 65426 5788 65432 5800
rect 65484 5788 65490 5840
rect 89441 5831 89499 5837
rect 89441 5797 89453 5831
rect 89487 5828 89499 5831
rect 93044 5828 93072 6072
rect 100938 6060 100944 6072
rect 100996 6060 101002 6112
rect 107746 6060 107752 6112
rect 107804 6100 107810 6112
rect 117682 6100 117688 6112
rect 107804 6072 117688 6100
rect 107804 6060 107810 6072
rect 117682 6060 117688 6072
rect 117740 6060 117746 6112
rect 124122 6060 124128 6112
rect 124180 6060 124186 6112
rect 143460 6100 143488 6140
rect 143644 6140 148876 6168
rect 143644 6100 143672 6140
rect 148870 6128 148876 6140
rect 148928 6128 148934 6180
rect 150250 6128 150256 6180
rect 150308 6168 150314 6180
rect 154669 6171 154727 6177
rect 154669 6168 154681 6171
rect 150308 6140 154681 6168
rect 150308 6128 150314 6140
rect 154669 6137 154681 6140
rect 154715 6137 154727 6171
rect 154669 6131 154727 6137
rect 157426 6128 157432 6180
rect 157484 6168 157490 6180
rect 164878 6168 164884 6180
rect 157484 6140 164884 6168
rect 157484 6128 157490 6140
rect 164878 6128 164884 6140
rect 164936 6128 164942 6180
rect 165154 6168 165160 6180
rect 165115 6140 165160 6168
rect 165154 6128 165160 6140
rect 165212 6128 165218 6180
rect 156322 6100 156328 6112
rect 143460 6072 143672 6100
rect 156283 6072 156328 6100
rect 156322 6060 156328 6072
rect 156380 6060 156386 6112
rect 163590 6100 163596 6112
rect 163551 6072 163596 6100
rect 163590 6060 163596 6072
rect 163648 6060 163654 6112
rect 102028 6010 169556 6032
rect 93210 5924 93216 5976
rect 93268 5964 93274 5976
rect 93268 5936 101444 5964
rect 102028 5958 141299 6010
rect 141351 5958 141363 6010
rect 141415 5958 141427 6010
rect 141479 5958 141491 6010
rect 141543 5958 169556 6010
rect 102028 5936 169556 5958
rect 93268 5924 93274 5936
rect 101416 5896 101444 5936
rect 116118 5896 116124 5908
rect 101416 5868 116124 5896
rect 116118 5856 116124 5868
rect 116176 5856 116182 5908
rect 116210 5856 116216 5908
rect 116268 5896 116274 5908
rect 116305 5899 116363 5905
rect 116305 5896 116317 5899
rect 116268 5868 116317 5896
rect 116268 5856 116274 5868
rect 116305 5865 116317 5868
rect 116351 5865 116363 5899
rect 128906 5896 128912 5908
rect 116305 5859 116363 5865
rect 121472 5868 123892 5896
rect 128867 5868 128912 5896
rect 89487 5800 93072 5828
rect 95053 5831 95111 5837
rect 89487 5797 89499 5800
rect 89441 5791 89499 5797
rect 95053 5797 95065 5831
rect 95099 5828 95111 5831
rect 106642 5828 106648 5840
rect 95099 5800 106648 5828
rect 95099 5797 95111 5800
rect 95053 5791 95111 5797
rect 58437 5763 58495 5769
rect 58437 5760 58449 5763
rect 56045 5723 56103 5729
rect 56152 5732 57652 5760
rect 57808 5732 58449 5760
rect 56152 5692 56180 5732
rect 56594 5692 56600 5704
rect 55232 5664 56180 5692
rect 56244 5664 56600 5692
rect 55309 5627 55367 5633
rect 55309 5624 55321 5627
rect 54956 5596 55321 5624
rect 55309 5593 55321 5596
rect 55355 5593 55367 5627
rect 55309 5587 55367 5593
rect 55490 5584 55496 5636
rect 55548 5624 55554 5636
rect 56244 5624 56272 5664
rect 56594 5652 56600 5664
rect 56652 5652 56658 5704
rect 56689 5695 56747 5701
rect 56689 5661 56701 5695
rect 56735 5692 56747 5695
rect 57149 5695 57207 5701
rect 57149 5692 57161 5695
rect 56735 5664 57161 5692
rect 56735 5661 56747 5664
rect 56689 5655 56747 5661
rect 57149 5661 57161 5664
rect 57195 5692 57207 5695
rect 57514 5692 57520 5704
rect 57195 5664 57520 5692
rect 57195 5661 57207 5664
rect 57149 5655 57207 5661
rect 57514 5652 57520 5664
rect 57572 5652 57578 5704
rect 57701 5695 57759 5701
rect 57701 5661 57713 5695
rect 57747 5692 57759 5695
rect 57808 5692 57836 5732
rect 58437 5729 58449 5732
rect 58483 5729 58495 5763
rect 58437 5723 58495 5729
rect 59814 5720 59820 5772
rect 59872 5760 59878 5772
rect 66806 5760 66812 5772
rect 59872 5732 66812 5760
rect 59872 5720 59878 5732
rect 66806 5720 66812 5732
rect 66864 5720 66870 5772
rect 87506 5760 87512 5772
rect 87467 5732 87512 5760
rect 87506 5720 87512 5732
rect 87564 5720 87570 5772
rect 88702 5760 88708 5772
rect 88663 5732 88708 5760
rect 88702 5720 88708 5732
rect 88760 5720 88766 5772
rect 63310 5692 63316 5704
rect 57747 5664 57836 5692
rect 57900 5664 63316 5692
rect 57747 5661 57759 5664
rect 57701 5655 57759 5661
rect 57900 5624 57928 5664
rect 63310 5652 63316 5664
rect 63368 5652 63374 5704
rect 89073 5695 89131 5701
rect 89073 5661 89085 5695
rect 89119 5692 89131 5695
rect 89456 5692 89484 5791
rect 106642 5788 106648 5800
rect 106700 5788 106706 5840
rect 106734 5788 106740 5840
rect 106792 5828 106798 5840
rect 121472 5828 121500 5868
rect 106792 5800 121500 5828
rect 106792 5788 106798 5800
rect 94961 5763 95019 5769
rect 94961 5729 94973 5763
rect 95007 5760 95019 5763
rect 107654 5760 107660 5772
rect 95007 5732 107660 5760
rect 95007 5729 95019 5732
rect 94961 5723 95019 5729
rect 107654 5720 107660 5732
rect 107712 5720 107718 5772
rect 112714 5760 112720 5772
rect 110432 5732 112720 5760
rect 89119 5664 89484 5692
rect 102321 5695 102379 5701
rect 89119 5661 89131 5664
rect 89073 5655 89131 5661
rect 102321 5661 102333 5695
rect 102367 5692 102379 5695
rect 102597 5695 102655 5701
rect 102597 5692 102609 5695
rect 102367 5664 102609 5692
rect 102367 5661 102379 5664
rect 102321 5655 102379 5661
rect 102597 5661 102609 5664
rect 102643 5661 102655 5695
rect 102597 5655 102655 5661
rect 104434 5652 104440 5704
rect 104492 5692 104498 5704
rect 110432 5692 110460 5732
rect 112714 5720 112720 5732
rect 112772 5720 112778 5772
rect 115201 5763 115259 5769
rect 115201 5760 115213 5763
rect 114572 5732 115213 5760
rect 104492 5664 110460 5692
rect 110877 5695 110935 5701
rect 104492 5652 104498 5664
rect 110877 5661 110889 5695
rect 110923 5692 110935 5695
rect 111153 5695 111211 5701
rect 111153 5692 111165 5695
rect 110923 5664 111165 5692
rect 110923 5661 110935 5664
rect 110877 5655 110935 5661
rect 111153 5661 111165 5664
rect 111199 5661 111211 5695
rect 114572 5692 114600 5732
rect 115201 5729 115213 5732
rect 115247 5760 115259 5763
rect 118326 5760 118332 5772
rect 115247 5732 118332 5760
rect 115247 5729 115259 5732
rect 115201 5723 115259 5729
rect 118326 5720 118332 5732
rect 118384 5720 118390 5772
rect 123864 5769 123892 5868
rect 128906 5856 128912 5868
rect 128964 5856 128970 5908
rect 148410 5896 148416 5908
rect 148371 5868 148416 5896
rect 148410 5856 148416 5868
rect 148468 5856 148474 5908
rect 152921 5899 152979 5905
rect 152921 5865 152933 5899
rect 152967 5896 152979 5899
rect 153378 5896 153384 5908
rect 152967 5868 153384 5896
rect 152967 5865 152979 5868
rect 152921 5859 152979 5865
rect 153378 5856 153384 5868
rect 153436 5856 153442 5908
rect 157426 5896 157432 5908
rect 153488 5868 157432 5896
rect 123849 5763 123907 5769
rect 123849 5729 123861 5763
rect 123895 5729 123907 5763
rect 128924 5760 128952 5856
rect 129001 5763 129059 5769
rect 129001 5760 129013 5763
rect 128924 5732 129013 5760
rect 123849 5723 123907 5729
rect 129001 5729 129013 5732
rect 129047 5729 129059 5763
rect 130010 5760 130016 5772
rect 129971 5732 130016 5760
rect 129001 5723 129059 5729
rect 130010 5720 130016 5732
rect 130068 5720 130074 5772
rect 148428 5760 148456 5856
rect 148870 5788 148876 5840
rect 148928 5828 148934 5840
rect 153488 5828 153516 5868
rect 157426 5856 157432 5868
rect 157484 5856 157490 5908
rect 157518 5856 157524 5908
rect 157576 5896 157582 5908
rect 158257 5899 158315 5905
rect 158257 5896 158269 5899
rect 157576 5868 158269 5896
rect 157576 5856 157582 5868
rect 158257 5865 158269 5868
rect 158303 5865 158315 5899
rect 159266 5896 159272 5908
rect 159227 5868 159272 5896
rect 158257 5859 158315 5865
rect 159266 5856 159272 5868
rect 159324 5856 159330 5908
rect 163498 5896 163504 5908
rect 163459 5868 163504 5896
rect 163498 5856 163504 5868
rect 163556 5856 163562 5908
rect 148928 5800 153516 5828
rect 154485 5831 154543 5837
rect 148928 5788 148934 5800
rect 154485 5797 154497 5831
rect 154531 5828 154543 5831
rect 154666 5828 154672 5840
rect 154531 5800 154672 5828
rect 154531 5797 154543 5800
rect 154485 5791 154543 5797
rect 154666 5788 154672 5800
rect 154724 5788 154730 5840
rect 148781 5763 148839 5769
rect 148781 5760 148793 5763
rect 148428 5732 148793 5760
rect 148781 5729 148793 5732
rect 148827 5729 148839 5763
rect 148781 5723 148839 5729
rect 150989 5763 151047 5769
rect 150989 5729 151001 5763
rect 151035 5760 151047 5763
rect 153838 5760 153844 5772
rect 151035 5732 153844 5760
rect 151035 5729 151047 5732
rect 150989 5723 151047 5729
rect 153838 5720 153844 5732
rect 153896 5720 153902 5772
rect 156414 5720 156420 5772
rect 156472 5760 156478 5772
rect 156785 5763 156843 5769
rect 156785 5760 156797 5763
rect 156472 5732 156797 5760
rect 156472 5720 156478 5732
rect 156785 5729 156797 5732
rect 156831 5729 156843 5763
rect 156785 5723 156843 5729
rect 162581 5763 162639 5769
rect 162581 5729 162593 5763
rect 162627 5760 162639 5763
rect 163590 5760 163596 5772
rect 162627 5732 163596 5760
rect 162627 5729 162639 5732
rect 162581 5723 162639 5729
rect 163590 5720 163596 5732
rect 163648 5720 163654 5772
rect 164694 5760 164700 5772
rect 164655 5732 164700 5760
rect 164694 5720 164700 5732
rect 164752 5720 164758 5772
rect 114649 5695 114707 5701
rect 114649 5692 114661 5695
rect 114572 5664 114661 5692
rect 111153 5655 111211 5661
rect 114649 5661 114661 5664
rect 114695 5661 114707 5695
rect 114649 5655 114707 5661
rect 116213 5695 116271 5701
rect 116213 5661 116225 5695
rect 116259 5661 116271 5695
rect 116213 5655 116271 5661
rect 120997 5695 121055 5701
rect 120997 5661 121009 5695
rect 121043 5692 121055 5695
rect 121454 5692 121460 5704
rect 121043 5664 121460 5692
rect 121043 5661 121055 5664
rect 120997 5655 121055 5661
rect 55548 5596 56272 5624
rect 56336 5596 57928 5624
rect 55548 5584 55554 5596
rect 21232 5528 22692 5556
rect 22741 5559 22799 5565
rect 21232 5516 21238 5528
rect 22741 5525 22753 5559
rect 22787 5556 22799 5559
rect 23017 5559 23075 5565
rect 23017 5556 23029 5559
rect 22787 5528 23029 5556
rect 22787 5525 22799 5528
rect 22741 5519 22799 5525
rect 23017 5525 23029 5528
rect 23063 5556 23075 5559
rect 26510 5556 26516 5568
rect 23063 5528 26516 5556
rect 23063 5525 23075 5528
rect 23017 5519 23075 5525
rect 26510 5516 26516 5528
rect 26568 5516 26574 5568
rect 30374 5516 30380 5568
rect 30432 5556 30438 5568
rect 36446 5556 36452 5568
rect 30432 5528 36452 5556
rect 30432 5516 30438 5528
rect 36446 5516 36452 5528
rect 36504 5516 36510 5568
rect 38194 5516 38200 5568
rect 38252 5556 38258 5568
rect 41874 5556 41880 5568
rect 38252 5528 41880 5556
rect 38252 5516 38258 5528
rect 41874 5516 41880 5528
rect 41932 5516 41938 5568
rect 41966 5516 41972 5568
rect 42024 5556 42030 5568
rect 42334 5556 42340 5568
rect 42024 5528 42340 5556
rect 42024 5516 42030 5528
rect 42334 5516 42340 5528
rect 42392 5516 42398 5568
rect 42426 5516 42432 5568
rect 42484 5556 42490 5568
rect 46842 5556 46848 5568
rect 42484 5528 46848 5556
rect 42484 5516 42490 5528
rect 46842 5516 46848 5528
rect 46900 5516 46906 5568
rect 47029 5559 47087 5565
rect 47029 5525 47041 5559
rect 47075 5556 47087 5559
rect 47210 5556 47216 5568
rect 47075 5528 47216 5556
rect 47075 5525 47087 5528
rect 47029 5519 47087 5525
rect 47210 5516 47216 5528
rect 47268 5556 47274 5568
rect 55030 5556 55036 5568
rect 47268 5528 55036 5556
rect 47268 5516 47274 5528
rect 55030 5516 55036 5528
rect 55088 5516 55094 5568
rect 55122 5516 55128 5568
rect 55180 5556 55186 5568
rect 55585 5559 55643 5565
rect 55585 5556 55597 5559
rect 55180 5528 55597 5556
rect 55180 5516 55186 5528
rect 55585 5525 55597 5528
rect 55631 5556 55643 5559
rect 55950 5556 55956 5568
rect 55631 5528 55956 5556
rect 55631 5525 55643 5528
rect 55585 5519 55643 5525
rect 55950 5516 55956 5528
rect 56008 5516 56014 5568
rect 56134 5516 56140 5568
rect 56192 5556 56198 5568
rect 56336 5556 56364 5596
rect 58342 5584 58348 5636
rect 58400 5624 58406 5636
rect 69106 5624 69112 5636
rect 58400 5596 69112 5624
rect 58400 5584 58406 5596
rect 69106 5584 69112 5596
rect 69164 5584 69170 5636
rect 91278 5584 91284 5636
rect 91336 5624 91342 5636
rect 91741 5627 91799 5633
rect 91741 5624 91753 5627
rect 91336 5596 91753 5624
rect 91336 5584 91342 5596
rect 91741 5593 91753 5596
rect 91787 5593 91799 5627
rect 101398 5624 101404 5636
rect 91741 5587 91799 5593
rect 94056 5596 101404 5624
rect 56192 5528 56364 5556
rect 56873 5559 56931 5565
rect 56192 5516 56198 5528
rect 56873 5525 56885 5559
rect 56919 5556 56931 5559
rect 58986 5556 58992 5568
rect 56919 5528 58992 5556
rect 56919 5525 56931 5528
rect 56873 5519 56931 5525
rect 58986 5516 58992 5528
rect 59044 5516 59050 5568
rect 59081 5559 59139 5565
rect 59081 5525 59093 5559
rect 59127 5556 59139 5559
rect 59262 5556 59268 5568
rect 59127 5528 59268 5556
rect 59127 5525 59139 5528
rect 59081 5519 59139 5525
rect 59262 5516 59268 5528
rect 59320 5556 59326 5568
rect 64414 5556 64420 5568
rect 59320 5528 64420 5556
rect 59320 5516 59326 5528
rect 64414 5516 64420 5528
rect 64472 5516 64478 5568
rect 65889 5559 65947 5565
rect 65889 5525 65901 5559
rect 65935 5556 65947 5559
rect 66070 5556 66076 5568
rect 65935 5528 66076 5556
rect 65935 5525 65947 5528
rect 65889 5519 65947 5525
rect 66070 5516 66076 5528
rect 66128 5556 66134 5568
rect 71038 5556 71044 5568
rect 66128 5528 71044 5556
rect 66128 5516 66134 5528
rect 71038 5516 71044 5528
rect 71096 5516 71102 5568
rect 71317 5559 71375 5565
rect 71317 5525 71329 5559
rect 71363 5556 71375 5559
rect 71774 5556 71780 5568
rect 71363 5528 71780 5556
rect 71363 5525 71375 5528
rect 71317 5519 71375 5525
rect 71774 5516 71780 5528
rect 71832 5516 71838 5568
rect 90726 5556 90732 5568
rect 90687 5528 90732 5556
rect 90726 5516 90732 5528
rect 90784 5516 90790 5568
rect 91649 5559 91707 5565
rect 91649 5525 91661 5559
rect 91695 5556 91707 5559
rect 91830 5556 91836 5568
rect 91695 5528 91836 5556
rect 91695 5525 91707 5528
rect 91649 5519 91707 5525
rect 91830 5516 91836 5528
rect 91888 5556 91894 5568
rect 94056 5556 94084 5596
rect 101398 5584 101404 5596
rect 101456 5584 101462 5636
rect 101493 5627 101551 5633
rect 101493 5593 101505 5627
rect 101539 5624 101551 5627
rect 104066 5624 104072 5636
rect 101539 5596 104072 5624
rect 101539 5593 101551 5596
rect 101493 5587 101551 5593
rect 104066 5584 104072 5596
rect 104124 5584 104130 5636
rect 108758 5624 108764 5636
rect 104360 5596 108764 5624
rect 91888 5528 94084 5556
rect 94961 5559 95019 5565
rect 91888 5516 91894 5528
rect 94961 5525 94973 5559
rect 95007 5556 95019 5559
rect 99009 5559 99067 5565
rect 99009 5556 99021 5559
rect 95007 5528 99021 5556
rect 95007 5525 95019 5528
rect 94961 5519 95019 5525
rect 99009 5525 99021 5528
rect 99055 5525 99067 5559
rect 99009 5519 99067 5525
rect 99098 5516 99104 5568
rect 99156 5556 99162 5568
rect 99156 5528 99512 5556
rect 99156 5516 99162 5528
rect 93121 5491 93179 5497
rect 368 5466 93012 5488
rect 368 5414 56667 5466
rect 56719 5414 56731 5466
rect 56783 5414 56795 5466
rect 56847 5414 56859 5466
rect 56911 5414 93012 5466
rect 93121 5457 93133 5491
rect 93167 5488 93179 5491
rect 99285 5491 99343 5497
rect 93167 5460 99236 5488
rect 93167 5457 93179 5460
rect 93121 5451 93179 5457
rect 99098 5420 99104 5432
rect 368 5392 93012 5414
rect 93044 5392 99104 5420
rect 7285 5355 7343 5361
rect 7285 5321 7297 5355
rect 7331 5352 7343 5355
rect 8018 5352 8024 5364
rect 7331 5324 8024 5352
rect 7331 5321 7343 5324
rect 7285 5315 7343 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 43530 5352 43536 5364
rect 14476 5324 43536 5352
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 14476 5284 14504 5324
rect 43530 5312 43536 5324
rect 43588 5312 43594 5364
rect 43622 5312 43628 5364
rect 43680 5352 43686 5364
rect 45646 5352 45652 5364
rect 43680 5324 45652 5352
rect 43680 5312 43686 5324
rect 45646 5312 45652 5324
rect 45704 5312 45710 5364
rect 45741 5355 45799 5361
rect 45741 5321 45753 5355
rect 45787 5352 45799 5355
rect 45830 5352 45836 5364
rect 45787 5324 45836 5352
rect 45787 5321 45799 5324
rect 45741 5315 45799 5321
rect 45830 5312 45836 5324
rect 45888 5312 45894 5364
rect 46106 5312 46112 5364
rect 46164 5352 46170 5364
rect 51074 5352 51080 5364
rect 46164 5324 51080 5352
rect 46164 5312 46170 5324
rect 51074 5312 51080 5324
rect 51132 5312 51138 5364
rect 51350 5312 51356 5364
rect 51408 5352 51414 5364
rect 57238 5352 57244 5364
rect 51408 5324 57244 5352
rect 51408 5312 51414 5324
rect 57238 5312 57244 5324
rect 57296 5312 57302 5364
rect 63862 5312 63868 5364
rect 63920 5352 63926 5364
rect 67082 5352 67088 5364
rect 63920 5324 67088 5352
rect 63920 5312 63926 5324
rect 67082 5312 67088 5324
rect 67140 5312 67146 5364
rect 92934 5312 92940 5364
rect 92992 5352 92998 5364
rect 93044 5352 93072 5392
rect 99098 5380 99104 5392
rect 99156 5380 99162 5432
rect 99208 5420 99236 5460
rect 99285 5457 99297 5491
rect 99331 5488 99343 5491
rect 99377 5491 99435 5497
rect 99377 5488 99389 5491
rect 99331 5460 99389 5488
rect 99331 5457 99343 5460
rect 99285 5451 99343 5457
rect 99377 5457 99389 5460
rect 99423 5457 99435 5491
rect 99484 5488 99512 5528
rect 102226 5516 102232 5568
rect 102284 5556 102290 5568
rect 102413 5559 102471 5565
rect 102413 5556 102425 5559
rect 102284 5528 102425 5556
rect 102284 5516 102290 5528
rect 102413 5525 102425 5528
rect 102459 5525 102471 5559
rect 102413 5519 102471 5525
rect 102597 5559 102655 5565
rect 102597 5525 102609 5559
rect 102643 5556 102655 5559
rect 102873 5559 102931 5565
rect 102873 5556 102885 5559
rect 102643 5528 102885 5556
rect 102643 5525 102655 5528
rect 102597 5519 102655 5525
rect 102873 5525 102885 5528
rect 102919 5556 102931 5559
rect 104360 5556 104388 5596
rect 108758 5584 108764 5596
rect 108816 5584 108822 5636
rect 114741 5627 114799 5633
rect 114741 5624 114753 5627
rect 110892 5596 114753 5624
rect 102919 5528 104388 5556
rect 102919 5525 102931 5528
rect 102873 5519 102931 5525
rect 104526 5516 104532 5568
rect 104584 5556 104590 5568
rect 110892 5556 110920 5596
rect 114741 5593 114753 5596
rect 114787 5593 114799 5627
rect 116228 5624 116256 5655
rect 121454 5652 121460 5664
rect 121512 5652 121518 5704
rect 121822 5692 121828 5704
rect 121783 5664 121828 5692
rect 121822 5652 121828 5664
rect 121880 5652 121886 5704
rect 122834 5692 122840 5704
rect 122795 5664 122840 5692
rect 122834 5652 122840 5664
rect 122892 5652 122898 5704
rect 124401 5695 124459 5701
rect 124401 5661 124413 5695
rect 124447 5692 124459 5695
rect 130565 5695 130623 5701
rect 124447 5664 124812 5692
rect 124447 5661 124459 5664
rect 124401 5655 124459 5661
rect 116765 5627 116823 5633
rect 116765 5624 116777 5627
rect 116228 5596 116777 5624
rect 114741 5587 114799 5593
rect 116765 5593 116777 5596
rect 116811 5624 116823 5627
rect 123110 5624 123116 5636
rect 116811 5596 123116 5624
rect 116811 5593 116823 5596
rect 116765 5587 116823 5593
rect 123110 5584 123116 5596
rect 123168 5584 123174 5636
rect 104584 5528 110920 5556
rect 104584 5516 104590 5528
rect 110966 5516 110972 5568
rect 111024 5556 111030 5568
rect 111153 5559 111211 5565
rect 111024 5528 111069 5556
rect 111024 5516 111030 5528
rect 111153 5525 111165 5559
rect 111199 5556 111211 5559
rect 111429 5559 111487 5565
rect 111429 5556 111441 5559
rect 111199 5528 111441 5556
rect 111199 5525 111211 5528
rect 111153 5519 111211 5525
rect 111429 5525 111441 5528
rect 111475 5556 111487 5559
rect 114646 5556 114652 5568
rect 111475 5528 114652 5556
rect 111475 5525 111487 5528
rect 111429 5519 111487 5525
rect 114646 5516 114652 5528
rect 114704 5516 114710 5568
rect 114830 5516 114836 5568
rect 114888 5556 114894 5568
rect 116854 5556 116860 5568
rect 114888 5528 116860 5556
rect 114888 5516 114894 5528
rect 116854 5516 116860 5528
rect 116912 5516 116918 5568
rect 122377 5559 122435 5565
rect 122377 5525 122389 5559
rect 122423 5556 122435 5559
rect 123018 5556 123024 5568
rect 122423 5528 123024 5556
rect 122423 5525 122435 5528
rect 122377 5519 122435 5525
rect 123018 5516 123024 5528
rect 123076 5556 123082 5568
rect 123754 5556 123760 5568
rect 123076 5528 123760 5556
rect 123076 5516 123082 5528
rect 123754 5516 123760 5528
rect 123812 5516 123818 5568
rect 124784 5565 124812 5664
rect 130565 5661 130577 5695
rect 130611 5692 130623 5695
rect 153013 5695 153071 5701
rect 130611 5664 130976 5692
rect 130611 5661 130623 5664
rect 130565 5655 130623 5661
rect 130948 5568 130976 5664
rect 153013 5661 153025 5695
rect 153059 5692 153071 5695
rect 153470 5692 153476 5704
rect 153059 5664 153476 5692
rect 153059 5661 153071 5664
rect 153013 5655 153071 5661
rect 153470 5652 153476 5664
rect 153528 5652 153534 5704
rect 154577 5695 154635 5701
rect 154577 5661 154589 5695
rect 154623 5692 154635 5695
rect 155773 5695 155831 5701
rect 154623 5664 155356 5692
rect 154623 5661 154635 5664
rect 154577 5655 154635 5661
rect 124769 5559 124827 5565
rect 124769 5525 124781 5559
rect 124815 5556 124827 5559
rect 126054 5556 126060 5568
rect 124815 5528 126060 5556
rect 124815 5525 124827 5528
rect 124769 5519 124827 5525
rect 126054 5516 126060 5528
rect 126112 5516 126118 5568
rect 130930 5556 130936 5568
rect 130891 5528 130936 5556
rect 130930 5516 130936 5528
rect 130988 5516 130994 5568
rect 150066 5556 150072 5568
rect 150027 5528 150072 5556
rect 150066 5516 150072 5528
rect 150124 5516 150130 5568
rect 151998 5556 152004 5568
rect 151959 5528 152004 5556
rect 151998 5516 152004 5528
rect 152056 5516 152062 5568
rect 154574 5516 154580 5568
rect 154632 5556 154638 5568
rect 154850 5556 154856 5568
rect 154632 5528 154856 5556
rect 154632 5516 154638 5528
rect 154850 5516 154856 5528
rect 154908 5516 154914 5568
rect 155328 5565 155356 5664
rect 155773 5661 155785 5695
rect 155819 5692 155831 5695
rect 156322 5692 156328 5704
rect 155819 5664 156328 5692
rect 155819 5661 155831 5664
rect 155773 5655 155831 5661
rect 156322 5652 156328 5664
rect 156380 5652 156386 5704
rect 157334 5652 157340 5704
rect 157392 5692 157398 5704
rect 157613 5695 157671 5701
rect 157613 5692 157625 5695
rect 157392 5664 157625 5692
rect 157392 5652 157398 5664
rect 157613 5661 157625 5664
rect 157659 5661 157671 5695
rect 157613 5655 157671 5661
rect 158070 5652 158076 5704
rect 158128 5692 158134 5704
rect 158165 5695 158223 5701
rect 158165 5692 158177 5695
rect 158128 5664 158177 5692
rect 158128 5652 158134 5664
rect 158165 5661 158177 5664
rect 158211 5692 158223 5695
rect 158625 5695 158683 5701
rect 158625 5692 158637 5695
rect 158211 5664 158637 5692
rect 158211 5661 158223 5664
rect 158165 5655 158223 5661
rect 158625 5661 158637 5664
rect 158671 5661 158683 5695
rect 159174 5692 159180 5704
rect 159135 5664 159180 5692
rect 158625 5655 158683 5661
rect 159174 5652 159180 5664
rect 159232 5692 159238 5704
rect 159637 5695 159695 5701
rect 159637 5692 159649 5695
rect 159232 5664 159649 5692
rect 159232 5652 159238 5664
rect 159637 5661 159649 5664
rect 159683 5661 159695 5695
rect 165062 5692 165068 5704
rect 165023 5664 165068 5692
rect 159637 5655 159695 5661
rect 165062 5652 165068 5664
rect 165120 5692 165126 5704
rect 165433 5695 165491 5701
rect 165433 5692 165445 5695
rect 165120 5664 165445 5692
rect 165120 5652 165126 5664
rect 165433 5661 165445 5664
rect 165479 5661 165491 5695
rect 165433 5655 165491 5661
rect 155313 5559 155371 5565
rect 155313 5525 155325 5559
rect 155359 5556 155371 5559
rect 155770 5556 155776 5568
rect 155359 5528 155776 5556
rect 155359 5525 155371 5528
rect 155313 5519 155371 5525
rect 155770 5516 155776 5528
rect 155828 5516 155834 5568
rect 164970 5516 164976 5568
rect 165028 5556 165034 5568
rect 165801 5559 165859 5565
rect 165801 5556 165813 5559
rect 165028 5528 165813 5556
rect 165028 5516 165034 5528
rect 165801 5525 165813 5528
rect 165847 5525 165859 5559
rect 165801 5519 165859 5525
rect 99484 5460 101996 5488
rect 99377 5451 99435 5457
rect 99208 5392 100156 5420
rect 92992 5324 93072 5352
rect 92992 5312 92998 5324
rect 18874 5284 18880 5296
rect 6512 5256 14504 5284
rect 18432 5256 18880 5284
rect 6512 5244 6518 5256
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3292 5188 3433 5216
rect 3292 5176 3298 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5350 5216 5356 5228
rect 5031 5188 5356 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 16022 5176 16028 5228
rect 16080 5216 16086 5228
rect 16209 5219 16267 5225
rect 16209 5216 16221 5219
rect 16080 5188 16221 5216
rect 16080 5176 16086 5188
rect 16209 5185 16221 5188
rect 16255 5216 16267 5219
rect 18046 5216 18052 5228
rect 16255 5188 18052 5216
rect 16255 5185 16267 5188
rect 16209 5179 16267 5185
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 18432 5225 18460 5256
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 20257 5287 20315 5293
rect 20257 5253 20269 5287
rect 20303 5284 20315 5287
rect 21266 5284 21272 5296
rect 20303 5256 21272 5284
rect 20303 5253 20315 5256
rect 20257 5247 20315 5253
rect 21266 5244 21272 5256
rect 21324 5244 21330 5296
rect 23290 5244 23296 5296
rect 23348 5284 23354 5296
rect 26237 5287 26295 5293
rect 23348 5256 26188 5284
rect 23348 5244 23354 5256
rect 18417 5219 18475 5225
rect 18417 5185 18429 5219
rect 18463 5185 18475 5219
rect 21450 5216 21456 5228
rect 21411 5188 21456 5216
rect 18417 5179 18475 5185
rect 21450 5176 21456 5188
rect 21508 5176 21514 5228
rect 24489 5219 24547 5225
rect 24489 5185 24501 5219
rect 24535 5216 24547 5219
rect 26160 5216 26188 5256
rect 26237 5253 26249 5287
rect 26283 5284 26295 5287
rect 26418 5284 26424 5296
rect 26283 5256 26424 5284
rect 26283 5253 26295 5256
rect 26237 5247 26295 5253
rect 26418 5244 26424 5256
rect 26476 5244 26482 5296
rect 34422 5244 34428 5296
rect 34480 5284 34486 5296
rect 46014 5284 46020 5296
rect 34480 5256 46020 5284
rect 34480 5244 34486 5256
rect 46014 5244 46020 5256
rect 46072 5244 46078 5296
rect 46124 5256 46612 5284
rect 29178 5216 29184 5228
rect 24535 5188 24900 5216
rect 26160 5188 29184 5216
rect 24535 5185 24547 5188
rect 24489 5179 24547 5185
rect 4430 5148 4436 5160
rect 4391 5120 4436 5148
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 15010 5108 15016 5160
rect 15068 5148 15074 5160
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 15068 5120 15577 5148
rect 15068 5108 15074 5120
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 21269 5151 21327 5157
rect 21269 5148 21281 5151
rect 20772 5120 21281 5148
rect 20772 5108 20778 5120
rect 21269 5117 21281 5120
rect 21315 5117 21327 5151
rect 21269 5111 21327 5117
rect 22554 5108 22560 5160
rect 22612 5148 22618 5160
rect 22925 5151 22983 5157
rect 22925 5148 22937 5151
rect 22612 5120 22937 5148
rect 22612 5108 22618 5120
rect 22925 5117 22937 5120
rect 22971 5117 22983 5151
rect 22925 5111 22983 5117
rect 23937 5151 23995 5157
rect 23937 5117 23949 5151
rect 23983 5117 23995 5151
rect 23937 5111 23995 5117
rect 8202 5040 8208 5092
rect 8260 5080 8266 5092
rect 23952 5080 23980 5111
rect 24872 5089 24900 5188
rect 29178 5176 29184 5188
rect 29236 5176 29242 5228
rect 29270 5176 29276 5228
rect 29328 5216 29334 5228
rect 34793 5219 34851 5225
rect 29328 5188 34192 5216
rect 29328 5176 29334 5188
rect 25314 5148 25320 5160
rect 25275 5120 25320 5148
rect 25314 5108 25320 5120
rect 25372 5108 25378 5160
rect 29638 5108 29644 5160
rect 29696 5148 29702 5160
rect 34054 5148 34060 5160
rect 29696 5120 34060 5148
rect 29696 5108 29702 5120
rect 34054 5108 34060 5120
rect 34112 5108 34118 5160
rect 34164 5148 34192 5188
rect 34793 5185 34805 5219
rect 34839 5216 34851 5219
rect 34882 5216 34888 5228
rect 34839 5188 34888 5216
rect 34839 5185 34851 5188
rect 34793 5179 34851 5185
rect 34882 5176 34888 5188
rect 34940 5176 34946 5228
rect 34974 5176 34980 5228
rect 35032 5216 35038 5228
rect 40770 5216 40776 5228
rect 35032 5188 40776 5216
rect 35032 5176 35038 5188
rect 40770 5176 40776 5188
rect 40828 5176 40834 5228
rect 40862 5176 40868 5228
rect 40920 5216 40926 5228
rect 41322 5216 41328 5228
rect 40920 5188 41328 5216
rect 40920 5176 40926 5188
rect 41322 5176 41328 5188
rect 41380 5176 41386 5228
rect 41414 5176 41420 5228
rect 41472 5216 41478 5228
rect 43070 5216 43076 5228
rect 41472 5188 43076 5216
rect 41472 5176 41478 5188
rect 43070 5176 43076 5188
rect 43128 5176 43134 5228
rect 46124 5216 46152 5256
rect 46382 5216 46388 5228
rect 43180 5188 46152 5216
rect 46343 5188 46388 5216
rect 43180 5148 43208 5188
rect 46382 5176 46388 5188
rect 46440 5176 46446 5228
rect 46584 5216 46612 5256
rect 46658 5244 46664 5296
rect 46716 5284 46722 5296
rect 67634 5284 67640 5296
rect 46716 5256 67640 5284
rect 46716 5244 46722 5256
rect 67634 5244 67640 5256
rect 67692 5244 67698 5296
rect 89717 5287 89775 5293
rect 89717 5284 89729 5287
rect 89364 5256 89729 5284
rect 47673 5219 47731 5225
rect 47673 5216 47685 5219
rect 46584 5188 47685 5216
rect 47673 5185 47685 5188
rect 47719 5185 47731 5219
rect 47673 5179 47731 5185
rect 48038 5176 48044 5228
rect 48096 5216 48102 5228
rect 48317 5219 48375 5225
rect 48317 5216 48329 5219
rect 48096 5188 48329 5216
rect 48096 5176 48102 5188
rect 48317 5185 48329 5188
rect 48363 5216 48375 5219
rect 48498 5216 48504 5228
rect 48363 5188 48504 5216
rect 48363 5185 48375 5188
rect 48317 5179 48375 5185
rect 48498 5176 48504 5188
rect 48556 5176 48562 5228
rect 49694 5176 49700 5228
rect 49752 5216 49758 5228
rect 49881 5219 49939 5225
rect 49881 5216 49893 5219
rect 49752 5188 49893 5216
rect 49752 5176 49758 5188
rect 49881 5185 49893 5188
rect 49927 5216 49939 5219
rect 52822 5216 52828 5228
rect 49927 5188 52828 5216
rect 49927 5185 49939 5188
rect 49881 5179 49939 5185
rect 52822 5176 52828 5188
rect 52880 5176 52886 5228
rect 53650 5176 53656 5228
rect 53708 5216 53714 5228
rect 54113 5219 54171 5225
rect 54113 5216 54125 5219
rect 53708 5188 54125 5216
rect 53708 5176 53714 5188
rect 54113 5185 54125 5188
rect 54159 5216 54171 5219
rect 55398 5216 55404 5228
rect 54159 5188 55404 5216
rect 54159 5185 54171 5188
rect 54113 5179 54171 5185
rect 55398 5176 55404 5188
rect 55456 5176 55462 5228
rect 55766 5176 55772 5228
rect 55824 5216 55830 5228
rect 57054 5216 57060 5228
rect 55824 5188 57060 5216
rect 55824 5176 55830 5188
rect 57054 5176 57060 5188
rect 57112 5176 57118 5228
rect 57241 5219 57299 5225
rect 57241 5185 57253 5219
rect 57287 5216 57299 5219
rect 57330 5216 57336 5228
rect 57287 5188 57336 5216
rect 57287 5185 57299 5188
rect 57241 5179 57299 5185
rect 57330 5176 57336 5188
rect 57388 5216 57394 5228
rect 59538 5216 59544 5228
rect 57388 5188 59544 5216
rect 57388 5176 57394 5188
rect 59538 5176 59544 5188
rect 59596 5176 59602 5228
rect 63310 5176 63316 5228
rect 63368 5216 63374 5228
rect 66530 5216 66536 5228
rect 63368 5188 66536 5216
rect 63368 5176 63374 5188
rect 66530 5176 66536 5188
rect 66588 5176 66594 5228
rect 89364 5225 89392 5256
rect 89717 5253 89729 5256
rect 89763 5284 89775 5287
rect 93121 5287 93179 5293
rect 93121 5284 93133 5287
rect 89763 5256 93133 5284
rect 89763 5253 89775 5256
rect 89717 5247 89775 5253
rect 93121 5253 93133 5256
rect 93167 5253 93179 5287
rect 93121 5247 93179 5253
rect 89349 5219 89407 5225
rect 89349 5185 89361 5219
rect 89395 5185 89407 5219
rect 89349 5179 89407 5185
rect 90729 5219 90787 5225
rect 90729 5185 90741 5219
rect 90775 5216 90787 5219
rect 91094 5216 91100 5228
rect 90775 5188 91100 5216
rect 90775 5185 90787 5188
rect 90729 5179 90787 5185
rect 91094 5176 91100 5188
rect 91152 5176 91158 5228
rect 91741 5219 91799 5225
rect 91741 5185 91753 5219
rect 91787 5216 91799 5219
rect 92290 5216 92296 5228
rect 91787 5188 92296 5216
rect 91787 5185 91799 5188
rect 91741 5179 91799 5185
rect 92290 5176 92296 5188
rect 92348 5176 92354 5228
rect 34164 5120 43208 5148
rect 43346 5108 43352 5160
rect 43404 5148 43410 5160
rect 46109 5151 46167 5157
rect 46109 5148 46121 5151
rect 43404 5120 46121 5148
rect 43404 5108 43410 5120
rect 46109 5117 46121 5120
rect 46155 5117 46167 5151
rect 46109 5111 46167 5117
rect 46198 5108 46204 5160
rect 46256 5148 46262 5160
rect 49237 5151 49295 5157
rect 49237 5148 49249 5151
rect 46256 5120 49249 5148
rect 46256 5108 46262 5120
rect 49237 5117 49249 5120
rect 49283 5117 49295 5151
rect 49237 5111 49295 5117
rect 49326 5108 49332 5160
rect 49384 5148 49390 5160
rect 53469 5151 53527 5157
rect 53469 5148 53481 5151
rect 49384 5120 53481 5148
rect 49384 5108 49390 5120
rect 53469 5117 53481 5120
rect 53515 5117 53527 5151
rect 62666 5148 62672 5160
rect 53469 5111 53527 5117
rect 53576 5120 62672 5148
rect 8260 5052 23980 5080
rect 24857 5083 24915 5089
rect 8260 5040 8266 5052
rect 24857 5049 24869 5083
rect 24903 5080 24915 5083
rect 53576 5080 53604 5120
rect 62666 5108 62672 5120
rect 62724 5108 62730 5160
rect 63402 5108 63408 5160
rect 63460 5148 63466 5160
rect 70486 5148 70492 5160
rect 63460 5120 70492 5148
rect 63460 5108 63466 5120
rect 70486 5108 70492 5120
rect 70544 5108 70550 5160
rect 86770 5148 86776 5160
rect 86731 5120 86776 5148
rect 86770 5108 86776 5120
rect 86828 5108 86834 5160
rect 87782 5148 87788 5160
rect 87743 5120 87788 5148
rect 87782 5108 87788 5120
rect 87840 5108 87846 5160
rect 89257 5151 89315 5157
rect 89257 5117 89269 5151
rect 89303 5148 89315 5151
rect 89438 5148 89444 5160
rect 89303 5120 89444 5148
rect 89303 5117 89315 5120
rect 89257 5111 89315 5117
rect 89438 5108 89444 5120
rect 89496 5108 89502 5160
rect 90818 5148 90824 5160
rect 90779 5120 90824 5148
rect 90818 5108 90824 5120
rect 90876 5108 90882 5160
rect 24903 5052 53604 5080
rect 53668 5052 57008 5080
rect 24903 5049 24915 5052
rect 24857 5043 24915 5049
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 23382 4972 23388 5024
rect 23440 5012 23446 5024
rect 31570 5012 31576 5024
rect 23440 4984 31576 5012
rect 23440 4972 23446 4984
rect 31570 4972 31576 4984
rect 31628 4972 31634 5024
rect 31662 4972 31668 5024
rect 31720 5012 31726 5024
rect 34425 5015 34483 5021
rect 34425 5012 34437 5015
rect 31720 4984 34437 5012
rect 31720 4972 31726 4984
rect 34425 4981 34437 4984
rect 34471 4981 34483 5015
rect 34425 4975 34483 4981
rect 35066 4972 35072 5024
rect 35124 5012 35130 5024
rect 36446 5012 36452 5024
rect 35124 4984 36452 5012
rect 35124 4972 35130 4984
rect 36446 4972 36452 4984
rect 36504 4972 36510 5024
rect 36538 4972 36544 5024
rect 36596 5012 36602 5024
rect 43346 5012 43352 5024
rect 36596 4984 43352 5012
rect 36596 4972 36602 4984
rect 43346 4972 43352 4984
rect 43404 4972 43410 5024
rect 43530 4972 43536 5024
rect 43588 5012 43594 5024
rect 50982 5012 50988 5024
rect 43588 4984 50988 5012
rect 43588 4972 43594 4984
rect 50982 4972 50988 4984
rect 51040 4972 51046 5024
rect 51258 4972 51264 5024
rect 51316 5012 51322 5024
rect 53668 5012 53696 5052
rect 51316 4984 53696 5012
rect 51316 4972 51322 4984
rect 53742 4972 53748 5024
rect 53800 5012 53806 5024
rect 56042 5012 56048 5024
rect 53800 4984 56048 5012
rect 53800 4972 53806 4984
rect 56042 4972 56048 4984
rect 56100 4972 56106 5024
rect 56318 4972 56324 5024
rect 56376 5012 56382 5024
rect 56873 5015 56931 5021
rect 56873 5012 56885 5015
rect 56376 4984 56885 5012
rect 56376 4972 56382 4984
rect 56873 4981 56885 4984
rect 56919 4981 56931 5015
rect 56980 5012 57008 5052
rect 57054 5040 57060 5092
rect 57112 5080 57118 5092
rect 57974 5080 57980 5092
rect 57112 5052 57980 5080
rect 57112 5040 57118 5052
rect 57974 5040 57980 5052
rect 58032 5040 58038 5092
rect 58986 5040 58992 5092
rect 59044 5080 59050 5092
rect 65058 5080 65064 5092
rect 59044 5052 65064 5080
rect 59044 5040 59050 5052
rect 65058 5040 65064 5052
rect 65116 5040 65122 5092
rect 90358 5040 90364 5092
rect 90416 5080 90422 5092
rect 90545 5083 90603 5089
rect 90545 5080 90557 5083
rect 90416 5052 90557 5080
rect 90416 5040 90422 5052
rect 90545 5049 90557 5052
rect 90591 5080 90603 5083
rect 94961 5083 95019 5089
rect 94961 5080 94973 5083
rect 90591 5052 94973 5080
rect 90591 5049 90603 5052
rect 90545 5043 90603 5049
rect 94961 5049 94973 5052
rect 95007 5049 95019 5083
rect 100128 5080 100156 5392
rect 101968 5352 101996 5460
rect 102028 5466 169556 5488
rect 102028 5414 113088 5466
rect 113140 5414 113152 5466
rect 113204 5414 113216 5466
rect 113268 5414 113280 5466
rect 113332 5414 169556 5466
rect 102028 5392 169556 5414
rect 102134 5352 102140 5364
rect 101968 5324 102140 5352
rect 102134 5312 102140 5324
rect 102192 5312 102198 5364
rect 105909 5355 105967 5361
rect 105909 5352 105921 5355
rect 102244 5324 105921 5352
rect 100754 5176 100760 5228
rect 100812 5216 100818 5228
rect 102244 5216 102272 5324
rect 105909 5321 105921 5324
rect 105955 5321 105967 5355
rect 105909 5315 105967 5321
rect 106016 5324 106228 5352
rect 106016 5284 106044 5324
rect 100812 5188 102272 5216
rect 102520 5256 106044 5284
rect 106200 5284 106228 5324
rect 106458 5312 106464 5364
rect 106516 5352 106522 5364
rect 121914 5352 121920 5364
rect 106516 5324 121920 5352
rect 106516 5312 106522 5324
rect 121914 5312 121920 5324
rect 121972 5312 121978 5364
rect 127618 5312 127624 5364
rect 127676 5352 127682 5364
rect 127805 5355 127863 5361
rect 127805 5352 127817 5355
rect 127676 5324 127817 5352
rect 127676 5312 127682 5324
rect 127805 5321 127817 5324
rect 127851 5321 127863 5355
rect 145834 5352 145840 5364
rect 145795 5324 145840 5352
rect 127805 5315 127863 5321
rect 145834 5312 145840 5324
rect 145892 5312 145898 5364
rect 164697 5355 164755 5361
rect 164697 5321 164709 5355
rect 164743 5352 164755 5355
rect 166902 5352 166908 5364
rect 164743 5324 166908 5352
rect 164743 5321 164755 5324
rect 164697 5315 164755 5321
rect 166902 5312 166908 5324
rect 166960 5312 166966 5364
rect 109770 5284 109776 5296
rect 106200 5256 109776 5284
rect 100812 5176 100818 5188
rect 100205 5151 100263 5157
rect 100205 5117 100217 5151
rect 100251 5148 100263 5151
rect 102520 5148 102548 5256
rect 109770 5244 109776 5256
rect 109828 5244 109834 5296
rect 112898 5284 112904 5296
rect 110064 5256 112904 5284
rect 104434 5176 104440 5228
rect 104492 5216 104498 5228
rect 104621 5219 104679 5225
rect 104621 5216 104633 5219
rect 104492 5188 104633 5216
rect 104492 5176 104498 5188
rect 104621 5185 104633 5188
rect 104667 5216 104679 5219
rect 105630 5216 105636 5228
rect 104667 5188 105636 5216
rect 104667 5185 104679 5188
rect 104621 5179 104679 5185
rect 105630 5176 105636 5188
rect 105688 5176 105694 5228
rect 105814 5216 105820 5228
rect 105775 5188 105820 5216
rect 105814 5176 105820 5188
rect 105872 5176 105878 5228
rect 106182 5176 106188 5228
rect 106240 5216 106246 5228
rect 107930 5216 107936 5228
rect 106240 5188 107936 5216
rect 106240 5176 106246 5188
rect 107930 5176 107936 5188
rect 107988 5176 107994 5228
rect 103054 5148 103060 5160
rect 100251 5120 102548 5148
rect 103015 5120 103060 5148
rect 100251 5117 100263 5120
rect 100205 5111 100263 5117
rect 103054 5108 103060 5120
rect 103112 5108 103118 5160
rect 104066 5148 104072 5160
rect 104027 5120 104072 5148
rect 104066 5108 104072 5120
rect 104124 5108 104130 5160
rect 105998 5108 106004 5160
rect 106056 5148 106062 5160
rect 110064 5148 110092 5256
rect 112898 5244 112904 5256
rect 112956 5244 112962 5296
rect 110230 5216 110236 5228
rect 110191 5188 110236 5216
rect 110230 5176 110236 5188
rect 110288 5176 110294 5228
rect 115293 5219 115351 5225
rect 115293 5185 115305 5219
rect 115339 5216 115351 5219
rect 115382 5216 115388 5228
rect 115339 5188 115388 5216
rect 115339 5185 115351 5188
rect 115293 5179 115351 5185
rect 115382 5176 115388 5188
rect 115440 5176 115446 5228
rect 117130 5176 117136 5228
rect 117188 5216 117194 5228
rect 124674 5216 124680 5228
rect 117188 5188 124680 5216
rect 117188 5176 117194 5188
rect 124674 5176 124680 5188
rect 124732 5176 124738 5228
rect 127713 5219 127771 5225
rect 127713 5185 127725 5219
rect 127759 5216 127771 5219
rect 128354 5216 128360 5228
rect 127759 5188 128360 5216
rect 127759 5185 127771 5188
rect 127713 5179 127771 5185
rect 128354 5176 128360 5188
rect 128412 5176 128418 5228
rect 145745 5219 145803 5225
rect 145745 5185 145757 5219
rect 145791 5216 145803 5219
rect 146294 5216 146300 5228
rect 145791 5188 146300 5216
rect 145791 5185 145803 5188
rect 145745 5179 145803 5185
rect 146294 5176 146300 5188
rect 146352 5176 146358 5228
rect 151998 5176 152004 5228
rect 152056 5216 152062 5228
rect 152918 5216 152924 5228
rect 152056 5188 152924 5216
rect 152056 5176 152062 5188
rect 152918 5176 152924 5188
rect 152976 5176 152982 5228
rect 154485 5219 154543 5225
rect 154485 5185 154497 5219
rect 154531 5216 154543 5219
rect 154850 5216 154856 5228
rect 154531 5188 154856 5216
rect 154531 5185 154543 5188
rect 154485 5179 154543 5185
rect 154850 5176 154856 5188
rect 154908 5176 154914 5228
rect 156598 5216 156604 5228
rect 156559 5188 156604 5216
rect 156598 5176 156604 5188
rect 156656 5176 156662 5228
rect 158254 5216 158260 5228
rect 158215 5188 158260 5216
rect 158254 5176 158260 5188
rect 158312 5176 158318 5228
rect 159542 5216 159548 5228
rect 159503 5188 159548 5216
rect 159542 5176 159548 5188
rect 159600 5176 159606 5228
rect 164605 5219 164663 5225
rect 164605 5185 164617 5219
rect 164651 5216 164663 5219
rect 164694 5216 164700 5228
rect 164651 5188 164700 5216
rect 164651 5185 164663 5188
rect 164605 5179 164663 5185
rect 164694 5176 164700 5188
rect 164752 5176 164758 5228
rect 110322 5148 110328 5160
rect 106056 5120 110092 5148
rect 110283 5120 110328 5148
rect 106056 5108 106062 5120
rect 110322 5108 110328 5120
rect 110380 5108 110386 5160
rect 153930 5148 153936 5160
rect 153891 5120 153936 5148
rect 153930 5108 153936 5120
rect 153988 5108 153994 5160
rect 155310 5148 155316 5160
rect 155271 5120 155316 5148
rect 155310 5108 155316 5120
rect 155368 5108 155374 5160
rect 156506 5148 156512 5160
rect 156467 5120 156512 5148
rect 156506 5108 156512 5120
rect 156564 5108 156570 5160
rect 158806 5108 158812 5160
rect 158864 5148 158870 5160
rect 159269 5151 159327 5157
rect 159269 5148 159281 5151
rect 158864 5120 159281 5148
rect 158864 5108 158870 5120
rect 159269 5117 159281 5120
rect 159315 5117 159327 5151
rect 159269 5111 159327 5117
rect 103790 5080 103796 5092
rect 100128 5052 103796 5080
rect 94961 5043 95019 5049
rect 103790 5040 103796 5052
rect 103848 5040 103854 5092
rect 106090 5040 106096 5092
rect 106148 5080 106154 5092
rect 110414 5080 110420 5092
rect 106148 5052 110420 5080
rect 106148 5040 106154 5052
rect 110414 5040 110420 5052
rect 110472 5040 110478 5092
rect 115290 5040 115296 5092
rect 115348 5080 115354 5092
rect 115385 5083 115443 5089
rect 115385 5080 115397 5083
rect 115348 5052 115397 5080
rect 115348 5040 115354 5052
rect 115385 5049 115397 5052
rect 115431 5049 115443 5083
rect 115385 5043 115443 5049
rect 62482 5012 62488 5024
rect 56980 4984 62488 5012
rect 56873 4975 56931 4981
rect 62482 4972 62488 4984
rect 62540 4972 62546 5024
rect 64414 4972 64420 5024
rect 64472 5012 64478 5024
rect 70670 5012 70676 5024
rect 64472 4984 70676 5012
rect 64472 4972 64478 4984
rect 70670 4972 70676 4984
rect 70728 4972 70734 5024
rect 91830 5012 91836 5024
rect 91791 4984 91836 5012
rect 91830 4972 91836 4984
rect 91888 4972 91894 5024
rect 106182 4972 106188 5024
rect 106240 5012 106246 5024
rect 116210 5012 116216 5024
rect 106240 4984 116216 5012
rect 106240 4972 106246 4984
rect 116210 4972 116216 4984
rect 116268 4972 116274 5024
rect 368 4922 93012 4944
rect 368 4870 28456 4922
rect 28508 4870 28520 4922
rect 28572 4870 28584 4922
rect 28636 4870 28648 4922
rect 28700 4870 84878 4922
rect 84930 4870 84942 4922
rect 84994 4870 85006 4922
rect 85058 4870 85070 4922
rect 85122 4870 93012 4922
rect 368 4848 93012 4870
rect 102028 4922 169556 4944
rect 102028 4870 141299 4922
rect 141351 4870 141363 4922
rect 141415 4870 141427 4922
rect 141479 4870 141491 4922
rect 141543 4870 169556 4922
rect 102028 4848 169556 4870
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 3513 4811 3571 4817
rect 3513 4808 3525 4811
rect 3292 4780 3525 4808
rect 3292 4768 3298 4780
rect 3513 4777 3525 4780
rect 3559 4777 3571 4811
rect 3513 4771 3571 4777
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 7374 4808 7380 4820
rect 3752 4780 7380 4808
rect 3752 4768 3758 4780
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 16022 4808 16028 4820
rect 15983 4780 16028 4808
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 17313 4811 17371 4817
rect 17313 4777 17325 4811
rect 17359 4808 17371 4811
rect 17402 4808 17408 4820
rect 17359 4780 17408 4808
rect 17359 4777 17371 4780
rect 17313 4771 17371 4777
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4212 4644 4997 4672
rect 4212 4632 4218 4644
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 4985 4635 5043 4641
rect 3970 4604 3976 4616
rect 3931 4576 3976 4604
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 17328 4604 17356 4771
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 21450 4768 21456 4820
rect 21508 4808 21514 4820
rect 21637 4811 21695 4817
rect 21637 4808 21649 4811
rect 21508 4780 21649 4808
rect 21508 4768 21514 4780
rect 21637 4777 21649 4780
rect 21683 4777 21695 4811
rect 22554 4808 22560 4820
rect 21637 4771 21695 4777
rect 22020 4780 22560 4808
rect 20993 4675 21051 4681
rect 20993 4641 21005 4675
rect 21039 4672 21051 4675
rect 21358 4672 21364 4684
rect 21039 4644 21364 4672
rect 21039 4641 21051 4644
rect 20993 4635 21051 4641
rect 21358 4632 21364 4644
rect 21416 4632 21422 4684
rect 22020 4681 22048 4780
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 22925 4811 22983 4817
rect 22925 4777 22937 4811
rect 22971 4808 22983 4811
rect 25314 4808 25320 4820
rect 22971 4780 25320 4808
rect 22971 4777 22983 4780
rect 22925 4771 22983 4777
rect 23032 4681 23060 4780
rect 25314 4768 25320 4780
rect 25372 4768 25378 4820
rect 26605 4811 26663 4817
rect 26605 4777 26617 4811
rect 26651 4808 26663 4811
rect 26881 4811 26939 4817
rect 26881 4808 26893 4811
rect 26651 4780 26893 4808
rect 26651 4777 26663 4780
rect 26605 4771 26663 4777
rect 26881 4777 26893 4780
rect 26927 4808 26939 4811
rect 27890 4808 27896 4820
rect 26927 4780 27896 4808
rect 26927 4777 26939 4780
rect 26881 4771 26939 4777
rect 27890 4768 27896 4780
rect 27948 4768 27954 4820
rect 29730 4768 29736 4820
rect 29788 4808 29794 4820
rect 36538 4808 36544 4820
rect 29788 4780 36544 4808
rect 29788 4768 29794 4780
rect 36538 4768 36544 4780
rect 36596 4768 36602 4820
rect 36832 4780 46336 4808
rect 36832 4752 36860 4780
rect 26142 4700 26148 4752
rect 26200 4740 26206 4752
rect 30374 4740 30380 4752
rect 26200 4712 30380 4740
rect 26200 4700 26206 4712
rect 30374 4700 30380 4712
rect 30432 4700 30438 4752
rect 30561 4743 30619 4749
rect 30561 4709 30573 4743
rect 30607 4740 30619 4743
rect 33137 4743 33195 4749
rect 33137 4740 33149 4743
rect 30607 4712 33149 4740
rect 30607 4709 30619 4712
rect 30561 4703 30619 4709
rect 33137 4709 33149 4712
rect 33183 4709 33195 4743
rect 33137 4703 33195 4709
rect 33229 4743 33287 4749
rect 33229 4709 33241 4743
rect 33275 4740 33287 4743
rect 33413 4743 33471 4749
rect 33413 4740 33425 4743
rect 33275 4712 33425 4740
rect 33275 4709 33287 4712
rect 33229 4703 33287 4709
rect 33413 4709 33425 4712
rect 33459 4740 33471 4743
rect 34514 4740 34520 4752
rect 33459 4712 34520 4740
rect 33459 4709 33471 4712
rect 33413 4703 33471 4709
rect 22005 4675 22063 4681
rect 22005 4641 22017 4675
rect 22051 4641 22063 4675
rect 22005 4635 22063 4641
rect 23017 4675 23075 4681
rect 23017 4641 23029 4675
rect 23063 4641 23075 4675
rect 23017 4635 23075 4641
rect 24029 4675 24087 4681
rect 24029 4641 24041 4675
rect 24075 4641 24087 4675
rect 25777 4675 25835 4681
rect 25777 4672 25789 4675
rect 24029 4635 24087 4641
rect 24136 4644 25789 4672
rect 17954 4604 17960 4616
rect 16899 4576 17356 4604
rect 17915 4576 17960 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 5552 4536 5580 4567
rect 17954 4564 17960 4576
rect 18012 4604 18018 4616
rect 18785 4607 18843 4613
rect 18785 4604 18797 4607
rect 18012 4576 18797 4604
rect 18012 4564 18018 4576
rect 18785 4573 18797 4576
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 5902 4536 5908 4548
rect 5552 4508 5908 4536
rect 5902 4496 5908 4508
rect 5960 4496 5966 4548
rect 12250 4496 12256 4548
rect 12308 4536 12314 4548
rect 24044 4536 24072 4635
rect 12308 4508 24072 4536
rect 12308 4496 12314 4508
rect 3878 4428 3884 4480
rect 3936 4468 3942 4480
rect 5810 4468 5816 4480
rect 3936 4440 5816 4468
rect 3936 4428 3942 4440
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 7193 4471 7251 4477
rect 7193 4437 7205 4471
rect 7239 4468 7251 4471
rect 8478 4468 8484 4480
rect 7239 4440 8484 4468
rect 7239 4437 7251 4440
rect 7193 4431 7251 4437
rect 8478 4428 8484 4440
rect 8536 4428 8542 4480
rect 16666 4468 16672 4480
rect 16627 4440 16672 4468
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18049 4471 18107 4477
rect 18049 4468 18061 4471
rect 18012 4440 18061 4468
rect 18012 4428 18018 4440
rect 18049 4437 18061 4440
rect 18095 4437 18107 4471
rect 18049 4431 18107 4437
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 24136 4468 24164 4644
rect 25777 4641 25789 4644
rect 25823 4641 25835 4675
rect 25777 4635 25835 4641
rect 26970 4632 26976 4684
rect 27028 4672 27034 4684
rect 30466 4672 30472 4684
rect 27028 4644 30472 4672
rect 27028 4632 27034 4644
rect 30466 4632 30472 4644
rect 30524 4632 30530 4684
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 26329 4607 26387 4613
rect 24627 4576 24992 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 24964 4480 24992 4576
rect 26329 4573 26341 4607
rect 26375 4604 26387 4607
rect 26605 4607 26663 4613
rect 26605 4604 26617 4607
rect 26375 4576 26617 4604
rect 26375 4573 26387 4576
rect 26329 4567 26387 4573
rect 26605 4573 26617 4576
rect 26651 4573 26663 4607
rect 26605 4567 26663 4573
rect 28166 4564 28172 4616
rect 28224 4604 28230 4616
rect 30101 4607 30159 4613
rect 28224 4576 30052 4604
rect 28224 4564 28230 4576
rect 26418 4496 26424 4548
rect 26476 4536 26482 4548
rect 29457 4539 29515 4545
rect 29457 4536 29469 4539
rect 26476 4508 29469 4536
rect 26476 4496 26482 4508
rect 29457 4505 29469 4508
rect 29503 4505 29515 4539
rect 30024 4536 30052 4576
rect 30101 4573 30113 4607
rect 30147 4604 30159 4607
rect 30576 4604 30604 4703
rect 34514 4700 34520 4712
rect 34572 4700 34578 4752
rect 34609 4743 34667 4749
rect 34609 4709 34621 4743
rect 34655 4740 34667 4743
rect 34882 4740 34888 4752
rect 34655 4712 34888 4740
rect 34655 4709 34667 4712
rect 34609 4703 34667 4709
rect 34882 4700 34888 4712
rect 34940 4700 34946 4752
rect 35158 4700 35164 4752
rect 35216 4740 35222 4752
rect 36446 4740 36452 4752
rect 35216 4712 36452 4740
rect 35216 4700 35222 4712
rect 36446 4700 36452 4712
rect 36504 4700 36510 4752
rect 36556 4712 36768 4740
rect 36556 4672 36584 4712
rect 30147 4576 30604 4604
rect 30668 4644 36584 4672
rect 36740 4672 36768 4712
rect 36814 4700 36820 4752
rect 36872 4700 36878 4752
rect 36998 4700 37004 4752
rect 37056 4740 37062 4752
rect 38930 4740 38936 4752
rect 37056 4712 38936 4740
rect 37056 4700 37062 4712
rect 38930 4700 38936 4712
rect 38988 4700 38994 4752
rect 39206 4700 39212 4752
rect 39264 4740 39270 4752
rect 46198 4740 46204 4752
rect 39264 4712 46204 4740
rect 39264 4700 39270 4712
rect 46198 4700 46204 4712
rect 46256 4700 46262 4752
rect 46308 4740 46336 4780
rect 46382 4768 46388 4820
rect 46440 4808 46446 4820
rect 49513 4811 49571 4817
rect 49513 4808 49525 4811
rect 46440 4780 49525 4808
rect 46440 4768 46446 4780
rect 49513 4777 49525 4780
rect 49559 4777 49571 4811
rect 49694 4808 49700 4820
rect 49655 4780 49700 4808
rect 49513 4771 49571 4777
rect 49694 4768 49700 4780
rect 49752 4768 49758 4820
rect 50062 4768 50068 4820
rect 50120 4808 50126 4820
rect 50120 4780 50476 4808
rect 50120 4768 50126 4780
rect 49326 4740 49332 4752
rect 46308 4712 49332 4740
rect 49326 4700 49332 4712
rect 49384 4700 49390 4752
rect 50448 4740 50476 4780
rect 50522 4768 50528 4820
rect 50580 4808 50586 4820
rect 52822 4808 52828 4820
rect 50580 4780 52828 4808
rect 50580 4768 50586 4780
rect 52822 4768 52828 4780
rect 52880 4768 52886 4820
rect 53650 4808 53656 4820
rect 53611 4780 53656 4808
rect 53650 4768 53656 4780
rect 53708 4768 53714 4820
rect 54665 4811 54723 4817
rect 54665 4777 54677 4811
rect 54711 4808 54723 4811
rect 54941 4811 54999 4817
rect 54941 4808 54953 4811
rect 54711 4780 54953 4808
rect 54711 4777 54723 4780
rect 54665 4771 54723 4777
rect 54941 4777 54953 4780
rect 54987 4808 54999 4811
rect 55214 4808 55220 4820
rect 54987 4780 55220 4808
rect 54987 4777 54999 4780
rect 54941 4771 54999 4777
rect 55214 4768 55220 4780
rect 55272 4768 55278 4820
rect 55490 4768 55496 4820
rect 55548 4808 55554 4820
rect 57422 4808 57428 4820
rect 55548 4780 57428 4808
rect 55548 4768 55554 4780
rect 57422 4768 57428 4780
rect 57480 4768 57486 4820
rect 57606 4768 57612 4820
rect 57664 4808 57670 4820
rect 81618 4808 81624 4820
rect 57664 4780 81624 4808
rect 57664 4768 57670 4780
rect 81618 4768 81624 4780
rect 81676 4768 81682 4820
rect 86770 4768 86776 4820
rect 86828 4808 86834 4820
rect 88613 4811 88671 4817
rect 88613 4808 88625 4811
rect 86828 4780 88625 4808
rect 86828 4768 86834 4780
rect 88613 4777 88625 4780
rect 88659 4808 88671 4811
rect 91833 4811 91891 4817
rect 88659 4780 88840 4808
rect 88659 4777 88671 4780
rect 88613 4771 88671 4777
rect 55953 4743 56011 4749
rect 55953 4740 55965 4743
rect 50448 4712 55965 4740
rect 55953 4709 55965 4712
rect 55999 4709 56011 4743
rect 55953 4703 56011 4709
rect 56781 4743 56839 4749
rect 56781 4709 56793 4743
rect 56827 4740 56839 4743
rect 56962 4740 56968 4752
rect 56827 4712 56968 4740
rect 56827 4709 56839 4712
rect 56781 4703 56839 4709
rect 56962 4700 56968 4712
rect 57020 4700 57026 4752
rect 57149 4743 57207 4749
rect 57149 4709 57161 4743
rect 57195 4740 57207 4743
rect 57330 4740 57336 4752
rect 57195 4712 57336 4740
rect 57195 4709 57207 4712
rect 57149 4703 57207 4709
rect 57330 4700 57336 4712
rect 57388 4700 57394 4752
rect 60458 4700 60464 4752
rect 60516 4740 60522 4752
rect 60734 4740 60740 4752
rect 60516 4712 60740 4740
rect 60516 4700 60522 4712
rect 60734 4700 60740 4712
rect 60792 4700 60798 4752
rect 39761 4675 39819 4681
rect 39761 4672 39773 4675
rect 36740 4644 39773 4672
rect 30147 4573 30159 4576
rect 30101 4567 30159 4573
rect 30668 4536 30696 4644
rect 39761 4641 39773 4644
rect 39807 4641 39819 4675
rect 39761 4635 39819 4641
rect 39850 4632 39856 4684
rect 39908 4672 39914 4684
rect 41506 4672 41512 4684
rect 39908 4644 41512 4672
rect 39908 4632 39914 4644
rect 41506 4632 41512 4644
rect 41564 4632 41570 4684
rect 41598 4632 41604 4684
rect 41656 4672 41662 4684
rect 45646 4672 45652 4684
rect 41656 4644 45652 4672
rect 41656 4632 41662 4644
rect 45646 4632 45652 4644
rect 45704 4632 45710 4684
rect 45756 4644 46060 4672
rect 30742 4564 30748 4616
rect 30800 4604 30806 4616
rect 31478 4604 31484 4616
rect 30800 4576 31484 4604
rect 30800 4564 30806 4576
rect 31478 4564 31484 4576
rect 31536 4564 31542 4616
rect 32953 4607 33011 4613
rect 31588 4576 32628 4604
rect 30024 4508 30696 4536
rect 29457 4499 29515 4505
rect 30834 4496 30840 4548
rect 30892 4536 30898 4548
rect 31588 4536 31616 4576
rect 30892 4508 31616 4536
rect 30892 4496 30898 4508
rect 31846 4496 31852 4548
rect 31904 4536 31910 4548
rect 32309 4539 32367 4545
rect 32309 4536 32321 4539
rect 31904 4508 32321 4536
rect 31904 4496 31910 4508
rect 32309 4505 32321 4508
rect 32355 4505 32367 4539
rect 32309 4499 32367 4505
rect 24946 4468 24952 4480
rect 22336 4440 24164 4468
rect 24907 4440 24952 4468
rect 22336 4428 22342 4440
rect 24946 4428 24952 4440
rect 25004 4428 25010 4480
rect 25038 4428 25044 4480
rect 25096 4468 25102 4480
rect 32490 4468 32496 4480
rect 25096 4440 32496 4468
rect 25096 4428 25102 4440
rect 32490 4428 32496 4440
rect 32548 4428 32554 4480
rect 32600 4468 32628 4576
rect 32953 4573 32965 4607
rect 32999 4604 33011 4607
rect 33229 4607 33287 4613
rect 33229 4604 33241 4607
rect 32999 4576 33241 4604
rect 32999 4573 33011 4576
rect 32953 4567 33011 4573
rect 33229 4573 33241 4576
rect 33275 4573 33287 4607
rect 33229 4567 33287 4573
rect 34422 4564 34428 4616
rect 34480 4604 34486 4616
rect 36814 4604 36820 4616
rect 34480 4576 36820 4604
rect 34480 4564 34486 4576
rect 36814 4564 36820 4576
rect 36872 4564 36878 4616
rect 36906 4564 36912 4616
rect 36964 4604 36970 4616
rect 40034 4604 40040 4616
rect 36964 4576 40040 4604
rect 36964 4564 36970 4576
rect 40034 4564 40040 4576
rect 40092 4564 40098 4616
rect 40218 4604 40224 4616
rect 40179 4576 40224 4604
rect 40218 4564 40224 4576
rect 40276 4604 40282 4616
rect 40773 4607 40831 4613
rect 40773 4604 40785 4607
rect 40276 4576 40785 4604
rect 40276 4564 40282 4576
rect 40773 4573 40785 4576
rect 40819 4573 40831 4607
rect 40773 4567 40831 4573
rect 40862 4564 40868 4616
rect 40920 4604 40926 4616
rect 45554 4604 45560 4616
rect 40920 4576 45560 4604
rect 40920 4564 40926 4576
rect 45554 4564 45560 4576
rect 45612 4564 45618 4616
rect 33137 4539 33195 4545
rect 33137 4505 33149 4539
rect 33183 4536 33195 4539
rect 36630 4536 36636 4548
rect 33183 4508 36636 4536
rect 33183 4505 33195 4508
rect 33137 4499 33195 4505
rect 36630 4496 36636 4508
rect 36688 4496 36694 4548
rect 36722 4496 36728 4548
rect 36780 4536 36786 4548
rect 41414 4536 41420 4548
rect 36780 4508 41420 4536
rect 36780 4496 36786 4508
rect 41414 4496 41420 4508
rect 41472 4496 41478 4548
rect 41506 4496 41512 4548
rect 41564 4536 41570 4548
rect 44910 4536 44916 4548
rect 41564 4508 44916 4536
rect 41564 4496 41570 4508
rect 44910 4496 44916 4508
rect 44968 4496 44974 4548
rect 45186 4496 45192 4548
rect 45244 4536 45250 4548
rect 45756 4536 45784 4644
rect 45244 4508 45784 4536
rect 45244 4496 45250 4508
rect 33962 4468 33968 4480
rect 32600 4440 33968 4468
rect 33962 4428 33968 4440
rect 34020 4428 34026 4480
rect 34054 4428 34060 4480
rect 34112 4468 34118 4480
rect 45738 4468 45744 4480
rect 34112 4440 45744 4468
rect 34112 4428 34118 4440
rect 45738 4428 45744 4440
rect 45796 4428 45802 4480
rect 46032 4468 46060 4644
rect 46106 4632 46112 4684
rect 46164 4672 46170 4684
rect 46382 4672 46388 4684
rect 46164 4644 46388 4672
rect 46164 4632 46170 4644
rect 46382 4632 46388 4644
rect 46440 4632 46446 4684
rect 46566 4672 46572 4684
rect 46527 4644 46572 4672
rect 46566 4632 46572 4644
rect 46624 4632 46630 4684
rect 46842 4632 46848 4684
rect 46900 4672 46906 4684
rect 47670 4672 47676 4684
rect 46900 4644 47676 4672
rect 46900 4632 46906 4644
rect 47670 4632 47676 4644
rect 47728 4632 47734 4684
rect 47857 4675 47915 4681
rect 47857 4641 47869 4675
rect 47903 4672 47915 4675
rect 56318 4672 56324 4684
rect 47903 4644 56324 4672
rect 47903 4641 47915 4644
rect 47857 4635 47915 4641
rect 56318 4632 56324 4644
rect 56376 4632 56382 4684
rect 57606 4632 57612 4684
rect 57664 4672 57670 4684
rect 63678 4672 63684 4684
rect 57664 4644 63684 4672
rect 57664 4632 57670 4644
rect 63678 4632 63684 4644
rect 63736 4632 63742 4684
rect 87782 4672 87788 4684
rect 87743 4644 87788 4672
rect 87782 4632 87788 4644
rect 87840 4672 87846 4684
rect 88812 4681 88840 4780
rect 91833 4777 91845 4811
rect 91879 4808 91891 4811
rect 92750 4808 92756 4820
rect 91879 4780 92756 4808
rect 91879 4777 91891 4780
rect 91833 4771 91891 4777
rect 92750 4768 92756 4780
rect 92808 4768 92814 4820
rect 104434 4808 104440 4820
rect 104395 4780 104440 4808
rect 104434 4768 104440 4780
rect 104492 4768 104498 4820
rect 105725 4811 105783 4817
rect 105725 4777 105737 4811
rect 105771 4808 105783 4811
rect 118878 4808 118884 4820
rect 105771 4780 118884 4808
rect 105771 4777 105783 4780
rect 105725 4771 105783 4777
rect 118878 4768 118884 4780
rect 118936 4768 118942 4820
rect 121914 4808 121920 4820
rect 121875 4780 121920 4808
rect 121914 4768 121920 4780
rect 121972 4768 121978 4820
rect 129182 4808 129188 4820
rect 129143 4780 129188 4808
rect 129182 4768 129188 4780
rect 129240 4768 129246 4820
rect 130194 4808 130200 4820
rect 130155 4780 130200 4808
rect 130194 4768 130200 4780
rect 130252 4768 130258 4820
rect 131209 4811 131267 4817
rect 131209 4777 131221 4811
rect 131255 4808 131267 4811
rect 131298 4808 131304 4820
rect 131255 4780 131304 4808
rect 131255 4777 131267 4780
rect 131209 4771 131267 4777
rect 131298 4768 131304 4780
rect 131356 4768 131362 4820
rect 146662 4768 146668 4820
rect 146720 4808 146726 4820
rect 147309 4811 147367 4817
rect 147309 4808 147321 4811
rect 146720 4780 147321 4808
rect 146720 4768 146726 4780
rect 147309 4777 147321 4780
rect 147355 4777 147367 4811
rect 150158 4808 150164 4820
rect 150119 4780 150164 4808
rect 147309 4771 147367 4777
rect 150158 4768 150164 4780
rect 150216 4768 150222 4820
rect 151722 4808 151728 4820
rect 151683 4780 151728 4808
rect 151722 4768 151728 4780
rect 151780 4768 151786 4820
rect 152918 4768 152924 4820
rect 152976 4808 152982 4820
rect 153381 4811 153439 4817
rect 153381 4808 153393 4811
rect 152976 4780 153393 4808
rect 152976 4768 152982 4780
rect 153381 4777 153393 4780
rect 153427 4777 153439 4811
rect 153381 4771 153439 4777
rect 153654 4768 153660 4820
rect 153712 4808 153718 4820
rect 154025 4811 154083 4817
rect 154025 4808 154037 4811
rect 153712 4780 154037 4808
rect 153712 4768 153718 4780
rect 154025 4777 154037 4780
rect 154071 4777 154083 4811
rect 154025 4771 154083 4777
rect 155865 4811 155923 4817
rect 155865 4777 155877 4811
rect 155911 4808 155923 4811
rect 156046 4808 156052 4820
rect 155911 4780 156052 4808
rect 155911 4777 155923 4780
rect 155865 4771 155923 4777
rect 156046 4768 156052 4780
rect 156104 4768 156110 4820
rect 156598 4808 156604 4820
rect 156559 4780 156604 4808
rect 156598 4768 156604 4780
rect 156656 4768 156662 4820
rect 158254 4808 158260 4820
rect 158215 4780 158260 4808
rect 158254 4768 158260 4780
rect 158312 4768 158318 4820
rect 163225 4811 163283 4817
rect 163225 4777 163237 4811
rect 163271 4808 163283 4811
rect 163958 4808 163964 4820
rect 163271 4780 163964 4808
rect 163271 4777 163283 4780
rect 163225 4771 163283 4777
rect 163958 4768 163964 4780
rect 164016 4768 164022 4820
rect 90269 4743 90327 4749
rect 90269 4709 90281 4743
rect 90315 4740 90327 4743
rect 90542 4740 90548 4752
rect 90315 4712 90548 4740
rect 90315 4709 90327 4712
rect 90269 4703 90327 4709
rect 90542 4700 90548 4712
rect 90600 4700 90606 4752
rect 92661 4743 92719 4749
rect 92661 4709 92673 4743
rect 92707 4740 92719 4743
rect 94869 4743 94927 4749
rect 94869 4740 94881 4743
rect 92707 4712 94881 4740
rect 92707 4709 92719 4712
rect 92661 4703 92719 4709
rect 94869 4709 94881 4712
rect 94915 4709 94927 4743
rect 94869 4703 94927 4709
rect 88245 4675 88303 4681
rect 88245 4672 88257 4675
rect 87840 4644 88257 4672
rect 87840 4632 87846 4644
rect 88245 4641 88257 4644
rect 88291 4641 88303 4675
rect 88245 4635 88303 4641
rect 88797 4675 88855 4681
rect 88797 4641 88809 4675
rect 88843 4641 88855 4675
rect 88797 4635 88855 4641
rect 46474 4564 46480 4616
rect 46532 4604 46538 4616
rect 48869 4607 48927 4613
rect 46532 4576 48360 4604
rect 46532 4564 46538 4576
rect 46198 4496 46204 4548
rect 46256 4536 46262 4548
rect 46256 4508 46612 4536
rect 46256 4496 46262 4508
rect 46474 4468 46480 4480
rect 46032 4440 46480 4468
rect 46474 4428 46480 4440
rect 46532 4428 46538 4480
rect 46584 4468 46612 4508
rect 46658 4496 46664 4548
rect 46716 4536 46722 4548
rect 47857 4539 47915 4545
rect 47857 4536 47869 4539
rect 46716 4508 47869 4536
rect 46716 4496 46722 4508
rect 47857 4505 47869 4508
rect 47903 4505 47915 4539
rect 48038 4536 48044 4548
rect 47999 4508 48044 4536
rect 47857 4499 47915 4505
rect 48038 4496 48044 4508
rect 48096 4496 48102 4548
rect 48222 4536 48228 4548
rect 48183 4508 48228 4536
rect 48222 4496 48228 4508
rect 48280 4496 48286 4548
rect 48332 4536 48360 4576
rect 48869 4573 48881 4607
rect 48915 4604 48927 4607
rect 48958 4604 48964 4616
rect 48915 4576 48964 4604
rect 48915 4573 48927 4576
rect 48869 4567 48927 4573
rect 48958 4564 48964 4576
rect 49016 4564 49022 4616
rect 49053 4607 49111 4613
rect 49053 4573 49065 4607
rect 49099 4604 49111 4607
rect 53837 4607 53895 4613
rect 53837 4604 53849 4607
rect 49099 4576 53849 4604
rect 49099 4573 49111 4576
rect 49053 4567 49111 4573
rect 53837 4573 53849 4576
rect 53883 4573 53895 4607
rect 53837 4567 53895 4573
rect 54481 4607 54539 4613
rect 54481 4573 54493 4607
rect 54527 4604 54539 4607
rect 54665 4607 54723 4613
rect 54665 4604 54677 4607
rect 54527 4576 54677 4604
rect 54527 4573 54539 4576
rect 54481 4567 54539 4573
rect 54665 4573 54677 4576
rect 54711 4573 54723 4607
rect 54665 4567 54723 4573
rect 54754 4564 54760 4616
rect 54812 4604 54818 4616
rect 55582 4604 55588 4616
rect 54812 4576 55588 4604
rect 54812 4564 54818 4576
rect 55582 4564 55588 4576
rect 55640 4564 55646 4616
rect 55766 4604 55772 4616
rect 55727 4576 55772 4604
rect 55766 4564 55772 4576
rect 55824 4564 55830 4616
rect 61286 4604 61292 4616
rect 55876 4576 61292 4604
rect 49513 4539 49571 4545
rect 48332 4508 49464 4536
rect 49053 4471 49111 4477
rect 49053 4468 49065 4471
rect 46584 4440 49065 4468
rect 49053 4437 49065 4440
rect 49099 4437 49111 4471
rect 49234 4468 49240 4480
rect 49195 4440 49240 4468
rect 49053 4431 49111 4437
rect 49234 4428 49240 4440
rect 49292 4428 49298 4480
rect 49436 4468 49464 4508
rect 49513 4505 49525 4539
rect 49559 4536 49571 4539
rect 55876 4536 55904 4576
rect 61286 4564 61292 4576
rect 61344 4564 61350 4616
rect 90358 4604 90364 4616
rect 90319 4576 90364 4604
rect 90358 4564 90364 4576
rect 90416 4564 90422 4616
rect 91741 4607 91799 4613
rect 91741 4573 91753 4607
rect 91787 4604 91799 4607
rect 92676 4604 92704 4703
rect 100386 4700 100392 4752
rect 100444 4740 100450 4752
rect 100444 4712 103468 4740
rect 100444 4700 100450 4712
rect 102873 4675 102931 4681
rect 102873 4641 102885 4675
rect 102919 4672 102931 4675
rect 103054 4672 103060 4684
rect 102919 4644 103060 4672
rect 102919 4641 102931 4644
rect 102873 4635 102931 4641
rect 103054 4632 103060 4644
rect 103112 4672 103118 4684
rect 103333 4675 103391 4681
rect 103333 4672 103345 4675
rect 103112 4644 103345 4672
rect 103112 4632 103118 4644
rect 103333 4641 103345 4644
rect 103379 4641 103391 4675
rect 103440 4672 103468 4712
rect 103790 4700 103796 4752
rect 103848 4740 103854 4752
rect 110782 4740 110788 4752
rect 103848 4712 110788 4740
rect 103848 4700 103854 4712
rect 110782 4700 110788 4712
rect 110840 4700 110846 4752
rect 107010 4672 107016 4684
rect 103440 4644 107016 4672
rect 103333 4635 103391 4641
rect 107010 4632 107016 4644
rect 107068 4632 107074 4684
rect 109586 4632 109592 4684
rect 109644 4672 109650 4684
rect 117038 4672 117044 4684
rect 109644 4644 117044 4672
rect 109644 4632 109650 4644
rect 117038 4632 117044 4644
rect 117096 4632 117102 4684
rect 150621 4675 150679 4681
rect 150621 4672 150633 4675
rect 147140 4644 147812 4672
rect 91787 4576 92704 4604
rect 91787 4573 91799 4576
rect 91741 4567 91799 4573
rect 100570 4564 100576 4616
rect 100628 4604 100634 4616
rect 110322 4604 110328 4616
rect 100628 4576 110328 4604
rect 100628 4564 100634 4576
rect 110322 4564 110328 4576
rect 110380 4564 110386 4616
rect 121825 4607 121883 4613
rect 121825 4573 121837 4607
rect 121871 4604 121883 4607
rect 129093 4607 129151 4613
rect 121871 4576 122420 4604
rect 121871 4573 121883 4576
rect 121825 4567 121883 4573
rect 57514 4536 57520 4548
rect 49559 4508 55904 4536
rect 55968 4508 57520 4536
rect 49559 4505 49571 4508
rect 49513 4499 49571 4505
rect 49970 4468 49976 4480
rect 49436 4440 49976 4468
rect 49970 4428 49976 4440
rect 50028 4428 50034 4480
rect 50614 4428 50620 4480
rect 50672 4468 50678 4480
rect 51626 4468 51632 4480
rect 50672 4440 51632 4468
rect 50672 4428 50678 4440
rect 51626 4428 51632 4440
rect 51684 4428 51690 4480
rect 52086 4428 52092 4480
rect 52144 4468 52150 4480
rect 55122 4468 55128 4480
rect 52144 4440 55128 4468
rect 52144 4428 52150 4440
rect 55122 4428 55128 4440
rect 55180 4428 55186 4480
rect 55490 4428 55496 4480
rect 55548 4468 55554 4480
rect 55968 4468 55996 4508
rect 57514 4496 57520 4508
rect 57572 4496 57578 4548
rect 60642 4496 60648 4548
rect 60700 4536 60706 4548
rect 61378 4536 61384 4548
rect 60700 4508 61384 4536
rect 60700 4496 60706 4508
rect 61378 4496 61384 4508
rect 61436 4496 61442 4548
rect 90821 4539 90879 4545
rect 90821 4505 90833 4539
rect 90867 4536 90879 4539
rect 91094 4536 91100 4548
rect 90867 4508 91100 4536
rect 90867 4505 90879 4508
rect 90821 4499 90879 4505
rect 91094 4496 91100 4508
rect 91152 4536 91158 4548
rect 92198 4536 92204 4548
rect 91152 4508 92204 4536
rect 91152 4496 91158 4508
rect 92198 4496 92204 4508
rect 92256 4496 92262 4548
rect 100021 4539 100079 4545
rect 100021 4505 100033 4539
rect 100067 4536 100079 4539
rect 113450 4536 113456 4548
rect 100067 4508 113456 4536
rect 100067 4505 100079 4508
rect 100021 4499 100079 4505
rect 113450 4496 113456 4508
rect 113508 4496 113514 4548
rect 113542 4496 113548 4548
rect 113600 4536 113606 4548
rect 117130 4536 117136 4548
rect 113600 4508 117136 4536
rect 113600 4496 113606 4508
rect 117130 4496 117136 4508
rect 117188 4496 117194 4548
rect 55548 4440 55996 4468
rect 55548 4428 55554 4440
rect 56042 4428 56048 4480
rect 56100 4468 56106 4480
rect 57606 4468 57612 4480
rect 56100 4440 57612 4468
rect 56100 4428 56106 4440
rect 57606 4428 57612 4440
rect 57664 4428 57670 4480
rect 57698 4428 57704 4480
rect 57756 4468 57762 4480
rect 66438 4468 66444 4480
rect 57756 4440 66444 4468
rect 57756 4428 57762 4440
rect 66438 4428 66444 4440
rect 66496 4428 66502 4480
rect 92290 4468 92296 4480
rect 92203 4440 92296 4468
rect 92290 4428 92296 4440
rect 92348 4468 92354 4480
rect 94958 4468 94964 4480
rect 92348 4440 94964 4468
rect 92348 4428 92354 4440
rect 94958 4428 94964 4440
rect 95016 4428 95022 4480
rect 100386 4428 100392 4480
rect 100444 4468 100450 4480
rect 105725 4471 105783 4477
rect 105725 4468 105737 4471
rect 100444 4440 105737 4468
rect 100444 4428 100450 4440
rect 105725 4437 105737 4440
rect 105771 4437 105783 4471
rect 105906 4468 105912 4480
rect 105867 4440 105912 4468
rect 105725 4431 105783 4437
rect 105906 4428 105912 4440
rect 105964 4428 105970 4480
rect 110230 4468 110236 4480
rect 110191 4440 110236 4468
rect 110230 4428 110236 4440
rect 110288 4428 110294 4480
rect 115382 4468 115388 4480
rect 115343 4440 115388 4468
rect 115382 4428 115388 4440
rect 115440 4428 115446 4480
rect 122392 4477 122420 4576
rect 129093 4573 129105 4607
rect 129139 4573 129151 4607
rect 129093 4567 129151 4573
rect 130105 4607 130163 4613
rect 130105 4573 130117 4607
rect 130151 4604 130163 4607
rect 131117 4607 131175 4613
rect 130151 4576 130700 4604
rect 130151 4573 130163 4576
rect 130105 4567 130163 4573
rect 129108 4536 129136 4567
rect 129645 4539 129703 4545
rect 129645 4536 129657 4539
rect 129108 4508 129657 4536
rect 129645 4505 129657 4508
rect 129691 4536 129703 4539
rect 130470 4536 130476 4548
rect 129691 4508 130476 4536
rect 129691 4505 129703 4508
rect 129645 4499 129703 4505
rect 130470 4496 130476 4508
rect 130528 4496 130534 4548
rect 122377 4471 122435 4477
rect 122377 4437 122389 4471
rect 122423 4468 122435 4471
rect 122742 4468 122748 4480
rect 122423 4440 122748 4468
rect 122423 4437 122435 4440
rect 122377 4431 122435 4437
rect 122742 4428 122748 4440
rect 122800 4428 122806 4480
rect 127805 4471 127863 4477
rect 127805 4437 127817 4471
rect 127851 4468 127863 4471
rect 128354 4468 128360 4480
rect 127851 4440 128360 4468
rect 127851 4437 127863 4440
rect 127805 4431 127863 4437
rect 128354 4428 128360 4440
rect 128412 4468 128418 4480
rect 129366 4468 129372 4480
rect 128412 4440 129372 4468
rect 128412 4428 128418 4440
rect 129366 4428 129372 4440
rect 129424 4428 129430 4480
rect 130672 4477 130700 4576
rect 131117 4573 131129 4607
rect 131163 4604 131175 4607
rect 147140 4604 147168 4644
rect 147209 4607 147267 4613
rect 147209 4604 147221 4607
rect 131163 4576 131712 4604
rect 147140 4576 147221 4604
rect 131163 4573 131175 4576
rect 131117 4567 131175 4573
rect 130657 4471 130715 4477
rect 130657 4437 130669 4471
rect 130703 4468 130715 4471
rect 130838 4468 130844 4480
rect 130703 4440 130844 4468
rect 130703 4437 130715 4440
rect 130657 4431 130715 4437
rect 130838 4428 130844 4440
rect 130896 4428 130902 4480
rect 131684 4477 131712 4576
rect 147209 4573 147221 4576
rect 147255 4573 147267 4607
rect 147209 4567 147267 4573
rect 145837 4539 145895 4545
rect 145837 4505 145849 4539
rect 145883 4536 145895 4539
rect 146294 4536 146300 4548
rect 145883 4508 146300 4536
rect 145883 4505 145895 4508
rect 145837 4499 145895 4505
rect 146294 4496 146300 4508
rect 146352 4536 146358 4548
rect 147398 4536 147404 4548
rect 146352 4508 147404 4536
rect 146352 4496 146358 4508
rect 147398 4496 147404 4508
rect 147456 4496 147462 4548
rect 147784 4545 147812 4644
rect 150084 4644 150633 4672
rect 150084 4613 150112 4644
rect 150621 4641 150633 4644
rect 150667 4672 150679 4675
rect 152182 4672 152188 4684
rect 150667 4644 152188 4672
rect 150667 4641 150679 4644
rect 150621 4635 150679 4641
rect 152182 4632 152188 4644
rect 152240 4632 152246 4684
rect 152921 4675 152979 4681
rect 152921 4641 152933 4675
rect 152967 4672 152979 4675
rect 155221 4675 155279 4681
rect 155221 4672 155233 4675
rect 152967 4644 155233 4672
rect 152967 4641 152979 4644
rect 152921 4635 152979 4641
rect 155221 4641 155233 4644
rect 155267 4672 155279 4675
rect 155310 4672 155316 4684
rect 155267 4644 155316 4672
rect 155267 4641 155279 4644
rect 155221 4635 155279 4641
rect 155310 4632 155316 4644
rect 155368 4632 155374 4684
rect 156322 4632 156328 4684
rect 156380 4672 156386 4684
rect 156785 4675 156843 4681
rect 156785 4672 156797 4675
rect 156380 4644 156797 4672
rect 156380 4632 156386 4644
rect 156785 4641 156797 4644
rect 156831 4641 156843 4675
rect 156785 4635 156843 4641
rect 150069 4607 150127 4613
rect 150069 4573 150081 4607
rect 150115 4573 150127 4607
rect 150069 4567 150127 4573
rect 151633 4607 151691 4613
rect 151633 4573 151645 4607
rect 151679 4604 151691 4607
rect 153933 4607 153991 4613
rect 151679 4576 152228 4604
rect 151679 4573 151691 4576
rect 151633 4567 151691 4573
rect 147769 4539 147827 4545
rect 147769 4505 147781 4539
rect 147815 4536 147827 4539
rect 149606 4536 149612 4548
rect 147815 4508 149612 4536
rect 147815 4505 147827 4508
rect 147769 4499 147827 4505
rect 149606 4496 149612 4508
rect 149664 4496 149670 4548
rect 131669 4471 131727 4477
rect 131669 4437 131681 4471
rect 131715 4468 131727 4471
rect 132678 4468 132684 4480
rect 131715 4440 132684 4468
rect 131715 4437 131727 4440
rect 131669 4431 131727 4437
rect 132678 4428 132684 4440
rect 132736 4428 132742 4480
rect 152200 4477 152228 4576
rect 153933 4573 153945 4607
rect 153979 4604 153991 4607
rect 155773 4607 155831 4613
rect 153979 4576 154528 4604
rect 153979 4573 153991 4576
rect 153933 4567 153991 4573
rect 154500 4545 154528 4576
rect 155773 4573 155785 4607
rect 155819 4604 155831 4607
rect 163133 4607 163191 4613
rect 155819 4576 156368 4604
rect 155819 4573 155831 4576
rect 155773 4567 155831 4573
rect 154485 4539 154543 4545
rect 154485 4505 154497 4539
rect 154531 4536 154543 4539
rect 155126 4536 155132 4548
rect 154531 4508 155132 4536
rect 154531 4505 154543 4508
rect 154485 4499 154543 4505
rect 155126 4496 155132 4508
rect 155184 4496 155190 4548
rect 152185 4471 152243 4477
rect 152185 4437 152197 4471
rect 152231 4468 152243 4471
rect 153286 4468 153292 4480
rect 152231 4440 153292 4468
rect 152231 4437 152243 4440
rect 152185 4431 152243 4437
rect 153286 4428 153292 4440
rect 153344 4428 153350 4480
rect 154850 4468 154856 4480
rect 154811 4440 154856 4468
rect 154850 4428 154856 4440
rect 154908 4428 154914 4480
rect 156340 4477 156368 4576
rect 163133 4573 163145 4607
rect 163179 4604 163191 4607
rect 163179 4576 163636 4604
rect 163179 4573 163191 4576
rect 163133 4567 163191 4573
rect 163608 4480 163636 4576
rect 156325 4471 156383 4477
rect 156325 4437 156337 4471
rect 156371 4468 156383 4471
rect 156414 4468 156420 4480
rect 156371 4440 156420 4468
rect 156371 4437 156383 4440
rect 156325 4431 156383 4437
rect 156414 4428 156420 4440
rect 156472 4428 156478 4480
rect 159542 4468 159548 4480
rect 159503 4440 159548 4468
rect 159542 4428 159548 4440
rect 159600 4428 159606 4480
rect 163590 4468 163596 4480
rect 163551 4440 163596 4468
rect 163590 4428 163596 4440
rect 163648 4428 163654 4480
rect 164694 4468 164700 4480
rect 164655 4440 164700 4468
rect 164694 4428 164700 4440
rect 164752 4428 164758 4480
rect 368 4378 93012 4400
rect 368 4326 56667 4378
rect 56719 4326 56731 4378
rect 56783 4326 56795 4378
rect 56847 4326 56859 4378
rect 56911 4326 93012 4378
rect 368 4304 93012 4326
rect 102028 4378 169556 4400
rect 102028 4326 113088 4378
rect 113140 4326 113152 4378
rect 113204 4326 113216 4378
rect 113268 4326 113280 4378
rect 113332 4326 169556 4378
rect 102028 4304 169556 4326
rect 3513 4267 3571 4273
rect 3513 4233 3525 4267
rect 3559 4264 3571 4267
rect 3970 4264 3976 4276
rect 3559 4236 3976 4264
rect 3559 4233 3571 4236
rect 3513 4227 3571 4233
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 9858 4264 9864 4276
rect 4120 4236 9864 4264
rect 4120 4224 4126 4236
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 12066 4224 12072 4276
rect 12124 4264 12130 4276
rect 31570 4264 31576 4276
rect 12124 4236 31576 4264
rect 12124 4224 12130 4236
rect 31570 4224 31576 4236
rect 31628 4224 31634 4276
rect 31662 4224 31668 4276
rect 31720 4264 31726 4276
rect 31846 4264 31852 4276
rect 31720 4236 31852 4264
rect 31720 4224 31726 4236
rect 31846 4224 31852 4236
rect 31904 4224 31910 4276
rect 32214 4224 32220 4276
rect 32272 4264 32278 4276
rect 34974 4264 34980 4276
rect 32272 4236 34980 4264
rect 32272 4224 32278 4236
rect 34974 4224 34980 4236
rect 35032 4224 35038 4276
rect 35158 4224 35164 4276
rect 35216 4264 35222 4276
rect 35216 4236 36492 4264
rect 35216 4224 35222 4236
rect 9214 4156 9220 4208
rect 9272 4196 9278 4208
rect 9585 4199 9643 4205
rect 9585 4196 9597 4199
rect 9272 4168 9597 4196
rect 9272 4156 9278 4168
rect 9585 4165 9597 4168
rect 9631 4165 9643 4199
rect 29822 4196 29828 4208
rect 9585 4159 9643 4165
rect 24596 4168 25544 4196
rect 1302 4088 1308 4140
rect 1360 4128 1366 4140
rect 7653 4131 7711 4137
rect 1360 4100 7604 4128
rect 1360 4088 1366 4100
rect 4522 4060 4528 4072
rect 4483 4032 4528 4060
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 7006 4060 7012 4072
rect 6135 4032 7012 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4029 7159 4063
rect 7576 4060 7604 4100
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 8018 4128 8024 4140
rect 7699 4100 8024 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 10134 4128 10140 4140
rect 8128 4100 10140 4128
rect 8128 4060 8156 4100
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 18877 4131 18935 4137
rect 14424 4100 18368 4128
rect 14424 4088 14430 4100
rect 7576 4032 8156 4060
rect 7101 4023 7159 4029
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 7116 3992 7144 4023
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 16298 4060 16304 4072
rect 8444 4032 16304 4060
rect 8444 4020 8450 4032
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 18233 4063 18291 4069
rect 18233 4060 18245 4063
rect 16448 4032 18245 4060
rect 16448 4020 16454 4032
rect 18233 4029 18245 4032
rect 18279 4029 18291 4063
rect 18340 4060 18368 4100
rect 18877 4097 18889 4131
rect 18923 4128 18935 4131
rect 19610 4128 19616 4140
rect 18923 4100 19616 4128
rect 18923 4097 18935 4100
rect 18877 4091 18935 4097
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 19720 4100 21312 4128
rect 19720 4060 19748 4100
rect 21082 4060 21088 4072
rect 18340 4032 19748 4060
rect 20995 4032 21088 4060
rect 18233 4023 18291 4029
rect 21082 4020 21088 4032
rect 21140 4060 21146 4072
rect 21177 4063 21235 4069
rect 21177 4060 21189 4063
rect 21140 4032 21189 4060
rect 21140 4020 21146 4032
rect 21177 4029 21189 4032
rect 21223 4029 21235 4063
rect 21284 4060 21312 4100
rect 21358 4088 21364 4140
rect 21416 4128 21422 4140
rect 24029 4131 24087 4137
rect 24029 4128 24041 4131
rect 21416 4100 24041 4128
rect 21416 4088 21422 4100
rect 24029 4097 24041 4100
rect 24075 4097 24087 4131
rect 24029 4091 24087 4097
rect 24118 4088 24124 4140
rect 24176 4128 24182 4140
rect 24596 4128 24624 4168
rect 24176 4100 24624 4128
rect 24673 4131 24731 4137
rect 24176 4088 24182 4100
rect 24673 4097 24685 4131
rect 24719 4128 24731 4131
rect 25133 4131 25191 4137
rect 25133 4128 25145 4131
rect 24719 4100 25145 4128
rect 24719 4097 24731 4100
rect 24673 4091 24731 4097
rect 25133 4097 25145 4100
rect 25179 4128 25191 4131
rect 25406 4128 25412 4140
rect 25179 4100 25412 4128
rect 25179 4097 25191 4100
rect 25133 4091 25191 4097
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 25516 4128 25544 4168
rect 26160 4168 29828 4196
rect 26160 4128 26188 4168
rect 29822 4156 29828 4168
rect 29880 4156 29886 4208
rect 31110 4156 31116 4208
rect 31168 4196 31174 4208
rect 36354 4196 36360 4208
rect 31168 4168 36360 4196
rect 31168 4156 31174 4168
rect 36354 4156 36360 4168
rect 36412 4156 36418 4208
rect 36464 4196 36492 4236
rect 36630 4224 36636 4276
rect 36688 4264 36694 4276
rect 48222 4264 48228 4276
rect 36688 4236 48228 4264
rect 36688 4224 36694 4236
rect 48222 4224 48228 4236
rect 48280 4224 48286 4276
rect 48516 4236 49924 4264
rect 36722 4196 36728 4208
rect 36464 4168 36728 4196
rect 36722 4156 36728 4168
rect 36780 4156 36786 4208
rect 36814 4156 36820 4208
rect 36872 4196 36878 4208
rect 39666 4196 39672 4208
rect 36872 4168 39672 4196
rect 36872 4156 36878 4168
rect 39666 4156 39672 4168
rect 39724 4156 39730 4208
rect 40034 4156 40040 4208
rect 40092 4196 40098 4208
rect 41506 4196 41512 4208
rect 40092 4168 41512 4196
rect 40092 4156 40098 4168
rect 41506 4156 41512 4168
rect 41564 4156 41570 4208
rect 42794 4196 42800 4208
rect 41616 4168 42800 4196
rect 25516 4100 26188 4128
rect 26237 4131 26295 4137
rect 26237 4097 26249 4131
rect 26283 4128 26295 4131
rect 26326 4128 26332 4140
rect 26283 4100 26332 4128
rect 26283 4097 26295 4100
rect 26237 4091 26295 4097
rect 26326 4088 26332 4100
rect 26384 4088 26390 4140
rect 27798 4088 27804 4140
rect 27856 4128 27862 4140
rect 32674 4128 32680 4140
rect 27856 4100 32536 4128
rect 32635 4100 32680 4128
rect 27856 4088 27862 4100
rect 25498 4060 25504 4072
rect 21284 4032 25504 4060
rect 21177 4023 21235 4029
rect 25498 4020 25504 4032
rect 25556 4020 25562 4072
rect 25593 4063 25651 4069
rect 25593 4029 25605 4063
rect 25639 4029 25651 4063
rect 25593 4023 25651 4029
rect 9306 3992 9312 4004
rect 5408 3964 7144 3992
rect 7208 3964 9312 3992
rect 5408 3952 5414 3964
rect 3142 3884 3148 3936
rect 3200 3924 3206 3936
rect 7208 3924 7236 3964
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 9456 3964 24164 3992
rect 9456 3952 9462 3964
rect 3200 3896 7236 3924
rect 3200 3884 3206 3896
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 16574 3924 16580 3936
rect 7984 3896 16580 3924
rect 7984 3884 7990 3896
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 18046 3924 18052 3936
rect 16816 3896 18052 3924
rect 16816 3884 16822 3896
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18414 3884 18420 3936
rect 18472 3924 18478 3936
rect 20254 3924 20260 3936
rect 18472 3896 20260 3924
rect 18472 3884 18478 3896
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 21358 3924 21364 3936
rect 20496 3896 21364 3924
rect 20496 3884 20502 3896
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 22002 3884 22008 3936
rect 22060 3924 22066 3936
rect 23934 3924 23940 3936
rect 22060 3896 23940 3924
rect 22060 3884 22066 3896
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 24136 3924 24164 3964
rect 24210 3952 24216 4004
rect 24268 3992 24274 4004
rect 25608 3992 25636 4023
rect 25682 4020 25688 4072
rect 25740 4060 25746 4072
rect 32309 4063 32367 4069
rect 32309 4060 32321 4063
rect 25740 4032 32321 4060
rect 25740 4020 25746 4032
rect 32309 4029 32321 4032
rect 32355 4029 32367 4063
rect 32508 4060 32536 4100
rect 32674 4088 32680 4100
rect 32732 4088 32738 4140
rect 33226 4088 33232 4140
rect 33284 4128 33290 4140
rect 41616 4128 41644 4168
rect 42794 4156 42800 4168
rect 42852 4156 42858 4208
rect 45922 4196 45928 4208
rect 42904 4168 45928 4196
rect 33284 4100 41644 4128
rect 41693 4131 41751 4137
rect 33284 4088 33290 4100
rect 41693 4097 41705 4131
rect 41739 4128 41751 4131
rect 41966 4128 41972 4140
rect 41739 4100 41972 4128
rect 41739 4097 41751 4100
rect 41693 4091 41751 4097
rect 41966 4088 41972 4100
rect 42024 4128 42030 4140
rect 42518 4128 42524 4140
rect 42024 4100 42524 4128
rect 42024 4088 42030 4100
rect 42518 4088 42524 4100
rect 42576 4088 42582 4140
rect 42610 4088 42616 4140
rect 42668 4128 42674 4140
rect 42904 4128 42932 4168
rect 45922 4156 45928 4168
rect 45980 4156 45986 4208
rect 46014 4156 46020 4208
rect 46072 4196 46078 4208
rect 48516 4196 48544 4236
rect 46072 4168 48544 4196
rect 46072 4156 46078 4168
rect 48590 4156 48596 4208
rect 48648 4196 48654 4208
rect 49786 4196 49792 4208
rect 48648 4168 49792 4196
rect 48648 4156 48654 4168
rect 49786 4156 49792 4168
rect 49844 4156 49850 4208
rect 49896 4196 49924 4236
rect 49970 4224 49976 4276
rect 50028 4264 50034 4276
rect 53190 4264 53196 4276
rect 50028 4236 53196 4264
rect 50028 4224 50034 4236
rect 53190 4224 53196 4236
rect 53248 4224 53254 4276
rect 55030 4264 55036 4276
rect 53300 4236 55036 4264
rect 51258 4196 51264 4208
rect 49896 4168 51264 4196
rect 51258 4156 51264 4168
rect 51316 4156 51322 4208
rect 51534 4156 51540 4208
rect 51592 4196 51598 4208
rect 53300 4196 53328 4236
rect 55030 4224 55036 4236
rect 55088 4224 55094 4276
rect 55122 4224 55128 4276
rect 55180 4264 55186 4276
rect 55180 4236 55720 4264
rect 55180 4224 55186 4236
rect 51592 4168 53328 4196
rect 53653 4199 53711 4205
rect 51592 4156 51598 4168
rect 53653 4165 53665 4199
rect 53699 4196 53711 4199
rect 55582 4196 55588 4208
rect 53699 4168 55588 4196
rect 53699 4165 53711 4168
rect 53653 4159 53711 4165
rect 55582 4156 55588 4168
rect 55640 4156 55646 4208
rect 55692 4196 55720 4236
rect 55766 4224 55772 4276
rect 55824 4264 55830 4276
rect 56962 4264 56968 4276
rect 55824 4236 56968 4264
rect 55824 4224 55830 4236
rect 56962 4224 56968 4236
rect 57020 4224 57026 4276
rect 57054 4224 57060 4276
rect 57112 4264 57118 4276
rect 61197 4267 61255 4273
rect 61197 4264 61209 4267
rect 57112 4236 61209 4264
rect 57112 4224 57118 4236
rect 61197 4233 61209 4236
rect 61243 4233 61255 4267
rect 61197 4227 61255 4233
rect 61470 4224 61476 4276
rect 61528 4264 61534 4276
rect 62301 4267 62359 4273
rect 62301 4264 62313 4267
rect 61528 4236 62313 4264
rect 61528 4224 61534 4236
rect 62301 4233 62313 4236
rect 62347 4233 62359 4267
rect 62301 4227 62359 4233
rect 64598 4224 64604 4276
rect 64656 4264 64662 4276
rect 68465 4267 68523 4273
rect 68465 4264 68477 4267
rect 64656 4236 68477 4264
rect 64656 4224 64662 4236
rect 68465 4233 68477 4236
rect 68511 4233 68523 4267
rect 68465 4227 68523 4233
rect 70504 4236 76144 4264
rect 57698 4196 57704 4208
rect 55692 4168 57704 4196
rect 57698 4156 57704 4168
rect 57756 4156 57762 4208
rect 68278 4196 68284 4208
rect 60936 4168 68284 4196
rect 42668 4100 42932 4128
rect 42668 4088 42674 4100
rect 43346 4088 43352 4140
rect 43404 4128 43410 4140
rect 44542 4128 44548 4140
rect 43404 4100 44548 4128
rect 43404 4088 43410 4100
rect 44542 4088 44548 4100
rect 44600 4088 44606 4140
rect 44818 4088 44824 4140
rect 44876 4128 44882 4140
rect 47486 4128 47492 4140
rect 44876 4100 47492 4128
rect 44876 4088 44882 4100
rect 47486 4088 47492 4100
rect 47544 4088 47550 4140
rect 47946 4128 47952 4140
rect 47907 4100 47952 4128
rect 47946 4088 47952 4100
rect 48004 4088 48010 4140
rect 48222 4088 48228 4140
rect 48280 4128 48286 4140
rect 49602 4128 49608 4140
rect 48280 4100 49372 4128
rect 49563 4100 49608 4128
rect 48280 4088 48286 4100
rect 40770 4060 40776 4072
rect 32508 4032 40776 4060
rect 32309 4023 32367 4029
rect 40770 4020 40776 4032
rect 40828 4020 40834 4072
rect 41046 4060 41052 4072
rect 41007 4032 41052 4060
rect 41046 4020 41052 4032
rect 41104 4020 41110 4072
rect 49237 4063 49295 4069
rect 49237 4060 49249 4063
rect 41432 4032 49249 4060
rect 24268 3964 25636 3992
rect 24268 3952 24274 3964
rect 26694 3952 26700 4004
rect 26752 3992 26758 4004
rect 26752 3964 30880 3992
rect 26752 3952 26758 3964
rect 30742 3924 30748 3936
rect 24136 3896 30748 3924
rect 30742 3884 30748 3896
rect 30800 3884 30806 3936
rect 30852 3924 30880 3964
rect 31294 3952 31300 4004
rect 31352 3992 31358 4004
rect 41432 3992 41460 4032
rect 49237 4029 49249 4032
rect 49283 4029 49295 4063
rect 49344 4060 49372 4100
rect 49602 4088 49608 4100
rect 49660 4088 49666 4140
rect 49694 4088 49700 4140
rect 49752 4128 49758 4140
rect 49752 4100 51580 4128
rect 49752 4088 49758 4100
rect 51442 4060 51448 4072
rect 49344 4032 51448 4060
rect 49237 4023 49295 4029
rect 51442 4020 51448 4032
rect 51500 4020 51506 4072
rect 51552 4060 51580 4100
rect 51626 4088 51632 4140
rect 51684 4128 51690 4140
rect 51684 4100 52132 4128
rect 51684 4088 51690 4100
rect 51810 4060 51816 4072
rect 51552 4032 51816 4060
rect 51810 4020 51816 4032
rect 51868 4020 51874 4072
rect 51994 4060 52000 4072
rect 51955 4032 52000 4060
rect 51994 4020 52000 4032
rect 52052 4020 52058 4072
rect 52104 4060 52132 4100
rect 52362 4088 52368 4140
rect 52420 4128 52426 4140
rect 52641 4131 52699 4137
rect 52641 4128 52653 4131
rect 52420 4100 52653 4128
rect 52420 4088 52426 4100
rect 52641 4097 52653 4100
rect 52687 4128 52699 4131
rect 54294 4128 54300 4140
rect 52687 4100 54300 4128
rect 52687 4097 52699 4100
rect 52641 4091 52699 4097
rect 54294 4088 54300 4100
rect 54352 4088 54358 4140
rect 55306 4128 55312 4140
rect 55267 4100 55312 4128
rect 55306 4088 55312 4100
rect 55364 4088 55370 4140
rect 55490 4088 55496 4140
rect 55548 4128 55554 4140
rect 56226 4128 56232 4140
rect 55548 4100 56232 4128
rect 55548 4088 55554 4100
rect 56226 4088 56232 4100
rect 56284 4088 56290 4140
rect 56318 4088 56324 4140
rect 56376 4128 56382 4140
rect 60550 4128 60556 4140
rect 56376 4100 60556 4128
rect 56376 4088 56382 4100
rect 60550 4088 60556 4100
rect 60608 4088 60614 4140
rect 54665 4063 54723 4069
rect 54665 4060 54677 4063
rect 52104 4032 54677 4060
rect 54665 4029 54677 4032
rect 54711 4029 54723 4063
rect 54665 4023 54723 4029
rect 54754 4020 54760 4072
rect 54812 4060 54818 4072
rect 55766 4060 55772 4072
rect 54812 4032 55772 4060
rect 54812 4020 54818 4032
rect 55766 4020 55772 4032
rect 55824 4020 55830 4072
rect 60936 4060 60964 4168
rect 68278 4156 68284 4168
rect 68336 4156 68342 4208
rect 61102 4128 61108 4140
rect 61063 4100 61108 4128
rect 61102 4088 61108 4100
rect 61160 4088 61166 4140
rect 62206 4128 62212 4140
rect 62167 4100 62212 4128
rect 62206 4088 62212 4100
rect 62264 4088 62270 4140
rect 62758 4128 62764 4140
rect 62719 4100 62764 4128
rect 62758 4088 62764 4100
rect 62816 4128 62822 4140
rect 62942 4128 62948 4140
rect 62816 4100 62948 4128
rect 62816 4088 62822 4100
rect 62942 4088 62948 4100
rect 63000 4088 63006 4140
rect 63218 4128 63224 4140
rect 63179 4100 63224 4128
rect 63218 4088 63224 4100
rect 63276 4088 63282 4140
rect 63310 4088 63316 4140
rect 63368 4128 63374 4140
rect 68373 4131 68431 4137
rect 63368 4100 63413 4128
rect 63368 4088 63374 4100
rect 68373 4097 68385 4131
rect 68419 4128 68431 4131
rect 68738 4128 68744 4140
rect 68419 4100 68744 4128
rect 68419 4097 68431 4100
rect 68373 4091 68431 4097
rect 68738 4088 68744 4100
rect 68796 4088 68802 4140
rect 69937 4131 69995 4137
rect 69937 4097 69949 4131
rect 69983 4097 69995 4131
rect 69937 4091 69995 4097
rect 64414 4060 64420 4072
rect 55876 4032 60964 4060
rect 61212 4032 64420 4060
rect 31352 3964 41460 3992
rect 31352 3952 31358 3964
rect 41506 3952 41512 4004
rect 41564 3992 41570 4004
rect 45278 3992 45284 4004
rect 41564 3964 45284 3992
rect 41564 3952 41570 3964
rect 45278 3952 45284 3964
rect 45336 3952 45342 4004
rect 49418 3992 49424 4004
rect 45388 3964 49424 3992
rect 39942 3924 39948 3936
rect 30852 3896 39948 3924
rect 39942 3884 39948 3896
rect 40000 3884 40006 3936
rect 40034 3884 40040 3936
rect 40092 3924 40098 3936
rect 45388 3924 45416 3964
rect 49418 3952 49424 3964
rect 49476 3952 49482 4004
rect 50062 3952 50068 4004
rect 50120 3992 50126 4004
rect 55876 3992 55904 4032
rect 50120 3964 55904 3992
rect 50120 3952 50126 3964
rect 56042 3952 56048 4004
rect 56100 3992 56106 4004
rect 61212 3992 61240 4032
rect 64414 4020 64420 4032
rect 64472 4020 64478 4072
rect 69952 4060 69980 4091
rect 70026 4088 70032 4140
rect 70084 4128 70090 4140
rect 70084 4100 70129 4128
rect 70084 4088 70090 4100
rect 70210 4088 70216 4140
rect 70268 4128 70274 4140
rect 70504 4128 70532 4236
rect 70780 4168 71268 4196
rect 70268 4100 70532 4128
rect 70268 4088 70274 4100
rect 70578 4088 70584 4140
rect 70636 4128 70642 4140
rect 70780 4128 70808 4168
rect 70946 4128 70952 4140
rect 70636 4100 70808 4128
rect 70907 4100 70952 4128
rect 70636 4088 70642 4100
rect 70946 4088 70952 4100
rect 71004 4088 71010 4140
rect 71038 4088 71044 4140
rect 71096 4128 71102 4140
rect 71240 4128 71268 4168
rect 71792 4168 72280 4196
rect 71792 4128 71820 4168
rect 71958 4128 71964 4140
rect 71096 4100 71141 4128
rect 71240 4100 71820 4128
rect 71919 4100 71964 4128
rect 71096 4088 71102 4100
rect 71958 4088 71964 4100
rect 72016 4088 72022 4140
rect 72050 4088 72056 4140
rect 72108 4128 72114 4140
rect 72252 4128 72280 4168
rect 76006 4128 76012 4140
rect 72108 4100 72153 4128
rect 72252 4100 76012 4128
rect 72108 4088 72114 4100
rect 76006 4088 76012 4100
rect 76064 4088 76070 4140
rect 76116 4128 76144 4236
rect 105906 4224 105912 4276
rect 105964 4264 105970 4276
rect 113542 4264 113548 4276
rect 105964 4236 113548 4264
rect 105964 4224 105970 4236
rect 113542 4224 113548 4236
rect 113600 4224 113606 4276
rect 114002 4224 114008 4276
rect 114060 4264 114066 4276
rect 114833 4267 114891 4273
rect 114833 4264 114845 4267
rect 114060 4236 114845 4264
rect 114060 4224 114066 4236
rect 114833 4233 114845 4236
rect 114879 4233 114891 4267
rect 114833 4227 114891 4233
rect 115382 4224 115388 4276
rect 115440 4264 115446 4276
rect 125870 4264 125876 4276
rect 115440 4236 125876 4264
rect 115440 4224 115446 4236
rect 125870 4224 125876 4236
rect 125928 4224 125934 4276
rect 153470 4264 153476 4276
rect 153431 4236 153476 4264
rect 153470 4224 153476 4236
rect 153528 4224 153534 4276
rect 88153 4199 88211 4205
rect 88153 4165 88165 4199
rect 88199 4196 88211 4199
rect 88886 4196 88892 4208
rect 88199 4168 88892 4196
rect 88199 4165 88211 4168
rect 88153 4159 88211 4165
rect 88886 4156 88892 4168
rect 88944 4156 88950 4208
rect 115937 4199 115995 4205
rect 115937 4196 115949 4199
rect 102152 4168 102456 4196
rect 76374 4128 76380 4140
rect 76116 4100 76380 4128
rect 76374 4088 76380 4100
rect 76432 4088 76438 4140
rect 89162 4128 89168 4140
rect 89123 4100 89168 4128
rect 89162 4088 89168 4100
rect 89220 4088 89226 4140
rect 90269 4131 90327 4137
rect 90269 4097 90281 4131
rect 90315 4128 90327 4131
rect 91094 4128 91100 4140
rect 90315 4100 91100 4128
rect 90315 4097 90327 4100
rect 90269 4091 90327 4097
rect 91094 4088 91100 4100
rect 91152 4088 91158 4140
rect 91741 4131 91799 4137
rect 91741 4097 91753 4131
rect 91787 4128 91799 4131
rect 92290 4128 92296 4140
rect 91787 4100 92296 4128
rect 91787 4097 91799 4100
rect 91741 4091 91799 4097
rect 92290 4088 92296 4100
rect 92348 4088 92354 4140
rect 100478 4088 100484 4140
rect 100536 4128 100542 4140
rect 102152 4128 102180 4168
rect 100536 4100 102180 4128
rect 100536 4088 100542 4100
rect 102226 4088 102232 4140
rect 102284 4128 102290 4140
rect 102321 4131 102379 4137
rect 102321 4128 102333 4131
rect 102284 4100 102333 4128
rect 102284 4088 102290 4100
rect 102321 4097 102333 4100
rect 102367 4097 102379 4131
rect 102428 4128 102456 4168
rect 106384 4168 106872 4196
rect 106384 4128 106412 4168
rect 102428 4100 106412 4128
rect 102321 4091 102379 4097
rect 106458 4088 106464 4140
rect 106516 4128 106522 4140
rect 106553 4131 106611 4137
rect 106553 4128 106565 4131
rect 106516 4100 106565 4128
rect 106516 4088 106522 4100
rect 106553 4097 106565 4100
rect 106599 4097 106611 4131
rect 106553 4091 106611 4097
rect 106642 4088 106648 4140
rect 106700 4128 106706 4140
rect 106844 4128 106872 4168
rect 107580 4168 108068 4196
rect 107580 4128 107608 4168
rect 107746 4128 107752 4140
rect 106700 4100 106745 4128
rect 106844 4100 107608 4128
rect 107707 4100 107752 4128
rect 106700 4088 106706 4100
rect 107746 4088 107752 4100
rect 107804 4088 107810 4140
rect 107838 4088 107844 4140
rect 107896 4128 107902 4140
rect 108040 4128 108068 4168
rect 113560 4168 113864 4196
rect 109034 4128 109040 4140
rect 107896 4100 107941 4128
rect 108040 4100 109040 4128
rect 107896 4088 107902 4100
rect 109034 4088 109040 4100
rect 109092 4088 109098 4140
rect 113560 4128 113588 4168
rect 109236 4100 113588 4128
rect 70394 4060 70400 4072
rect 69952 4032 70400 4060
rect 70394 4020 70400 4032
rect 70452 4060 70458 4072
rect 71222 4060 71228 4072
rect 70452 4032 71228 4060
rect 70452 4020 70458 4032
rect 71222 4020 71228 4032
rect 71280 4020 71286 4072
rect 71314 4020 71320 4072
rect 71372 4060 71378 4072
rect 77846 4060 77852 4072
rect 71372 4032 77852 4060
rect 71372 4020 71378 4032
rect 77846 4020 77852 4032
rect 77904 4020 77910 4072
rect 89990 4020 89996 4072
rect 90048 4060 90054 4072
rect 90361 4063 90419 4069
rect 90361 4060 90373 4063
rect 90048 4032 90373 4060
rect 90048 4020 90054 4032
rect 90361 4029 90373 4032
rect 90407 4029 90419 4063
rect 90361 4023 90419 4029
rect 91833 4063 91891 4069
rect 91833 4029 91845 4063
rect 91879 4060 91891 4063
rect 91922 4060 91928 4072
rect 91879 4032 91928 4060
rect 91879 4029 91891 4032
rect 91833 4023 91891 4029
rect 91922 4020 91928 4032
rect 91980 4020 91986 4072
rect 100294 4020 100300 4072
rect 100352 4060 100358 4072
rect 108206 4060 108212 4072
rect 100352 4032 108212 4060
rect 100352 4020 100358 4032
rect 108206 4020 108212 4032
rect 108264 4020 108270 4072
rect 108390 4020 108396 4072
rect 108448 4060 108454 4072
rect 109236 4060 109264 4100
rect 113634 4088 113640 4140
rect 113692 4128 113698 4140
rect 113737 4131 113795 4137
rect 113737 4128 113749 4131
rect 113692 4100 113749 4128
rect 113692 4088 113698 4100
rect 113737 4097 113749 4100
rect 113783 4097 113795 4131
rect 113836 4128 113864 4168
rect 114664 4168 114968 4196
rect 114664 4128 114692 4168
rect 113836 4100 114692 4128
rect 114741 4131 114799 4137
rect 113737 4091 113795 4097
rect 114741 4097 114753 4131
rect 114787 4128 114799 4131
rect 114830 4128 114836 4140
rect 114787 4100 114836 4128
rect 114787 4097 114799 4100
rect 114741 4091 114799 4097
rect 114830 4088 114836 4100
rect 114888 4088 114894 4140
rect 114940 4128 114968 4168
rect 115768 4168 115949 4196
rect 115768 4128 115796 4168
rect 115937 4165 115949 4168
rect 115983 4165 115995 4199
rect 115937 4159 115995 4165
rect 117038 4156 117044 4208
rect 117096 4196 117102 4208
rect 124677 4199 124735 4205
rect 124677 4196 124689 4199
rect 117096 4168 124689 4196
rect 117096 4156 117102 4168
rect 124677 4165 124689 4168
rect 124723 4165 124735 4199
rect 124677 4159 124735 4165
rect 137925 4199 137983 4205
rect 137925 4165 137937 4199
rect 137971 4196 137983 4199
rect 138658 4196 138664 4208
rect 137971 4168 138664 4196
rect 137971 4165 137983 4168
rect 137925 4159 137983 4165
rect 138658 4156 138664 4168
rect 138716 4156 138722 4208
rect 114940 4100 115796 4128
rect 115842 4088 115848 4140
rect 115900 4128 115906 4140
rect 119525 4131 119583 4137
rect 115900 4100 115945 4128
rect 115900 4088 115906 4100
rect 119525 4097 119537 4131
rect 119571 4128 119583 4131
rect 120074 4128 120080 4140
rect 119571 4100 120080 4128
rect 119571 4097 119583 4100
rect 119525 4091 119583 4097
rect 120074 4088 120080 4100
rect 120132 4088 120138 4140
rect 121549 4131 121607 4137
rect 121549 4097 121561 4131
rect 121595 4128 121607 4131
rect 121638 4128 121644 4140
rect 121595 4100 121644 4128
rect 121595 4097 121607 4100
rect 121549 4091 121607 4097
rect 121638 4088 121644 4100
rect 121696 4088 121702 4140
rect 124582 4128 124588 4140
rect 124543 4100 124588 4128
rect 124582 4088 124588 4100
rect 124640 4088 124646 4140
rect 125594 4128 125600 4140
rect 125555 4100 125600 4128
rect 125594 4088 125600 4100
rect 125652 4088 125658 4140
rect 125689 4131 125747 4137
rect 125689 4097 125701 4131
rect 125735 4128 125747 4131
rect 125962 4128 125968 4140
rect 125735 4100 125968 4128
rect 125735 4097 125747 4100
rect 125689 4091 125747 4097
rect 125962 4088 125968 4100
rect 126020 4088 126026 4140
rect 126882 4128 126888 4140
rect 126843 4100 126888 4128
rect 126882 4088 126888 4100
rect 126940 4088 126946 4140
rect 126977 4131 127035 4137
rect 126977 4097 126989 4131
rect 127023 4128 127035 4131
rect 127158 4128 127164 4140
rect 127023 4100 127164 4128
rect 127023 4097 127035 4100
rect 126977 4091 127035 4097
rect 127158 4088 127164 4100
rect 127216 4088 127222 4140
rect 130194 4128 130200 4140
rect 130155 4100 130200 4128
rect 130194 4088 130200 4100
rect 130252 4088 130258 4140
rect 130286 4088 130292 4140
rect 130344 4128 130350 4140
rect 131298 4128 131304 4140
rect 130344 4100 130389 4128
rect 131259 4100 131304 4128
rect 130344 4088 130350 4100
rect 131298 4088 131304 4100
rect 131356 4088 131362 4140
rect 131390 4088 131396 4140
rect 131448 4128 131454 4140
rect 148137 4131 148195 4137
rect 131448 4100 131493 4128
rect 131448 4088 131454 4100
rect 148137 4097 148149 4131
rect 148183 4097 148195 4131
rect 148137 4091 148195 4097
rect 108448 4032 109264 4060
rect 108448 4020 108454 4032
rect 109310 4020 109316 4072
rect 109368 4060 109374 4072
rect 109368 4032 121684 4060
rect 109368 4020 109374 4032
rect 56100 3964 61240 3992
rect 56100 3952 56106 3964
rect 61378 3952 61384 4004
rect 61436 3992 61442 4004
rect 61436 3964 74488 3992
rect 61436 3952 61442 3964
rect 40092 3896 45416 3924
rect 40092 3884 40098 3896
rect 45646 3884 45652 3936
rect 45704 3924 45710 3936
rect 46017 3927 46075 3933
rect 46017 3924 46029 3927
rect 45704 3896 46029 3924
rect 45704 3884 45710 3896
rect 46017 3893 46029 3896
rect 46063 3924 46075 3927
rect 47762 3924 47768 3936
rect 46063 3896 47768 3924
rect 46063 3893 46075 3896
rect 46017 3887 46075 3893
rect 47762 3884 47768 3896
rect 47820 3884 47826 3936
rect 47946 3924 47952 3936
rect 47907 3896 47952 3924
rect 47946 3884 47952 3896
rect 48004 3884 48010 3936
rect 48498 3884 48504 3936
rect 48556 3924 48562 3936
rect 55490 3924 55496 3936
rect 48556 3896 55496 3924
rect 48556 3884 48562 3896
rect 55490 3884 55496 3896
rect 55548 3884 55554 3936
rect 55766 3884 55772 3936
rect 55824 3924 55830 3936
rect 58526 3924 58532 3936
rect 55824 3896 58532 3924
rect 55824 3884 55830 3896
rect 58526 3884 58532 3896
rect 58584 3884 58590 3936
rect 58710 3884 58716 3936
rect 58768 3924 58774 3936
rect 64046 3924 64052 3936
rect 58768 3896 64052 3924
rect 58768 3884 58774 3896
rect 64046 3884 64052 3896
rect 64104 3884 64110 3936
rect 64598 3884 64604 3936
rect 64656 3924 64662 3936
rect 70118 3924 70124 3936
rect 64656 3896 70124 3924
rect 64656 3884 64662 3896
rect 70118 3884 70124 3896
rect 70176 3884 70182 3936
rect 70302 3884 70308 3936
rect 70360 3924 70366 3936
rect 70578 3924 70584 3936
rect 70360 3896 70584 3924
rect 70360 3884 70366 3896
rect 70578 3884 70584 3896
rect 70636 3884 70642 3936
rect 74460 3924 74488 3964
rect 74534 3952 74540 4004
rect 74592 3992 74598 4004
rect 84654 3992 84660 4004
rect 74592 3964 84660 3992
rect 74592 3952 74598 3964
rect 84654 3952 84660 3964
rect 84712 3952 84718 4004
rect 100478 3952 100484 4004
rect 100536 3992 100542 4004
rect 100536 3964 102548 3992
rect 100536 3952 100542 3964
rect 82998 3924 83004 3936
rect 74460 3896 83004 3924
rect 82998 3884 83004 3896
rect 83056 3884 83062 3936
rect 89254 3924 89260 3936
rect 89215 3896 89260 3924
rect 89254 3884 89260 3896
rect 89312 3884 89318 3936
rect 100202 3884 100208 3936
rect 100260 3924 100266 3936
rect 102413 3927 102471 3933
rect 102413 3924 102425 3927
rect 100260 3896 102425 3924
rect 100260 3884 100266 3896
rect 102413 3893 102425 3896
rect 102459 3893 102471 3927
rect 102520 3924 102548 3964
rect 104250 3952 104256 4004
rect 104308 3992 104314 4004
rect 107562 3992 107568 4004
rect 104308 3964 107568 3992
rect 104308 3952 104314 3964
rect 107562 3952 107568 3964
rect 107620 3952 107626 4004
rect 109218 3952 109224 4004
rect 109276 3992 109282 4004
rect 111610 3992 111616 4004
rect 109276 3964 111616 3992
rect 109276 3952 109282 3964
rect 111610 3952 111616 3964
rect 111668 3952 111674 4004
rect 114738 3992 114744 4004
rect 113468 3964 114744 3992
rect 108850 3924 108856 3936
rect 102520 3896 108856 3924
rect 102413 3887 102471 3893
rect 108850 3884 108856 3896
rect 108908 3884 108914 3936
rect 108942 3884 108948 3936
rect 109000 3924 109006 3936
rect 113468 3924 113496 3964
rect 114738 3952 114744 3964
rect 114796 3952 114802 4004
rect 114922 3952 114928 4004
rect 114980 3992 114986 4004
rect 121656 4001 121684 4032
rect 121730 4020 121736 4072
rect 121788 4060 121794 4072
rect 129826 4060 129832 4072
rect 121788 4032 129832 4060
rect 121788 4020 121794 4032
rect 129826 4020 129832 4032
rect 129884 4020 129890 4072
rect 148152 4060 148180 4091
rect 148226 4088 148232 4140
rect 148284 4128 148290 4140
rect 150069 4131 150127 4137
rect 148284 4100 148329 4128
rect 148284 4088 148290 4100
rect 150069 4097 150081 4131
rect 150115 4128 150127 4131
rect 150158 4128 150164 4140
rect 150115 4100 150164 4128
rect 150115 4097 150127 4100
rect 150069 4091 150127 4097
rect 150158 4088 150164 4100
rect 150216 4088 150222 4140
rect 155034 4128 155040 4140
rect 154995 4100 155040 4128
rect 155034 4088 155040 4100
rect 155092 4088 155098 4140
rect 156046 4128 156052 4140
rect 156007 4100 156052 4128
rect 156046 4088 156052 4100
rect 156104 4088 156110 4140
rect 156141 4131 156199 4137
rect 156141 4097 156153 4131
rect 156187 4128 156199 4131
rect 156230 4128 156236 4140
rect 156187 4100 156236 4128
rect 156187 4097 156199 4100
rect 156141 4091 156199 4097
rect 156230 4088 156236 4100
rect 156288 4088 156294 4140
rect 158441 4131 158499 4137
rect 158441 4097 158453 4131
rect 158487 4097 158499 4131
rect 158441 4091 158499 4097
rect 149054 4060 149060 4072
rect 148152 4032 149060 4060
rect 149054 4020 149060 4032
rect 149112 4020 149118 4072
rect 155129 4063 155187 4069
rect 155129 4029 155141 4063
rect 155175 4060 155187 4063
rect 155954 4060 155960 4072
rect 155175 4032 155960 4060
rect 155175 4029 155187 4032
rect 155129 4023 155187 4029
rect 155954 4020 155960 4032
rect 156012 4020 156018 4072
rect 158456 4060 158484 4091
rect 158530 4088 158536 4140
rect 158588 4128 158594 4140
rect 160189 4131 160247 4137
rect 158588 4100 158633 4128
rect 158588 4088 158594 4100
rect 160189 4097 160201 4131
rect 160235 4128 160247 4131
rect 160554 4128 160560 4140
rect 160235 4100 160560 4128
rect 160235 4097 160247 4100
rect 160189 4091 160247 4097
rect 160554 4088 160560 4100
rect 160612 4088 160618 4140
rect 161201 4131 161259 4137
rect 161201 4097 161213 4131
rect 161247 4128 161259 4131
rect 161750 4128 161756 4140
rect 161247 4100 161756 4128
rect 161247 4097 161259 4100
rect 161201 4091 161259 4097
rect 161750 4088 161756 4100
rect 161808 4088 161814 4140
rect 162213 4131 162271 4137
rect 162213 4097 162225 4131
rect 162259 4128 162271 4131
rect 162486 4128 162492 4140
rect 162259 4100 162492 4128
rect 162259 4097 162271 4100
rect 162213 4091 162271 4097
rect 162486 4088 162492 4100
rect 162544 4088 162550 4140
rect 164878 4088 164884 4140
rect 164936 4128 164942 4140
rect 165522 4128 165528 4140
rect 164936 4100 165528 4128
rect 164936 4088 164942 4100
rect 165522 4088 165528 4100
rect 165580 4088 165586 4140
rect 165614 4088 165620 4140
rect 165672 4128 165678 4140
rect 165672 4100 165717 4128
rect 165672 4088 165678 4100
rect 158714 4060 158720 4072
rect 158456 4032 158720 4060
rect 158714 4020 158720 4032
rect 158772 4020 158778 4072
rect 160278 4060 160284 4072
rect 160239 4032 160284 4060
rect 160278 4020 160284 4032
rect 160336 4020 160342 4072
rect 161293 4063 161351 4069
rect 161293 4029 161305 4063
rect 161339 4060 161351 4063
rect 161566 4060 161572 4072
rect 161339 4032 161572 4060
rect 161339 4029 161351 4032
rect 161293 4023 161351 4029
rect 161566 4020 161572 4032
rect 161624 4020 161630 4072
rect 162302 4060 162308 4072
rect 162263 4032 162308 4060
rect 162302 4020 162308 4032
rect 162360 4020 162366 4072
rect 119617 3995 119675 4001
rect 119617 3992 119629 3995
rect 114980 3964 119629 3992
rect 114980 3952 114986 3964
rect 119617 3961 119629 3964
rect 119663 3961 119675 3995
rect 119617 3955 119675 3961
rect 121641 3995 121699 4001
rect 121641 3961 121653 3995
rect 121687 3961 121699 3995
rect 134886 3992 134892 4004
rect 121641 3955 121699 3961
rect 124784 3964 134892 3992
rect 109000 3896 113496 3924
rect 109000 3884 109006 3896
rect 113542 3884 113548 3936
rect 113600 3924 113606 3936
rect 113821 3927 113879 3933
rect 113821 3924 113833 3927
rect 113600 3896 113833 3924
rect 113600 3884 113606 3896
rect 113821 3893 113833 3896
rect 113867 3893 113879 3927
rect 113821 3887 113879 3893
rect 114830 3884 114836 3936
rect 114888 3924 114894 3936
rect 115014 3924 115020 3936
rect 114888 3896 115020 3924
rect 114888 3884 114894 3896
rect 115014 3884 115020 3896
rect 115072 3924 115078 3936
rect 117590 3924 117596 3936
rect 115072 3896 117596 3924
rect 115072 3884 115078 3896
rect 117590 3884 117596 3896
rect 117648 3884 117654 3936
rect 122282 3884 122288 3936
rect 122340 3924 122346 3936
rect 124784 3924 124812 3964
rect 134886 3952 134892 3964
rect 134944 3952 134950 4004
rect 144086 3952 144092 4004
rect 144144 3992 144150 4004
rect 158162 3992 158168 4004
rect 144144 3964 158168 3992
rect 144144 3952 144150 3964
rect 158162 3952 158168 3964
rect 158220 3952 158226 4004
rect 126422 3924 126428 3936
rect 122340 3896 124812 3924
rect 126383 3896 126428 3924
rect 122340 3884 122346 3896
rect 126422 3884 126428 3896
rect 126480 3884 126486 3936
rect 150161 3927 150219 3933
rect 150161 3893 150173 3927
rect 150207 3924 150219 3927
rect 151078 3924 151084 3936
rect 150207 3896 151084 3924
rect 150207 3893 150219 3896
rect 150161 3887 150219 3893
rect 151078 3884 151084 3896
rect 151136 3884 151142 3936
rect 368 3834 93012 3856
rect 368 3782 28456 3834
rect 28508 3782 28520 3834
rect 28572 3782 28584 3834
rect 28636 3782 28648 3834
rect 28700 3782 84878 3834
rect 84930 3782 84942 3834
rect 84994 3782 85006 3834
rect 85058 3782 85070 3834
rect 85122 3782 93012 3834
rect 368 3760 93012 3782
rect 102028 3834 169556 3856
rect 102028 3782 141299 3834
rect 141351 3782 141363 3834
rect 141415 3782 141427 3834
rect 141479 3782 141491 3834
rect 141543 3782 169556 3834
rect 102028 3760 169556 3782
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 6362 3720 6368 3732
rect 3660 3692 6368 3720
rect 3660 3680 3666 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 6638 3720 6644 3732
rect 6599 3692 6644 3720
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7190 3720 7196 3732
rect 7151 3692 7196 3720
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 9272 3692 9413 3720
rect 9272 3680 9278 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 9401 3683 9459 3689
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 11698 3720 11704 3732
rect 9732 3692 11704 3720
rect 9732 3680 9738 3692
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 18693 3723 18751 3729
rect 16356 3692 17172 3720
rect 16356 3680 16362 3692
rect 4062 3612 4068 3664
rect 4120 3652 4126 3664
rect 7377 3655 7435 3661
rect 7377 3652 7389 3655
rect 4120 3624 7389 3652
rect 4120 3612 4126 3624
rect 7377 3621 7389 3624
rect 7423 3621 7435 3655
rect 7377 3615 7435 3621
rect 8662 3612 8668 3664
rect 8720 3652 8726 3664
rect 8720 3624 14504 3652
rect 8720 3612 8726 3624
rect 5718 3584 5724 3596
rect 5679 3556 5724 3584
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 7116 3556 7573 3584
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4540 3488 4721 3516
rect 4540 3457 4568 3488
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3516 6331 3519
rect 6638 3516 6644 3528
rect 6319 3488 6644 3516
rect 6319 3485 6331 3488
rect 6273 3479 6331 3485
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 7116 3525 7144 3556
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 9272 3556 9597 3584
rect 9272 3544 9278 3556
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 10597 3587 10655 3593
rect 10597 3553 10609 3587
rect 10643 3553 10655 3587
rect 14366 3584 14372 3596
rect 10597 3547 10655 3553
rect 11072 3556 14372 3584
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 6748 3488 7113 3516
rect 3697 3451 3755 3457
rect 3697 3417 3709 3451
rect 3743 3448 3755 3451
rect 4525 3451 4583 3457
rect 4525 3448 4537 3451
rect 3743 3420 4537 3448
rect 3743 3417 3755 3420
rect 3697 3411 3755 3417
rect 4525 3417 4537 3420
rect 4571 3417 4583 3451
rect 4525 3411 4583 3417
rect 4890 3408 4896 3460
rect 4948 3448 4954 3460
rect 6748 3448 6776 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3516 7435 3519
rect 10612 3516 10640 3547
rect 7423 3488 10640 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 7006 3448 7012 3460
rect 4948 3420 6776 3448
rect 6919 3420 7012 3448
rect 4948 3408 4954 3420
rect 7006 3408 7012 3420
rect 7064 3448 7070 3460
rect 7742 3448 7748 3460
rect 7064 3420 7748 3448
rect 7064 3408 7070 3420
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 11072 3448 11100 3556
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 10100 3420 11100 3448
rect 11164 3448 11192 3479
rect 11514 3448 11520 3460
rect 11164 3420 11520 3448
rect 10100 3408 10106 3420
rect 11514 3408 11520 3420
rect 11572 3408 11578 3460
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 10686 3380 10692 3392
rect 4028 3352 10692 3380
rect 4028 3340 4034 3352
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 11974 3380 11980 3392
rect 11935 3352 11980 3380
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 14476 3380 14504 3624
rect 15286 3612 15292 3664
rect 15344 3652 15350 3664
rect 16666 3652 16672 3664
rect 15344 3624 16672 3652
rect 15344 3612 15350 3624
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 17144 3652 17172 3692
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 19610 3720 19616 3732
rect 18739 3692 19616 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 24213 3723 24271 3729
rect 24213 3720 24225 3723
rect 19944 3692 24225 3720
rect 19944 3680 19950 3692
rect 24213 3689 24225 3692
rect 24259 3689 24271 3723
rect 25038 3720 25044 3732
rect 24999 3692 25044 3720
rect 24213 3683 24271 3689
rect 25038 3680 25044 3692
rect 25096 3680 25102 3732
rect 26145 3723 26203 3729
rect 26145 3720 26157 3723
rect 25148 3692 26157 3720
rect 24026 3652 24032 3664
rect 17144 3624 24032 3652
rect 24026 3612 24032 3624
rect 24084 3612 24090 3664
rect 24118 3612 24124 3664
rect 24176 3652 24182 3664
rect 24854 3652 24860 3664
rect 24176 3624 24860 3652
rect 24176 3612 24182 3624
rect 24854 3612 24860 3624
rect 24912 3612 24918 3664
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 17954 3584 17960 3596
rect 15712 3556 17960 3584
rect 15712 3544 15718 3556
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 19334 3584 19340 3596
rect 18279 3556 19340 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 18248 3516 18276 3547
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 21910 3584 21916 3596
rect 21560 3556 21916 3584
rect 17819 3488 18276 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 20714 3516 20720 3528
rect 18380 3488 20720 3516
rect 18380 3476 18386 3488
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 21082 3516 21088 3528
rect 21043 3488 21088 3516
rect 21082 3476 21088 3488
rect 21140 3476 21146 3528
rect 21560 3525 21588 3556
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 24486 3544 24492 3596
rect 24544 3584 24550 3596
rect 25148 3584 25176 3692
rect 26145 3689 26157 3692
rect 26191 3689 26203 3723
rect 26326 3720 26332 3732
rect 26287 3692 26332 3720
rect 26145 3683 26203 3689
rect 26326 3680 26332 3692
rect 26384 3680 26390 3732
rect 27982 3720 27988 3732
rect 27943 3692 27988 3720
rect 27982 3680 27988 3692
rect 28040 3680 28046 3732
rect 28074 3680 28080 3732
rect 28132 3720 28138 3732
rect 28902 3720 28908 3732
rect 28132 3692 28908 3720
rect 28132 3680 28138 3692
rect 28902 3680 28908 3692
rect 28960 3680 28966 3732
rect 29365 3723 29423 3729
rect 29365 3689 29377 3723
rect 29411 3720 29423 3723
rect 29638 3720 29644 3732
rect 29411 3692 29644 3720
rect 29411 3689 29423 3692
rect 29365 3683 29423 3689
rect 29638 3680 29644 3692
rect 29696 3680 29702 3732
rect 30006 3680 30012 3732
rect 30064 3720 30070 3732
rect 47670 3720 47676 3732
rect 30064 3692 47676 3720
rect 30064 3680 30070 3692
rect 47670 3680 47676 3692
rect 47728 3680 47734 3732
rect 48038 3720 48044 3732
rect 47999 3692 48044 3720
rect 48038 3680 48044 3692
rect 48096 3680 48102 3732
rect 48130 3680 48136 3732
rect 48188 3720 48194 3732
rect 49513 3723 49571 3729
rect 49513 3720 49525 3723
rect 48188 3692 49525 3720
rect 48188 3680 48194 3692
rect 49513 3689 49525 3692
rect 49559 3689 49571 3723
rect 49513 3683 49571 3689
rect 49602 3680 49608 3732
rect 49660 3720 49666 3732
rect 49660 3692 49705 3720
rect 49660 3680 49666 3692
rect 50154 3680 50160 3732
rect 50212 3720 50218 3732
rect 51077 3723 51135 3729
rect 51077 3720 51089 3723
rect 50212 3692 51089 3720
rect 50212 3680 50218 3692
rect 51077 3689 51089 3692
rect 51123 3689 51135 3723
rect 51077 3683 51135 3689
rect 51718 3680 51724 3732
rect 51776 3720 51782 3732
rect 51813 3723 51871 3729
rect 51813 3720 51825 3723
rect 51776 3692 51825 3720
rect 51776 3680 51782 3692
rect 51813 3689 51825 3692
rect 51859 3689 51871 3723
rect 51813 3683 51871 3689
rect 51902 3680 51908 3732
rect 51960 3720 51966 3732
rect 51960 3692 55168 3720
rect 51960 3680 51966 3692
rect 25406 3612 25412 3664
rect 25464 3652 25470 3664
rect 26970 3652 26976 3664
rect 25464 3624 26976 3652
rect 25464 3612 25470 3624
rect 26970 3612 26976 3624
rect 27028 3612 27034 3664
rect 27246 3612 27252 3664
rect 27304 3652 27310 3664
rect 32490 3652 32496 3664
rect 27304 3624 32496 3652
rect 27304 3612 27310 3624
rect 32490 3612 32496 3624
rect 32548 3612 32554 3664
rect 32674 3652 32680 3664
rect 32635 3624 32680 3652
rect 32674 3612 32680 3624
rect 32732 3612 32738 3664
rect 32950 3612 32956 3664
rect 33008 3652 33014 3664
rect 41230 3652 41236 3664
rect 33008 3624 41236 3652
rect 33008 3612 33014 3624
rect 41230 3612 41236 3624
rect 41288 3612 41294 3664
rect 41340 3624 45600 3652
rect 24544 3556 25176 3584
rect 24544 3544 24550 3556
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 35802 3584 35808 3596
rect 25556 3556 35808 3584
rect 25556 3544 25562 3556
rect 35802 3544 35808 3556
rect 35860 3544 35866 3596
rect 35894 3544 35900 3596
rect 35952 3584 35958 3596
rect 36354 3584 36360 3596
rect 35952 3556 36360 3584
rect 35952 3544 35958 3556
rect 36354 3544 36360 3556
rect 36412 3544 36418 3596
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 41340 3584 41368 3624
rect 37424 3556 41368 3584
rect 41509 3587 41567 3593
rect 37424 3544 37430 3556
rect 41509 3553 41521 3587
rect 41555 3584 41567 3587
rect 41966 3584 41972 3596
rect 41555 3556 41972 3584
rect 41555 3553 41567 3556
rect 41509 3547 41567 3553
rect 41966 3544 41972 3556
rect 42024 3544 42030 3596
rect 42058 3544 42064 3596
rect 42116 3584 42122 3596
rect 42978 3584 42984 3596
rect 42116 3556 42984 3584
rect 42116 3544 42122 3556
rect 42978 3544 42984 3556
rect 43036 3544 43042 3596
rect 43070 3544 43076 3596
rect 43128 3584 43134 3596
rect 43349 3587 43407 3593
rect 43349 3584 43361 3587
rect 43128 3556 43361 3584
rect 43128 3544 43134 3556
rect 43349 3553 43361 3556
rect 43395 3553 43407 3587
rect 44450 3584 44456 3596
rect 43349 3547 43407 3553
rect 43916 3556 44456 3584
rect 21177 3519 21235 3525
rect 21177 3485 21189 3519
rect 21223 3485 21235 3519
rect 21177 3479 21235 3485
rect 21545 3519 21603 3525
rect 21545 3485 21557 3519
rect 21591 3485 21603 3519
rect 21545 3479 21603 3485
rect 23017 3519 23075 3525
rect 23017 3485 23029 3519
rect 23063 3516 23075 3519
rect 24581 3519 24639 3525
rect 23063 3488 23520 3516
rect 23063 3485 23075 3488
rect 23017 3479 23075 3485
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 17129 3451 17187 3457
rect 17129 3448 17141 3451
rect 14608 3420 17141 3448
rect 14608 3408 14614 3420
rect 17129 3417 17141 3420
rect 17175 3417 17187 3451
rect 17129 3411 17187 3417
rect 17310 3408 17316 3460
rect 17368 3448 17374 3460
rect 20898 3448 20904 3460
rect 17368 3420 20904 3448
rect 17368 3408 17374 3420
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 21082 3380 21088 3392
rect 14476 3352 21088 3380
rect 21082 3340 21088 3352
rect 21140 3340 21146 3392
rect 21192 3380 21220 3479
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 22373 3451 22431 3457
rect 22373 3448 22385 3451
rect 21876 3420 22385 3448
rect 21876 3408 21882 3420
rect 22373 3417 22385 3420
rect 22419 3417 22431 3451
rect 22373 3411 22431 3417
rect 22002 3380 22008 3392
rect 21192 3352 22008 3380
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 23492 3389 23520 3488
rect 24581 3485 24593 3519
rect 24627 3516 24639 3519
rect 25038 3516 25044 3528
rect 24627 3488 25044 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 25038 3476 25044 3488
rect 25096 3476 25102 3528
rect 27525 3519 27583 3525
rect 27525 3485 27537 3519
rect 27571 3516 27583 3519
rect 27982 3516 27988 3528
rect 27571 3488 27988 3516
rect 27571 3485 27583 3488
rect 27525 3479 27583 3485
rect 27982 3476 27988 3488
rect 28040 3476 28046 3528
rect 29181 3519 29239 3525
rect 29181 3485 29193 3519
rect 29227 3516 29239 3519
rect 29365 3519 29423 3525
rect 29365 3516 29377 3519
rect 29227 3488 29377 3516
rect 29227 3485 29239 3488
rect 29181 3479 29239 3485
rect 29365 3485 29377 3488
rect 29411 3485 29423 3519
rect 37001 3519 37059 3525
rect 37001 3516 37013 3519
rect 29365 3479 29423 3485
rect 29472 3488 37013 3516
rect 25498 3408 25504 3460
rect 25556 3448 25562 3460
rect 26881 3451 26939 3457
rect 26881 3448 26893 3451
rect 25556 3420 26893 3448
rect 25556 3408 25562 3420
rect 26881 3417 26893 3420
rect 26927 3417 26939 3451
rect 26881 3411 26939 3417
rect 27062 3408 27068 3460
rect 27120 3448 27126 3460
rect 28537 3451 28595 3457
rect 28537 3448 28549 3451
rect 27120 3420 28549 3448
rect 27120 3408 27126 3420
rect 28537 3417 28549 3420
rect 28583 3417 28595 3451
rect 28537 3411 28595 3417
rect 23477 3383 23535 3389
rect 23477 3349 23489 3383
rect 23523 3380 23535 3383
rect 25682 3380 25688 3392
rect 23523 3352 25688 3380
rect 23523 3349 23535 3352
rect 23477 3343 23535 3349
rect 25682 3340 25688 3352
rect 25740 3340 25746 3392
rect 25866 3380 25872 3392
rect 25827 3352 25872 3380
rect 25866 3340 25872 3352
rect 25924 3340 25930 3392
rect 26145 3383 26203 3389
rect 26145 3349 26157 3383
rect 26191 3380 26203 3383
rect 29472 3380 29500 3488
rect 37001 3485 37013 3488
rect 37047 3485 37059 3519
rect 37458 3516 37464 3528
rect 37419 3488 37464 3516
rect 37001 3479 37059 3485
rect 37458 3476 37464 3488
rect 37516 3516 37522 3528
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 37516 3488 38025 3516
rect 37516 3476 37522 3488
rect 38013 3485 38025 3488
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 38102 3476 38108 3528
rect 38160 3516 38166 3528
rect 39850 3516 39856 3528
rect 38160 3488 39856 3516
rect 38160 3476 38166 3488
rect 39850 3476 39856 3488
rect 39908 3476 39914 3528
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40000 3488 41552 3516
rect 40000 3476 40006 3488
rect 29546 3408 29552 3460
rect 29604 3448 29610 3460
rect 41046 3448 41052 3460
rect 29604 3420 41052 3448
rect 29604 3408 29610 3420
rect 41046 3408 41052 3420
rect 41104 3408 41110 3460
rect 41414 3448 41420 3460
rect 41156 3420 41420 3448
rect 26191 3352 29500 3380
rect 26191 3349 26203 3352
rect 26145 3343 26203 3349
rect 29638 3340 29644 3392
rect 29696 3380 29702 3392
rect 34606 3380 34612 3392
rect 29696 3352 34612 3380
rect 29696 3340 29702 3352
rect 34606 3340 34612 3352
rect 34664 3340 34670 3392
rect 34698 3340 34704 3392
rect 34756 3380 34762 3392
rect 41156 3380 41184 3420
rect 41414 3408 41420 3420
rect 41472 3408 41478 3460
rect 41524 3448 41552 3488
rect 41598 3476 41604 3528
rect 41656 3516 41662 3528
rect 43530 3516 43536 3528
rect 41656 3488 43536 3516
rect 41656 3476 41662 3488
rect 43530 3476 43536 3488
rect 43588 3476 43594 3528
rect 43916 3525 43944 3556
rect 44450 3544 44456 3556
rect 44508 3544 44514 3596
rect 44542 3544 44548 3596
rect 44600 3584 44606 3596
rect 45462 3584 45468 3596
rect 44600 3556 45468 3584
rect 44600 3544 44606 3556
rect 45462 3544 45468 3556
rect 45520 3544 45526 3596
rect 45572 3584 45600 3624
rect 45646 3612 45652 3664
rect 45704 3652 45710 3664
rect 46290 3652 46296 3664
rect 45704 3624 46296 3652
rect 45704 3612 45710 3624
rect 46290 3612 46296 3624
rect 46348 3612 46354 3664
rect 49053 3655 49111 3661
rect 49053 3652 49065 3655
rect 46400 3624 49065 3652
rect 46400 3584 46428 3624
rect 49053 3621 49065 3624
rect 49099 3621 49111 3655
rect 49053 3615 49111 3621
rect 49418 3612 49424 3664
rect 49476 3652 49482 3664
rect 51994 3652 52000 3664
rect 49476 3624 52000 3652
rect 49476 3612 49482 3624
rect 51994 3612 52000 3624
rect 52052 3612 52058 3664
rect 54754 3652 54760 3664
rect 52104 3624 54760 3652
rect 46845 3587 46903 3593
rect 46845 3584 46857 3587
rect 45572 3556 46428 3584
rect 46676 3556 46857 3584
rect 43901 3519 43959 3525
rect 43901 3485 43913 3519
rect 43947 3485 43959 3519
rect 45649 3519 45707 3525
rect 45649 3516 45661 3519
rect 43901 3479 43959 3485
rect 44008 3488 45661 3516
rect 41874 3448 41880 3460
rect 41524 3420 41880 3448
rect 41874 3408 41880 3420
rect 41932 3408 41938 3460
rect 42334 3408 42340 3460
rect 42392 3448 42398 3460
rect 44008 3448 44036 3488
rect 45649 3485 45661 3488
rect 45695 3485 45707 3519
rect 45830 3516 45836 3528
rect 45791 3488 45836 3516
rect 45649 3479 45707 3485
rect 45830 3476 45836 3488
rect 45888 3476 45894 3528
rect 46106 3516 46112 3528
rect 46067 3488 46112 3516
rect 46106 3476 46112 3488
rect 46164 3476 46170 3528
rect 46477 3519 46535 3525
rect 46477 3485 46489 3519
rect 46523 3516 46535 3519
rect 46676 3516 46704 3556
rect 46845 3553 46857 3556
rect 46891 3584 46903 3587
rect 51074 3584 51080 3596
rect 46891 3556 51080 3584
rect 46891 3553 46903 3556
rect 46845 3547 46903 3553
rect 51074 3544 51080 3556
rect 51132 3544 51138 3596
rect 52104 3584 52132 3624
rect 54754 3612 54760 3624
rect 54812 3612 54818 3664
rect 55140 3652 55168 3692
rect 55306 3680 55312 3732
rect 55364 3720 55370 3732
rect 55401 3723 55459 3729
rect 55401 3720 55413 3723
rect 55364 3692 55413 3720
rect 55364 3680 55370 3692
rect 55401 3689 55413 3692
rect 55447 3689 55459 3723
rect 57238 3720 57244 3732
rect 55401 3683 55459 3689
rect 55508 3692 57244 3720
rect 55508 3652 55536 3692
rect 57238 3680 57244 3692
rect 57296 3680 57302 3732
rect 58250 3720 58256 3732
rect 58211 3692 58256 3720
rect 58250 3680 58256 3692
rect 58308 3680 58314 3732
rect 58437 3723 58495 3729
rect 58437 3689 58449 3723
rect 58483 3720 58495 3723
rect 58710 3720 58716 3732
rect 58483 3692 58716 3720
rect 58483 3689 58495 3692
rect 58437 3683 58495 3689
rect 58710 3680 58716 3692
rect 58768 3680 58774 3732
rect 60642 3720 60648 3732
rect 58820 3692 60648 3720
rect 55140 3624 55536 3652
rect 55674 3612 55680 3664
rect 55732 3652 55738 3664
rect 56045 3655 56103 3661
rect 56045 3652 56057 3655
rect 55732 3624 56057 3652
rect 55732 3612 55738 3624
rect 56045 3621 56057 3624
rect 56091 3621 56103 3655
rect 56045 3615 56103 3621
rect 56410 3612 56416 3664
rect 56468 3652 56474 3664
rect 58820 3652 58848 3692
rect 60642 3680 60648 3692
rect 60700 3680 60706 3732
rect 60734 3680 60740 3732
rect 60792 3720 60798 3732
rect 61289 3723 61347 3729
rect 61289 3720 61301 3723
rect 60792 3692 61301 3720
rect 60792 3680 60798 3692
rect 61289 3689 61301 3692
rect 61335 3689 61347 3723
rect 61289 3683 61347 3689
rect 61841 3723 61899 3729
rect 61841 3689 61853 3723
rect 61887 3720 61899 3723
rect 83734 3720 83740 3732
rect 61887 3692 83740 3720
rect 61887 3689 61899 3692
rect 61841 3683 61899 3689
rect 83734 3680 83740 3692
rect 83792 3680 83798 3732
rect 89162 3720 89168 3732
rect 89123 3692 89168 3720
rect 89162 3680 89168 3692
rect 89220 3720 89226 3732
rect 92566 3720 92572 3732
rect 89220 3692 92572 3720
rect 89220 3680 89226 3692
rect 92566 3680 92572 3692
rect 92624 3680 92630 3732
rect 92661 3723 92719 3729
rect 92661 3689 92673 3723
rect 92707 3720 92719 3723
rect 93210 3720 93216 3732
rect 92707 3692 93216 3720
rect 92707 3689 92719 3692
rect 92661 3683 92719 3689
rect 56468 3624 58848 3652
rect 56468 3612 56474 3624
rect 61102 3612 61108 3664
rect 61160 3652 61166 3664
rect 61749 3655 61807 3661
rect 61749 3652 61761 3655
rect 61160 3624 61761 3652
rect 61160 3612 61166 3624
rect 61749 3621 61761 3624
rect 61795 3652 61807 3655
rect 63586 3652 63592 3664
rect 61795 3624 63592 3652
rect 61795 3621 61807 3624
rect 61749 3615 61807 3621
rect 63586 3612 63592 3624
rect 63644 3612 63650 3664
rect 63862 3652 63868 3664
rect 63823 3624 63868 3652
rect 63862 3612 63868 3624
rect 63920 3612 63926 3664
rect 64049 3655 64107 3661
rect 64049 3621 64061 3655
rect 64095 3652 64107 3655
rect 68830 3652 68836 3664
rect 64095 3624 68836 3652
rect 64095 3621 64107 3624
rect 64049 3615 64107 3621
rect 68830 3612 68836 3624
rect 68888 3612 68894 3664
rect 69477 3655 69535 3661
rect 69477 3621 69489 3655
rect 69523 3652 69535 3655
rect 70578 3652 70584 3664
rect 69523 3624 70584 3652
rect 69523 3621 69535 3624
rect 69477 3615 69535 3621
rect 52362 3584 52368 3596
rect 51184 3556 52132 3584
rect 52323 3556 52368 3584
rect 46523 3488 46704 3516
rect 46523 3485 46535 3488
rect 46477 3479 46535 3485
rect 46750 3476 46756 3528
rect 46808 3516 46814 3528
rect 48866 3516 48872 3528
rect 46808 3488 48728 3516
rect 48827 3488 48872 3516
rect 46808 3476 46814 3488
rect 42392 3420 44036 3448
rect 42392 3408 42398 3420
rect 44082 3408 44088 3460
rect 44140 3448 44146 3460
rect 45462 3448 45468 3460
rect 44140 3420 45468 3448
rect 44140 3408 44146 3420
rect 45462 3408 45468 3420
rect 45520 3408 45526 3460
rect 46198 3448 46204 3460
rect 45572 3420 46204 3448
rect 34756 3352 41184 3380
rect 34756 3340 34762 3352
rect 41230 3340 41236 3392
rect 41288 3380 41294 3392
rect 43438 3380 43444 3392
rect 41288 3352 43444 3380
rect 41288 3340 41294 3352
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 43530 3340 43536 3392
rect 43588 3380 43594 3392
rect 45572 3380 45600 3420
rect 46198 3408 46204 3420
rect 46256 3408 46262 3460
rect 46290 3408 46296 3460
rect 46348 3448 46354 3460
rect 48225 3451 48283 3457
rect 48225 3448 48237 3451
rect 46348 3420 48237 3448
rect 46348 3408 46354 3420
rect 48225 3417 48237 3420
rect 48271 3417 48283 3451
rect 48590 3448 48596 3460
rect 48225 3411 48283 3417
rect 48332 3420 48596 3448
rect 43588 3352 45600 3380
rect 45649 3383 45707 3389
rect 43588 3340 43594 3352
rect 45649 3349 45661 3383
rect 45695 3380 45707 3383
rect 48332 3380 48360 3420
rect 48590 3408 48596 3420
rect 48648 3408 48654 3460
rect 48700 3448 48728 3488
rect 48866 3476 48872 3488
rect 48924 3516 48930 3528
rect 49237 3519 49295 3525
rect 49237 3516 49249 3519
rect 48924 3488 49249 3516
rect 48924 3476 48930 3488
rect 49237 3485 49249 3488
rect 49283 3485 49295 3519
rect 49237 3479 49295 3485
rect 49513 3519 49571 3525
rect 49513 3485 49525 3519
rect 49559 3516 49571 3519
rect 51184 3516 51212 3556
rect 52362 3544 52368 3556
rect 52420 3544 52426 3596
rect 57146 3584 57152 3596
rect 55048 3556 57152 3584
rect 49559 3488 51212 3516
rect 51445 3519 51503 3525
rect 49559 3485 49571 3488
rect 49513 3479 49571 3485
rect 51445 3485 51457 3519
rect 51491 3516 51503 3519
rect 51721 3519 51779 3525
rect 51721 3516 51733 3519
rect 51491 3488 51733 3516
rect 51491 3485 51503 3488
rect 51445 3479 51503 3485
rect 51721 3485 51733 3488
rect 51767 3485 51779 3519
rect 51721 3479 51779 3485
rect 51810 3476 51816 3528
rect 51868 3516 51874 3528
rect 54018 3516 54024 3528
rect 51868 3488 54024 3516
rect 51868 3476 51874 3488
rect 54018 3476 54024 3488
rect 54076 3476 54082 3528
rect 55048 3525 55076 3556
rect 57146 3544 57152 3556
rect 57204 3544 57210 3596
rect 60550 3544 60556 3596
rect 60608 3584 60614 3596
rect 63034 3584 63040 3596
rect 60608 3556 63040 3584
rect 60608 3544 60614 3556
rect 63034 3544 63040 3556
rect 63092 3544 63098 3596
rect 63218 3544 63224 3596
rect 63276 3584 63282 3596
rect 63313 3587 63371 3593
rect 63313 3584 63325 3587
rect 63276 3556 63325 3584
rect 63276 3544 63282 3556
rect 63313 3553 63325 3556
rect 63359 3584 63371 3587
rect 65242 3584 65248 3596
rect 63359 3556 65248 3584
rect 63359 3553 63371 3556
rect 63313 3547 63371 3553
rect 65242 3544 65248 3556
rect 65300 3544 65306 3596
rect 68097 3587 68155 3593
rect 68097 3584 68109 3587
rect 67560 3556 68109 3584
rect 54297 3519 54355 3525
rect 54297 3485 54309 3519
rect 54343 3516 54355 3519
rect 55033 3519 55091 3525
rect 55033 3516 55045 3519
rect 54343 3488 55045 3516
rect 54343 3485 54355 3488
rect 54297 3479 54355 3485
rect 55033 3485 55045 3488
rect 55079 3485 55091 3519
rect 55033 3479 55091 3485
rect 55953 3519 56011 3525
rect 55953 3485 55965 3519
rect 55999 3516 56011 3519
rect 56318 3516 56324 3528
rect 55999 3488 56324 3516
rect 55999 3485 56011 3488
rect 55953 3479 56011 3485
rect 56318 3476 56324 3488
rect 56376 3516 56382 3528
rect 56413 3519 56471 3525
rect 56413 3516 56425 3519
rect 56376 3488 56425 3516
rect 56376 3476 56382 3488
rect 56413 3485 56425 3488
rect 56459 3485 56471 3519
rect 56413 3479 56471 3485
rect 58161 3519 58219 3525
rect 58161 3485 58173 3519
rect 58207 3516 58219 3519
rect 58437 3519 58495 3525
rect 58437 3516 58449 3519
rect 58207 3488 58449 3516
rect 58207 3485 58219 3488
rect 58161 3479 58219 3485
rect 58437 3485 58449 3488
rect 58483 3485 58495 3519
rect 60090 3516 60096 3528
rect 58437 3479 58495 3485
rect 58820 3488 60096 3516
rect 48958 3448 48964 3460
rect 48700 3420 48964 3448
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 49053 3451 49111 3457
rect 49053 3417 49065 3451
rect 49099 3448 49111 3451
rect 54389 3451 54447 3457
rect 54389 3448 54401 3451
rect 49099 3420 54401 3448
rect 49099 3417 49111 3420
rect 49053 3411 49111 3417
rect 54389 3417 54401 3420
rect 54435 3417 54447 3451
rect 54389 3411 54447 3417
rect 54478 3408 54484 3460
rect 54536 3448 54542 3460
rect 55858 3448 55864 3460
rect 54536 3420 55864 3448
rect 54536 3408 54542 3420
rect 55858 3408 55864 3420
rect 55916 3408 55922 3460
rect 56686 3408 56692 3460
rect 56744 3448 56750 3460
rect 58820 3448 58848 3488
rect 60090 3476 60096 3488
rect 60148 3476 60154 3528
rect 61105 3519 61163 3525
rect 61105 3485 61117 3519
rect 61151 3516 61163 3519
rect 61197 3519 61255 3525
rect 61197 3516 61209 3519
rect 61151 3488 61209 3516
rect 61151 3485 61163 3488
rect 61105 3479 61163 3485
rect 61197 3485 61209 3488
rect 61243 3516 61255 3519
rect 62758 3516 62764 3528
rect 61243 3488 62764 3516
rect 61243 3485 61255 3488
rect 61197 3479 61255 3485
rect 62758 3476 62764 3488
rect 62816 3476 62822 3528
rect 62853 3519 62911 3525
rect 62853 3485 62865 3519
rect 62899 3516 62911 3519
rect 62942 3516 62948 3528
rect 62899 3488 62948 3516
rect 62899 3485 62911 3488
rect 62853 3479 62911 3485
rect 62942 3476 62948 3488
rect 63000 3476 63006 3528
rect 67560 3525 67588 3556
rect 68097 3553 68109 3556
rect 68143 3584 68155 3587
rect 69014 3584 69020 3596
rect 68143 3556 69020 3584
rect 68143 3553 68155 3556
rect 68097 3547 68155 3553
rect 69014 3544 69020 3556
rect 69072 3544 69078 3596
rect 63773 3519 63831 3525
rect 63773 3485 63785 3519
rect 63819 3516 63831 3519
rect 67545 3519 67603 3525
rect 63819 3488 64368 3516
rect 63819 3485 63831 3488
rect 63773 3479 63831 3485
rect 62022 3448 62028 3460
rect 56744 3420 58848 3448
rect 58912 3420 62028 3448
rect 56744 3408 56750 3420
rect 45695 3352 48360 3380
rect 45695 3349 45707 3352
rect 45649 3343 45707 3349
rect 48406 3340 48412 3392
rect 48464 3380 48470 3392
rect 52178 3380 52184 3392
rect 48464 3352 52184 3380
rect 48464 3340 48470 3352
rect 52178 3340 52184 3352
rect 52236 3340 52242 3392
rect 53282 3340 53288 3392
rect 53340 3380 53346 3392
rect 55950 3380 55956 3392
rect 53340 3352 55956 3380
rect 53340 3340 53346 3352
rect 55950 3340 55956 3352
rect 56008 3340 56014 3392
rect 56962 3380 56968 3392
rect 56923 3352 56968 3380
rect 56962 3340 56968 3352
rect 57020 3340 57026 3392
rect 57054 3340 57060 3392
rect 57112 3380 57118 3392
rect 58912 3380 58940 3420
rect 62022 3408 62028 3420
rect 62080 3408 62086 3460
rect 62117 3451 62175 3457
rect 62117 3417 62129 3451
rect 62163 3448 62175 3451
rect 62206 3448 62212 3460
rect 62163 3420 62212 3448
rect 62163 3417 62175 3420
rect 62117 3411 62175 3417
rect 62206 3408 62212 3420
rect 62264 3448 62270 3460
rect 64230 3448 64236 3460
rect 62264 3420 64236 3448
rect 62264 3408 62270 3420
rect 64230 3408 64236 3420
rect 64288 3408 64294 3460
rect 57112 3352 58940 3380
rect 59449 3383 59507 3389
rect 57112 3340 57118 3352
rect 59449 3349 59461 3383
rect 59495 3380 59507 3383
rect 60366 3380 60372 3392
rect 59495 3352 60372 3380
rect 59495 3349 59507 3352
rect 59449 3343 59507 3349
rect 60366 3340 60372 3352
rect 60424 3340 60430 3392
rect 60458 3340 60464 3392
rect 60516 3380 60522 3392
rect 61841 3383 61899 3389
rect 61841 3380 61853 3383
rect 60516 3352 61853 3380
rect 60516 3340 60522 3352
rect 61841 3349 61853 3352
rect 61887 3349 61899 3383
rect 62482 3380 62488 3392
rect 62443 3352 62488 3380
rect 61841 3343 61899 3349
rect 62482 3340 62488 3352
rect 62540 3340 62546 3392
rect 62758 3340 62764 3392
rect 62816 3380 62822 3392
rect 64340 3389 64368 3488
rect 67545 3485 67557 3519
rect 67591 3485 67603 3519
rect 67545 3479 67603 3485
rect 67634 3476 67640 3528
rect 67692 3516 67698 3528
rect 68925 3519 68983 3525
rect 67692 3488 67737 3516
rect 67692 3476 67698 3488
rect 68925 3485 68937 3519
rect 68971 3516 68983 3519
rect 69492 3516 69520 3615
rect 70578 3612 70584 3624
rect 70636 3612 70642 3664
rect 71774 3652 71780 3664
rect 71735 3624 71780 3652
rect 71774 3612 71780 3624
rect 71832 3612 71838 3664
rect 71958 3612 71964 3664
rect 72016 3652 72022 3664
rect 72237 3655 72295 3661
rect 72237 3652 72249 3655
rect 72016 3624 72249 3652
rect 72016 3612 72022 3624
rect 72237 3621 72249 3624
rect 72283 3652 72295 3655
rect 72694 3652 72700 3664
rect 72283 3624 72700 3652
rect 72283 3621 72295 3624
rect 72237 3615 72295 3621
rect 72694 3612 72700 3624
rect 72752 3612 72758 3664
rect 72878 3652 72884 3664
rect 72804 3624 72884 3652
rect 72142 3584 72148 3596
rect 68971 3488 69520 3516
rect 69584 3556 72148 3584
rect 68971 3485 68983 3488
rect 68925 3479 68983 3485
rect 67450 3408 67456 3460
rect 67508 3448 67514 3460
rect 69584 3448 69612 3556
rect 72142 3544 72148 3556
rect 72200 3544 72206 3596
rect 72804 3593 72832 3624
rect 72878 3612 72884 3624
rect 72936 3612 72942 3664
rect 72970 3612 72976 3664
rect 73028 3652 73034 3664
rect 78214 3652 78220 3664
rect 73028 3624 78220 3652
rect 73028 3612 73034 3624
rect 78214 3612 78220 3624
rect 78272 3612 78278 3664
rect 89438 3652 89444 3664
rect 89399 3624 89444 3652
rect 89438 3612 89444 3624
rect 89496 3612 89502 3664
rect 90269 3655 90327 3661
rect 90269 3621 90281 3655
rect 90315 3652 90327 3655
rect 91094 3652 91100 3664
rect 90315 3624 91100 3652
rect 90315 3621 90327 3624
rect 90269 3615 90327 3621
rect 91094 3612 91100 3624
rect 91152 3652 91158 3664
rect 91738 3652 91744 3664
rect 91152 3624 91744 3652
rect 91152 3612 91158 3624
rect 91738 3612 91744 3624
rect 91796 3612 91802 3664
rect 72789 3587 72847 3593
rect 72789 3553 72801 3587
rect 72835 3553 72847 3587
rect 72789 3547 72847 3553
rect 73062 3544 73068 3596
rect 73120 3584 73126 3596
rect 88426 3584 88432 3596
rect 73120 3556 88432 3584
rect 73120 3544 73126 3556
rect 88426 3544 88432 3556
rect 88484 3544 88490 3596
rect 70673 3519 70731 3525
rect 70673 3485 70685 3519
rect 70719 3485 70731 3519
rect 71130 3516 71136 3528
rect 70673 3479 70731 3485
rect 70780 3488 71136 3516
rect 67508 3420 69612 3448
rect 67508 3408 67514 3420
rect 64049 3383 64107 3389
rect 64049 3380 64061 3383
rect 62816 3352 64061 3380
rect 62816 3340 62822 3352
rect 64049 3349 64061 3352
rect 64095 3349 64107 3383
rect 64049 3343 64107 3349
rect 64325 3383 64383 3389
rect 64325 3349 64337 3383
rect 64371 3380 64383 3383
rect 66070 3380 66076 3392
rect 64371 3352 66076 3380
rect 64371 3349 64383 3352
rect 64325 3343 64383 3349
rect 66070 3340 66076 3352
rect 66128 3340 66134 3392
rect 66346 3340 66352 3392
rect 66404 3380 66410 3392
rect 66533 3383 66591 3389
rect 66533 3380 66545 3383
rect 66404 3352 66545 3380
rect 66404 3340 66410 3352
rect 66533 3349 66545 3352
rect 66579 3349 66591 3383
rect 66533 3343 66591 3349
rect 68465 3383 68523 3389
rect 68465 3349 68477 3383
rect 68511 3380 68523 3383
rect 68738 3380 68744 3392
rect 68511 3352 68744 3380
rect 68511 3349 68523 3352
rect 68465 3343 68523 3349
rect 68738 3340 68744 3352
rect 68796 3340 68802 3392
rect 69017 3383 69075 3389
rect 69017 3349 69029 3383
rect 69063 3380 69075 3383
rect 69106 3380 69112 3392
rect 69063 3352 69112 3380
rect 69063 3349 69075 3352
rect 69017 3343 69075 3349
rect 69106 3340 69112 3352
rect 69164 3340 69170 3392
rect 70029 3383 70087 3389
rect 70029 3349 70041 3383
rect 70075 3380 70087 3383
rect 70394 3380 70400 3392
rect 70075 3352 70400 3380
rect 70075 3349 70087 3352
rect 70029 3343 70087 3349
rect 70394 3340 70400 3352
rect 70452 3340 70458 3392
rect 70688 3380 70716 3479
rect 70780 3457 70808 3488
rect 71130 3476 71136 3488
rect 71188 3476 71194 3528
rect 71685 3519 71743 3525
rect 71685 3485 71697 3519
rect 71731 3516 71743 3519
rect 71961 3519 72019 3525
rect 71961 3516 71973 3519
rect 71731 3488 71973 3516
rect 71731 3485 71743 3488
rect 71685 3479 71743 3485
rect 71961 3485 71973 3488
rect 72007 3485 72019 3519
rect 71961 3479 72019 3485
rect 72326 3476 72332 3528
rect 72384 3516 72390 3528
rect 72697 3519 72755 3525
rect 72697 3516 72709 3519
rect 72384 3488 72709 3516
rect 72384 3476 72390 3488
rect 72697 3485 72709 3488
rect 72743 3516 72755 3519
rect 73157 3519 73215 3525
rect 73157 3516 73169 3519
rect 72743 3488 73169 3516
rect 72743 3485 72755 3488
rect 72697 3479 72755 3485
rect 73157 3485 73169 3488
rect 73203 3485 73215 3519
rect 73157 3479 73215 3485
rect 73338 3476 73344 3528
rect 73396 3516 73402 3528
rect 78950 3516 78956 3528
rect 73396 3488 78956 3516
rect 73396 3476 73402 3488
rect 78950 3476 78956 3488
rect 79008 3476 79014 3528
rect 88245 3519 88303 3525
rect 88245 3485 88257 3519
rect 88291 3516 88303 3519
rect 89349 3519 89407 3525
rect 88291 3488 88840 3516
rect 88291 3485 88303 3488
rect 88245 3479 88303 3485
rect 70765 3451 70823 3457
rect 70765 3417 70777 3451
rect 70811 3417 70823 3451
rect 70765 3411 70823 3417
rect 70946 3408 70952 3460
rect 71004 3448 71010 3460
rect 71225 3451 71283 3457
rect 71225 3448 71237 3451
rect 71004 3420 71237 3448
rect 71004 3408 71010 3420
rect 71225 3417 71237 3420
rect 71271 3448 71283 3451
rect 71590 3448 71596 3460
rect 71271 3420 71596 3448
rect 71271 3417 71283 3420
rect 71225 3411 71283 3417
rect 71590 3408 71596 3420
rect 71648 3408 71654 3460
rect 72050 3448 72056 3460
rect 71884 3420 72056 3448
rect 71501 3383 71559 3389
rect 71501 3380 71513 3383
rect 70688 3352 71513 3380
rect 71501 3349 71513 3352
rect 71547 3380 71559 3383
rect 71884 3380 71912 3420
rect 72050 3408 72056 3420
rect 72108 3408 72114 3460
rect 72418 3408 72424 3460
rect 72476 3448 72482 3460
rect 81894 3448 81900 3460
rect 72476 3420 81900 3448
rect 72476 3408 72482 3420
rect 81894 3408 81900 3420
rect 81952 3408 81958 3460
rect 88812 3392 88840 3488
rect 89349 3485 89361 3519
rect 89395 3485 89407 3519
rect 89349 3479 89407 3485
rect 90361 3519 90419 3525
rect 90361 3485 90373 3519
rect 90407 3516 90419 3519
rect 91741 3519 91799 3525
rect 90407 3488 90956 3516
rect 90407 3485 90419 3488
rect 90361 3479 90419 3485
rect 89364 3448 89392 3479
rect 89364 3420 89944 3448
rect 71547 3352 71912 3380
rect 71961 3383 72019 3389
rect 71547 3349 71559 3352
rect 71501 3343 71559 3349
rect 71961 3349 71973 3383
rect 72007 3380 72019 3383
rect 72605 3383 72663 3389
rect 72605 3380 72617 3383
rect 72007 3352 72617 3380
rect 72007 3349 72019 3352
rect 71961 3343 72019 3349
rect 72605 3349 72617 3352
rect 72651 3380 72663 3383
rect 73338 3380 73344 3392
rect 72651 3352 73344 3380
rect 72651 3349 72663 3352
rect 72605 3343 72663 3349
rect 73338 3340 73344 3352
rect 73396 3340 73402 3392
rect 73706 3380 73712 3392
rect 73667 3352 73712 3380
rect 73706 3340 73712 3352
rect 73764 3340 73770 3392
rect 73798 3340 73804 3392
rect 73856 3380 73862 3392
rect 85942 3380 85948 3392
rect 73856 3352 85948 3380
rect 73856 3340 73862 3352
rect 85942 3340 85948 3352
rect 86000 3340 86006 3392
rect 88334 3380 88340 3392
rect 88295 3352 88340 3380
rect 88334 3340 88340 3352
rect 88392 3340 88398 3392
rect 88794 3380 88800 3392
rect 88755 3352 88800 3380
rect 88794 3340 88800 3352
rect 88852 3340 88858 3392
rect 89916 3389 89944 3420
rect 89901 3383 89959 3389
rect 89901 3349 89913 3383
rect 89947 3380 89959 3383
rect 89990 3380 89996 3392
rect 89947 3352 89996 3380
rect 89947 3349 89959 3352
rect 89901 3343 89959 3349
rect 89990 3340 89996 3352
rect 90048 3340 90054 3392
rect 90450 3380 90456 3392
rect 90411 3352 90456 3380
rect 90450 3340 90456 3352
rect 90508 3340 90514 3392
rect 90928 3389 90956 3488
rect 91741 3485 91753 3519
rect 91787 3516 91799 3519
rect 92676 3516 92704 3683
rect 93210 3680 93216 3692
rect 93268 3680 93274 3732
rect 100570 3680 100576 3732
rect 100628 3720 100634 3732
rect 100628 3692 108344 3720
rect 100628 3680 100634 3692
rect 100018 3612 100024 3664
rect 100076 3652 100082 3664
rect 107930 3652 107936 3664
rect 100076 3624 107936 3652
rect 100076 3612 100082 3624
rect 107930 3612 107936 3624
rect 107988 3612 107994 3664
rect 100294 3544 100300 3596
rect 100352 3584 100358 3596
rect 108114 3584 108120 3596
rect 100352 3556 108120 3584
rect 100352 3544 100358 3556
rect 108114 3544 108120 3556
rect 108172 3544 108178 3596
rect 108316 3584 108344 3692
rect 108390 3680 108396 3732
rect 108448 3720 108454 3732
rect 113542 3720 113548 3732
rect 108448 3692 113548 3720
rect 108448 3680 108454 3692
rect 113542 3680 113548 3692
rect 113600 3680 113606 3732
rect 113634 3680 113640 3732
rect 113692 3720 113698 3732
rect 113821 3723 113879 3729
rect 113821 3720 113833 3723
rect 113692 3692 113833 3720
rect 113692 3680 113698 3692
rect 113821 3689 113833 3692
rect 113867 3720 113879 3723
rect 115750 3720 115756 3732
rect 113867 3692 115756 3720
rect 113867 3689 113879 3692
rect 113821 3683 113879 3689
rect 115750 3680 115756 3692
rect 115808 3680 115814 3732
rect 117498 3680 117504 3732
rect 117556 3720 117562 3732
rect 121917 3723 121975 3729
rect 121917 3720 121929 3723
rect 117556 3692 121929 3720
rect 117556 3680 117562 3692
rect 121917 3689 121929 3692
rect 121963 3689 121975 3723
rect 124950 3720 124956 3732
rect 124911 3692 124956 3720
rect 121917 3683 121975 3689
rect 124950 3680 124956 3692
rect 125008 3680 125014 3732
rect 125686 3680 125692 3732
rect 125744 3720 125750 3732
rect 126425 3723 126483 3729
rect 126425 3720 126437 3723
rect 125744 3692 126437 3720
rect 125744 3680 125750 3692
rect 126425 3689 126437 3692
rect 126471 3689 126483 3723
rect 126425 3683 126483 3689
rect 130841 3723 130899 3729
rect 130841 3689 130853 3723
rect 130887 3720 130899 3723
rect 131022 3720 131028 3732
rect 130887 3692 131028 3720
rect 130887 3689 130899 3692
rect 130841 3683 130899 3689
rect 131022 3680 131028 3692
rect 131080 3680 131086 3732
rect 133506 3720 133512 3732
rect 133467 3692 133512 3720
rect 133506 3680 133512 3692
rect 133564 3680 133570 3732
rect 143350 3680 143356 3732
rect 143408 3720 143414 3732
rect 164237 3723 164295 3729
rect 143408 3692 162164 3720
rect 143408 3680 143414 3692
rect 108942 3612 108948 3664
rect 109000 3652 109006 3664
rect 139946 3652 139952 3664
rect 109000 3624 139952 3652
rect 109000 3612 109006 3624
rect 139946 3612 139952 3624
rect 140004 3612 140010 3664
rect 146018 3652 146024 3664
rect 145979 3624 146024 3652
rect 146018 3612 146024 3624
rect 146076 3612 146082 3664
rect 149974 3652 149980 3664
rect 149935 3624 149980 3652
rect 149974 3612 149980 3624
rect 150032 3612 150038 3664
rect 150158 3612 150164 3664
rect 150216 3652 150222 3664
rect 150805 3655 150863 3661
rect 150805 3652 150817 3655
rect 150216 3624 150817 3652
rect 150216 3612 150222 3624
rect 150805 3621 150817 3624
rect 150851 3652 150863 3655
rect 152550 3652 152556 3664
rect 150851 3624 152556 3652
rect 150851 3621 150863 3624
rect 150805 3615 150863 3621
rect 152550 3612 152556 3624
rect 152608 3612 152614 3664
rect 162136 3652 162164 3692
rect 164237 3689 164249 3723
rect 164283 3720 164295 3723
rect 164418 3720 164424 3732
rect 164283 3692 164424 3720
rect 164283 3689 164295 3692
rect 164237 3683 164295 3689
rect 164418 3680 164424 3692
rect 164476 3680 164482 3732
rect 165522 3720 165528 3732
rect 165483 3692 165528 3720
rect 165522 3680 165528 3692
rect 165580 3680 165586 3732
rect 166718 3652 166724 3664
rect 162136 3624 166724 3652
rect 166718 3612 166724 3624
rect 166776 3612 166782 3664
rect 126606 3584 126612 3596
rect 108316 3556 126612 3584
rect 126606 3544 126612 3556
rect 126664 3544 126670 3596
rect 130194 3544 130200 3596
rect 130252 3584 130258 3596
rect 130289 3587 130347 3593
rect 130289 3584 130301 3587
rect 130252 3556 130301 3584
rect 130252 3544 130258 3556
rect 130289 3553 130301 3556
rect 130335 3584 130347 3587
rect 131574 3584 131580 3596
rect 130335 3556 131580 3584
rect 130335 3553 130347 3556
rect 130289 3547 130347 3553
rect 131574 3544 131580 3556
rect 131632 3544 131638 3596
rect 144730 3544 144736 3596
rect 144788 3584 144794 3596
rect 162302 3584 162308 3596
rect 144788 3556 162308 3584
rect 144788 3544 144794 3556
rect 162302 3544 162308 3556
rect 162360 3544 162366 3596
rect 102318 3516 102324 3528
rect 91787 3488 92704 3516
rect 102231 3488 102324 3516
rect 91787 3485 91799 3488
rect 91741 3479 91799 3485
rect 102318 3476 102324 3488
rect 102376 3516 102382 3528
rect 102781 3519 102839 3525
rect 102781 3516 102793 3519
rect 102376 3488 102793 3516
rect 102376 3476 102382 3488
rect 102781 3485 102793 3488
rect 102827 3485 102839 3519
rect 102781 3479 102839 3485
rect 102962 3476 102968 3528
rect 103020 3516 103026 3528
rect 108022 3516 108028 3528
rect 103020 3488 108028 3516
rect 103020 3476 103026 3488
rect 108022 3476 108028 3488
rect 108080 3476 108086 3528
rect 108206 3476 108212 3528
rect 108264 3516 108270 3528
rect 109218 3516 109224 3528
rect 108264 3488 109224 3516
rect 108264 3476 108270 3488
rect 109218 3476 109224 3488
rect 109276 3476 109282 3528
rect 109402 3476 109408 3528
rect 109460 3516 109466 3528
rect 114002 3516 114008 3528
rect 109460 3488 114008 3516
rect 109460 3476 109466 3488
rect 114002 3476 114008 3488
rect 114060 3476 114066 3528
rect 121730 3516 121736 3528
rect 114112 3488 121736 3516
rect 91833 3451 91891 3457
rect 91833 3417 91845 3451
rect 91879 3448 91891 3451
rect 94222 3448 94228 3460
rect 91879 3420 94228 3448
rect 91879 3417 91891 3420
rect 91833 3411 91891 3417
rect 94222 3408 94228 3420
rect 94280 3408 94286 3460
rect 100849 3451 100907 3457
rect 100849 3417 100861 3451
rect 100895 3448 100907 3451
rect 102226 3448 102232 3460
rect 100895 3420 102232 3448
rect 100895 3417 100907 3420
rect 100849 3411 100907 3417
rect 102226 3408 102232 3420
rect 102284 3448 102290 3460
rect 103149 3451 103207 3457
rect 103149 3448 103161 3451
rect 102284 3420 103161 3448
rect 102284 3408 102290 3420
rect 103149 3417 103161 3420
rect 103195 3417 103207 3451
rect 103149 3411 103207 3417
rect 106458 3408 106464 3460
rect 106516 3448 106522 3460
rect 106645 3451 106703 3457
rect 106645 3448 106657 3451
rect 106516 3420 106657 3448
rect 106516 3408 106522 3420
rect 106645 3417 106657 3420
rect 106691 3448 106703 3451
rect 106734 3448 106740 3460
rect 106691 3420 106740 3448
rect 106691 3417 106703 3420
rect 106645 3411 106703 3417
rect 106734 3408 106740 3420
rect 106792 3408 106798 3460
rect 107930 3408 107936 3460
rect 107988 3448 107994 3460
rect 108850 3448 108856 3460
rect 107988 3420 108856 3448
rect 107988 3408 107994 3420
rect 108850 3408 108856 3420
rect 108908 3408 108914 3460
rect 108942 3408 108948 3460
rect 109000 3448 109006 3460
rect 114112 3448 114140 3488
rect 121730 3476 121736 3488
rect 121788 3476 121794 3528
rect 121825 3519 121883 3525
rect 121825 3485 121837 3519
rect 121871 3516 121883 3519
rect 122101 3519 122159 3525
rect 122101 3516 122113 3519
rect 121871 3488 122113 3516
rect 121871 3485 121883 3488
rect 121825 3479 121883 3485
rect 122101 3485 122113 3488
rect 122147 3485 122159 3519
rect 122101 3479 122159 3485
rect 124861 3519 124919 3525
rect 124861 3485 124873 3519
rect 124907 3516 124919 3519
rect 124950 3516 124956 3528
rect 124907 3488 124956 3516
rect 124907 3485 124919 3488
rect 124861 3479 124919 3485
rect 124950 3476 124956 3488
rect 125008 3516 125014 3528
rect 125321 3519 125379 3525
rect 125321 3516 125333 3519
rect 125008 3488 125333 3516
rect 125008 3476 125014 3488
rect 125321 3485 125333 3488
rect 125367 3485 125379 3519
rect 125321 3479 125379 3485
rect 126333 3519 126391 3525
rect 126333 3485 126345 3519
rect 126379 3516 126391 3519
rect 126422 3516 126428 3528
rect 126379 3488 126428 3516
rect 126379 3485 126391 3488
rect 126333 3479 126391 3485
rect 126422 3476 126428 3488
rect 126480 3516 126486 3528
rect 129734 3516 129740 3528
rect 126480 3488 129740 3516
rect 126480 3476 126486 3488
rect 129734 3476 129740 3488
rect 129792 3476 129798 3528
rect 130749 3519 130807 3525
rect 130749 3485 130761 3519
rect 130795 3516 130807 3519
rect 131301 3519 131359 3525
rect 131301 3516 131313 3519
rect 130795 3488 131313 3516
rect 130795 3485 130807 3488
rect 130749 3479 130807 3485
rect 131301 3485 131313 3488
rect 131347 3516 131359 3519
rect 131942 3516 131948 3528
rect 131347 3488 131948 3516
rect 131347 3485 131359 3488
rect 131301 3479 131359 3485
rect 131942 3476 131948 3488
rect 132000 3476 132006 3528
rect 133417 3519 133475 3525
rect 133417 3485 133429 3519
rect 133463 3516 133475 3519
rect 133782 3516 133788 3528
rect 133463 3488 133788 3516
rect 133463 3485 133475 3488
rect 133417 3479 133475 3485
rect 133782 3476 133788 3488
rect 133840 3516 133846 3528
rect 133877 3519 133935 3525
rect 133877 3516 133889 3519
rect 133840 3488 133889 3516
rect 133840 3476 133846 3488
rect 133877 3485 133889 3488
rect 133923 3485 133935 3519
rect 133877 3479 133935 3485
rect 137094 3476 137100 3528
rect 137152 3516 137158 3528
rect 138661 3519 138719 3525
rect 138661 3516 138673 3519
rect 137152 3488 138673 3516
rect 137152 3476 137158 3488
rect 138661 3485 138673 3488
rect 138707 3516 138719 3519
rect 139121 3519 139179 3525
rect 139121 3516 139133 3519
rect 138707 3488 139133 3516
rect 138707 3485 138719 3488
rect 138661 3479 138719 3485
rect 139121 3485 139133 3488
rect 139167 3485 139179 3519
rect 139121 3479 139179 3485
rect 145929 3519 145987 3525
rect 145929 3485 145941 3519
rect 145975 3516 145987 3519
rect 146481 3519 146539 3525
rect 146481 3516 146493 3519
rect 145975 3488 146493 3516
rect 145975 3485 145987 3488
rect 145929 3479 145987 3485
rect 146481 3485 146493 3488
rect 146527 3516 146539 3519
rect 148134 3516 148140 3528
rect 146527 3488 148140 3516
rect 146527 3485 146539 3488
rect 146481 3479 146539 3485
rect 148134 3476 148140 3488
rect 148192 3476 148198 3528
rect 149885 3519 149943 3525
rect 149885 3485 149897 3519
rect 149931 3485 149943 3519
rect 149885 3479 149943 3485
rect 151541 3519 151599 3525
rect 151541 3485 151553 3519
rect 151587 3516 151599 3519
rect 151587 3488 152136 3516
rect 151587 3485 151599 3488
rect 151541 3479 151599 3485
rect 109000 3420 114140 3448
rect 109000 3408 109006 3420
rect 115014 3408 115020 3460
rect 115072 3448 115078 3460
rect 115072 3420 141464 3448
rect 115072 3408 115078 3420
rect 90913 3383 90971 3389
rect 90913 3349 90925 3383
rect 90959 3380 90971 3383
rect 91462 3380 91468 3392
rect 90959 3352 91468 3380
rect 90959 3349 90971 3352
rect 90913 3343 90971 3349
rect 91462 3340 91468 3352
rect 91520 3340 91526 3392
rect 92290 3380 92296 3392
rect 92251 3352 92296 3380
rect 92290 3340 92296 3352
rect 92348 3340 92354 3392
rect 100018 3340 100024 3392
rect 100076 3380 100082 3392
rect 102413 3383 102471 3389
rect 102413 3380 102425 3383
rect 100076 3352 102425 3380
rect 100076 3340 100082 3352
rect 102413 3349 102425 3352
rect 102459 3349 102471 3383
rect 103330 3380 103336 3392
rect 103291 3352 103336 3380
rect 102413 3343 102471 3349
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 103422 3340 103428 3392
rect 103480 3380 103486 3392
rect 107562 3380 107568 3392
rect 103480 3352 107568 3380
rect 103480 3340 103486 3352
rect 107562 3340 107568 3352
rect 107620 3340 107626 3392
rect 107746 3340 107752 3392
rect 107804 3380 107810 3392
rect 107841 3383 107899 3389
rect 107841 3380 107853 3383
rect 107804 3352 107853 3380
rect 107804 3340 107810 3352
rect 107841 3349 107853 3352
rect 107887 3380 107899 3383
rect 109862 3380 109868 3392
rect 107887 3352 109868 3380
rect 107887 3349 107899 3352
rect 107841 3343 107899 3349
rect 109862 3340 109868 3352
rect 109920 3340 109926 3392
rect 114830 3380 114836 3392
rect 114791 3352 114836 3380
rect 114830 3340 114836 3352
rect 114888 3340 114894 3392
rect 115842 3340 115848 3392
rect 115900 3380 115906 3392
rect 115937 3383 115995 3389
rect 115937 3380 115949 3383
rect 115900 3352 115949 3380
rect 115900 3340 115906 3352
rect 115937 3349 115949 3352
rect 115983 3380 115995 3383
rect 117958 3380 117964 3392
rect 115983 3352 117964 3380
rect 115983 3349 115995 3352
rect 115937 3343 115995 3349
rect 117958 3340 117964 3352
rect 118016 3340 118022 3392
rect 119617 3383 119675 3389
rect 119617 3349 119629 3383
rect 119663 3380 119675 3383
rect 120074 3380 120080 3392
rect 119663 3352 120080 3380
rect 119663 3349 119675 3352
rect 119617 3343 119675 3349
rect 120074 3340 120080 3352
rect 120132 3380 120138 3392
rect 121270 3380 121276 3392
rect 120132 3352 121276 3380
rect 120132 3340 120138 3352
rect 121270 3340 121276 3352
rect 121328 3340 121334 3392
rect 121638 3380 121644 3392
rect 121599 3352 121644 3380
rect 121638 3340 121644 3352
rect 121696 3340 121702 3392
rect 122101 3383 122159 3389
rect 122101 3349 122113 3383
rect 122147 3380 122159 3383
rect 122377 3383 122435 3389
rect 122377 3380 122389 3383
rect 122147 3352 122389 3380
rect 122147 3349 122159 3352
rect 122101 3343 122159 3349
rect 122377 3349 122389 3352
rect 122423 3380 122435 3383
rect 123478 3380 123484 3392
rect 122423 3352 123484 3380
rect 122423 3349 122435 3352
rect 122377 3343 122435 3349
rect 123478 3340 123484 3352
rect 123536 3340 123542 3392
rect 124582 3380 124588 3392
rect 124543 3352 124588 3380
rect 124582 3340 124588 3352
rect 124640 3340 124646 3392
rect 125594 3340 125600 3392
rect 125652 3380 125658 3392
rect 125781 3383 125839 3389
rect 125781 3380 125793 3383
rect 125652 3352 125793 3380
rect 125652 3340 125658 3352
rect 125781 3349 125793 3352
rect 125827 3380 125839 3383
rect 126330 3380 126336 3392
rect 125827 3352 126336 3380
rect 125827 3349 125839 3352
rect 125781 3343 125839 3349
rect 126330 3340 126336 3352
rect 126388 3340 126394 3392
rect 126882 3340 126888 3392
rect 126940 3380 126946 3392
rect 126977 3383 127035 3389
rect 126977 3380 126989 3383
rect 126940 3352 126989 3380
rect 126940 3340 126946 3352
rect 126977 3349 126989 3352
rect 127023 3380 127035 3383
rect 128630 3380 128636 3392
rect 127023 3352 128636 3380
rect 127023 3349 127035 3352
rect 126977 3343 127035 3349
rect 128630 3340 128636 3352
rect 128688 3340 128694 3392
rect 131298 3340 131304 3392
rect 131356 3380 131362 3392
rect 131669 3383 131727 3389
rect 131669 3380 131681 3383
rect 131356 3352 131681 3380
rect 131356 3340 131362 3352
rect 131669 3349 131681 3352
rect 131715 3380 131727 3383
rect 132310 3380 132316 3392
rect 131715 3352 132316 3380
rect 131715 3349 131727 3352
rect 131669 3343 131727 3349
rect 132310 3340 132316 3352
rect 132368 3340 132374 3392
rect 137278 3380 137284 3392
rect 137239 3352 137284 3380
rect 137278 3340 137284 3352
rect 137336 3340 137342 3392
rect 138750 3380 138756 3392
rect 138711 3352 138756 3380
rect 138750 3340 138756 3352
rect 138808 3340 138814 3392
rect 141436 3380 141464 3420
rect 142982 3408 142988 3460
rect 143040 3448 143046 3460
rect 149900 3448 149928 3479
rect 150437 3451 150495 3457
rect 150437 3448 150449 3451
rect 143040 3420 149836 3448
rect 149900 3420 150449 3448
rect 143040 3408 143046 3420
rect 144822 3380 144828 3392
rect 141436 3352 144828 3380
rect 144822 3340 144828 3352
rect 144880 3340 144886 3392
rect 148229 3383 148287 3389
rect 148229 3349 148241 3383
rect 148275 3380 148287 3383
rect 149054 3380 149060 3392
rect 148275 3352 149060 3380
rect 148275 3349 148287 3352
rect 148229 3343 148287 3349
rect 149054 3340 149060 3352
rect 149112 3340 149118 3392
rect 149808 3380 149836 3420
rect 150437 3417 150449 3420
rect 150483 3448 150495 3451
rect 151078 3448 151084 3460
rect 150483 3420 151084 3448
rect 150483 3417 150495 3420
rect 150437 3411 150495 3417
rect 151078 3408 151084 3420
rect 151136 3408 151142 3460
rect 151630 3448 151636 3460
rect 151591 3420 151636 3448
rect 151630 3408 151636 3420
rect 151688 3408 151694 3460
rect 151998 3380 152004 3392
rect 149808 3352 152004 3380
rect 151998 3340 152004 3352
rect 152056 3340 152062 3392
rect 152108 3389 152136 3488
rect 163222 3476 163228 3528
rect 163280 3516 163286 3528
rect 164145 3519 164203 3525
rect 164145 3516 164157 3519
rect 163280 3488 164157 3516
rect 163280 3476 163286 3488
rect 164145 3485 164157 3488
rect 164191 3516 164203 3519
rect 164605 3519 164663 3525
rect 164605 3516 164617 3519
rect 164191 3488 164617 3516
rect 164191 3485 164203 3488
rect 164145 3479 164203 3485
rect 164605 3485 164617 3488
rect 164651 3485 164663 3519
rect 164605 3479 164663 3485
rect 155034 3408 155040 3460
rect 155092 3448 155098 3460
rect 155129 3451 155187 3457
rect 155129 3448 155141 3451
rect 155092 3420 155141 3448
rect 155092 3408 155098 3420
rect 155129 3417 155141 3420
rect 155175 3448 155187 3451
rect 157242 3448 157248 3460
rect 155175 3420 157248 3448
rect 155175 3417 155187 3420
rect 155129 3411 155187 3417
rect 157242 3408 157248 3420
rect 157300 3408 157306 3460
rect 158533 3451 158591 3457
rect 158533 3417 158545 3451
rect 158579 3448 158591 3451
rect 158714 3448 158720 3460
rect 158579 3420 158720 3448
rect 158579 3417 158591 3420
rect 158533 3411 158591 3417
rect 158714 3408 158720 3420
rect 158772 3448 158778 3460
rect 159910 3448 159916 3460
rect 158772 3420 159916 3448
rect 158772 3408 158778 3420
rect 159910 3408 159916 3420
rect 159968 3408 159974 3460
rect 152093 3383 152151 3389
rect 152093 3349 152105 3383
rect 152139 3380 152151 3383
rect 153562 3380 153568 3392
rect 152139 3352 153568 3380
rect 152139 3349 152151 3352
rect 152093 3343 152151 3349
rect 153562 3340 153568 3352
rect 153620 3340 153626 3392
rect 156046 3340 156052 3392
rect 156104 3380 156110 3392
rect 156141 3383 156199 3389
rect 156141 3380 156153 3383
rect 156104 3352 156153 3380
rect 156104 3340 156110 3352
rect 156141 3349 156153 3352
rect 156187 3380 156199 3383
rect 156966 3380 156972 3392
rect 156187 3352 156972 3380
rect 156187 3349 156199 3352
rect 156141 3343 156199 3349
rect 156966 3340 156972 3352
rect 157024 3340 157030 3392
rect 159450 3340 159456 3392
rect 159508 3380 159514 3392
rect 159637 3383 159695 3389
rect 159637 3380 159649 3383
rect 159508 3352 159649 3380
rect 159508 3340 159514 3352
rect 159637 3349 159649 3352
rect 159683 3349 159695 3383
rect 159637 3343 159695 3349
rect 160281 3383 160339 3389
rect 160281 3349 160293 3383
rect 160327 3380 160339 3383
rect 160554 3380 160560 3392
rect 160327 3352 160560 3380
rect 160327 3349 160339 3352
rect 160281 3343 160339 3349
rect 160554 3340 160560 3352
rect 160612 3340 160618 3392
rect 161385 3383 161443 3389
rect 161385 3349 161397 3383
rect 161431 3380 161443 3383
rect 161750 3380 161756 3392
rect 161431 3352 161756 3380
rect 161431 3349 161443 3352
rect 161385 3343 161443 3349
rect 161750 3340 161756 3352
rect 161808 3340 161814 3392
rect 162305 3383 162363 3389
rect 162305 3349 162317 3383
rect 162351 3380 162363 3383
rect 162486 3380 162492 3392
rect 162351 3352 162492 3380
rect 162351 3349 162363 3352
rect 162305 3343 162363 3349
rect 162486 3340 162492 3352
rect 162544 3340 162550 3392
rect 164418 3340 164424 3392
rect 164476 3380 164482 3392
rect 164602 3380 164608 3392
rect 164476 3352 164608 3380
rect 164476 3340 164482 3352
rect 164602 3340 164608 3352
rect 164660 3340 164666 3392
rect 368 3290 93012 3312
rect 368 3238 56667 3290
rect 56719 3238 56731 3290
rect 56783 3238 56795 3290
rect 56847 3238 56859 3290
rect 56911 3238 93012 3290
rect 368 3216 93012 3238
rect 102028 3290 169556 3312
rect 102028 3238 113088 3290
rect 113140 3238 113152 3290
rect 113204 3238 113216 3290
rect 113268 3238 113280 3290
rect 113332 3238 169556 3290
rect 102028 3216 169556 3238
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 11606 3176 11612 3188
rect 3936 3148 11612 3176
rect 3936 3136 3942 3148
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 21634 3176 21640 3188
rect 11756 3148 21640 3176
rect 11756 3136 11762 3148
rect 21634 3136 21640 3148
rect 21692 3136 21698 3188
rect 21913 3179 21971 3185
rect 21913 3145 21925 3179
rect 21959 3176 21971 3179
rect 22462 3176 22468 3188
rect 21959 3148 22468 3176
rect 21959 3145 21971 3148
rect 21913 3139 21971 3145
rect 22462 3136 22468 3148
rect 22520 3136 22526 3188
rect 23216 3148 25084 3176
rect 6362 3068 6368 3120
rect 6420 3108 6426 3120
rect 6420 3080 9904 3108
rect 6420 3068 6426 3080
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 3694 3040 3700 3052
rect 3651 3012 3700 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3694 3000 3700 3012
rect 3752 3040 3758 3052
rect 4522 3040 4528 3052
rect 3752 3012 4528 3040
rect 3752 3000 3758 3012
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4706 3040 4712 3052
rect 4667 3012 4712 3040
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7834 3040 7840 3052
rect 7699 3012 7840 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 8478 3040 8484 3052
rect 8439 3012 8484 3040
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 9766 3040 9772 3052
rect 9727 3012 9772 3040
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 9876 3040 9904 3080
rect 10134 3068 10140 3120
rect 10192 3108 10198 3120
rect 17310 3108 17316 3120
rect 10192 3080 17316 3108
rect 10192 3068 10198 3080
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 17862 3068 17868 3120
rect 17920 3108 17926 3120
rect 19889 3111 19947 3117
rect 19889 3108 19901 3111
rect 17920 3080 19901 3108
rect 17920 3068 17926 3080
rect 19889 3077 19901 3080
rect 19935 3077 19947 3111
rect 23216 3108 23244 3148
rect 19889 3071 19947 3077
rect 19996 3080 23244 3108
rect 23293 3111 23351 3117
rect 10226 3040 10232 3052
rect 9876 3012 10232 3040
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3040 11759 3043
rect 11974 3040 11980 3052
rect 11747 3012 11980 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 13262 3040 13268 3052
rect 13223 3012 13268 3040
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 16022 3000 16028 3052
rect 16080 3040 16086 3052
rect 17954 3040 17960 3052
rect 16080 3012 17960 3040
rect 16080 3000 16086 3012
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 18414 3040 18420 3052
rect 18340 3012 18420 3040
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 6089 2975 6147 2981
rect 6089 2972 6101 2975
rect 2639 2944 6101 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 6089 2941 6101 2944
rect 6135 2941 6147 2975
rect 6089 2935 6147 2941
rect 750 2864 756 2916
rect 808 2904 814 2916
rect 4890 2904 4896 2916
rect 808 2876 4896 2904
rect 808 2864 814 2876
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 4982 2864 4988 2916
rect 5040 2904 5046 2916
rect 6104 2904 6132 2935
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 12713 2975 12771 2981
rect 12713 2972 12725 2975
rect 6236 2944 12725 2972
rect 6236 2932 6242 2944
rect 12713 2941 12725 2944
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 17126 2932 17132 2984
rect 17184 2972 17190 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17184 2944 18061 2972
rect 17184 2932 17190 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 6270 2904 6276 2916
rect 5040 2876 5672 2904
rect 6104 2876 6276 2904
rect 5040 2864 5046 2876
rect 5534 2836 5540 2848
rect 5495 2808 5540 2836
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 5644 2836 5672 2876
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 7374 2904 7380 2916
rect 7335 2876 7380 2904
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 7466 2864 7472 2916
rect 7524 2904 7530 2916
rect 7524 2876 9812 2904
rect 7524 2864 7530 2876
rect 9674 2836 9680 2848
rect 5644 2808 9680 2836
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9784 2836 9812 2876
rect 9858 2864 9864 2916
rect 9916 2904 9922 2916
rect 9953 2907 10011 2913
rect 9953 2904 9965 2907
rect 9916 2876 9965 2904
rect 9916 2864 9922 2876
rect 9953 2873 9965 2876
rect 9999 2873 10011 2907
rect 15378 2904 15384 2916
rect 9953 2867 10011 2873
rect 10060 2876 15384 2904
rect 10060 2836 10088 2876
rect 15378 2864 15384 2876
rect 15436 2864 15442 2916
rect 18340 2848 18368 3012
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 19996 3040 20024 3080
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24949 3111 25007 3117
rect 24949 3108 24961 3111
rect 23339 3080 24961 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24949 3077 24961 3080
rect 24995 3077 25007 3111
rect 25056 3108 25084 3148
rect 25314 3136 25320 3188
rect 25372 3176 25378 3188
rect 25372 3148 28672 3176
rect 25372 3136 25378 3148
rect 25056 3080 25912 3108
rect 24949 3071 25007 3077
rect 20530 3040 20536 3052
rect 18656 3012 20024 3040
rect 20443 3012 20536 3040
rect 18656 3000 18662 3012
rect 20530 3000 20536 3012
rect 20588 3040 20594 3052
rect 21542 3040 21548 3052
rect 20588 3012 21548 3040
rect 20588 3000 20594 3012
rect 21542 3000 21548 3012
rect 21600 3000 21606 3052
rect 21726 3000 21732 3052
rect 21784 3040 21790 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21784 3012 21833 3040
rect 21784 3000 21790 3012
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 24029 3043 24087 3049
rect 23164 3012 23612 3040
rect 23164 3000 23170 3012
rect 18966 2932 18972 2984
rect 19024 2972 19030 2984
rect 19024 2944 19840 2972
rect 19024 2932 19030 2944
rect 18690 2864 18696 2916
rect 18748 2904 18754 2916
rect 19702 2904 19708 2916
rect 18748 2876 19708 2904
rect 18748 2864 18754 2876
rect 19702 2864 19708 2876
rect 19760 2864 19766 2916
rect 19812 2904 19840 2944
rect 20346 2932 20352 2984
rect 20404 2972 20410 2984
rect 23293 2975 23351 2981
rect 23293 2972 23305 2975
rect 20404 2944 23305 2972
rect 20404 2932 20410 2944
rect 23293 2941 23305 2944
rect 23339 2941 23351 2975
rect 23293 2935 23351 2941
rect 23385 2975 23443 2981
rect 23385 2941 23397 2975
rect 23431 2941 23443 2975
rect 23385 2935 23443 2941
rect 23400 2904 23428 2935
rect 19812 2876 23428 2904
rect 9784 2808 10088 2836
rect 10226 2796 10232 2848
rect 10284 2836 10290 2848
rect 12434 2836 12440 2848
rect 10284 2808 12440 2836
rect 10284 2796 10290 2808
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 17954 2836 17960 2848
rect 14240 2808 17960 2836
rect 14240 2796 14246 2808
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18322 2796 18328 2848
rect 18380 2796 18386 2848
rect 18506 2796 18512 2848
rect 18564 2836 18570 2848
rect 19061 2839 19119 2845
rect 19061 2836 19073 2839
rect 18564 2808 19073 2836
rect 18564 2796 18570 2808
rect 19061 2805 19073 2808
rect 19107 2805 19119 2839
rect 19061 2799 19119 2805
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 23474 2836 23480 2848
rect 19392 2808 23480 2836
rect 19392 2796 19398 2808
rect 23474 2796 23480 2808
rect 23532 2796 23538 2848
rect 23584 2836 23612 3012
rect 24029 3009 24041 3043
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 23750 2932 23756 2984
rect 23808 2972 23814 2984
rect 24044 2972 24072 3003
rect 25406 3000 25412 3052
rect 25464 3040 25470 3052
rect 25593 3043 25651 3049
rect 25593 3040 25605 3043
rect 25464 3012 25605 3040
rect 25464 3000 25470 3012
rect 25593 3009 25605 3012
rect 25639 3040 25651 3043
rect 25639 3012 25820 3040
rect 25639 3009 25651 3012
rect 25593 3003 25651 3009
rect 25222 2972 25228 2984
rect 23808 2944 25228 2972
rect 23808 2932 23814 2944
rect 25222 2932 25228 2944
rect 25280 2932 25286 2984
rect 25792 2904 25820 3012
rect 25884 2972 25912 3080
rect 25958 3068 25964 3120
rect 26016 3108 26022 3120
rect 28537 3111 28595 3117
rect 28537 3108 28549 3111
rect 26016 3080 28549 3108
rect 26016 3068 26022 3080
rect 28537 3077 28549 3080
rect 28583 3077 28595 3111
rect 28644 3108 28672 3148
rect 28902 3136 28908 3188
rect 28960 3176 28966 3188
rect 29546 3176 29552 3188
rect 28960 3148 29552 3176
rect 28960 3136 28966 3148
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 30374 3136 30380 3188
rect 30432 3176 30438 3188
rect 33226 3176 33232 3188
rect 30432 3148 33232 3176
rect 30432 3136 30438 3148
rect 33226 3136 33232 3148
rect 33284 3136 33290 3188
rect 33318 3136 33324 3188
rect 33376 3176 33382 3188
rect 39482 3176 39488 3188
rect 33376 3148 39488 3176
rect 33376 3136 33382 3148
rect 39482 3136 39488 3148
rect 39540 3136 39546 3188
rect 39574 3136 39580 3188
rect 39632 3176 39638 3188
rect 41506 3176 41512 3188
rect 39632 3148 41512 3176
rect 39632 3136 39638 3148
rect 41506 3136 41512 3148
rect 41564 3136 41570 3188
rect 41598 3136 41604 3188
rect 41656 3176 41662 3188
rect 44082 3176 44088 3188
rect 41656 3148 44088 3176
rect 41656 3136 41662 3148
rect 44082 3136 44088 3148
rect 44140 3136 44146 3188
rect 44818 3176 44824 3188
rect 44779 3148 44824 3176
rect 44818 3136 44824 3148
rect 44876 3136 44882 3188
rect 44910 3136 44916 3188
rect 44968 3176 44974 3188
rect 46290 3176 46296 3188
rect 44968 3148 46296 3176
rect 44968 3136 44974 3148
rect 46290 3136 46296 3148
rect 46348 3136 46354 3188
rect 46474 3176 46480 3188
rect 46435 3148 46480 3176
rect 46474 3136 46480 3148
rect 46532 3136 46538 3188
rect 46658 3136 46664 3188
rect 46716 3176 46722 3188
rect 47118 3176 47124 3188
rect 46716 3148 47124 3176
rect 46716 3136 46722 3148
rect 47118 3136 47124 3148
rect 47176 3136 47182 3188
rect 47578 3176 47584 3188
rect 47539 3148 47584 3176
rect 47578 3136 47584 3148
rect 47636 3136 47642 3188
rect 49326 3176 49332 3188
rect 47688 3148 49332 3176
rect 28644 3080 30696 3108
rect 28537 3071 28595 3077
rect 27430 3040 27436 3052
rect 27391 3012 27436 3040
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 29181 3043 29239 3049
rect 29181 3009 29193 3043
rect 29227 3040 29239 3043
rect 29638 3040 29644 3052
rect 29227 3012 29644 3040
rect 29227 3009 29239 3012
rect 29181 3003 29239 3009
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 25884 2944 28028 2972
rect 26142 2904 26148 2916
rect 25792 2876 26148 2904
rect 26142 2864 26148 2876
rect 26200 2864 26206 2916
rect 27338 2864 27344 2916
rect 27396 2904 27402 2916
rect 27893 2907 27951 2913
rect 27893 2904 27905 2907
rect 27396 2876 27905 2904
rect 27396 2864 27402 2876
rect 27893 2873 27905 2876
rect 27939 2873 27951 2907
rect 28000 2904 28028 2944
rect 28166 2932 28172 2984
rect 28224 2972 28230 2984
rect 30561 2975 30619 2981
rect 30561 2972 30573 2975
rect 28224 2944 30573 2972
rect 28224 2932 28230 2944
rect 30561 2941 30573 2944
rect 30607 2941 30619 2975
rect 30561 2935 30619 2941
rect 30282 2904 30288 2916
rect 28000 2876 30288 2904
rect 27893 2867 27951 2873
rect 30282 2864 30288 2876
rect 30340 2864 30346 2916
rect 30668 2904 30696 3080
rect 30742 3068 30748 3120
rect 30800 3108 30806 3120
rect 36538 3108 36544 3120
rect 30800 3080 36544 3108
rect 30800 3068 30806 3080
rect 36538 3068 36544 3080
rect 36596 3068 36602 3120
rect 36648 3080 36952 3108
rect 30926 3040 30932 3052
rect 30887 3012 30932 3040
rect 30926 3000 30932 3012
rect 30984 3000 30990 3052
rect 31202 3000 31208 3052
rect 31260 3040 31266 3052
rect 31938 3040 31944 3052
rect 31260 3012 31944 3040
rect 31260 3000 31266 3012
rect 31938 3000 31944 3012
rect 31996 3000 32002 3052
rect 33686 3000 33692 3052
rect 33744 3040 33750 3052
rect 36648 3040 36676 3080
rect 33744 3012 36676 3040
rect 33744 3000 33750 3012
rect 36722 3000 36728 3052
rect 36780 3040 36786 3052
rect 36924 3040 36952 3080
rect 36998 3068 37004 3120
rect 37056 3108 37062 3120
rect 39022 3108 39028 3120
rect 37056 3080 39028 3108
rect 37056 3068 37062 3080
rect 39022 3068 39028 3080
rect 39080 3068 39086 3120
rect 39942 3108 39948 3120
rect 39316 3080 39948 3108
rect 37826 3040 37832 3052
rect 36780 3012 36825 3040
rect 36924 3012 37832 3040
rect 36780 3000 36786 3012
rect 37826 3000 37832 3012
rect 37884 3000 37890 3052
rect 39316 3040 39344 3080
rect 39942 3068 39948 3080
rect 40000 3068 40006 3120
rect 40034 3068 40040 3120
rect 40092 3108 40098 3120
rect 41046 3108 41052 3120
rect 40092 3080 41052 3108
rect 40092 3068 40098 3080
rect 41046 3068 41052 3080
rect 41104 3068 41110 3120
rect 43070 3108 43076 3120
rect 41156 3080 43076 3108
rect 37936 3012 39344 3040
rect 31662 2932 31668 2984
rect 31720 2972 31726 2984
rect 31846 2972 31852 2984
rect 31720 2944 31852 2972
rect 31720 2932 31726 2944
rect 31846 2932 31852 2944
rect 31904 2932 31910 2984
rect 32582 2932 32588 2984
rect 32640 2972 32646 2984
rect 36173 2975 36231 2981
rect 36173 2972 36185 2975
rect 32640 2944 36185 2972
rect 32640 2932 32646 2944
rect 36173 2941 36185 2944
rect 36219 2941 36231 2975
rect 36173 2935 36231 2941
rect 36354 2932 36360 2984
rect 36412 2972 36418 2984
rect 37936 2972 37964 3012
rect 39666 3000 39672 3052
rect 39724 3040 39730 3052
rect 39724 3012 39896 3040
rect 39724 3000 39730 3012
rect 36412 2944 37964 2972
rect 36412 2932 36418 2944
rect 38010 2932 38016 2984
rect 38068 2972 38074 2984
rect 38746 2972 38752 2984
rect 38068 2944 38752 2972
rect 38068 2932 38074 2944
rect 38746 2932 38752 2944
rect 38804 2932 38810 2984
rect 38930 2972 38936 2984
rect 38891 2944 38936 2972
rect 38930 2932 38936 2944
rect 38988 2932 38994 2984
rect 39022 2932 39028 2984
rect 39080 2972 39086 2984
rect 39574 2972 39580 2984
rect 39080 2944 39580 2972
rect 39080 2932 39086 2944
rect 39574 2932 39580 2944
rect 39632 2932 39638 2984
rect 39761 2975 39819 2981
rect 39761 2941 39773 2975
rect 39807 2941 39819 2975
rect 39761 2935 39819 2941
rect 39776 2904 39804 2935
rect 30668 2876 39804 2904
rect 39868 2904 39896 3012
rect 40126 3000 40132 3052
rect 40184 3040 40190 3052
rect 40310 3040 40316 3052
rect 40184 3012 40316 3040
rect 40184 3000 40190 3012
rect 40310 3000 40316 3012
rect 40368 3000 40374 3052
rect 40770 3000 40776 3052
rect 40828 3040 40834 3052
rect 41156 3040 41184 3080
rect 43070 3068 43076 3080
rect 43128 3068 43134 3120
rect 43438 3068 43444 3120
rect 43496 3108 43502 3120
rect 45373 3111 45431 3117
rect 45373 3108 45385 3111
rect 43496 3080 45385 3108
rect 43496 3068 43502 3080
rect 45373 3077 45385 3080
rect 45419 3077 45431 3111
rect 47688 3108 47716 3148
rect 49326 3136 49332 3148
rect 49384 3136 49390 3188
rect 49510 3136 49516 3188
rect 49568 3176 49574 3188
rect 49568 3148 54524 3176
rect 49568 3136 49574 3148
rect 45373 3071 45431 3077
rect 45480 3080 47716 3108
rect 40828 3012 41184 3040
rect 41325 3043 41383 3049
rect 40828 3000 40834 3012
rect 41325 3009 41337 3043
rect 41371 3040 41383 3043
rect 41690 3040 41696 3052
rect 41371 3012 41696 3040
rect 41371 3009 41383 3012
rect 41325 3003 41383 3009
rect 41690 3000 41696 3012
rect 41748 3040 41754 3052
rect 42334 3040 42340 3052
rect 41748 3012 42340 3040
rect 41748 3000 41754 3012
rect 42334 3000 42340 3012
rect 42392 3000 42398 3052
rect 43346 3040 43352 3052
rect 42444 3012 43352 3040
rect 39942 2932 39948 2984
rect 40000 2972 40006 2984
rect 42444 2972 42472 3012
rect 43346 3000 43352 3012
rect 43404 3000 43410 3052
rect 43530 3000 43536 3052
rect 43588 3040 43594 3052
rect 43717 3043 43775 3049
rect 43717 3040 43729 3043
rect 43588 3012 43729 3040
rect 43588 3000 43594 3012
rect 43717 3009 43729 3012
rect 43763 3009 43775 3043
rect 43717 3003 43775 3009
rect 43806 3000 43812 3052
rect 43864 3040 43870 3052
rect 44085 3043 44143 3049
rect 44085 3040 44097 3043
rect 43864 3012 44097 3040
rect 43864 3000 43870 3012
rect 44085 3009 44097 3012
rect 44131 3009 44143 3043
rect 44085 3003 44143 3009
rect 44453 3043 44511 3049
rect 44453 3009 44465 3043
rect 44499 3040 44511 3043
rect 44818 3040 44824 3052
rect 44499 3012 44824 3040
rect 44499 3009 44511 3012
rect 44453 3003 44511 3009
rect 44818 3000 44824 3012
rect 44876 3000 44882 3052
rect 44910 3000 44916 3052
rect 44968 3040 44974 3052
rect 45480 3040 45508 3080
rect 48038 3068 48044 3120
rect 48096 3108 48102 3120
rect 53098 3108 53104 3120
rect 48096 3080 53104 3108
rect 48096 3068 48102 3080
rect 53098 3068 53104 3080
rect 53156 3068 53162 3120
rect 53190 3068 53196 3120
rect 53248 3108 53254 3120
rect 53561 3111 53619 3117
rect 53561 3108 53573 3111
rect 53248 3080 53573 3108
rect 53248 3068 53254 3080
rect 53561 3077 53573 3080
rect 53607 3077 53619 3111
rect 54496 3108 54524 3148
rect 55214 3136 55220 3188
rect 55272 3176 55278 3188
rect 55272 3148 55812 3176
rect 55272 3136 55278 3148
rect 55674 3108 55680 3120
rect 54496 3080 55680 3108
rect 53561 3071 53619 3077
rect 55674 3068 55680 3080
rect 55732 3068 55738 3120
rect 55784 3108 55812 3148
rect 56134 3136 56140 3188
rect 56192 3176 56198 3188
rect 56689 3179 56747 3185
rect 56689 3176 56701 3179
rect 56192 3148 56701 3176
rect 56192 3136 56198 3148
rect 56689 3145 56701 3148
rect 56735 3145 56747 3179
rect 56689 3139 56747 3145
rect 56962 3136 56968 3188
rect 57020 3176 57026 3188
rect 57333 3179 57391 3185
rect 57333 3176 57345 3179
rect 57020 3148 57345 3176
rect 57020 3136 57026 3148
rect 57333 3145 57345 3148
rect 57379 3145 57391 3179
rect 60458 3176 60464 3188
rect 57333 3139 57391 3145
rect 57440 3148 60464 3176
rect 57440 3108 57468 3148
rect 60458 3136 60464 3148
rect 60516 3136 60522 3188
rect 60550 3136 60556 3188
rect 60608 3176 60614 3188
rect 61102 3176 61108 3188
rect 60608 3148 61108 3176
rect 60608 3136 60614 3148
rect 61102 3136 61108 3148
rect 61160 3176 61166 3188
rect 61381 3179 61439 3185
rect 61381 3176 61393 3179
rect 61160 3148 61393 3176
rect 61160 3136 61166 3148
rect 61381 3145 61393 3148
rect 61427 3145 61439 3179
rect 62298 3176 62304 3188
rect 62259 3148 62304 3176
rect 61381 3139 61439 3145
rect 62298 3136 62304 3148
rect 62356 3136 62362 3188
rect 62666 3136 62672 3188
rect 62724 3176 62730 3188
rect 63405 3179 63463 3185
rect 63405 3176 63417 3179
rect 62724 3148 63417 3176
rect 62724 3136 62730 3148
rect 63405 3145 63417 3148
rect 63451 3145 63463 3179
rect 64414 3176 64420 3188
rect 64375 3148 64420 3176
rect 63405 3139 63463 3145
rect 64414 3136 64420 3148
rect 64472 3136 64478 3188
rect 64506 3136 64512 3188
rect 64564 3176 64570 3188
rect 70118 3176 70124 3188
rect 64564 3148 70124 3176
rect 64564 3136 64570 3148
rect 70118 3136 70124 3148
rect 70176 3136 70182 3188
rect 70394 3136 70400 3188
rect 70452 3176 70458 3188
rect 71774 3176 71780 3188
rect 70452 3148 71780 3176
rect 70452 3136 70458 3148
rect 71774 3136 71780 3148
rect 71832 3136 71838 3188
rect 73522 3176 73528 3188
rect 73483 3148 73528 3176
rect 73522 3136 73528 3148
rect 73580 3136 73586 3188
rect 88426 3176 88432 3188
rect 88387 3148 88432 3176
rect 88426 3136 88432 3148
rect 88484 3136 88490 3188
rect 88794 3136 88800 3188
rect 88852 3176 88858 3188
rect 93302 3176 93308 3188
rect 88852 3148 93308 3176
rect 88852 3136 88858 3148
rect 93302 3136 93308 3148
rect 93360 3136 93366 3188
rect 104434 3136 104440 3188
rect 104492 3176 104498 3188
rect 108942 3176 108948 3188
rect 104492 3148 108948 3176
rect 104492 3136 104498 3148
rect 108942 3136 108948 3148
rect 109000 3136 109006 3188
rect 109034 3136 109040 3188
rect 109092 3176 109098 3188
rect 133230 3176 133236 3188
rect 109092 3148 132356 3176
rect 133191 3148 133236 3176
rect 109092 3136 109098 3148
rect 55784 3080 57468 3108
rect 57974 3068 57980 3120
rect 58032 3108 58038 3120
rect 58713 3111 58771 3117
rect 58713 3108 58725 3111
rect 58032 3080 58725 3108
rect 58032 3068 58038 3080
rect 58713 3077 58725 3080
rect 58759 3077 58771 3111
rect 58713 3071 58771 3077
rect 58986 3068 58992 3120
rect 59044 3108 59050 3120
rect 65702 3108 65708 3120
rect 59044 3080 65708 3108
rect 59044 3068 59050 3080
rect 65702 3068 65708 3080
rect 65760 3068 65766 3120
rect 65978 3068 65984 3120
rect 66036 3108 66042 3120
rect 66036 3080 71820 3108
rect 66036 3068 66042 3080
rect 44968 3012 45508 3040
rect 44968 3000 44974 3012
rect 45554 3000 45560 3052
rect 45612 3040 45618 3052
rect 45612 3012 45657 3040
rect 45612 3000 45618 3012
rect 45738 3000 45744 3052
rect 45796 3040 45802 3052
rect 45796 3012 46704 3040
rect 45796 3000 45802 3012
rect 42702 2972 42708 2984
rect 40000 2944 42472 2972
rect 42663 2944 42708 2972
rect 40000 2932 40006 2944
rect 42702 2932 42708 2944
rect 42760 2932 42766 2984
rect 46566 2972 46572 2984
rect 42812 2944 46572 2972
rect 39868 2876 41552 2904
rect 25682 2836 25688 2848
rect 23584 2808 25688 2836
rect 25682 2796 25688 2808
rect 25740 2796 25746 2848
rect 25774 2796 25780 2848
rect 25832 2836 25838 2848
rect 25961 2839 26019 2845
rect 25961 2836 25973 2839
rect 25832 2808 25973 2836
rect 25832 2796 25838 2808
rect 25961 2805 25973 2808
rect 26007 2805 26019 2839
rect 25961 2799 26019 2805
rect 26510 2796 26516 2848
rect 26568 2836 26574 2848
rect 27525 2839 27583 2845
rect 27525 2836 27537 2839
rect 26568 2808 27537 2836
rect 26568 2796 26574 2808
rect 27525 2805 27537 2808
rect 27571 2805 27583 2839
rect 27525 2799 27583 2805
rect 27614 2796 27620 2848
rect 27672 2836 27678 2848
rect 34698 2836 34704 2848
rect 27672 2808 34704 2836
rect 27672 2796 27678 2808
rect 34698 2796 34704 2808
rect 34756 2796 34762 2848
rect 34790 2796 34796 2848
rect 34848 2836 34854 2848
rect 35618 2836 35624 2848
rect 34848 2808 35624 2836
rect 34848 2796 34854 2808
rect 35618 2796 35624 2808
rect 35676 2796 35682 2848
rect 36354 2796 36360 2848
rect 36412 2836 36418 2848
rect 36722 2836 36728 2848
rect 36412 2808 36728 2836
rect 36412 2796 36418 2808
rect 36722 2796 36728 2808
rect 36780 2836 36786 2848
rect 38194 2836 38200 2848
rect 36780 2808 38200 2836
rect 36780 2796 36786 2808
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 38286 2796 38292 2848
rect 38344 2836 38350 2848
rect 39850 2836 39856 2848
rect 38344 2808 39856 2836
rect 38344 2796 38350 2808
rect 39850 2796 39856 2808
rect 39908 2796 39914 2848
rect 40494 2796 40500 2848
rect 40552 2836 40558 2848
rect 41417 2839 41475 2845
rect 41417 2836 41429 2839
rect 40552 2808 41429 2836
rect 40552 2796 40558 2808
rect 41417 2805 41429 2808
rect 41463 2805 41475 2839
rect 41524 2836 41552 2876
rect 41690 2864 41696 2916
rect 41748 2904 41754 2916
rect 41874 2904 41880 2916
rect 41748 2876 41880 2904
rect 41748 2864 41754 2876
rect 41874 2864 41880 2876
rect 41932 2864 41938 2916
rect 41966 2864 41972 2916
rect 42024 2904 42030 2916
rect 42812 2904 42840 2944
rect 46566 2932 46572 2944
rect 46624 2932 46630 2984
rect 46676 2972 46704 3012
rect 47210 3000 47216 3052
rect 47268 3040 47274 3052
rect 47489 3043 47547 3049
rect 47489 3040 47501 3043
rect 47268 3012 47501 3040
rect 47268 3000 47274 3012
rect 47489 3009 47501 3012
rect 47535 3009 47547 3043
rect 47489 3003 47547 3009
rect 47578 3000 47584 3052
rect 47636 3040 47642 3052
rect 48222 3040 48228 3052
rect 47636 3012 48228 3040
rect 47636 3000 47642 3012
rect 48222 3000 48228 3012
rect 48280 3000 48286 3052
rect 48774 3040 48780 3052
rect 48735 3012 48780 3040
rect 48774 3000 48780 3012
rect 48832 3040 48838 3052
rect 49050 3040 49056 3052
rect 48832 3012 49056 3040
rect 48832 3000 48838 3012
rect 49050 3000 49056 3012
rect 49108 3000 49114 3052
rect 49142 3000 49148 3052
rect 49200 3040 49206 3052
rect 50706 3040 50712 3052
rect 49200 3012 50712 3040
rect 49200 3000 49206 3012
rect 50706 3000 50712 3012
rect 50764 3000 50770 3052
rect 50798 3000 50804 3052
rect 50856 3040 50862 3052
rect 53466 3040 53472 3052
rect 50856 3012 53472 3040
rect 50856 3000 50862 3012
rect 53466 3000 53472 3012
rect 53524 3000 53530 3052
rect 53650 3000 53656 3052
rect 53708 3040 53714 3052
rect 54205 3043 54263 3049
rect 54205 3040 54217 3043
rect 53708 3012 54217 3040
rect 53708 3000 53714 3012
rect 54205 3009 54217 3012
rect 54251 3040 54263 3043
rect 54938 3040 54944 3052
rect 54251 3012 54944 3040
rect 54251 3009 54263 3012
rect 54205 3003 54263 3009
rect 54938 3000 54944 3012
rect 54996 3000 55002 3052
rect 55122 3040 55128 3052
rect 55083 3012 55128 3040
rect 55122 3000 55128 3012
rect 55180 3000 55186 3052
rect 55858 3000 55864 3052
rect 55916 3040 55922 3052
rect 56318 3040 56324 3052
rect 55916 3012 56324 3040
rect 55916 3000 55922 3012
rect 56318 3000 56324 3012
rect 56376 3000 56382 3052
rect 56597 3043 56655 3049
rect 56597 3009 56609 3043
rect 56643 3040 56655 3043
rect 57054 3040 57060 3052
rect 56643 3012 57060 3040
rect 56643 3009 56655 3012
rect 56597 3003 56655 3009
rect 57054 3000 57060 3012
rect 57112 3000 57118 3052
rect 57238 3000 57244 3052
rect 57296 3040 57302 3052
rect 58621 3043 58679 3049
rect 57296 3012 58572 3040
rect 57296 3000 57302 3012
rect 46676 2944 49280 2972
rect 45646 2904 45652 2916
rect 42024 2876 42840 2904
rect 42904 2876 45652 2904
rect 42024 2864 42030 2876
rect 42904 2836 42932 2876
rect 45646 2864 45652 2876
rect 45704 2864 45710 2916
rect 45830 2864 45836 2916
rect 45888 2904 45894 2916
rect 49142 2904 49148 2916
rect 45888 2876 49148 2904
rect 45888 2864 45894 2876
rect 49142 2864 49148 2876
rect 49200 2864 49206 2916
rect 49252 2904 49280 2944
rect 49326 2932 49332 2984
rect 49384 2972 49390 2984
rect 49384 2944 51212 2972
rect 49384 2932 49390 2944
rect 51074 2904 51080 2916
rect 49252 2876 51080 2904
rect 51074 2864 51080 2876
rect 51132 2864 51138 2916
rect 51184 2904 51212 2944
rect 51258 2932 51264 2984
rect 51316 2972 51322 2984
rect 51316 2944 55444 2972
rect 51316 2932 51322 2944
rect 51718 2904 51724 2916
rect 51184 2876 51724 2904
rect 51718 2864 51724 2876
rect 51776 2864 51782 2916
rect 52178 2864 52184 2916
rect 52236 2904 52242 2916
rect 55306 2904 55312 2916
rect 52236 2876 55312 2904
rect 52236 2864 52242 2876
rect 55306 2864 55312 2876
rect 55364 2864 55370 2916
rect 55416 2904 55444 2944
rect 55490 2932 55496 2984
rect 55548 2972 55554 2984
rect 57422 2972 57428 2984
rect 55548 2944 57428 2972
rect 55548 2932 55554 2944
rect 57422 2932 57428 2944
rect 57480 2932 57486 2984
rect 57609 2975 57667 2981
rect 57609 2941 57621 2975
rect 57655 2972 57667 2975
rect 58434 2972 58440 2984
rect 57655 2944 58440 2972
rect 57655 2941 57667 2944
rect 57609 2935 57667 2941
rect 58434 2932 58440 2944
rect 58492 2932 58498 2984
rect 58544 2972 58572 3012
rect 58621 3009 58633 3043
rect 58667 3040 58679 3043
rect 58802 3040 58808 3052
rect 58667 3012 58808 3040
rect 58667 3009 58679 3012
rect 58621 3003 58679 3009
rect 58802 3000 58808 3012
rect 58860 3000 58866 3052
rect 58894 3000 58900 3052
rect 58952 3040 58958 3052
rect 60277 3043 60335 3049
rect 58952 3012 60228 3040
rect 58952 3000 58958 3012
rect 59630 2972 59636 2984
rect 58544 2944 59636 2972
rect 59630 2932 59636 2944
rect 59688 2932 59694 2984
rect 60200 2972 60228 3012
rect 60277 3009 60289 3043
rect 60323 3040 60335 3043
rect 60369 3043 60427 3049
rect 60369 3040 60381 3043
rect 60323 3012 60381 3040
rect 60323 3009 60335 3012
rect 60277 3003 60335 3009
rect 60369 3009 60381 3012
rect 60415 3040 60427 3043
rect 60458 3040 60464 3052
rect 60415 3012 60464 3040
rect 60415 3009 60427 3012
rect 60369 3003 60427 3009
rect 60458 3000 60464 3012
rect 60516 3000 60522 3052
rect 60550 3000 60556 3052
rect 60608 3040 60614 3052
rect 60737 3043 60795 3049
rect 60737 3040 60749 3043
rect 60608 3012 60749 3040
rect 60608 3000 60614 3012
rect 60737 3009 60749 3012
rect 60783 3009 60795 3043
rect 60737 3003 60795 3009
rect 61105 3043 61163 3049
rect 61105 3009 61117 3043
rect 61151 3040 61163 3043
rect 62209 3043 62267 3049
rect 61151 3012 61240 3040
rect 61151 3009 61163 3012
rect 61105 3003 61163 3009
rect 60642 2972 60648 2984
rect 60200 2944 60648 2972
rect 60642 2932 60648 2944
rect 60700 2932 60706 2984
rect 60918 2932 60924 2984
rect 60976 2972 60982 2984
rect 61212 2972 61240 3012
rect 62209 3009 62221 3043
rect 62255 3040 62267 3043
rect 62390 3040 62396 3052
rect 62255 3012 62396 3040
rect 62255 3009 62267 3012
rect 62209 3003 62267 3009
rect 62390 3000 62396 3012
rect 62448 3000 62454 3052
rect 63313 3043 63371 3049
rect 63313 3009 63325 3043
rect 63359 3040 63371 3043
rect 63494 3040 63500 3052
rect 63359 3012 63500 3040
rect 63359 3009 63371 3012
rect 63313 3003 63371 3009
rect 63494 3000 63500 3012
rect 63552 3000 63558 3052
rect 63770 3000 63776 3052
rect 63828 3040 63834 3052
rect 64325 3043 64383 3049
rect 63828 3012 64092 3040
rect 63828 3000 63834 3012
rect 60976 2944 61240 2972
rect 61289 2975 61347 2981
rect 60976 2932 60982 2944
rect 61289 2941 61301 2975
rect 61335 2972 61347 2975
rect 63954 2972 63960 2984
rect 61335 2944 63960 2972
rect 61335 2941 61347 2944
rect 61289 2935 61347 2941
rect 63954 2932 63960 2944
rect 64012 2932 64018 2984
rect 64064 2972 64092 3012
rect 64325 3009 64337 3043
rect 64371 3040 64383 3043
rect 64506 3040 64512 3052
rect 64371 3012 64512 3040
rect 64371 3009 64383 3012
rect 64325 3003 64383 3009
rect 64506 3000 64512 3012
rect 64564 3000 64570 3052
rect 68370 3040 68376 3052
rect 64616 3012 68376 3040
rect 64616 2972 64644 3012
rect 68370 3000 68376 3012
rect 68428 3000 68434 3052
rect 68465 3043 68523 3049
rect 68465 3009 68477 3043
rect 68511 3009 68523 3043
rect 68465 3003 68523 3009
rect 69477 3043 69535 3049
rect 69477 3009 69489 3043
rect 69523 3040 69535 3043
rect 70210 3040 70216 3052
rect 69523 3012 70216 3040
rect 69523 3009 69535 3012
rect 69477 3003 69535 3009
rect 65334 2972 65340 2984
rect 64064 2944 64644 2972
rect 65295 2944 65340 2972
rect 65334 2932 65340 2944
rect 65392 2932 65398 2984
rect 66714 2972 66720 2984
rect 66675 2944 66720 2972
rect 66714 2932 66720 2944
rect 66772 2932 66778 2984
rect 68480 2972 68508 3003
rect 70210 3000 70216 3012
rect 70268 3000 70274 3052
rect 70489 3043 70547 3049
rect 70489 3009 70501 3043
rect 70535 3040 70547 3043
rect 70578 3040 70584 3052
rect 70535 3012 70584 3040
rect 70535 3009 70547 3012
rect 70489 3003 70547 3009
rect 70578 3000 70584 3012
rect 70636 3000 70642 3052
rect 71130 3000 71136 3052
rect 71188 3040 71194 3052
rect 71501 3043 71559 3049
rect 71501 3040 71513 3043
rect 71188 3012 71513 3040
rect 71188 3000 71194 3012
rect 71501 3009 71513 3012
rect 71547 3009 71559 3043
rect 71501 3003 71559 3009
rect 71593 3043 71651 3049
rect 71593 3009 71605 3043
rect 71639 3040 71651 3043
rect 71682 3040 71688 3052
rect 71639 3012 71688 3040
rect 71639 3009 71651 3012
rect 71593 3003 71651 3009
rect 71682 3000 71688 3012
rect 71740 3000 71746 3052
rect 71792 3040 71820 3080
rect 72050 3068 72056 3120
rect 72108 3108 72114 3120
rect 86678 3108 86684 3120
rect 72108 3080 86684 3108
rect 72108 3068 72114 3080
rect 86678 3068 86684 3080
rect 86736 3068 86742 3120
rect 101582 3068 101588 3120
rect 101640 3108 101646 3120
rect 101640 3080 103468 3108
rect 101640 3068 101646 3080
rect 73249 3043 73307 3049
rect 73249 3040 73261 3043
rect 71792 3012 73261 3040
rect 73249 3009 73261 3012
rect 73295 3009 73307 3043
rect 73249 3003 73307 3009
rect 73433 3043 73491 3049
rect 73433 3009 73445 3043
rect 73479 3040 73491 3043
rect 74258 3040 74264 3052
rect 73479 3012 74264 3040
rect 73479 3009 73491 3012
rect 73433 3003 73491 3009
rect 74258 3000 74264 3012
rect 74316 3000 74322 3052
rect 87322 3040 87328 3052
rect 87283 3012 87328 3040
rect 87322 3000 87328 3012
rect 87380 3000 87386 3052
rect 88337 3043 88395 3049
rect 88337 3009 88349 3043
rect 88383 3040 88395 3043
rect 88426 3040 88432 3052
rect 88383 3012 88432 3040
rect 88383 3009 88395 3012
rect 88337 3003 88395 3009
rect 88426 3000 88432 3012
rect 88484 3000 88490 3052
rect 90266 3000 90272 3052
rect 90324 3040 90330 3052
rect 90361 3043 90419 3049
rect 90361 3040 90373 3043
rect 90324 3012 90373 3040
rect 90324 3000 90330 3012
rect 90361 3009 90373 3012
rect 90407 3040 90419 3043
rect 90726 3040 90732 3052
rect 90407 3012 90732 3040
rect 90407 3009 90419 3012
rect 90361 3003 90419 3009
rect 90726 3000 90732 3012
rect 90784 3000 90790 3052
rect 91830 3040 91836 3052
rect 91791 3012 91836 3040
rect 91830 3000 91836 3012
rect 91888 3040 91894 3052
rect 92201 3043 92259 3049
rect 92201 3040 92213 3043
rect 91888 3012 92213 3040
rect 91888 3000 91894 3012
rect 92201 3009 92213 3012
rect 92247 3009 92259 3043
rect 92201 3003 92259 3009
rect 102134 3000 102140 3052
rect 102192 3040 102198 3052
rect 102321 3043 102379 3049
rect 102321 3040 102333 3043
rect 102192 3012 102333 3040
rect 102192 3000 102198 3012
rect 102321 3009 102333 3012
rect 102367 3040 102379 3043
rect 102781 3043 102839 3049
rect 102781 3040 102793 3043
rect 102367 3012 102793 3040
rect 102367 3009 102379 3012
rect 102321 3003 102379 3009
rect 102781 3009 102793 3012
rect 102827 3009 102839 3043
rect 103325 3043 103383 3049
rect 103325 3040 103337 3043
rect 102781 3003 102839 3009
rect 103256 3012 103337 3040
rect 68554 2972 68560 2984
rect 68467 2944 68560 2972
rect 68554 2932 68560 2944
rect 68612 2972 68618 2984
rect 71314 2972 71320 2984
rect 68612 2944 71320 2972
rect 68612 2932 68618 2944
rect 71314 2932 71320 2944
rect 71372 2932 71378 2984
rect 73614 2932 73620 2984
rect 73672 2972 73678 2984
rect 74445 2975 74503 2981
rect 74445 2972 74457 2975
rect 73672 2944 74457 2972
rect 73672 2932 73678 2944
rect 74445 2941 74457 2944
rect 74491 2941 74503 2975
rect 74445 2935 74503 2941
rect 76098 2932 76104 2984
rect 76156 2972 76162 2984
rect 76193 2975 76251 2981
rect 76193 2972 76205 2975
rect 76156 2944 76205 2972
rect 76156 2932 76162 2944
rect 76193 2941 76205 2944
rect 76239 2941 76251 2975
rect 76193 2935 76251 2941
rect 76558 2932 76564 2984
rect 76616 2972 76622 2984
rect 76745 2975 76803 2981
rect 76745 2972 76757 2975
rect 76616 2944 76757 2972
rect 76616 2932 76622 2944
rect 76745 2941 76757 2944
rect 76791 2972 76803 2975
rect 77205 2975 77263 2981
rect 77205 2972 77217 2975
rect 76791 2944 77217 2972
rect 76791 2941 76803 2944
rect 76745 2935 76803 2941
rect 77205 2941 77217 2944
rect 77251 2941 77263 2975
rect 77205 2935 77263 2941
rect 80885 2975 80943 2981
rect 80885 2941 80897 2975
rect 80931 2972 80943 2975
rect 80974 2972 80980 2984
rect 80931 2944 80980 2972
rect 80931 2941 80943 2944
rect 80885 2935 80943 2941
rect 80974 2932 80980 2944
rect 81032 2932 81038 2984
rect 83090 2972 83096 2984
rect 83051 2944 83096 2972
rect 83090 2932 83096 2944
rect 83148 2932 83154 2984
rect 86310 2972 86316 2984
rect 86271 2944 86316 2972
rect 86310 2932 86316 2944
rect 86368 2932 86374 2984
rect 88150 2932 88156 2984
rect 88208 2972 88214 2984
rect 91373 2975 91431 2981
rect 91373 2972 91385 2975
rect 88208 2944 91385 2972
rect 88208 2932 88214 2944
rect 91373 2941 91385 2944
rect 91419 2941 91431 2975
rect 91373 2935 91431 2941
rect 103054 2932 103060 2984
rect 103112 2972 103118 2984
rect 103256 2972 103284 3012
rect 103325 3009 103337 3012
rect 103371 3009 103383 3043
rect 103440 3040 103468 3080
rect 103514 3068 103520 3120
rect 103572 3108 103578 3120
rect 107565 3111 107623 3117
rect 107565 3108 107577 3111
rect 103572 3080 107577 3108
rect 103572 3068 103578 3080
rect 107565 3077 107577 3080
rect 107611 3077 107623 3111
rect 107838 3108 107844 3120
rect 107799 3080 107844 3108
rect 107565 3071 107623 3077
rect 107838 3068 107844 3080
rect 107896 3068 107902 3120
rect 108114 3068 108120 3120
rect 108172 3108 108178 3120
rect 108172 3080 108804 3108
rect 108172 3068 108178 3080
rect 107470 3040 107476 3052
rect 103440 3012 107476 3040
rect 103325 3003 103383 3009
rect 107470 3000 107476 3012
rect 107528 3000 107534 3052
rect 107746 3040 107752 3052
rect 107707 3012 107752 3040
rect 107746 3000 107752 3012
rect 107804 3000 107810 3052
rect 108776 3040 108804 3080
rect 108850 3068 108856 3120
rect 108908 3108 108914 3120
rect 130013 3111 130071 3117
rect 130013 3108 130025 3111
rect 108908 3080 130025 3108
rect 108908 3068 108914 3080
rect 130013 3077 130025 3080
rect 130059 3077 130071 3111
rect 130013 3071 130071 3077
rect 109402 3040 109408 3052
rect 108776 3012 109408 3040
rect 109402 3000 109408 3012
rect 109460 3000 109466 3052
rect 109586 3040 109592 3052
rect 109547 3012 109592 3040
rect 109586 3000 109592 3012
rect 109644 3000 109650 3052
rect 109681 3043 109739 3049
rect 109681 3009 109693 3043
rect 109727 3040 109739 3043
rect 109770 3040 109776 3052
rect 109727 3012 109776 3040
rect 109727 3009 109739 3012
rect 109681 3003 109739 3009
rect 109770 3000 109776 3012
rect 109828 3000 109834 3052
rect 110877 3043 110935 3049
rect 110877 3009 110889 3043
rect 110923 3040 110935 3043
rect 111518 3040 111524 3052
rect 110923 3012 111524 3040
rect 110923 3009 110935 3012
rect 110877 3003 110935 3009
rect 111518 3000 111524 3012
rect 111576 3040 111582 3052
rect 112806 3040 112812 3052
rect 111576 3012 112812 3040
rect 111576 3000 111582 3012
rect 112806 3000 112812 3012
rect 112864 3000 112870 3052
rect 113637 3043 113695 3049
rect 113637 3009 113649 3043
rect 113683 3040 113695 3043
rect 114554 3040 114560 3052
rect 113683 3012 114560 3040
rect 113683 3009 113695 3012
rect 113637 3003 113695 3009
rect 114554 3000 114560 3012
rect 114612 3000 114618 3052
rect 117133 3043 117191 3049
rect 117133 3009 117145 3043
rect 117179 3040 117191 3043
rect 117222 3040 117228 3052
rect 117179 3012 117228 3040
rect 117179 3009 117191 3012
rect 117133 3003 117191 3009
rect 117222 3000 117228 3012
rect 117280 3040 117286 3052
rect 119430 3040 119436 3052
rect 117280 3012 119436 3040
rect 117280 3000 117286 3012
rect 119430 3000 119436 3012
rect 119488 3000 119494 3052
rect 122377 3043 122435 3049
rect 122377 3009 122389 3043
rect 122423 3009 122435 3043
rect 122377 3003 122435 3009
rect 104158 2972 104164 2984
rect 103112 2944 104164 2972
rect 103112 2932 103118 2944
rect 104158 2932 104164 2944
rect 104216 2932 104222 2984
rect 104342 2972 104348 2984
rect 104303 2944 104348 2972
rect 104342 2932 104348 2944
rect 104400 2932 104406 2984
rect 105446 2932 105452 2984
rect 105504 2972 105510 2984
rect 108574 2972 108580 2984
rect 105504 2944 108580 2972
rect 105504 2932 105510 2944
rect 108574 2932 108580 2944
rect 108632 2932 108638 2984
rect 109126 2932 109132 2984
rect 109184 2972 109190 2984
rect 120074 2972 120080 2984
rect 109184 2944 120080 2972
rect 109184 2932 109190 2944
rect 120074 2932 120080 2944
rect 120132 2932 120138 2984
rect 122392 2916 122420 3003
rect 122466 3000 122472 3052
rect 122524 3040 122530 3052
rect 126333 3043 126391 3049
rect 122524 3012 122569 3040
rect 122524 3000 122530 3012
rect 126333 3009 126345 3043
rect 126379 3040 126391 3043
rect 126882 3040 126888 3052
rect 126379 3012 126888 3040
rect 126379 3009 126391 3012
rect 126333 3003 126391 3009
rect 126882 3000 126888 3012
rect 126940 3000 126946 3052
rect 127897 3043 127955 3049
rect 127897 3009 127909 3043
rect 127943 3040 127955 3043
rect 128170 3040 128176 3052
rect 127943 3012 128176 3040
rect 127943 3009 127955 3012
rect 127897 3003 127955 3009
rect 128170 3000 128176 3012
rect 128228 3000 128234 3052
rect 125778 2932 125784 2984
rect 125836 2972 125842 2984
rect 126425 2975 126483 2981
rect 126425 2972 126437 2975
rect 125836 2944 126437 2972
rect 125836 2932 125842 2944
rect 126425 2941 126437 2944
rect 126471 2941 126483 2975
rect 127986 2972 127992 2984
rect 127947 2944 127992 2972
rect 126425 2935 126483 2941
rect 127986 2932 127992 2944
rect 128044 2932 128050 2984
rect 132328 2972 132356 3148
rect 133230 3136 133236 3148
rect 133288 3136 133294 3188
rect 134242 3176 134248 3188
rect 134203 3148 134248 3176
rect 134242 3136 134248 3148
rect 134300 3136 134306 3188
rect 138566 3136 138572 3188
rect 138624 3176 138630 3188
rect 144914 3176 144920 3188
rect 138624 3148 144920 3176
rect 138624 3136 138630 3148
rect 144914 3136 144920 3148
rect 144972 3136 144978 3188
rect 145374 3176 145380 3188
rect 145335 3148 145380 3176
rect 145374 3136 145380 3148
rect 145432 3136 145438 3188
rect 149054 3136 149060 3188
rect 149112 3176 149118 3188
rect 150342 3176 150348 3188
rect 149112 3148 150348 3176
rect 149112 3136 149118 3148
rect 150342 3136 150348 3148
rect 150400 3136 150406 3188
rect 154298 3176 154304 3188
rect 154259 3148 154304 3176
rect 154298 3136 154304 3148
rect 154356 3136 154362 3188
rect 154942 3136 154948 3188
rect 155000 3176 155006 3188
rect 155313 3179 155371 3185
rect 155313 3176 155325 3179
rect 155000 3148 155325 3176
rect 155000 3136 155006 3148
rect 155313 3145 155325 3148
rect 155359 3145 155371 3179
rect 155313 3139 155371 3145
rect 156325 3179 156383 3185
rect 156325 3145 156337 3179
rect 156371 3176 156383 3179
rect 156598 3176 156604 3188
rect 156371 3148 156604 3176
rect 156371 3145 156383 3148
rect 156325 3139 156383 3145
rect 156598 3136 156604 3148
rect 156656 3136 156662 3188
rect 159545 3179 159603 3185
rect 159545 3145 159557 3179
rect 159591 3176 159603 3179
rect 159726 3176 159732 3188
rect 159591 3148 159732 3176
rect 159591 3145 159603 3148
rect 159545 3139 159603 3145
rect 159726 3136 159732 3148
rect 159784 3136 159790 3188
rect 160738 3176 160744 3188
rect 160699 3148 160744 3176
rect 160738 3136 160744 3148
rect 160796 3136 160802 3188
rect 164053 3179 164111 3185
rect 164053 3145 164065 3179
rect 164099 3176 164111 3179
rect 164326 3176 164332 3188
rect 164099 3148 164332 3176
rect 164099 3145 164111 3148
rect 164053 3139 164111 3145
rect 164326 3136 164332 3148
rect 164384 3136 164390 3188
rect 165062 3176 165068 3188
rect 165023 3148 165068 3176
rect 165062 3136 165068 3148
rect 165120 3136 165126 3188
rect 144454 3068 144460 3120
rect 144512 3108 144518 3120
rect 161106 3108 161112 3120
rect 144512 3080 161112 3108
rect 144512 3068 144518 3080
rect 161106 3068 161112 3080
rect 161164 3068 161170 3120
rect 133046 3000 133052 3052
rect 133104 3040 133110 3052
rect 133141 3043 133199 3049
rect 133141 3040 133153 3043
rect 133104 3012 133153 3040
rect 133104 3000 133110 3012
rect 133141 3009 133153 3012
rect 133187 3009 133199 3043
rect 134150 3040 134156 3052
rect 134111 3012 134156 3040
rect 133141 3003 133199 3009
rect 134150 3000 134156 3012
rect 134208 3000 134214 3052
rect 136634 3040 136640 3052
rect 136595 3012 136640 3040
rect 136634 3000 136640 3012
rect 136692 3000 136698 3052
rect 136818 3000 136824 3052
rect 136876 3040 136882 3052
rect 137741 3043 137799 3049
rect 137741 3040 137753 3043
rect 136876 3012 137753 3040
rect 136876 3000 136882 3012
rect 137741 3009 137753 3012
rect 137787 3040 137799 3043
rect 138014 3040 138020 3052
rect 137787 3012 138020 3040
rect 137787 3009 137799 3012
rect 137741 3003 137799 3009
rect 138014 3000 138020 3012
rect 138072 3000 138078 3052
rect 138753 3043 138811 3049
rect 138753 3009 138765 3043
rect 138799 3040 138811 3043
rect 139029 3043 139087 3049
rect 139029 3040 139041 3043
rect 138799 3012 139041 3040
rect 138799 3009 138811 3012
rect 138753 3003 138811 3009
rect 139029 3009 139041 3012
rect 139075 3009 139087 3043
rect 139854 3040 139860 3052
rect 139029 3003 139087 3009
rect 139136 3012 139860 3040
rect 139136 2972 139164 3012
rect 139854 3000 139860 3012
rect 139912 3000 139918 3052
rect 145285 3043 145343 3049
rect 145285 3009 145297 3043
rect 145331 3040 145343 3043
rect 145558 3040 145564 3052
rect 145331 3012 145564 3040
rect 145331 3009 145343 3012
rect 145285 3003 145343 3009
rect 145558 3000 145564 3012
rect 145616 3000 145622 3052
rect 149054 3040 149060 3052
rect 149015 3012 149060 3040
rect 149054 3000 149060 3012
rect 149112 3000 149118 3052
rect 154209 3043 154267 3049
rect 149900 3012 151676 3040
rect 132328 2944 139164 2972
rect 139394 2932 139400 2984
rect 139452 2972 139458 2984
rect 139765 2975 139823 2981
rect 139765 2972 139777 2975
rect 139452 2944 139777 2972
rect 139452 2932 139458 2944
rect 139765 2941 139777 2944
rect 139811 2941 139823 2975
rect 139765 2935 139823 2941
rect 141142 2932 141148 2984
rect 141200 2972 141206 2984
rect 141421 2975 141479 2981
rect 141421 2972 141433 2975
rect 141200 2944 141433 2972
rect 141200 2932 141206 2944
rect 141421 2941 141433 2944
rect 141467 2941 141479 2975
rect 143166 2972 143172 2984
rect 143127 2944 143172 2972
rect 141421 2935 141479 2941
rect 143166 2932 143172 2944
rect 143224 2932 143230 2984
rect 143718 2932 143724 2984
rect 143776 2972 143782 2984
rect 149900 2972 149928 3012
rect 143776 2944 149928 2972
rect 151648 2972 151676 3012
rect 154209 3009 154221 3043
rect 154255 3040 154267 3043
rect 154390 3040 154396 3052
rect 154255 3012 154396 3040
rect 154255 3009 154267 3012
rect 154209 3003 154267 3009
rect 154390 3000 154396 3012
rect 154448 3000 154454 3052
rect 155218 3040 155224 3052
rect 155179 3012 155224 3040
rect 155218 3000 155224 3012
rect 155276 3000 155282 3052
rect 156230 3040 156236 3052
rect 156191 3012 156236 3040
rect 156230 3000 156236 3012
rect 156288 3000 156294 3052
rect 159453 3043 159511 3049
rect 159453 3009 159465 3043
rect 159499 3009 159511 3043
rect 160646 3040 160652 3052
rect 160607 3012 160652 3040
rect 159453 3003 159511 3009
rect 156690 2972 156696 2984
rect 151648 2944 156696 2972
rect 143776 2932 143782 2944
rect 156690 2932 156696 2944
rect 156748 2932 156754 2984
rect 158254 2972 158260 2984
rect 158215 2944 158260 2972
rect 158254 2932 158260 2944
rect 158312 2932 158318 2984
rect 55766 2904 55772 2916
rect 55416 2876 55772 2904
rect 55766 2864 55772 2876
rect 55824 2864 55830 2916
rect 56045 2907 56103 2913
rect 56045 2873 56057 2907
rect 56091 2904 56103 2907
rect 56134 2904 56140 2916
rect 56091 2876 56140 2904
rect 56091 2873 56103 2876
rect 56045 2867 56103 2873
rect 56134 2864 56140 2876
rect 56192 2904 56198 2916
rect 58066 2904 58072 2916
rect 56192 2876 58072 2904
rect 56192 2864 56198 2876
rect 58066 2864 58072 2876
rect 58124 2864 58130 2916
rect 58986 2904 58992 2916
rect 58176 2876 58992 2904
rect 41524 2808 42932 2836
rect 41417 2799 41475 2805
rect 42978 2796 42984 2848
rect 43036 2836 43042 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 43036 2808 48881 2836
rect 43036 2796 43042 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 48958 2796 48964 2848
rect 49016 2836 49022 2848
rect 54202 2836 54208 2848
rect 49016 2808 54208 2836
rect 49016 2796 49022 2808
rect 54202 2796 54208 2808
rect 54260 2796 54266 2848
rect 54570 2836 54576 2848
rect 54531 2808 54576 2836
rect 54570 2796 54576 2808
rect 54628 2796 54634 2848
rect 55217 2839 55275 2845
rect 55217 2805 55229 2839
rect 55263 2836 55275 2839
rect 55398 2836 55404 2848
rect 55263 2808 55404 2836
rect 55263 2805 55275 2808
rect 55217 2799 55275 2805
rect 55398 2796 55404 2808
rect 55456 2796 55462 2848
rect 55490 2796 55496 2848
rect 55548 2836 55554 2848
rect 57330 2836 57336 2848
rect 55548 2808 57336 2836
rect 55548 2796 55554 2808
rect 57330 2796 57336 2808
rect 57388 2796 57394 2848
rect 57698 2796 57704 2848
rect 57756 2836 57762 2848
rect 58176 2836 58204 2876
rect 58986 2864 58992 2876
rect 59044 2864 59050 2916
rect 59446 2864 59452 2916
rect 59504 2904 59510 2916
rect 61197 2907 61255 2913
rect 61197 2904 61209 2907
rect 59504 2876 61209 2904
rect 59504 2864 59510 2876
rect 61197 2873 61209 2876
rect 61243 2873 61255 2907
rect 62758 2904 62764 2916
rect 61197 2867 61255 2873
rect 61304 2876 62764 2904
rect 57756 2808 58204 2836
rect 57756 2796 57762 2808
rect 58802 2796 58808 2848
rect 58860 2836 58866 2848
rect 61304 2836 61332 2876
rect 62758 2864 62764 2876
rect 62816 2864 62822 2916
rect 63494 2864 63500 2916
rect 63552 2904 63558 2916
rect 67174 2904 67180 2916
rect 63552 2876 67180 2904
rect 63552 2864 63558 2876
rect 67174 2864 67180 2876
rect 67232 2864 67238 2916
rect 67358 2864 67364 2916
rect 67416 2904 67422 2916
rect 67416 2876 70440 2904
rect 67416 2864 67422 2876
rect 58860 2808 61332 2836
rect 58860 2796 58866 2808
rect 63218 2796 63224 2848
rect 63276 2836 63282 2848
rect 64598 2836 64604 2848
rect 63276 2808 64604 2836
rect 63276 2796 63282 2808
rect 64598 2796 64604 2808
rect 64656 2796 64662 2848
rect 67726 2796 67732 2848
rect 67784 2836 67790 2848
rect 68557 2839 68615 2845
rect 68557 2836 68569 2839
rect 67784 2808 68569 2836
rect 67784 2796 67790 2808
rect 68557 2805 68569 2808
rect 68603 2805 68615 2839
rect 69566 2836 69572 2848
rect 69527 2808 69572 2836
rect 68557 2799 68615 2805
rect 69566 2796 69572 2808
rect 69624 2796 69630 2848
rect 70412 2836 70440 2876
rect 70486 2864 70492 2916
rect 70544 2904 70550 2916
rect 70581 2907 70639 2913
rect 70581 2904 70593 2907
rect 70544 2876 70593 2904
rect 70544 2864 70550 2876
rect 70581 2873 70593 2876
rect 70627 2873 70639 2907
rect 70581 2867 70639 2873
rect 70946 2864 70952 2916
rect 71004 2904 71010 2916
rect 74902 2904 74908 2916
rect 71004 2876 74908 2904
rect 71004 2864 71010 2876
rect 74902 2864 74908 2876
rect 74960 2864 74966 2916
rect 103425 2907 103483 2913
rect 103425 2873 103437 2907
rect 103471 2904 103483 2907
rect 105262 2904 105268 2916
rect 103471 2876 105268 2904
rect 103471 2873 103483 2876
rect 103425 2867 103483 2873
rect 105262 2864 105268 2876
rect 105320 2864 105326 2916
rect 108850 2904 108856 2916
rect 105372 2876 108856 2904
rect 72418 2836 72424 2848
rect 70412 2808 72424 2836
rect 72418 2796 72424 2808
rect 72476 2796 72482 2848
rect 73249 2839 73307 2845
rect 73249 2805 73261 2839
rect 73295 2836 73307 2839
rect 73798 2836 73804 2848
rect 73295 2808 73804 2836
rect 73295 2805 73307 2808
rect 73249 2799 73307 2805
rect 73798 2796 73804 2808
rect 73856 2796 73862 2848
rect 74258 2796 74264 2848
rect 74316 2836 74322 2848
rect 77294 2836 77300 2848
rect 74316 2808 77300 2836
rect 74316 2796 74322 2808
rect 77294 2796 77300 2808
rect 77352 2796 77358 2848
rect 87414 2836 87420 2848
rect 87375 2808 87420 2836
rect 87414 2796 87420 2808
rect 87472 2796 87478 2848
rect 88518 2796 88524 2848
rect 88576 2836 88582 2848
rect 90358 2836 90364 2848
rect 88576 2808 90364 2836
rect 88576 2796 88582 2808
rect 90358 2796 90364 2808
rect 90416 2796 90422 2848
rect 100110 2796 100116 2848
rect 100168 2836 100174 2848
rect 102413 2839 102471 2845
rect 102413 2836 102425 2839
rect 100168 2808 102425 2836
rect 100168 2796 100174 2808
rect 102413 2805 102425 2808
rect 102459 2805 102471 2839
rect 103238 2836 103244 2848
rect 103199 2808 103244 2836
rect 102413 2799 102471 2805
rect 103238 2796 103244 2808
rect 103296 2796 103302 2848
rect 103882 2836 103888 2848
rect 103843 2808 103888 2836
rect 103882 2796 103888 2808
rect 103940 2796 103946 2848
rect 104250 2796 104256 2848
rect 104308 2836 104314 2848
rect 105372 2836 105400 2876
rect 108850 2864 108856 2876
rect 108908 2864 108914 2916
rect 109604 2876 109908 2904
rect 104308 2808 105400 2836
rect 107565 2839 107623 2845
rect 104308 2796 104314 2808
rect 107565 2805 107577 2839
rect 107611 2836 107623 2839
rect 109604 2836 109632 2876
rect 107611 2808 109632 2836
rect 109880 2836 109908 2876
rect 110322 2864 110328 2916
rect 110380 2904 110386 2916
rect 111426 2904 111432 2916
rect 110380 2876 111432 2904
rect 110380 2864 110386 2876
rect 111426 2864 111432 2876
rect 111484 2864 111490 2916
rect 111610 2864 111616 2916
rect 111668 2904 111674 2916
rect 113729 2907 113787 2913
rect 113729 2904 113741 2907
rect 111668 2876 113741 2904
rect 111668 2864 111674 2876
rect 113729 2873 113741 2876
rect 113775 2873 113787 2907
rect 113729 2867 113787 2873
rect 114554 2864 114560 2916
rect 114612 2904 114618 2916
rect 118694 2904 118700 2916
rect 114612 2876 118700 2904
rect 114612 2864 114618 2876
rect 118694 2864 118700 2876
rect 118752 2864 118758 2916
rect 122374 2864 122380 2916
rect 122432 2904 122438 2916
rect 123846 2904 123852 2916
rect 122432 2876 123852 2904
rect 122432 2864 122438 2876
rect 123846 2864 123852 2876
rect 123904 2864 123910 2916
rect 134518 2904 134524 2916
rect 124048 2876 134524 2904
rect 110690 2836 110696 2848
rect 109880 2808 110696 2836
rect 107611 2805 107623 2808
rect 107565 2799 107623 2805
rect 110690 2796 110696 2808
rect 110748 2796 110754 2848
rect 110874 2796 110880 2848
rect 110932 2836 110938 2848
rect 110969 2839 111027 2845
rect 110969 2836 110981 2839
rect 110932 2808 110981 2836
rect 110932 2796 110938 2808
rect 110969 2805 110981 2808
rect 111015 2805 111027 2839
rect 110969 2799 111027 2805
rect 111058 2796 111064 2848
rect 111116 2836 111122 2848
rect 116118 2836 116124 2848
rect 111116 2808 116124 2836
rect 111116 2796 111122 2808
rect 116118 2796 116124 2808
rect 116176 2796 116182 2848
rect 116210 2796 116216 2848
rect 116268 2836 116274 2848
rect 117225 2839 117283 2845
rect 117225 2836 117237 2839
rect 116268 2808 117237 2836
rect 116268 2796 116274 2808
rect 117225 2805 117237 2808
rect 117271 2805 117283 2839
rect 117225 2799 117283 2805
rect 122650 2796 122656 2848
rect 122708 2836 122714 2848
rect 124048 2836 124076 2876
rect 134518 2864 134524 2876
rect 134576 2864 134582 2916
rect 137833 2907 137891 2913
rect 137833 2873 137845 2907
rect 137879 2904 137891 2907
rect 139670 2904 139676 2916
rect 137879 2876 139676 2904
rect 137879 2873 137891 2876
rect 137833 2867 137891 2873
rect 139670 2864 139676 2876
rect 139728 2864 139734 2916
rect 142614 2864 142620 2916
rect 142672 2904 142678 2916
rect 151354 2904 151360 2916
rect 142672 2876 151360 2904
rect 142672 2864 142678 2876
rect 151354 2864 151360 2876
rect 151412 2864 151418 2916
rect 151998 2864 152004 2916
rect 152056 2904 152062 2916
rect 152056 2876 157288 2904
rect 152056 2864 152062 2876
rect 122708 2808 124076 2836
rect 122708 2796 122714 2808
rect 126882 2796 126888 2848
rect 126940 2836 126946 2848
rect 127894 2836 127900 2848
rect 126940 2808 127900 2836
rect 126940 2796 126946 2808
rect 127894 2796 127900 2808
rect 127952 2796 127958 2848
rect 130013 2839 130071 2845
rect 130013 2805 130025 2839
rect 130059 2836 130071 2839
rect 135438 2836 135444 2848
rect 130059 2808 135444 2836
rect 130059 2805 130071 2808
rect 130013 2799 130071 2805
rect 135438 2796 135444 2808
rect 135496 2796 135502 2848
rect 136726 2836 136732 2848
rect 136687 2808 136732 2836
rect 136726 2796 136732 2808
rect 136784 2796 136790 2848
rect 136910 2796 136916 2848
rect 136968 2836 136974 2848
rect 138845 2839 138903 2845
rect 138845 2836 138857 2839
rect 136968 2808 138857 2836
rect 136968 2796 136974 2808
rect 138845 2805 138857 2808
rect 138891 2805 138903 2839
rect 138845 2799 138903 2805
rect 139029 2839 139087 2845
rect 139029 2805 139041 2839
rect 139075 2836 139087 2839
rect 139305 2839 139363 2845
rect 139305 2836 139317 2839
rect 139075 2808 139317 2836
rect 139075 2805 139087 2808
rect 139029 2799 139087 2805
rect 139305 2805 139317 2808
rect 139351 2836 139363 2839
rect 140958 2836 140964 2848
rect 139351 2808 140964 2836
rect 139351 2805 139363 2808
rect 139305 2799 139363 2805
rect 140958 2796 140964 2808
rect 141016 2796 141022 2848
rect 142246 2796 142252 2848
rect 142304 2836 142310 2848
rect 145742 2836 145748 2848
rect 142304 2808 145748 2836
rect 142304 2796 142310 2808
rect 145742 2796 145748 2808
rect 145800 2796 145806 2848
rect 149146 2836 149152 2848
rect 149107 2808 149152 2836
rect 149146 2796 149152 2808
rect 149204 2796 149210 2848
rect 149238 2796 149244 2848
rect 149296 2836 149302 2848
rect 150894 2836 150900 2848
rect 149296 2808 150900 2836
rect 149296 2796 149302 2808
rect 150894 2796 150900 2808
rect 150952 2796 150958 2848
rect 157260 2836 157288 2876
rect 158806 2864 158812 2916
rect 158864 2904 158870 2916
rect 159468 2904 159496 3003
rect 160646 3000 160652 3012
rect 160704 3000 160710 3052
rect 163961 3043 164019 3049
rect 163961 3009 163973 3043
rect 164007 3040 164019 3043
rect 164142 3040 164148 3052
rect 164007 3012 164148 3040
rect 164007 3009 164019 3012
rect 163961 3003 164019 3009
rect 164142 3000 164148 3012
rect 164200 3000 164206 3052
rect 164973 3043 165031 3049
rect 164973 3009 164985 3043
rect 165019 3040 165031 3043
rect 165062 3040 165068 3052
rect 165019 3012 165068 3040
rect 165019 3009 165031 3012
rect 164973 3003 165031 3009
rect 165062 3000 165068 3012
rect 165120 3040 165126 3052
rect 165433 3043 165491 3049
rect 165433 3040 165445 3043
rect 165120 3012 165445 3040
rect 165120 3000 165126 3012
rect 165433 3009 165445 3012
rect 165479 3009 165491 3043
rect 165433 3003 165491 3009
rect 162026 2972 162032 2984
rect 161987 2944 162032 2972
rect 162026 2932 162032 2944
rect 162084 2932 162090 2984
rect 160186 2904 160192 2916
rect 158864 2876 160192 2904
rect 158864 2864 158870 2876
rect 160186 2864 160192 2876
rect 160244 2864 160250 2916
rect 159818 2836 159824 2848
rect 157260 2808 159824 2836
rect 159818 2796 159824 2808
rect 159876 2796 159882 2848
rect 164602 2796 164608 2848
rect 164660 2836 164666 2848
rect 164697 2839 164755 2845
rect 164697 2836 164709 2839
rect 164660 2808 164709 2836
rect 164660 2796 164666 2808
rect 164697 2805 164709 2808
rect 164743 2805 164755 2839
rect 164697 2799 164755 2805
rect 368 2746 93012 2768
rect 368 2694 28456 2746
rect 28508 2694 28520 2746
rect 28572 2694 28584 2746
rect 28636 2694 28648 2746
rect 28700 2694 84878 2746
rect 84930 2694 84942 2746
rect 84994 2694 85006 2746
rect 85058 2694 85070 2746
rect 85122 2694 93012 2746
rect 368 2672 93012 2694
rect 102028 2746 169556 2768
rect 102028 2694 141299 2746
rect 141351 2694 141363 2746
rect 141415 2694 141427 2746
rect 141479 2694 141491 2746
rect 141543 2694 169556 2746
rect 102028 2672 169556 2694
rect 3694 2632 3700 2644
rect 3655 2604 3700 2632
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 3881 2635 3939 2641
rect 3881 2601 3893 2635
rect 3927 2632 3939 2635
rect 4706 2632 4712 2644
rect 3927 2604 4712 2632
rect 3927 2601 3939 2604
rect 3881 2595 3939 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 22557 2635 22615 2641
rect 12216 2604 22508 2632
rect 12216 2592 12222 2604
rect 566 2524 572 2576
rect 624 2564 630 2576
rect 9490 2564 9496 2576
rect 624 2536 9496 2564
rect 624 2524 630 2536
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 18322 2564 18328 2576
rect 18283 2536 18328 2564
rect 18322 2524 18328 2536
rect 18380 2524 18386 2576
rect 19981 2567 20039 2573
rect 19981 2533 19993 2567
rect 20027 2564 20039 2567
rect 20530 2564 20536 2576
rect 20027 2536 20536 2564
rect 20027 2533 20039 2536
rect 19981 2527 20039 2533
rect 20530 2524 20536 2536
rect 20588 2524 20594 2576
rect 21637 2567 21695 2573
rect 21637 2533 21649 2567
rect 21683 2564 21695 2567
rect 21726 2564 21732 2576
rect 21683 2536 21732 2564
rect 21683 2533 21695 2536
rect 21637 2527 21695 2533
rect 21726 2524 21732 2536
rect 21784 2524 21790 2576
rect 22480 2564 22508 2604
rect 22557 2601 22569 2635
rect 22603 2632 22615 2635
rect 22833 2635 22891 2641
rect 22833 2632 22845 2635
rect 22603 2604 22845 2632
rect 22603 2601 22615 2604
rect 22557 2595 22615 2601
rect 22833 2601 22845 2604
rect 22879 2632 22891 2635
rect 23014 2632 23020 2644
rect 22879 2604 23020 2632
rect 22879 2601 22891 2604
rect 22833 2595 22891 2601
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 23750 2632 23756 2644
rect 23711 2604 23756 2632
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 24673 2635 24731 2641
rect 24673 2601 24685 2635
rect 24719 2632 24731 2635
rect 24949 2635 25007 2641
rect 24949 2632 24961 2635
rect 24719 2604 24961 2632
rect 24719 2601 24731 2604
rect 24673 2595 24731 2601
rect 24949 2601 24961 2604
rect 24995 2632 25007 2635
rect 25130 2632 25136 2644
rect 24995 2604 25136 2632
rect 24995 2601 25007 2604
rect 24949 2595 25007 2601
rect 25130 2592 25136 2604
rect 25188 2592 25194 2644
rect 25406 2632 25412 2644
rect 25367 2604 25412 2632
rect 25406 2592 25412 2604
rect 25464 2592 25470 2644
rect 27249 2635 27307 2641
rect 27249 2601 27261 2635
rect 27295 2632 27307 2635
rect 27430 2632 27436 2644
rect 27295 2604 27436 2632
rect 27295 2601 27307 2604
rect 27249 2595 27307 2601
rect 27430 2592 27436 2604
rect 27488 2592 27494 2644
rect 28258 2592 28264 2644
rect 28316 2632 28322 2644
rect 28810 2632 28816 2644
rect 28316 2604 28816 2632
rect 28316 2592 28322 2604
rect 28810 2592 28816 2604
rect 28868 2592 28874 2644
rect 29638 2632 29644 2644
rect 29599 2604 29644 2632
rect 29638 2592 29644 2604
rect 29696 2592 29702 2644
rect 30926 2632 30932 2644
rect 30887 2604 30932 2632
rect 30926 2592 30932 2604
rect 30984 2632 30990 2644
rect 35066 2632 35072 2644
rect 30984 2604 35072 2632
rect 30984 2592 30990 2604
rect 35066 2592 35072 2604
rect 35124 2592 35130 2644
rect 35342 2592 35348 2644
rect 35400 2632 35406 2644
rect 38010 2632 38016 2644
rect 35400 2604 38016 2632
rect 35400 2592 35406 2604
rect 38010 2592 38016 2604
rect 38068 2592 38074 2644
rect 38378 2592 38384 2644
rect 38436 2632 38442 2644
rect 39577 2635 39635 2641
rect 39577 2632 39589 2635
rect 38436 2604 39589 2632
rect 38436 2592 38442 2604
rect 39577 2601 39589 2604
rect 39623 2601 39635 2635
rect 39577 2595 39635 2601
rect 39666 2592 39672 2644
rect 39724 2632 39730 2644
rect 39724 2604 40080 2632
rect 39724 2592 39730 2604
rect 26050 2564 26056 2576
rect 22480 2536 26056 2564
rect 26050 2524 26056 2536
rect 26108 2524 26114 2576
rect 26510 2524 26516 2576
rect 26568 2564 26574 2576
rect 39942 2564 39948 2576
rect 26568 2536 37964 2564
rect 26568 2524 26574 2536
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 4801 2499 4859 2505
rect 4801 2496 4813 2499
rect 2271 2468 4813 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 4801 2465 4813 2468
rect 4847 2496 4859 2499
rect 5534 2496 5540 2508
rect 4847 2468 5540 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5810 2496 5816 2508
rect 5771 2468 5816 2496
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 9766 2496 9772 2508
rect 9631 2468 9772 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 10686 2496 10692 2508
rect 10647 2468 10692 2496
rect 10686 2456 10692 2468
rect 10744 2456 10750 2508
rect 11609 2499 11667 2505
rect 11609 2496 11621 2499
rect 11256 2468 11621 2496
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3786 2388 3792 2400
rect 3844 2428 3850 2440
rect 11256 2437 11284 2468
rect 11609 2465 11621 2468
rect 11655 2496 11667 2499
rect 11655 2468 20576 2496
rect 11655 2465 11667 2468
rect 11609 2459 11667 2465
rect 4249 2431 4307 2437
rect 4249 2428 4261 2431
rect 3844 2400 4261 2428
rect 3844 2388 3850 2400
rect 4249 2397 4261 2400
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 11241 2431 11299 2437
rect 11241 2397 11253 2431
rect 11287 2397 11299 2431
rect 18506 2428 18512 2440
rect 18467 2400 18512 2428
rect 11241 2391 11299 2397
rect 6380 2360 6408 2391
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 6380 2332 6745 2360
rect 6733 2329 6745 2332
rect 6779 2360 6791 2363
rect 9217 2363 9275 2369
rect 6779 2332 8340 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7190 2292 7196 2304
rect 7151 2264 7196 2292
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2292 7803 2295
rect 7834 2292 7840 2304
rect 7791 2264 7840 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 8312 2292 8340 2332
rect 9217 2329 9229 2363
rect 9263 2360 9275 2363
rect 9692 2360 9720 2391
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 18874 2428 18880 2440
rect 18835 2400 18880 2428
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 19610 2428 19616 2440
rect 19291 2400 19616 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 19610 2388 19616 2400
rect 19668 2388 19674 2440
rect 20254 2428 20260 2440
rect 20215 2400 20260 2428
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 20548 2428 20576 2468
rect 20732 2468 23428 2496
rect 20732 2428 20760 2468
rect 20548 2400 20760 2428
rect 21082 2388 21088 2440
rect 21140 2428 21146 2440
rect 21177 2431 21235 2437
rect 21177 2428 21189 2431
rect 21140 2400 21189 2428
rect 21140 2388 21146 2400
rect 21177 2397 21189 2400
rect 21223 2397 21235 2431
rect 21177 2391 21235 2397
rect 21453 2431 21511 2437
rect 21453 2397 21465 2431
rect 21499 2428 21511 2431
rect 22373 2431 22431 2437
rect 21499 2400 22324 2428
rect 21499 2397 21511 2400
rect 21453 2391 21511 2397
rect 12069 2363 12127 2369
rect 12069 2360 12081 2363
rect 9263 2332 12081 2360
rect 9263 2329 9275 2332
rect 9217 2323 9275 2329
rect 12069 2329 12081 2332
rect 12115 2329 12127 2363
rect 12069 2323 12127 2329
rect 13081 2363 13139 2369
rect 13081 2329 13093 2363
rect 13127 2360 13139 2363
rect 13262 2360 13268 2372
rect 13127 2332 13268 2360
rect 13127 2329 13139 2332
rect 13081 2323 13139 2329
rect 13262 2320 13268 2332
rect 13320 2360 13326 2372
rect 13320 2332 20668 2360
rect 13320 2320 13326 2332
rect 10318 2292 10324 2304
rect 8312 2264 10324 2292
rect 10318 2252 10324 2264
rect 10376 2252 10382 2304
rect 19610 2292 19616 2304
rect 19571 2264 19616 2292
rect 19610 2252 19616 2264
rect 19668 2252 19674 2304
rect 19702 2252 19708 2304
rect 19760 2292 19766 2304
rect 20441 2295 20499 2301
rect 20441 2292 20453 2295
rect 19760 2264 20453 2292
rect 19760 2252 19766 2264
rect 20441 2261 20453 2264
rect 20487 2261 20499 2295
rect 20640 2292 20668 2332
rect 21453 2295 21511 2301
rect 21453 2292 21465 2295
rect 20640 2264 21465 2292
rect 20441 2255 20499 2261
rect 21453 2261 21465 2264
rect 21499 2261 21511 2295
rect 22186 2292 22192 2304
rect 22147 2264 22192 2292
rect 21453 2255 21511 2261
rect 22186 2252 22192 2264
rect 22244 2252 22250 2304
rect 22296 2292 22324 2400
rect 22373 2397 22385 2431
rect 22419 2428 22431 2431
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 22419 2400 22569 2428
rect 22419 2397 22431 2400
rect 22373 2391 22431 2397
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 23400 2360 23428 2468
rect 23474 2456 23480 2508
rect 23532 2496 23538 2508
rect 23845 2499 23903 2505
rect 23845 2496 23857 2499
rect 23532 2468 23857 2496
rect 23532 2456 23538 2468
rect 23845 2465 23857 2468
rect 23891 2465 23903 2499
rect 23845 2459 23903 2465
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 28353 2499 28411 2505
rect 28353 2496 28365 2499
rect 23992 2468 28365 2496
rect 23992 2456 23998 2468
rect 28353 2465 28365 2468
rect 28399 2465 28411 2499
rect 29273 2499 29331 2505
rect 29273 2496 29285 2499
rect 28353 2459 28411 2465
rect 28920 2468 29285 2496
rect 24489 2431 24547 2437
rect 24489 2397 24501 2431
rect 24535 2428 24547 2431
rect 24673 2431 24731 2437
rect 24673 2428 24685 2431
rect 24535 2400 24685 2428
rect 24535 2397 24547 2400
rect 24489 2391 24547 2397
rect 24673 2397 24685 2400
rect 24719 2397 24731 2431
rect 25774 2428 25780 2440
rect 25735 2400 25780 2428
rect 24673 2391 24731 2397
rect 25774 2388 25780 2400
rect 25832 2388 25838 2440
rect 26142 2428 26148 2440
rect 26103 2400 26148 2428
rect 26142 2388 26148 2400
rect 26200 2388 26206 2440
rect 26513 2431 26571 2437
rect 26513 2397 26525 2431
rect 26559 2428 26571 2431
rect 26605 2431 26663 2437
rect 26605 2428 26617 2431
rect 26559 2400 26617 2428
rect 26559 2397 26571 2400
rect 26513 2391 26571 2397
rect 26605 2397 26617 2400
rect 26651 2397 26663 2431
rect 27338 2428 27344 2440
rect 27299 2400 27344 2428
rect 26605 2391 26663 2397
rect 27338 2388 27344 2400
rect 27396 2388 27402 2440
rect 28920 2437 28948 2468
rect 29273 2465 29285 2468
rect 29319 2496 29331 2499
rect 35710 2496 35716 2508
rect 29319 2468 35716 2496
rect 29319 2465 29331 2468
rect 29273 2459 29331 2465
rect 35710 2456 35716 2468
rect 35768 2456 35774 2508
rect 35802 2456 35808 2508
rect 35860 2496 35866 2508
rect 36998 2496 37004 2508
rect 35860 2468 37004 2496
rect 35860 2456 35866 2468
rect 36998 2456 37004 2468
rect 37056 2456 37062 2508
rect 37936 2496 37964 2536
rect 38672 2536 39948 2564
rect 38672 2496 38700 2536
rect 39942 2524 39948 2536
rect 40000 2524 40006 2576
rect 40052 2564 40080 2604
rect 40218 2592 40224 2644
rect 40276 2632 40282 2644
rect 41322 2632 41328 2644
rect 40276 2604 40321 2632
rect 40420 2604 41328 2632
rect 40276 2592 40282 2604
rect 40420 2564 40448 2604
rect 41322 2592 41328 2604
rect 41380 2592 41386 2644
rect 41417 2635 41475 2641
rect 41417 2601 41429 2635
rect 41463 2632 41475 2635
rect 41874 2632 41880 2644
rect 41463 2604 41880 2632
rect 41463 2601 41475 2604
rect 41417 2595 41475 2601
rect 41874 2592 41880 2604
rect 41932 2592 41938 2644
rect 42426 2592 42432 2644
rect 42484 2632 42490 2644
rect 43165 2635 43223 2641
rect 43165 2632 43177 2635
rect 42484 2604 43177 2632
rect 42484 2592 42490 2604
rect 43165 2601 43177 2604
rect 43211 2601 43223 2635
rect 43165 2595 43223 2601
rect 43349 2635 43407 2641
rect 43349 2601 43361 2635
rect 43395 2632 43407 2635
rect 43625 2635 43683 2641
rect 43625 2632 43637 2635
rect 43395 2604 43637 2632
rect 43395 2601 43407 2604
rect 43349 2595 43407 2601
rect 43625 2601 43637 2604
rect 43671 2632 43683 2635
rect 44082 2632 44088 2644
rect 43671 2604 44088 2632
rect 43671 2601 43683 2604
rect 43625 2595 43683 2601
rect 44082 2592 44088 2604
rect 44140 2592 44146 2644
rect 44174 2592 44180 2644
rect 44232 2632 44238 2644
rect 44913 2635 44971 2641
rect 44913 2632 44925 2635
rect 44232 2604 44925 2632
rect 44232 2592 44238 2604
rect 44913 2601 44925 2604
rect 44959 2601 44971 2635
rect 45554 2632 45560 2644
rect 45515 2604 45560 2632
rect 44913 2595 44971 2601
rect 45554 2592 45560 2604
rect 45612 2592 45618 2644
rect 45664 2604 45968 2632
rect 40052 2536 40448 2564
rect 40494 2524 40500 2576
rect 40552 2564 40558 2576
rect 45664 2564 45692 2604
rect 45830 2564 45836 2576
rect 40552 2536 45692 2564
rect 45756 2536 45836 2564
rect 40552 2524 40558 2536
rect 37936 2468 38700 2496
rect 38746 2456 38752 2508
rect 38804 2496 38810 2508
rect 39577 2499 39635 2505
rect 38804 2468 39436 2496
rect 38804 2456 38810 2468
rect 39408 2440 39436 2468
rect 39577 2465 39589 2499
rect 39623 2496 39635 2499
rect 39623 2468 40724 2496
rect 39623 2465 39635 2468
rect 39577 2459 39635 2465
rect 28905 2431 28963 2437
rect 28905 2397 28917 2431
rect 28951 2397 28963 2431
rect 32674 2428 32680 2440
rect 28905 2391 28963 2397
rect 29012 2400 32680 2428
rect 29012 2360 29040 2400
rect 32674 2388 32680 2400
rect 32732 2388 32738 2440
rect 32766 2388 32772 2440
rect 32824 2428 32830 2440
rect 35250 2428 35256 2440
rect 32824 2400 35256 2428
rect 32824 2388 32830 2400
rect 35250 2388 35256 2400
rect 35308 2388 35314 2440
rect 35526 2388 35532 2440
rect 35584 2428 35590 2440
rect 36262 2428 36268 2440
rect 35584 2400 36268 2428
rect 35584 2388 35590 2400
rect 36262 2388 36268 2400
rect 36320 2388 36326 2440
rect 36354 2388 36360 2440
rect 36412 2428 36418 2440
rect 36541 2431 36599 2437
rect 36541 2428 36553 2431
rect 36412 2400 36553 2428
rect 36412 2388 36418 2400
rect 36541 2397 36553 2400
rect 36587 2397 36599 2431
rect 36541 2391 36599 2397
rect 36630 2388 36636 2440
rect 36688 2428 36694 2440
rect 38654 2428 38660 2440
rect 36688 2400 38660 2428
rect 36688 2388 36694 2400
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 38930 2388 38936 2440
rect 38988 2428 38994 2440
rect 39114 2428 39120 2440
rect 38988 2400 39033 2428
rect 39075 2400 39120 2428
rect 38988 2388 38994 2400
rect 39114 2388 39120 2400
rect 39172 2388 39178 2440
rect 39390 2388 39396 2440
rect 39448 2388 39454 2440
rect 39485 2431 39543 2437
rect 39485 2397 39497 2431
rect 39531 2428 39543 2431
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39531 2400 39865 2428
rect 39531 2397 39543 2400
rect 39485 2391 39543 2397
rect 39853 2397 39865 2400
rect 39899 2428 39911 2431
rect 40494 2428 40500 2440
rect 39899 2400 40500 2428
rect 39899 2397 39911 2400
rect 39853 2391 39911 2397
rect 40494 2388 40500 2400
rect 40552 2388 40558 2440
rect 40696 2428 40724 2468
rect 40862 2456 40868 2508
rect 40920 2496 40926 2508
rect 41966 2496 41972 2508
rect 40920 2468 41972 2496
rect 40920 2456 40926 2468
rect 41966 2456 41972 2468
rect 42024 2456 42030 2508
rect 43898 2496 43904 2508
rect 42996 2468 43904 2496
rect 41138 2428 41144 2440
rect 40696 2400 41144 2428
rect 41138 2388 41144 2400
rect 41196 2388 41202 2440
rect 42996 2428 43024 2468
rect 43898 2456 43904 2468
rect 43956 2456 43962 2508
rect 44266 2496 44272 2508
rect 44008 2468 44272 2496
rect 42076 2400 43024 2428
rect 43073 2431 43131 2437
rect 42076 2360 42104 2400
rect 43073 2397 43085 2431
rect 43119 2428 43131 2431
rect 43349 2431 43407 2437
rect 43349 2428 43361 2431
rect 43119 2400 43361 2428
rect 43119 2397 43131 2400
rect 43073 2391 43131 2397
rect 43349 2397 43361 2400
rect 43395 2397 43407 2431
rect 44008 2428 44036 2468
rect 44266 2456 44272 2468
rect 44324 2456 44330 2508
rect 45189 2499 45247 2505
rect 45189 2496 45201 2499
rect 44744 2468 45201 2496
rect 43349 2391 43407 2397
rect 43456 2400 44036 2428
rect 44085 2431 44143 2437
rect 43456 2360 43484 2400
rect 44085 2397 44097 2431
rect 44131 2397 44143 2431
rect 44085 2391 44143 2397
rect 23400 2332 29040 2360
rect 29104 2332 42104 2360
rect 42536 2332 43484 2360
rect 43993 2363 44051 2369
rect 26510 2292 26516 2304
rect 22296 2264 26516 2292
rect 26510 2252 26516 2264
rect 26568 2252 26574 2304
rect 26605 2295 26663 2301
rect 26605 2261 26617 2295
rect 26651 2292 26663 2295
rect 26881 2295 26939 2301
rect 26881 2292 26893 2295
rect 26651 2264 26893 2292
rect 26651 2261 26663 2264
rect 26605 2255 26663 2261
rect 26881 2261 26893 2264
rect 26927 2292 26939 2295
rect 29104 2292 29132 2332
rect 26927 2264 29132 2292
rect 30285 2295 30343 2301
rect 26927 2261 26939 2264
rect 26881 2255 26939 2261
rect 30285 2261 30297 2295
rect 30331 2292 30343 2295
rect 30834 2292 30840 2304
rect 30331 2264 30840 2292
rect 30331 2261 30343 2264
rect 30285 2255 30343 2261
rect 30834 2252 30840 2264
rect 30892 2252 30898 2304
rect 31846 2252 31852 2304
rect 31904 2292 31910 2304
rect 35342 2292 35348 2304
rect 31904 2264 35348 2292
rect 31904 2252 31910 2264
rect 35342 2252 35348 2264
rect 35400 2252 35406 2304
rect 35618 2252 35624 2304
rect 35676 2292 35682 2304
rect 42536 2292 42564 2332
rect 43993 2329 44005 2363
rect 44039 2360 44051 2363
rect 44100 2360 44128 2391
rect 44174 2388 44180 2440
rect 44232 2428 44238 2440
rect 44744 2437 44772 2468
rect 45189 2465 45201 2468
rect 45235 2496 45247 2499
rect 45756 2496 45784 2536
rect 45830 2524 45836 2536
rect 45888 2524 45894 2576
rect 45940 2564 45968 2604
rect 46198 2592 46204 2644
rect 46256 2632 46262 2644
rect 46474 2632 46480 2644
rect 46256 2604 46480 2632
rect 46256 2592 46262 2604
rect 46474 2592 46480 2604
rect 46532 2592 46538 2644
rect 46566 2592 46572 2644
rect 46624 2632 46630 2644
rect 47026 2632 47032 2644
rect 46624 2604 47032 2632
rect 46624 2592 46630 2604
rect 47026 2592 47032 2604
rect 47084 2592 47090 2644
rect 47210 2592 47216 2644
rect 47268 2632 47274 2644
rect 47489 2635 47547 2641
rect 47489 2632 47501 2635
rect 47268 2604 47501 2632
rect 47268 2592 47274 2604
rect 47489 2601 47501 2604
rect 47535 2601 47547 2635
rect 47489 2595 47547 2601
rect 47762 2592 47768 2644
rect 47820 2632 47826 2644
rect 48866 2632 48872 2644
rect 47820 2604 48872 2632
rect 47820 2592 47826 2604
rect 48866 2592 48872 2604
rect 48924 2592 48930 2644
rect 49050 2632 49056 2644
rect 49011 2604 49056 2632
rect 49050 2592 49056 2604
rect 49108 2592 49114 2644
rect 49142 2592 49148 2644
rect 49200 2632 49206 2644
rect 50798 2632 50804 2644
rect 49200 2604 50804 2632
rect 49200 2592 49206 2604
rect 50798 2592 50804 2604
rect 50856 2592 50862 2644
rect 50890 2592 50896 2644
rect 50948 2632 50954 2644
rect 51718 2632 51724 2644
rect 50948 2604 51724 2632
rect 50948 2592 50954 2604
rect 51718 2592 51724 2604
rect 51776 2592 51782 2644
rect 52822 2632 52828 2644
rect 52783 2604 52828 2632
rect 52822 2592 52828 2604
rect 52880 2592 52886 2644
rect 53282 2632 53288 2644
rect 53243 2604 53288 2632
rect 53282 2592 53288 2604
rect 53340 2592 53346 2644
rect 53650 2632 53656 2644
rect 53611 2604 53656 2632
rect 53650 2592 53656 2604
rect 53708 2592 53714 2644
rect 55214 2632 55220 2644
rect 55175 2604 55220 2632
rect 55214 2592 55220 2604
rect 55272 2592 55278 2644
rect 55674 2592 55680 2644
rect 55732 2632 55738 2644
rect 56226 2632 56232 2644
rect 55732 2604 56232 2632
rect 55732 2592 55738 2604
rect 56226 2592 56232 2604
rect 56284 2592 56290 2644
rect 56689 2635 56747 2641
rect 56689 2601 56701 2635
rect 56735 2632 56747 2635
rect 57054 2632 57060 2644
rect 56735 2604 57060 2632
rect 56735 2601 56747 2604
rect 56689 2595 56747 2601
rect 57054 2592 57060 2604
rect 57112 2592 57118 2644
rect 57146 2592 57152 2644
rect 57204 2632 57210 2644
rect 57241 2635 57299 2641
rect 57241 2632 57253 2635
rect 57204 2604 57253 2632
rect 57204 2592 57210 2604
rect 57241 2601 57253 2604
rect 57287 2601 57299 2635
rect 57241 2595 57299 2601
rect 58713 2635 58771 2641
rect 58713 2601 58725 2635
rect 58759 2632 58771 2635
rect 58802 2632 58808 2644
rect 58759 2604 58808 2632
rect 58759 2601 58771 2604
rect 58713 2595 58771 2601
rect 58802 2592 58808 2604
rect 58860 2592 58866 2644
rect 60369 2635 60427 2641
rect 60369 2601 60381 2635
rect 60415 2632 60427 2635
rect 60734 2632 60740 2644
rect 60415 2604 60740 2632
rect 60415 2601 60427 2604
rect 60369 2595 60427 2601
rect 60734 2592 60740 2604
rect 60792 2592 60798 2644
rect 60918 2632 60924 2644
rect 60879 2604 60924 2632
rect 60918 2592 60924 2604
rect 60976 2592 60982 2644
rect 61286 2632 61292 2644
rect 61247 2604 61292 2632
rect 61286 2592 61292 2604
rect 61344 2592 61350 2644
rect 62574 2632 62580 2644
rect 61396 2604 62580 2632
rect 61396 2564 61424 2604
rect 62574 2592 62580 2604
rect 62632 2592 62638 2644
rect 62669 2635 62727 2641
rect 62669 2601 62681 2635
rect 62715 2632 62727 2635
rect 62850 2632 62856 2644
rect 62715 2604 62856 2632
rect 62715 2601 62727 2604
rect 62669 2595 62727 2601
rect 62850 2592 62856 2604
rect 62908 2592 62914 2644
rect 63494 2632 63500 2644
rect 63455 2604 63500 2632
rect 63494 2592 63500 2604
rect 63552 2592 63558 2644
rect 63678 2632 63684 2644
rect 63639 2604 63684 2632
rect 63678 2592 63684 2604
rect 63736 2592 63742 2644
rect 64506 2632 64512 2644
rect 64467 2604 64512 2632
rect 64506 2592 64512 2604
rect 64564 2592 64570 2644
rect 66530 2632 66536 2644
rect 66491 2604 66536 2632
rect 66530 2592 66536 2604
rect 66588 2592 66594 2644
rect 67542 2632 67548 2644
rect 67503 2604 67548 2632
rect 67542 2592 67548 2604
rect 67600 2592 67606 2644
rect 68554 2632 68560 2644
rect 68515 2604 68560 2632
rect 68554 2592 68560 2604
rect 68612 2592 68618 2644
rect 70121 2635 70179 2641
rect 70121 2601 70133 2635
rect 70167 2632 70179 2635
rect 70210 2632 70216 2644
rect 70167 2604 70216 2632
rect 70167 2601 70179 2604
rect 70121 2595 70179 2601
rect 70210 2592 70216 2604
rect 70268 2592 70274 2644
rect 70489 2635 70547 2641
rect 70489 2601 70501 2635
rect 70535 2632 70547 2635
rect 70578 2632 70584 2644
rect 70535 2604 70584 2632
rect 70535 2601 70547 2604
rect 70489 2595 70547 2601
rect 70578 2592 70584 2604
rect 70636 2592 70642 2644
rect 71130 2592 71136 2644
rect 71188 2632 71194 2644
rect 71593 2635 71651 2641
rect 71593 2632 71605 2635
rect 71188 2604 71605 2632
rect 71188 2592 71194 2604
rect 71593 2601 71605 2604
rect 71639 2632 71651 2635
rect 71682 2632 71688 2644
rect 71639 2604 71688 2632
rect 71639 2601 71651 2604
rect 71593 2595 71651 2601
rect 71682 2592 71688 2604
rect 71740 2592 71746 2644
rect 71866 2632 71872 2644
rect 71827 2604 71872 2632
rect 71866 2592 71872 2604
rect 71924 2592 71930 2644
rect 72142 2592 72148 2644
rect 72200 2632 72206 2644
rect 73525 2635 73583 2641
rect 73525 2632 73537 2635
rect 72200 2604 73537 2632
rect 72200 2592 72206 2604
rect 73525 2601 73537 2604
rect 73571 2601 73583 2635
rect 74258 2632 74264 2644
rect 74219 2604 74264 2632
rect 73525 2595 73583 2601
rect 74258 2592 74264 2604
rect 74316 2592 74322 2644
rect 74629 2635 74687 2641
rect 74629 2601 74641 2635
rect 74675 2632 74687 2635
rect 74718 2632 74724 2644
rect 74675 2604 74724 2632
rect 74675 2601 74687 2604
rect 74629 2595 74687 2601
rect 74718 2592 74724 2604
rect 74776 2592 74782 2644
rect 74813 2635 74871 2641
rect 74813 2601 74825 2635
rect 74859 2632 74871 2635
rect 75089 2635 75147 2641
rect 75089 2632 75101 2635
rect 74859 2604 75101 2632
rect 74859 2601 74871 2604
rect 74813 2595 74871 2601
rect 75089 2601 75101 2604
rect 75135 2632 75147 2635
rect 79686 2632 79692 2644
rect 75135 2604 79692 2632
rect 75135 2601 75147 2604
rect 75089 2595 75147 2601
rect 79686 2592 79692 2604
rect 79744 2592 79750 2644
rect 80793 2635 80851 2641
rect 80793 2601 80805 2635
rect 80839 2632 80851 2635
rect 80882 2632 80888 2644
rect 80839 2604 80888 2632
rect 80839 2601 80851 2604
rect 80793 2595 80851 2601
rect 80882 2592 80888 2604
rect 80940 2592 80946 2644
rect 81986 2632 81992 2644
rect 81947 2604 81992 2632
rect 81986 2592 81992 2604
rect 82044 2592 82050 2644
rect 83458 2632 83464 2644
rect 83419 2604 83464 2632
rect 83458 2592 83464 2604
rect 83516 2592 83522 2644
rect 83550 2592 83556 2644
rect 83608 2632 83614 2644
rect 86954 2632 86960 2644
rect 83608 2604 85896 2632
rect 86915 2604 86960 2632
rect 83608 2592 83614 2604
rect 45940 2536 61424 2564
rect 61470 2524 61476 2576
rect 61528 2564 61534 2576
rect 85758 2564 85764 2576
rect 61528 2536 85764 2564
rect 61528 2524 61534 2536
rect 85758 2524 85764 2536
rect 85816 2524 85822 2576
rect 85868 2564 85896 2604
rect 86954 2592 86960 2604
rect 87012 2592 87018 2644
rect 87322 2632 87328 2644
rect 87283 2604 87328 2632
rect 87322 2592 87328 2604
rect 87380 2592 87386 2644
rect 87598 2632 87604 2644
rect 87559 2604 87604 2632
rect 87598 2592 87604 2604
rect 87656 2592 87662 2644
rect 88426 2632 88432 2644
rect 88387 2604 88432 2632
rect 88426 2592 88432 2604
rect 88484 2592 88490 2644
rect 90266 2632 90272 2644
rect 90227 2604 90272 2632
rect 90266 2592 90272 2604
rect 90324 2592 90330 2644
rect 102134 2592 102140 2644
rect 102192 2632 102198 2644
rect 102962 2632 102968 2644
rect 102192 2604 102968 2632
rect 102192 2592 102198 2604
rect 102962 2592 102968 2604
rect 103020 2592 103026 2644
rect 103238 2592 103244 2644
rect 103296 2632 103302 2644
rect 103977 2635 104035 2641
rect 103977 2632 103989 2635
rect 103296 2604 103989 2632
rect 103296 2592 103302 2604
rect 103977 2601 103989 2604
rect 104023 2601 104035 2635
rect 104158 2632 104164 2644
rect 104119 2604 104164 2632
rect 103977 2595 104035 2601
rect 104158 2592 104164 2604
rect 104216 2592 104222 2644
rect 108482 2632 108488 2644
rect 108443 2604 108488 2632
rect 108482 2592 108488 2604
rect 108540 2592 108546 2644
rect 109494 2632 109500 2644
rect 109455 2604 109500 2632
rect 109494 2592 109500 2604
rect 109552 2592 109558 2644
rect 109586 2592 109592 2644
rect 109644 2632 109650 2644
rect 109865 2635 109923 2641
rect 109865 2632 109877 2635
rect 109644 2604 109877 2632
rect 109644 2592 109650 2604
rect 109865 2601 109877 2604
rect 109911 2632 109923 2635
rect 110322 2632 110328 2644
rect 109911 2604 110328 2632
rect 109911 2601 109923 2604
rect 109865 2595 109923 2601
rect 110322 2592 110328 2604
rect 110380 2592 110386 2644
rect 110414 2592 110420 2644
rect 110472 2632 110478 2644
rect 110693 2635 110751 2641
rect 110693 2632 110705 2635
rect 110472 2604 110705 2632
rect 110472 2592 110478 2604
rect 110693 2601 110705 2604
rect 110739 2601 110751 2635
rect 110693 2595 110751 2601
rect 110782 2592 110788 2644
rect 110840 2632 110846 2644
rect 111337 2635 111395 2641
rect 111337 2632 111349 2635
rect 110840 2604 111349 2632
rect 110840 2592 110846 2604
rect 111337 2601 111349 2604
rect 111383 2601 111395 2635
rect 111518 2632 111524 2644
rect 111479 2604 111524 2632
rect 111337 2595 111395 2601
rect 111518 2592 111524 2604
rect 111576 2592 111582 2644
rect 112714 2632 112720 2644
rect 112675 2604 112720 2632
rect 112714 2592 112720 2604
rect 112772 2592 112778 2644
rect 113450 2592 113456 2644
rect 113508 2632 113514 2644
rect 113729 2635 113787 2641
rect 113729 2632 113741 2635
rect 113508 2604 113741 2632
rect 113508 2592 113514 2604
rect 113729 2601 113741 2604
rect 113775 2601 113787 2635
rect 114554 2632 114560 2644
rect 114515 2604 114560 2632
rect 113729 2595 113787 2601
rect 114554 2592 114560 2604
rect 114612 2592 114618 2644
rect 117222 2632 117228 2644
rect 117183 2604 117228 2632
rect 117222 2592 117228 2604
rect 117280 2592 117286 2644
rect 117682 2592 117688 2644
rect 117740 2632 117746 2644
rect 118421 2635 118479 2641
rect 118421 2632 118433 2635
rect 117740 2604 118433 2632
rect 117740 2592 117746 2604
rect 118421 2601 118433 2604
rect 118467 2601 118479 2635
rect 118421 2595 118479 2601
rect 118510 2592 118516 2644
rect 118568 2632 118574 2644
rect 119798 2632 119804 2644
rect 118568 2604 119804 2632
rect 118568 2592 118574 2604
rect 119798 2592 119804 2604
rect 119856 2592 119862 2644
rect 120810 2632 120816 2644
rect 120771 2604 120816 2632
rect 120810 2592 120816 2604
rect 120868 2592 120874 2644
rect 122374 2632 122380 2644
rect 122335 2604 122380 2632
rect 122374 2592 122380 2604
rect 122432 2592 122438 2644
rect 123754 2632 123760 2644
rect 123715 2604 123760 2632
rect 123754 2592 123760 2604
rect 123812 2592 123818 2644
rect 124214 2592 124220 2644
rect 124272 2632 124278 2644
rect 124953 2635 125011 2641
rect 124953 2632 124965 2635
rect 124272 2604 124965 2632
rect 124272 2592 124278 2604
rect 124953 2601 124965 2604
rect 124999 2601 125011 2635
rect 126054 2632 126060 2644
rect 126015 2604 126060 2632
rect 124953 2595 125011 2601
rect 126054 2592 126060 2604
rect 126112 2592 126118 2644
rect 126882 2632 126888 2644
rect 126843 2604 126888 2632
rect 126882 2592 126888 2604
rect 126940 2592 126946 2644
rect 126974 2592 126980 2644
rect 127032 2632 127038 2644
rect 127529 2635 127587 2641
rect 127529 2632 127541 2635
rect 127032 2604 127541 2632
rect 127032 2592 127038 2604
rect 127529 2601 127541 2604
rect 127575 2601 127587 2635
rect 161566 2632 161572 2644
rect 127529 2595 127587 2601
rect 127636 2604 161572 2632
rect 88334 2564 88340 2576
rect 85868 2536 88340 2564
rect 88334 2524 88340 2536
rect 88392 2524 88398 2576
rect 100021 2567 100079 2573
rect 100021 2533 100033 2567
rect 100067 2564 100079 2567
rect 118050 2564 118056 2576
rect 100067 2536 118056 2564
rect 100067 2533 100079 2536
rect 100021 2527 100079 2533
rect 118050 2524 118056 2536
rect 118108 2524 118114 2576
rect 118160 2536 120672 2564
rect 45235 2468 45784 2496
rect 46017 2499 46075 2505
rect 45235 2465 45247 2468
rect 45189 2459 45247 2465
rect 46017 2465 46029 2499
rect 46063 2496 46075 2499
rect 46290 2496 46296 2508
rect 46063 2468 46296 2496
rect 46063 2465 46075 2468
rect 46017 2459 46075 2465
rect 46290 2456 46296 2468
rect 46348 2456 46354 2508
rect 46753 2499 46811 2505
rect 46753 2496 46765 2499
rect 46400 2468 46765 2496
rect 44453 2431 44511 2437
rect 44453 2428 44465 2431
rect 44232 2400 44465 2428
rect 44232 2388 44238 2400
rect 44453 2397 44465 2400
rect 44499 2397 44511 2431
rect 44453 2391 44511 2397
rect 44729 2431 44787 2437
rect 44729 2397 44741 2431
rect 44775 2397 44787 2431
rect 44729 2391 44787 2397
rect 44913 2431 44971 2437
rect 44913 2397 44925 2431
rect 44959 2428 44971 2431
rect 45738 2428 45744 2440
rect 44959 2400 45744 2428
rect 44959 2397 44971 2400
rect 44913 2391 44971 2397
rect 45738 2388 45744 2400
rect 45796 2388 45802 2440
rect 45925 2431 45983 2437
rect 45925 2397 45937 2431
rect 45971 2428 45983 2431
rect 46198 2428 46204 2440
rect 45971 2400 46204 2428
rect 45971 2397 45983 2400
rect 45925 2391 45983 2397
rect 46198 2388 46204 2400
rect 46256 2388 46262 2440
rect 46400 2437 46428 2468
rect 46753 2465 46765 2468
rect 46799 2496 46811 2499
rect 48406 2496 48412 2508
rect 46799 2468 48412 2496
rect 46799 2465 46811 2468
rect 46753 2459 46811 2465
rect 48406 2456 48412 2468
rect 48464 2456 48470 2508
rect 50614 2496 50620 2508
rect 48516 2468 50620 2496
rect 46385 2431 46443 2437
rect 46385 2397 46397 2431
rect 46431 2397 46443 2431
rect 46385 2391 46443 2397
rect 46474 2388 46480 2440
rect 46532 2428 46538 2440
rect 48516 2428 48544 2468
rect 50614 2456 50620 2468
rect 50672 2456 50678 2508
rect 50706 2456 50712 2508
rect 50764 2496 50770 2508
rect 52638 2496 52644 2508
rect 50764 2468 51120 2496
rect 50764 2456 50770 2468
rect 46532 2400 48544 2428
rect 46532 2388 46538 2400
rect 48590 2388 48596 2440
rect 48648 2428 48654 2440
rect 49881 2431 49939 2437
rect 49881 2428 49893 2431
rect 48648 2400 49893 2428
rect 48648 2388 48654 2400
rect 49881 2397 49893 2400
rect 49927 2397 49939 2431
rect 50246 2428 50252 2440
rect 50207 2400 50252 2428
rect 49881 2391 49939 2397
rect 50246 2388 50252 2400
rect 50304 2428 50310 2440
rect 50893 2431 50951 2437
rect 50893 2428 50905 2431
rect 50304 2400 50905 2428
rect 50304 2388 50310 2400
rect 50893 2397 50905 2400
rect 50939 2397 50951 2431
rect 50893 2391 50951 2397
rect 44818 2360 44824 2372
rect 44039 2332 44824 2360
rect 44039 2329 44051 2332
rect 43993 2323 44051 2329
rect 44818 2320 44824 2332
rect 44876 2320 44882 2372
rect 45370 2320 45376 2372
rect 45428 2360 45434 2372
rect 46842 2360 46848 2372
rect 45428 2332 46848 2360
rect 45428 2320 45434 2332
rect 46842 2320 46848 2332
rect 46900 2320 46906 2372
rect 47118 2320 47124 2372
rect 47176 2360 47182 2372
rect 47578 2360 47584 2372
rect 47176 2332 47584 2360
rect 47176 2320 47182 2332
rect 47578 2320 47584 2332
rect 47636 2320 47642 2372
rect 51092 2360 51120 2468
rect 51184 2468 52644 2496
rect 51184 2440 51212 2468
rect 52638 2456 52644 2468
rect 52696 2456 52702 2508
rect 54018 2496 54024 2508
rect 53979 2468 54024 2496
rect 54018 2456 54024 2468
rect 54076 2456 54082 2508
rect 54202 2456 54208 2508
rect 54260 2496 54266 2508
rect 54260 2468 54708 2496
rect 54260 2456 54266 2468
rect 51166 2388 51172 2440
rect 51224 2388 51230 2440
rect 51350 2388 51356 2440
rect 51408 2388 51414 2440
rect 51534 2388 51540 2440
rect 51592 2428 51598 2440
rect 52086 2428 52092 2440
rect 51592 2400 52092 2428
rect 51592 2388 51598 2400
rect 52086 2388 52092 2400
rect 52144 2388 52150 2440
rect 52733 2431 52791 2437
rect 52733 2397 52745 2431
rect 52779 2428 52791 2431
rect 53282 2428 53288 2440
rect 52779 2400 53288 2428
rect 52779 2397 52791 2400
rect 52733 2391 52791 2397
rect 53282 2388 53288 2400
rect 53340 2388 53346 2440
rect 54570 2428 54576 2440
rect 54531 2400 54576 2428
rect 54570 2388 54576 2400
rect 54628 2388 54634 2440
rect 54680 2428 54708 2468
rect 55674 2456 55680 2508
rect 55732 2496 55738 2508
rect 57238 2496 57244 2508
rect 55732 2468 57244 2496
rect 55732 2456 55738 2468
rect 57238 2456 57244 2468
rect 57296 2456 57302 2508
rect 57330 2456 57336 2508
rect 57388 2496 57394 2508
rect 59722 2496 59728 2508
rect 57388 2468 59728 2496
rect 57388 2456 57394 2468
rect 59722 2456 59728 2468
rect 59780 2456 59786 2508
rect 59814 2456 59820 2508
rect 59872 2496 59878 2508
rect 60550 2496 60556 2508
rect 59872 2468 60556 2496
rect 59872 2456 59878 2468
rect 60550 2456 60556 2468
rect 60608 2456 60614 2508
rect 61010 2456 61016 2508
rect 61068 2496 61074 2508
rect 61378 2496 61384 2508
rect 61068 2468 61384 2496
rect 61068 2456 61074 2468
rect 61378 2456 61384 2468
rect 61436 2456 61442 2508
rect 61746 2456 61752 2508
rect 61804 2496 61810 2508
rect 63218 2496 63224 2508
rect 61804 2468 63224 2496
rect 61804 2456 61810 2468
rect 63218 2456 63224 2468
rect 63276 2456 63282 2508
rect 63310 2456 63316 2508
rect 63368 2496 63374 2508
rect 65061 2499 65119 2505
rect 65061 2496 65073 2499
rect 63368 2468 65073 2496
rect 63368 2456 63374 2468
rect 65061 2465 65073 2468
rect 65107 2465 65119 2499
rect 68005 2499 68063 2505
rect 68005 2496 68017 2499
rect 65061 2459 65119 2465
rect 67468 2468 68017 2496
rect 56042 2428 56048 2440
rect 54680 2400 56048 2428
rect 56042 2388 56048 2400
rect 56100 2388 56106 2440
rect 56229 2431 56287 2437
rect 56229 2397 56241 2431
rect 56275 2428 56287 2431
rect 56502 2428 56508 2440
rect 56275 2400 56508 2428
rect 56275 2397 56287 2400
rect 56229 2391 56287 2397
rect 56502 2388 56508 2400
rect 56560 2388 56566 2440
rect 56962 2388 56968 2440
rect 57020 2428 57026 2440
rect 57149 2431 57207 2437
rect 57149 2428 57161 2431
rect 57020 2400 57161 2428
rect 57020 2388 57026 2400
rect 57149 2397 57161 2400
rect 57195 2397 57207 2431
rect 57149 2391 57207 2397
rect 57606 2388 57612 2440
rect 57664 2428 57670 2440
rect 57701 2431 57759 2437
rect 57701 2428 57713 2431
rect 57664 2400 57713 2428
rect 57664 2388 57670 2400
rect 57701 2397 57713 2400
rect 57747 2428 57759 2431
rect 58161 2431 58219 2437
rect 58161 2428 58173 2431
rect 57747 2400 58173 2428
rect 57747 2397 57759 2400
rect 57701 2391 57759 2397
rect 58161 2397 58173 2400
rect 58207 2397 58219 2431
rect 58161 2391 58219 2397
rect 59354 2388 59360 2440
rect 59412 2428 59418 2440
rect 60093 2431 60151 2437
rect 60093 2428 60105 2431
rect 59412 2400 60105 2428
rect 59412 2388 59418 2400
rect 60093 2397 60105 2400
rect 60139 2428 60151 2431
rect 60461 2431 60519 2437
rect 60461 2428 60473 2431
rect 60139 2400 60473 2428
rect 60139 2397 60151 2400
rect 60093 2391 60151 2397
rect 60461 2397 60473 2400
rect 60507 2397 60519 2431
rect 60461 2391 60519 2397
rect 61102 2388 61108 2440
rect 61160 2428 61166 2440
rect 61160 2400 61205 2428
rect 61160 2388 61166 2400
rect 61654 2388 61660 2440
rect 61712 2428 61718 2440
rect 62577 2431 62635 2437
rect 62577 2428 62589 2431
rect 61712 2400 62589 2428
rect 61712 2388 61718 2400
rect 62577 2397 62589 2400
rect 62623 2428 62635 2431
rect 63037 2431 63095 2437
rect 63037 2428 63049 2431
rect 62623 2400 63049 2428
rect 62623 2397 62635 2400
rect 62577 2391 62635 2397
rect 63037 2397 63049 2400
rect 63083 2397 63095 2431
rect 63037 2391 63095 2397
rect 63494 2388 63500 2440
rect 63552 2428 63558 2440
rect 67468 2437 67496 2468
rect 68005 2465 68017 2468
rect 68051 2496 68063 2499
rect 69750 2496 69756 2508
rect 68051 2468 69756 2496
rect 68051 2465 68063 2468
rect 68005 2459 68063 2465
rect 69750 2456 69756 2468
rect 69808 2456 69814 2508
rect 72878 2456 72884 2508
rect 72936 2496 72942 2508
rect 72936 2468 76880 2496
rect 72936 2456 72942 2468
rect 63589 2431 63647 2437
rect 63589 2428 63601 2431
rect 63552 2400 63601 2428
rect 63552 2388 63558 2400
rect 63589 2397 63601 2400
rect 63635 2397 63647 2431
rect 66441 2431 66499 2437
rect 63589 2391 63647 2397
rect 63696 2400 63908 2428
rect 51258 2360 51264 2372
rect 47780 2332 49556 2360
rect 51092 2332 51264 2360
rect 35676 2264 42564 2292
rect 35676 2252 35682 2264
rect 42610 2252 42616 2304
rect 42668 2292 42674 2304
rect 47780 2292 47808 2332
rect 42668 2264 47808 2292
rect 49528 2292 49556 2332
rect 51258 2320 51264 2332
rect 51316 2320 51322 2372
rect 51368 2360 51396 2388
rect 59449 2363 59507 2369
rect 59449 2360 59461 2363
rect 51368 2332 59461 2360
rect 59449 2329 59461 2332
rect 59495 2329 59507 2363
rect 59449 2323 59507 2329
rect 59998 2320 60004 2372
rect 60056 2360 60062 2372
rect 63696 2360 63724 2400
rect 60056 2332 63724 2360
rect 63880 2360 63908 2400
rect 66441 2397 66453 2431
rect 66487 2428 66499 2431
rect 66717 2431 66775 2437
rect 66717 2428 66729 2431
rect 66487 2400 66729 2428
rect 66487 2397 66499 2400
rect 66441 2391 66499 2397
rect 66717 2397 66729 2400
rect 66763 2397 66775 2431
rect 66717 2391 66775 2397
rect 67453 2431 67511 2437
rect 67453 2397 67465 2431
rect 67499 2397 67511 2431
rect 67453 2391 67511 2397
rect 69201 2431 69259 2437
rect 69201 2397 69213 2431
rect 69247 2428 69259 2431
rect 69477 2431 69535 2437
rect 69477 2428 69489 2431
rect 69247 2400 69489 2428
rect 69247 2397 69259 2400
rect 69201 2391 69259 2397
rect 69477 2397 69489 2400
rect 69523 2397 69535 2431
rect 69477 2391 69535 2397
rect 70673 2431 70731 2437
rect 70673 2397 70685 2431
rect 70719 2397 70731 2431
rect 70673 2391 70731 2397
rect 71777 2431 71835 2437
rect 71777 2397 71789 2431
rect 71823 2428 71835 2431
rect 73433 2431 73491 2437
rect 71823 2400 72372 2428
rect 71823 2397 71835 2400
rect 71777 2391 71835 2397
rect 70688 2360 70716 2391
rect 71225 2363 71283 2369
rect 71225 2360 71237 2363
rect 63880 2332 70624 2360
rect 70688 2332 71237 2360
rect 60056 2320 60062 2332
rect 51350 2292 51356 2304
rect 49528 2264 51356 2292
rect 42668 2252 42674 2264
rect 51350 2252 51356 2264
rect 51408 2252 51414 2304
rect 51442 2252 51448 2304
rect 51500 2292 51506 2304
rect 51810 2292 51816 2304
rect 51500 2264 51816 2292
rect 51500 2252 51506 2264
rect 51810 2252 51816 2264
rect 51868 2252 51874 2304
rect 51902 2252 51908 2304
rect 51960 2292 51966 2304
rect 55861 2295 55919 2301
rect 55861 2292 55873 2295
rect 51960 2264 55873 2292
rect 51960 2252 51966 2264
rect 55861 2261 55873 2264
rect 55907 2261 55919 2295
rect 55861 2255 55919 2261
rect 56042 2252 56048 2304
rect 56100 2292 56106 2304
rect 60369 2295 60427 2301
rect 60369 2292 60381 2295
rect 56100 2264 60381 2292
rect 56100 2252 56106 2264
rect 60369 2261 60381 2264
rect 60415 2261 60427 2295
rect 60369 2255 60427 2261
rect 60550 2252 60556 2304
rect 60608 2292 60614 2304
rect 62206 2292 62212 2304
rect 60608 2264 62212 2292
rect 60608 2252 60614 2264
rect 62206 2252 62212 2264
rect 62264 2252 62270 2304
rect 62301 2295 62359 2301
rect 62301 2261 62313 2295
rect 62347 2292 62359 2295
rect 62390 2292 62396 2304
rect 62347 2264 62396 2292
rect 62347 2261 62359 2264
rect 62301 2255 62359 2261
rect 62390 2252 62396 2264
rect 62448 2252 62454 2304
rect 63494 2252 63500 2304
rect 63552 2292 63558 2304
rect 64141 2295 64199 2301
rect 64141 2292 64153 2295
rect 63552 2264 64153 2292
rect 63552 2252 63558 2264
rect 64141 2261 64153 2264
rect 64187 2292 64199 2295
rect 64966 2292 64972 2304
rect 64187 2264 64972 2292
rect 64187 2261 64199 2264
rect 64141 2255 64199 2261
rect 64966 2252 64972 2264
rect 65024 2252 65030 2304
rect 66717 2295 66775 2301
rect 66717 2261 66729 2295
rect 66763 2292 66775 2295
rect 66993 2295 67051 2301
rect 66993 2292 67005 2295
rect 66763 2264 67005 2292
rect 66763 2261 66775 2264
rect 66717 2255 66775 2261
rect 66993 2261 67005 2264
rect 67039 2292 67051 2295
rect 67542 2292 67548 2304
rect 67039 2264 67548 2292
rect 67039 2261 67051 2264
rect 66993 2255 67051 2261
rect 67542 2252 67548 2264
rect 67600 2252 67606 2304
rect 68002 2252 68008 2304
rect 68060 2292 68066 2304
rect 69293 2295 69351 2301
rect 69293 2292 69305 2295
rect 68060 2264 69305 2292
rect 68060 2252 68066 2264
rect 69293 2261 69305 2264
rect 69339 2261 69351 2295
rect 69293 2255 69351 2261
rect 69477 2295 69535 2301
rect 69477 2261 69489 2295
rect 69523 2292 69535 2295
rect 69753 2295 69811 2301
rect 69753 2292 69765 2295
rect 69523 2264 69765 2292
rect 69523 2261 69535 2264
rect 69477 2255 69535 2261
rect 69753 2261 69765 2264
rect 69799 2292 69811 2295
rect 70394 2292 70400 2304
rect 69799 2264 70400 2292
rect 69799 2261 69811 2264
rect 69753 2255 69811 2261
rect 70394 2252 70400 2264
rect 70452 2252 70458 2304
rect 70596 2292 70624 2332
rect 71225 2329 71237 2332
rect 71271 2360 71283 2363
rect 71314 2360 71320 2372
rect 71271 2332 71320 2360
rect 71271 2329 71283 2332
rect 71225 2323 71283 2329
rect 71314 2320 71320 2332
rect 71372 2320 71378 2372
rect 72344 2301 72372 2400
rect 73433 2397 73445 2431
rect 73479 2428 73491 2431
rect 74537 2431 74595 2437
rect 73479 2400 74028 2428
rect 73479 2397 73491 2400
rect 73433 2391 73491 2397
rect 70765 2295 70823 2301
rect 70765 2292 70777 2295
rect 70596 2264 70777 2292
rect 70765 2261 70777 2264
rect 70811 2261 70823 2295
rect 70765 2255 70823 2261
rect 72329 2295 72387 2301
rect 72329 2261 72341 2295
rect 72375 2292 72387 2295
rect 73430 2292 73436 2304
rect 72375 2264 73436 2292
rect 72375 2261 72387 2264
rect 72329 2255 72387 2261
rect 73430 2252 73436 2264
rect 73488 2252 73494 2304
rect 74000 2301 74028 2400
rect 74537 2397 74549 2431
rect 74583 2397 74595 2431
rect 76558 2428 76564 2440
rect 76519 2400 76564 2428
rect 74537 2391 74595 2397
rect 74552 2360 74580 2391
rect 76558 2388 76564 2400
rect 76616 2388 76622 2440
rect 76650 2388 76656 2440
rect 76708 2428 76714 2440
rect 76852 2437 76880 2468
rect 80790 2456 80796 2508
rect 80848 2496 80854 2508
rect 85393 2499 85451 2505
rect 80848 2468 81940 2496
rect 80848 2456 80854 2468
rect 76837 2431 76895 2437
rect 76708 2400 76753 2428
rect 76708 2388 76714 2400
rect 76837 2397 76849 2431
rect 76883 2428 76895 2431
rect 77297 2431 77355 2437
rect 77297 2428 77309 2431
rect 76883 2400 77309 2428
rect 76883 2397 76895 2400
rect 76837 2391 76895 2397
rect 77297 2397 77309 2400
rect 77343 2397 77355 2431
rect 79318 2428 79324 2440
rect 79279 2400 79324 2428
rect 77297 2391 77355 2397
rect 79318 2388 79324 2400
rect 79376 2388 79382 2440
rect 80422 2388 80428 2440
rect 80480 2428 80486 2440
rect 81912 2437 81940 2468
rect 85393 2465 85405 2499
rect 85439 2496 85451 2499
rect 89809 2499 89867 2505
rect 89809 2496 89821 2499
rect 85439 2468 89821 2496
rect 85439 2465 85451 2468
rect 85393 2459 85451 2465
rect 89809 2465 89821 2468
rect 89855 2496 89867 2499
rect 90361 2499 90419 2505
rect 90361 2496 90373 2499
rect 89855 2468 90373 2496
rect 89855 2465 89867 2468
rect 89809 2459 89867 2465
rect 90361 2465 90373 2468
rect 90407 2465 90419 2499
rect 91370 2496 91376 2508
rect 91331 2468 91376 2496
rect 90361 2459 90419 2465
rect 91370 2456 91376 2468
rect 91428 2456 91434 2508
rect 102870 2456 102876 2508
rect 102928 2496 102934 2508
rect 103333 2499 103391 2505
rect 103333 2496 103345 2499
rect 102928 2468 103345 2496
rect 102928 2456 102934 2468
rect 103333 2465 103345 2468
rect 103379 2465 103391 2499
rect 103882 2496 103888 2508
rect 103333 2459 103391 2465
rect 103808 2468 103888 2496
rect 80701 2431 80759 2437
rect 80701 2428 80713 2431
rect 80480 2400 80713 2428
rect 80480 2388 80486 2400
rect 80701 2397 80713 2400
rect 80747 2428 80759 2431
rect 81161 2431 81219 2437
rect 81161 2428 81173 2431
rect 80747 2400 81173 2428
rect 80747 2397 80759 2400
rect 80701 2391 80759 2397
rect 81161 2397 81173 2400
rect 81207 2397 81219 2431
rect 81161 2391 81219 2397
rect 81897 2431 81955 2437
rect 81897 2397 81909 2431
rect 81943 2428 81955 2431
rect 82357 2431 82415 2437
rect 82357 2428 82369 2431
rect 81943 2400 82369 2428
rect 81943 2397 81955 2400
rect 81897 2391 81955 2397
rect 82357 2397 82369 2400
rect 82403 2397 82415 2431
rect 82357 2391 82415 2397
rect 83369 2431 83427 2437
rect 83369 2397 83381 2431
rect 83415 2428 83427 2431
rect 83645 2431 83703 2437
rect 83645 2428 83657 2431
rect 83415 2400 83657 2428
rect 83415 2397 83427 2400
rect 83369 2391 83427 2397
rect 83645 2397 83657 2400
rect 83691 2397 83703 2431
rect 83645 2391 83703 2397
rect 86405 2431 86463 2437
rect 86405 2397 86417 2431
rect 86451 2428 86463 2431
rect 86954 2428 86960 2440
rect 86451 2400 86960 2428
rect 86451 2397 86463 2400
rect 86405 2391 86463 2397
rect 86954 2388 86960 2400
rect 87012 2388 87018 2440
rect 87509 2431 87567 2437
rect 87509 2397 87521 2431
rect 87555 2397 87567 2431
rect 87509 2391 87567 2397
rect 88521 2431 88579 2437
rect 88521 2397 88533 2431
rect 88567 2428 88579 2431
rect 91925 2431 91983 2437
rect 88567 2400 89116 2428
rect 88567 2397 88579 2400
rect 88521 2391 88579 2397
rect 74813 2363 74871 2369
rect 74813 2360 74825 2363
rect 74552 2332 74825 2360
rect 74813 2329 74825 2332
rect 74859 2329 74871 2363
rect 74813 2323 74871 2329
rect 75730 2320 75736 2372
rect 75788 2360 75794 2372
rect 80882 2360 80888 2372
rect 75788 2332 80888 2360
rect 75788 2320 75794 2332
rect 80882 2320 80888 2332
rect 80940 2320 80946 2372
rect 86497 2363 86555 2369
rect 86497 2360 86509 2363
rect 81084 2332 86509 2360
rect 73985 2295 74043 2301
rect 73985 2261 73997 2295
rect 74031 2292 74043 2295
rect 74626 2292 74632 2304
rect 74031 2264 74632 2292
rect 74031 2261 74043 2264
rect 73985 2255 74043 2261
rect 74626 2252 74632 2264
rect 74684 2252 74690 2304
rect 74994 2252 75000 2304
rect 75052 2292 75058 2304
rect 81084 2292 81112 2332
rect 86497 2329 86509 2332
rect 86543 2329 86555 2363
rect 87524 2360 87552 2391
rect 88061 2363 88119 2369
rect 88061 2360 88073 2363
rect 87524 2332 88073 2360
rect 86497 2323 86555 2329
rect 88061 2329 88073 2332
rect 88107 2360 88119 2363
rect 88794 2360 88800 2372
rect 88107 2332 88800 2360
rect 88107 2329 88119 2332
rect 88061 2323 88119 2329
rect 88794 2320 88800 2332
rect 88852 2320 88858 2372
rect 75052 2264 81112 2292
rect 83645 2295 83703 2301
rect 75052 2252 75058 2264
rect 83645 2261 83657 2295
rect 83691 2292 83703 2295
rect 83921 2295 83979 2301
rect 83921 2292 83933 2295
rect 83691 2264 83933 2292
rect 83691 2261 83703 2264
rect 83645 2255 83703 2261
rect 83921 2261 83933 2264
rect 83967 2292 83979 2295
rect 84470 2292 84476 2304
rect 83967 2264 84476 2292
rect 83967 2261 83979 2264
rect 83921 2255 83979 2261
rect 84470 2252 84476 2264
rect 84528 2252 84534 2304
rect 88610 2292 88616 2304
rect 88571 2264 88616 2292
rect 88610 2252 88616 2264
rect 88668 2252 88674 2304
rect 89088 2301 89116 2400
rect 91925 2397 91937 2431
rect 91971 2428 91983 2431
rect 92014 2428 92020 2440
rect 91971 2400 92020 2428
rect 91971 2397 91983 2400
rect 91925 2391 91983 2397
rect 92014 2388 92020 2400
rect 92072 2428 92078 2440
rect 103808 2437 103836 2468
rect 103882 2456 103888 2468
rect 103940 2496 103946 2508
rect 103940 2468 108528 2496
rect 103940 2456 103946 2468
rect 92201 2431 92259 2437
rect 92201 2428 92213 2431
rect 92072 2400 92213 2428
rect 92072 2388 92078 2400
rect 92201 2397 92213 2400
rect 92247 2397 92259 2431
rect 92201 2391 92259 2397
rect 102321 2431 102379 2437
rect 102321 2397 102333 2431
rect 102367 2397 102379 2431
rect 102321 2391 102379 2397
rect 103793 2431 103851 2437
rect 103793 2397 103805 2431
rect 103839 2397 103851 2431
rect 108114 2428 108120 2440
rect 103793 2391 103851 2397
rect 104084 2400 108120 2428
rect 102336 2360 102364 2391
rect 103238 2360 103244 2372
rect 102336 2332 103244 2360
rect 103238 2320 103244 2332
rect 103296 2320 103302 2372
rect 104084 2360 104112 2400
rect 108114 2388 108120 2400
rect 108172 2388 108178 2440
rect 108393 2431 108451 2437
rect 108393 2397 108405 2431
rect 108439 2397 108451 2431
rect 108393 2391 108451 2397
rect 107838 2360 107844 2372
rect 103340 2332 104112 2360
rect 104176 2332 107844 2360
rect 89073 2295 89131 2301
rect 89073 2261 89085 2295
rect 89119 2292 89131 2295
rect 89898 2292 89904 2304
rect 89119 2264 89904 2292
rect 89119 2261 89131 2264
rect 89073 2255 89131 2261
rect 89898 2252 89904 2264
rect 89956 2252 89962 2304
rect 100754 2252 100760 2304
rect 100812 2292 100818 2304
rect 103340 2292 103368 2332
rect 100812 2264 103368 2292
rect 104069 2295 104127 2301
rect 100812 2252 100818 2264
rect 104069 2261 104081 2295
rect 104115 2292 104127 2295
rect 104176 2292 104204 2332
rect 107838 2320 107844 2332
rect 107896 2320 107902 2372
rect 104986 2292 104992 2304
rect 104115 2264 104204 2292
rect 104947 2264 104992 2292
rect 104115 2261 104127 2264
rect 104069 2255 104127 2261
rect 104986 2252 104992 2264
rect 105044 2252 105050 2304
rect 107746 2292 107752 2304
rect 107659 2264 107752 2292
rect 107746 2252 107752 2264
rect 107804 2292 107810 2304
rect 107930 2292 107936 2304
rect 107804 2264 107936 2292
rect 107804 2252 107810 2264
rect 107930 2252 107936 2264
rect 107988 2252 107994 2304
rect 108408 2292 108436 2391
rect 108500 2360 108528 2468
rect 108574 2456 108580 2508
rect 108632 2496 108638 2508
rect 118160 2496 118188 2536
rect 108632 2468 118188 2496
rect 108632 2456 108638 2468
rect 118234 2456 118240 2508
rect 118292 2496 118298 2508
rect 120644 2496 120672 2536
rect 120718 2524 120724 2576
rect 120776 2564 120782 2576
rect 127636 2564 127664 2604
rect 161566 2592 161572 2604
rect 161624 2592 161630 2644
rect 161753 2635 161811 2641
rect 161753 2601 161765 2635
rect 161799 2632 161811 2635
rect 161934 2632 161940 2644
rect 161799 2604 161940 2632
rect 161799 2601 161811 2604
rect 161753 2595 161811 2601
rect 161934 2592 161940 2604
rect 161992 2592 161998 2644
rect 162765 2635 162823 2641
rect 162765 2601 162777 2635
rect 162811 2632 162823 2635
rect 164326 2632 164332 2644
rect 162811 2604 164332 2632
rect 162811 2601 162823 2604
rect 162765 2595 162823 2601
rect 164326 2592 164332 2604
rect 164384 2592 164390 2644
rect 120776 2536 127664 2564
rect 127713 2567 127771 2573
rect 120776 2524 120782 2536
rect 127713 2533 127725 2567
rect 127759 2564 127771 2567
rect 151814 2564 151820 2576
rect 127759 2536 151820 2564
rect 127759 2533 127771 2536
rect 127713 2527 127771 2533
rect 151814 2524 151820 2536
rect 151872 2524 151878 2576
rect 155862 2564 155868 2576
rect 155823 2536 155868 2564
rect 155862 2524 155868 2536
rect 155920 2524 155926 2576
rect 157334 2564 157340 2576
rect 157295 2536 157340 2564
rect 157334 2524 157340 2536
rect 157392 2524 157398 2576
rect 158441 2567 158499 2573
rect 158441 2533 158453 2567
rect 158487 2564 158499 2567
rect 159542 2564 159548 2576
rect 158487 2536 159548 2564
rect 158487 2533 158499 2536
rect 158441 2527 158499 2533
rect 159542 2524 159548 2536
rect 159600 2524 159606 2576
rect 160186 2564 160192 2576
rect 160147 2536 160192 2564
rect 160186 2524 160192 2536
rect 160244 2524 160250 2576
rect 127805 2499 127863 2505
rect 127805 2496 127817 2499
rect 118292 2468 120396 2496
rect 120644 2468 127817 2496
rect 118292 2456 118298 2468
rect 109405 2431 109463 2437
rect 109405 2397 109417 2431
rect 109451 2428 109463 2431
rect 109681 2431 109739 2437
rect 109681 2428 109693 2431
rect 109451 2400 109693 2428
rect 109451 2397 109463 2400
rect 109405 2391 109463 2397
rect 109681 2397 109693 2400
rect 109727 2397 109739 2431
rect 109681 2391 109739 2397
rect 110601 2431 110659 2437
rect 110601 2397 110613 2431
rect 110647 2428 110659 2431
rect 111153 2431 111211 2437
rect 111153 2428 111165 2431
rect 110647 2400 111165 2428
rect 110647 2397 110659 2400
rect 110601 2391 110659 2397
rect 111153 2397 111165 2400
rect 111199 2428 111211 2431
rect 111518 2428 111524 2440
rect 111199 2400 111524 2428
rect 111199 2397 111211 2400
rect 111153 2391 111211 2397
rect 111518 2388 111524 2400
rect 111576 2388 111582 2440
rect 111613 2431 111671 2437
rect 111613 2397 111625 2431
rect 111659 2428 111671 2431
rect 111889 2431 111947 2437
rect 111889 2428 111901 2431
rect 111659 2400 111901 2428
rect 111659 2397 111671 2400
rect 111613 2391 111671 2397
rect 111889 2397 111901 2400
rect 111935 2397 111947 2431
rect 111889 2391 111947 2397
rect 112625 2431 112683 2437
rect 112625 2397 112637 2431
rect 112671 2428 112683 2431
rect 112901 2431 112959 2437
rect 112901 2428 112913 2431
rect 112671 2400 112913 2428
rect 112671 2397 112683 2400
rect 112625 2391 112683 2397
rect 112901 2397 112913 2400
rect 112947 2397 112959 2431
rect 112901 2391 112959 2397
rect 113637 2431 113695 2437
rect 113637 2397 113649 2431
rect 113683 2428 113695 2431
rect 114278 2428 114284 2440
rect 113683 2400 114284 2428
rect 113683 2397 113695 2400
rect 113637 2391 113695 2397
rect 114278 2388 114284 2400
rect 114336 2388 114342 2440
rect 116213 2431 116271 2437
rect 116213 2397 116225 2431
rect 116259 2428 116271 2431
rect 116762 2428 116768 2440
rect 116259 2400 116768 2428
rect 116259 2397 116271 2400
rect 116213 2391 116271 2397
rect 116762 2388 116768 2400
rect 116820 2388 116826 2440
rect 117317 2431 117375 2437
rect 117317 2397 117329 2431
rect 117363 2428 117375 2431
rect 117593 2431 117651 2437
rect 117593 2428 117605 2431
rect 117363 2400 117605 2428
rect 117363 2397 117375 2400
rect 117317 2391 117375 2397
rect 117593 2397 117605 2400
rect 117639 2397 117651 2431
rect 117593 2391 117651 2397
rect 118329 2431 118387 2437
rect 118329 2397 118341 2431
rect 118375 2428 118387 2431
rect 118881 2431 118939 2437
rect 118881 2428 118893 2431
rect 118375 2400 118893 2428
rect 118375 2397 118387 2400
rect 118329 2391 118387 2397
rect 118881 2397 118893 2400
rect 118927 2428 118939 2431
rect 118927 2400 119108 2428
rect 118927 2397 118939 2400
rect 118881 2391 118939 2397
rect 118970 2360 118976 2372
rect 108500 2332 118976 2360
rect 118970 2320 118976 2332
rect 119028 2320 119034 2372
rect 119080 2360 119108 2400
rect 120258 2360 120264 2372
rect 119080 2332 120264 2360
rect 120258 2320 120264 2332
rect 120316 2320 120322 2372
rect 120368 2360 120396 2468
rect 127805 2465 127817 2468
rect 127851 2465 127863 2499
rect 139673 2499 139731 2505
rect 139673 2496 139685 2499
rect 127805 2459 127863 2465
rect 128096 2468 139685 2496
rect 120721 2431 120779 2437
rect 120721 2397 120733 2431
rect 120767 2428 120779 2431
rect 120902 2428 120908 2440
rect 120767 2400 120908 2428
rect 120767 2397 120779 2400
rect 120721 2391 120779 2397
rect 120902 2388 120908 2400
rect 120960 2388 120966 2440
rect 123665 2431 123723 2437
rect 123665 2397 123677 2431
rect 123711 2428 123723 2431
rect 124214 2428 124220 2440
rect 123711 2400 124220 2428
rect 123711 2397 123723 2400
rect 123665 2391 123723 2397
rect 124214 2388 124220 2400
rect 124272 2388 124278 2440
rect 124861 2431 124919 2437
rect 124861 2397 124873 2431
rect 124907 2428 124919 2431
rect 125594 2428 125600 2440
rect 124907 2400 125600 2428
rect 124907 2397 124919 2400
rect 124861 2391 124919 2397
rect 125594 2388 125600 2400
rect 125652 2388 125658 2440
rect 125965 2431 126023 2437
rect 125965 2397 125977 2431
rect 126011 2428 126023 2431
rect 126241 2431 126299 2437
rect 126241 2428 126253 2431
rect 126011 2400 126253 2428
rect 126011 2397 126023 2400
rect 125965 2391 126023 2397
rect 126241 2397 126253 2400
rect 126287 2397 126299 2431
rect 126241 2391 126299 2397
rect 127437 2431 127495 2437
rect 127437 2397 127449 2431
rect 127483 2428 127495 2431
rect 127526 2428 127532 2440
rect 127483 2400 127532 2428
rect 127483 2397 127495 2400
rect 127437 2391 127495 2397
rect 127526 2388 127532 2400
rect 127584 2428 127590 2440
rect 127897 2431 127955 2437
rect 127897 2428 127909 2431
rect 127584 2400 127909 2428
rect 127584 2388 127590 2400
rect 127897 2397 127909 2400
rect 127943 2397 127955 2431
rect 127897 2391 127955 2397
rect 127713 2363 127771 2369
rect 127713 2360 127725 2363
rect 120368 2332 127725 2360
rect 127713 2329 127725 2332
rect 127759 2329 127771 2363
rect 127713 2323 127771 2329
rect 108945 2295 109003 2301
rect 108945 2292 108957 2295
rect 108408 2264 108957 2292
rect 108945 2261 108957 2264
rect 108991 2292 109003 2295
rect 109586 2292 109592 2304
rect 108991 2264 109592 2292
rect 108991 2261 109003 2264
rect 108945 2255 109003 2261
rect 109586 2252 109592 2264
rect 109644 2252 109650 2304
rect 109681 2295 109739 2301
rect 109681 2261 109693 2295
rect 109727 2292 109739 2295
rect 110325 2295 110383 2301
rect 110325 2292 110337 2295
rect 109727 2264 110337 2292
rect 109727 2261 109739 2264
rect 109681 2255 109739 2261
rect 110325 2261 110337 2264
rect 110371 2292 110383 2295
rect 111242 2292 111248 2304
rect 110371 2264 111248 2292
rect 110371 2261 110383 2264
rect 110325 2255 110383 2261
rect 111242 2252 111248 2264
rect 111300 2252 111306 2304
rect 111337 2295 111395 2301
rect 111337 2261 111349 2295
rect 111383 2292 111395 2295
rect 111705 2295 111763 2301
rect 111705 2292 111717 2295
rect 111383 2264 111717 2292
rect 111383 2261 111395 2264
rect 111337 2255 111395 2261
rect 111705 2261 111717 2264
rect 111751 2261 111763 2295
rect 111705 2255 111763 2261
rect 111889 2295 111947 2301
rect 111889 2261 111901 2295
rect 111935 2292 111947 2295
rect 112165 2295 112223 2301
rect 112165 2292 112177 2295
rect 111935 2264 112177 2292
rect 111935 2261 111947 2264
rect 111889 2255 111947 2261
rect 112165 2261 112177 2264
rect 112211 2292 112223 2295
rect 112254 2292 112260 2304
rect 112211 2264 112260 2292
rect 112211 2261 112223 2264
rect 112165 2255 112223 2261
rect 112254 2252 112260 2264
rect 112312 2252 112318 2304
rect 112901 2295 112959 2301
rect 112901 2261 112913 2295
rect 112947 2292 112959 2295
rect 113177 2295 113235 2301
rect 113177 2292 113189 2295
rect 112947 2264 113189 2292
rect 112947 2261 112959 2264
rect 112901 2255 112959 2261
rect 113177 2261 113189 2264
rect 113223 2292 113235 2295
rect 113910 2292 113916 2304
rect 113223 2264 113916 2292
rect 113223 2261 113235 2264
rect 113177 2255 113235 2261
rect 113910 2252 113916 2264
rect 113968 2252 113974 2304
rect 114189 2295 114247 2301
rect 114189 2261 114201 2295
rect 114235 2292 114247 2295
rect 114278 2292 114284 2304
rect 114235 2264 114284 2292
rect 114235 2261 114247 2264
rect 114189 2255 114247 2261
rect 114278 2252 114284 2264
rect 114336 2252 114342 2304
rect 114462 2252 114468 2304
rect 114520 2292 114526 2304
rect 115106 2292 115112 2304
rect 114520 2264 115112 2292
rect 114520 2252 114526 2264
rect 115106 2252 115112 2264
rect 115164 2252 115170 2304
rect 115934 2252 115940 2304
rect 115992 2292 115998 2304
rect 116305 2295 116363 2301
rect 116305 2292 116317 2295
rect 115992 2264 116317 2292
rect 115992 2252 115998 2264
rect 116305 2261 116317 2264
rect 116351 2261 116363 2295
rect 116762 2292 116768 2304
rect 116723 2264 116768 2292
rect 116305 2255 116363 2261
rect 116762 2252 116768 2264
rect 116820 2252 116826 2304
rect 117406 2292 117412 2304
rect 117367 2264 117412 2292
rect 117406 2252 117412 2264
rect 117464 2252 117470 2304
rect 117593 2295 117651 2301
rect 117593 2261 117605 2295
rect 117639 2292 117651 2295
rect 117869 2295 117927 2301
rect 117869 2292 117881 2295
rect 117639 2264 117881 2292
rect 117639 2261 117651 2264
rect 117593 2255 117651 2261
rect 117869 2261 117881 2264
rect 117915 2292 117927 2295
rect 118510 2292 118516 2304
rect 117915 2264 118516 2292
rect 117915 2261 117927 2264
rect 117869 2255 117927 2261
rect 118510 2252 118516 2264
rect 118568 2252 118574 2304
rect 118602 2252 118608 2304
rect 118660 2292 118666 2304
rect 119154 2292 119160 2304
rect 118660 2264 119160 2292
rect 118660 2252 118666 2264
rect 119154 2252 119160 2264
rect 119212 2252 119218 2304
rect 119338 2292 119344 2304
rect 119299 2264 119344 2292
rect 119338 2252 119344 2264
rect 119396 2252 119402 2304
rect 120902 2252 120908 2304
rect 120960 2292 120966 2304
rect 121181 2295 121239 2301
rect 121181 2292 121193 2295
rect 120960 2264 121193 2292
rect 120960 2252 120966 2264
rect 121181 2261 121193 2264
rect 121227 2261 121239 2295
rect 124214 2292 124220 2304
rect 124127 2264 124220 2292
rect 121181 2255 121239 2261
rect 124214 2252 124220 2264
rect 124272 2292 124278 2304
rect 125318 2292 125324 2304
rect 124272 2264 125324 2292
rect 124272 2252 124278 2264
rect 125318 2252 125324 2264
rect 125376 2252 125382 2304
rect 125413 2295 125471 2301
rect 125413 2261 125425 2295
rect 125459 2292 125471 2295
rect 125594 2292 125600 2304
rect 125459 2264 125600 2292
rect 125459 2261 125471 2264
rect 125413 2255 125471 2261
rect 125594 2252 125600 2264
rect 125652 2252 125658 2304
rect 126241 2295 126299 2301
rect 126241 2261 126253 2295
rect 126287 2292 126299 2295
rect 126517 2295 126575 2301
rect 126517 2292 126529 2295
rect 126287 2264 126529 2292
rect 126287 2261 126299 2264
rect 126241 2255 126299 2261
rect 126517 2261 126529 2264
rect 126563 2292 126575 2295
rect 127158 2292 127164 2304
rect 126563 2264 127164 2292
rect 126563 2261 126575 2264
rect 126517 2255 126575 2261
rect 127158 2252 127164 2264
rect 127216 2252 127222 2304
rect 127805 2295 127863 2301
rect 127805 2261 127817 2295
rect 127851 2292 127863 2295
rect 128096 2292 128124 2468
rect 139673 2465 139685 2468
rect 139719 2465 139731 2499
rect 142890 2496 142896 2508
rect 142851 2468 142896 2496
rect 139673 2459 139731 2465
rect 142890 2456 142896 2468
rect 142948 2456 142954 2508
rect 145190 2456 145196 2508
rect 145248 2496 145254 2508
rect 145377 2499 145435 2505
rect 145377 2496 145389 2499
rect 145248 2468 145389 2496
rect 145248 2456 145254 2468
rect 145377 2465 145389 2468
rect 145423 2465 145435 2499
rect 145377 2459 145435 2465
rect 146389 2499 146447 2505
rect 146389 2465 146401 2499
rect 146435 2496 146447 2499
rect 146478 2496 146484 2508
rect 146435 2468 146484 2496
rect 146435 2465 146447 2468
rect 146389 2459 146447 2465
rect 146478 2456 146484 2468
rect 146536 2456 146542 2508
rect 147766 2496 147772 2508
rect 147727 2468 147772 2496
rect 147766 2456 147772 2468
rect 147824 2456 147830 2508
rect 148781 2499 148839 2505
rect 148781 2465 148793 2499
rect 148827 2496 148839 2499
rect 149330 2496 149336 2508
rect 148827 2468 149336 2496
rect 148827 2465 148839 2468
rect 148781 2459 148839 2465
rect 149330 2456 149336 2468
rect 149388 2456 149394 2508
rect 149422 2456 149428 2508
rect 149480 2496 149486 2508
rect 149977 2499 150035 2505
rect 149977 2496 149989 2499
rect 149480 2468 149989 2496
rect 149480 2456 149486 2468
rect 149977 2465 149989 2468
rect 150023 2465 150035 2499
rect 149977 2459 150035 2465
rect 150989 2499 151047 2505
rect 150989 2465 151001 2499
rect 151035 2496 151047 2499
rect 152090 2496 152096 2508
rect 151035 2468 152096 2496
rect 151035 2465 151047 2468
rect 150989 2459 151047 2465
rect 152090 2456 152096 2468
rect 152148 2456 152154 2508
rect 159453 2499 159511 2505
rect 159453 2465 159465 2499
rect 159499 2496 159511 2499
rect 164510 2496 164516 2508
rect 159499 2468 164516 2496
rect 159499 2465 159511 2468
rect 159453 2459 159511 2465
rect 164510 2456 164516 2468
rect 164568 2456 164574 2508
rect 130102 2388 130108 2440
rect 130160 2428 130166 2440
rect 130197 2431 130255 2437
rect 130197 2428 130209 2431
rect 130160 2400 130209 2428
rect 130160 2388 130166 2400
rect 130197 2397 130209 2400
rect 130243 2397 130255 2431
rect 130197 2391 130255 2397
rect 130289 2431 130347 2437
rect 130289 2397 130301 2431
rect 130335 2428 130347 2431
rect 131114 2428 131120 2440
rect 130335 2400 131120 2428
rect 130335 2397 130347 2400
rect 130289 2391 130347 2397
rect 130212 2360 130240 2391
rect 131114 2388 131120 2400
rect 131172 2388 131178 2440
rect 134242 2388 134248 2440
rect 134300 2428 134306 2440
rect 134981 2431 135039 2437
rect 134981 2428 134993 2431
rect 134300 2400 134993 2428
rect 134300 2388 134306 2400
rect 134981 2397 134993 2400
rect 135027 2397 135039 2431
rect 134981 2391 135039 2397
rect 135073 2431 135131 2437
rect 135073 2397 135085 2431
rect 135119 2428 135131 2431
rect 135990 2428 135996 2440
rect 135119 2400 135996 2428
rect 135119 2397 135131 2400
rect 135073 2391 135131 2397
rect 130657 2363 130715 2369
rect 130657 2360 130669 2363
rect 130212 2332 130669 2360
rect 130657 2329 130669 2332
rect 130703 2329 130715 2363
rect 130657 2323 130715 2329
rect 131022 2320 131028 2372
rect 131080 2360 131086 2372
rect 134996 2360 135024 2391
rect 135990 2388 135996 2400
rect 136048 2388 136054 2440
rect 136361 2431 136419 2437
rect 136361 2397 136373 2431
rect 136407 2397 136419 2431
rect 136361 2391 136419 2397
rect 135441 2363 135499 2369
rect 135441 2360 135453 2363
rect 131080 2332 134288 2360
rect 134996 2332 135453 2360
rect 131080 2320 131086 2332
rect 127851 2264 128124 2292
rect 127851 2261 127863 2264
rect 127805 2255 127863 2261
rect 128170 2252 128176 2304
rect 128228 2292 128234 2304
rect 128357 2295 128415 2301
rect 128357 2292 128369 2295
rect 128228 2264 128369 2292
rect 128228 2252 128234 2264
rect 128357 2261 128369 2264
rect 128403 2292 128415 2295
rect 128998 2292 129004 2304
rect 128403 2264 129004 2292
rect 128403 2261 128415 2264
rect 128357 2255 128415 2261
rect 128998 2252 129004 2264
rect 129056 2252 129062 2304
rect 133046 2252 133052 2304
rect 133104 2292 133110 2304
rect 133233 2295 133291 2301
rect 133233 2292 133245 2295
rect 133104 2264 133245 2292
rect 133104 2252 133110 2264
rect 133233 2261 133245 2264
rect 133279 2261 133291 2295
rect 134150 2292 134156 2304
rect 134111 2264 134156 2292
rect 133233 2255 133291 2261
rect 134150 2252 134156 2264
rect 134208 2252 134214 2304
rect 134260 2292 134288 2332
rect 135441 2329 135453 2332
rect 135487 2329 135499 2363
rect 136376 2360 136404 2391
rect 137462 2388 137468 2440
rect 137520 2428 137526 2440
rect 137557 2431 137615 2437
rect 137557 2428 137569 2431
rect 137520 2400 137569 2428
rect 137520 2388 137526 2400
rect 137557 2397 137569 2400
rect 137603 2428 137615 2431
rect 138385 2431 138443 2437
rect 138385 2428 138397 2431
rect 137603 2400 138397 2428
rect 137603 2397 137615 2400
rect 137557 2391 137615 2397
rect 138385 2397 138397 2400
rect 138431 2397 138443 2431
rect 138658 2428 138664 2440
rect 138619 2400 138664 2428
rect 138385 2391 138443 2397
rect 138658 2388 138664 2400
rect 138716 2428 138722 2440
rect 139302 2428 139308 2440
rect 138716 2400 139308 2428
rect 138716 2388 138722 2400
rect 139302 2388 139308 2400
rect 139360 2388 139366 2440
rect 139578 2388 139584 2440
rect 139636 2428 139642 2440
rect 140225 2431 140283 2437
rect 140225 2428 140237 2431
rect 139636 2400 140237 2428
rect 139636 2388 139642 2400
rect 140225 2397 140237 2400
rect 140271 2428 140283 2431
rect 140501 2431 140559 2437
rect 140501 2428 140513 2431
rect 140271 2400 140513 2428
rect 140271 2397 140283 2400
rect 140225 2391 140283 2397
rect 140501 2397 140513 2400
rect 140547 2397 140559 2431
rect 140501 2391 140559 2397
rect 142801 2431 142859 2437
rect 142801 2397 142813 2431
rect 142847 2428 142859 2431
rect 145285 2431 145343 2437
rect 142847 2400 143396 2428
rect 142847 2397 142859 2400
rect 142801 2391 142859 2397
rect 137281 2363 137339 2369
rect 137281 2360 137293 2363
rect 136376 2332 137293 2360
rect 135441 2323 135499 2329
rect 137281 2329 137293 2332
rect 137327 2360 137339 2363
rect 138014 2360 138020 2372
rect 137327 2332 137784 2360
rect 137975 2332 138020 2360
rect 137327 2329 137339 2332
rect 137281 2323 137339 2329
rect 136453 2295 136511 2301
rect 136453 2292 136465 2295
rect 134260 2264 136465 2292
rect 136453 2261 136465 2264
rect 136499 2261 136511 2295
rect 136453 2255 136511 2261
rect 136634 2252 136640 2304
rect 136692 2292 136698 2304
rect 136821 2295 136879 2301
rect 136821 2292 136833 2295
rect 136692 2264 136833 2292
rect 136692 2252 136698 2264
rect 136821 2261 136833 2264
rect 136867 2261 136879 2295
rect 137646 2292 137652 2304
rect 137607 2264 137652 2292
rect 136821 2255 136879 2261
rect 137646 2252 137652 2264
rect 137704 2252 137710 2304
rect 137756 2292 137784 2332
rect 138014 2320 138020 2332
rect 138072 2320 138078 2372
rect 140866 2360 140872 2372
rect 138124 2332 140872 2360
rect 138124 2292 138152 2332
rect 140866 2320 140872 2332
rect 140924 2320 140930 2372
rect 137756 2264 138152 2292
rect 140774 2252 140780 2304
rect 140832 2292 140838 2304
rect 143368 2301 143396 2400
rect 145285 2397 145297 2431
rect 145331 2428 145343 2431
rect 146294 2428 146300 2440
rect 145331 2400 145972 2428
rect 146255 2400 146300 2428
rect 145331 2397 145343 2400
rect 145285 2391 145343 2397
rect 145944 2304 145972 2400
rect 146294 2388 146300 2400
rect 146352 2428 146358 2440
rect 146757 2431 146815 2437
rect 146757 2428 146769 2431
rect 146352 2400 146769 2428
rect 146352 2388 146358 2400
rect 146757 2397 146769 2400
rect 146803 2397 146815 2431
rect 146757 2391 146815 2397
rect 147030 2388 147036 2440
rect 147088 2428 147094 2440
rect 147677 2431 147735 2437
rect 147677 2428 147689 2431
rect 147088 2400 147689 2428
rect 147088 2388 147094 2400
rect 147677 2397 147689 2400
rect 147723 2428 147735 2431
rect 148137 2431 148195 2437
rect 148137 2428 148149 2431
rect 147723 2400 148149 2428
rect 147723 2397 147735 2400
rect 147677 2391 147735 2397
rect 148137 2397 148149 2400
rect 148183 2397 148195 2431
rect 148137 2391 148195 2397
rect 148689 2431 148747 2437
rect 148689 2397 148701 2431
rect 148735 2397 148747 2431
rect 148689 2391 148747 2397
rect 149885 2431 149943 2437
rect 149885 2397 149897 2431
rect 149931 2428 149943 2431
rect 150894 2428 150900 2440
rect 149931 2400 150480 2428
rect 150855 2400 150900 2428
rect 149931 2397 149943 2400
rect 149885 2391 149943 2397
rect 147766 2320 147772 2372
rect 147824 2360 147830 2372
rect 148704 2360 148732 2391
rect 149149 2363 149207 2369
rect 149149 2360 149161 2363
rect 147824 2332 149161 2360
rect 147824 2320 147830 2332
rect 149149 2329 149161 2332
rect 149195 2329 149207 2363
rect 149149 2323 149207 2329
rect 141053 2295 141111 2301
rect 141053 2292 141065 2295
rect 140832 2264 141065 2292
rect 140832 2252 140838 2264
rect 141053 2261 141065 2264
rect 141099 2261 141111 2295
rect 141053 2255 141111 2261
rect 143353 2295 143411 2301
rect 143353 2261 143365 2295
rect 143399 2292 143411 2295
rect 145190 2292 145196 2304
rect 143399 2264 145196 2292
rect 143399 2261 143411 2264
rect 143353 2255 143411 2261
rect 145190 2252 145196 2264
rect 145248 2252 145254 2304
rect 145558 2252 145564 2304
rect 145616 2292 145622 2304
rect 145745 2295 145803 2301
rect 145745 2292 145757 2295
rect 145616 2264 145757 2292
rect 145616 2252 145622 2264
rect 145745 2261 145757 2264
rect 145791 2261 145803 2295
rect 145745 2255 145803 2261
rect 145926 2252 145932 2304
rect 145984 2292 145990 2304
rect 146113 2295 146171 2301
rect 146113 2292 146125 2295
rect 145984 2264 146125 2292
rect 145984 2252 145990 2264
rect 146113 2261 146125 2264
rect 146159 2261 146171 2295
rect 146113 2255 146171 2261
rect 149054 2252 149060 2304
rect 149112 2292 149118 2304
rect 149609 2295 149667 2301
rect 149609 2292 149621 2295
rect 149112 2264 149621 2292
rect 149112 2252 149118 2264
rect 149609 2261 149621 2264
rect 149655 2292 149667 2295
rect 149882 2292 149888 2304
rect 149655 2264 149888 2292
rect 149655 2261 149667 2264
rect 149609 2255 149667 2261
rect 149882 2252 149888 2264
rect 149940 2252 149946 2304
rect 150452 2301 150480 2400
rect 150894 2388 150900 2400
rect 150952 2428 150958 2440
rect 151357 2431 151415 2437
rect 151357 2428 151369 2431
rect 150952 2400 151369 2428
rect 150952 2388 150958 2400
rect 151357 2397 151369 2400
rect 151403 2397 151415 2431
rect 151357 2391 151415 2397
rect 151814 2388 151820 2440
rect 151872 2428 151878 2440
rect 151909 2431 151967 2437
rect 151909 2428 151921 2431
rect 151872 2400 151921 2428
rect 151872 2388 151878 2400
rect 151909 2397 151921 2400
rect 151955 2428 151967 2431
rect 152369 2431 152427 2437
rect 152369 2428 152381 2431
rect 151955 2400 152381 2428
rect 151955 2397 151967 2400
rect 151909 2391 151967 2397
rect 152369 2397 152381 2400
rect 152415 2397 152427 2431
rect 152369 2391 152427 2397
rect 155494 2388 155500 2440
rect 155552 2428 155558 2440
rect 155773 2431 155831 2437
rect 155773 2428 155785 2431
rect 155552 2400 155785 2428
rect 155552 2388 155558 2400
rect 155773 2397 155785 2400
rect 155819 2397 155831 2431
rect 155773 2391 155831 2397
rect 151170 2320 151176 2372
rect 151228 2360 151234 2372
rect 152001 2363 152059 2369
rect 152001 2360 152013 2363
rect 151228 2332 152013 2360
rect 151228 2320 151234 2332
rect 152001 2329 152013 2332
rect 152047 2329 152059 2363
rect 155788 2360 155816 2391
rect 156230 2388 156236 2440
rect 156288 2428 156294 2440
rect 156601 2431 156659 2437
rect 156601 2428 156613 2431
rect 156288 2400 156613 2428
rect 156288 2388 156294 2400
rect 156601 2397 156613 2400
rect 156647 2397 156659 2431
rect 156601 2391 156659 2397
rect 157245 2431 157303 2437
rect 157245 2397 157257 2431
rect 157291 2428 157303 2431
rect 158349 2431 158407 2437
rect 157291 2400 157748 2428
rect 157291 2397 157303 2400
rect 157245 2391 157303 2397
rect 156325 2363 156383 2369
rect 156325 2360 156337 2363
rect 155788 2332 156337 2360
rect 152001 2323 152059 2329
rect 156325 2329 156337 2332
rect 156371 2329 156383 2363
rect 156325 2323 156383 2329
rect 157720 2304 157748 2400
rect 158349 2397 158361 2431
rect 158395 2428 158407 2431
rect 158438 2428 158444 2440
rect 158395 2400 158444 2428
rect 158395 2397 158407 2400
rect 158349 2391 158407 2397
rect 158438 2388 158444 2400
rect 158496 2428 158502 2440
rect 158809 2431 158867 2437
rect 158809 2428 158821 2431
rect 158496 2400 158821 2428
rect 158496 2388 158502 2400
rect 158809 2397 158821 2400
rect 158855 2397 158867 2431
rect 159358 2428 159364 2440
rect 159319 2400 159364 2428
rect 158809 2391 158867 2397
rect 159358 2388 159364 2400
rect 159416 2428 159422 2440
rect 159821 2431 159879 2437
rect 159821 2428 159833 2431
rect 159416 2400 159833 2428
rect 159416 2388 159422 2400
rect 159821 2397 159833 2400
rect 159867 2397 159879 2431
rect 159821 2391 159879 2397
rect 161014 2388 161020 2440
rect 161072 2428 161078 2440
rect 161661 2431 161719 2437
rect 161661 2428 161673 2431
rect 161072 2400 161673 2428
rect 161072 2388 161078 2400
rect 161661 2397 161673 2400
rect 161707 2428 161719 2431
rect 162121 2431 162179 2437
rect 162121 2428 162133 2431
rect 161707 2400 162133 2428
rect 161707 2397 161719 2400
rect 161661 2391 161719 2397
rect 162121 2397 162133 2400
rect 162167 2397 162179 2431
rect 162121 2391 162179 2397
rect 162210 2388 162216 2440
rect 162268 2428 162274 2440
rect 162673 2431 162731 2437
rect 162673 2428 162685 2431
rect 162268 2400 162685 2428
rect 162268 2388 162274 2400
rect 162673 2397 162685 2400
rect 162719 2428 162731 2431
rect 163133 2431 163191 2437
rect 163133 2428 163145 2431
rect 162719 2400 163145 2428
rect 162719 2397 162731 2400
rect 162673 2391 162731 2397
rect 163133 2397 163145 2400
rect 163179 2397 163191 2431
rect 164602 2428 164608 2440
rect 164515 2400 164608 2428
rect 163133 2391 163191 2397
rect 164602 2388 164608 2400
rect 164660 2388 164666 2440
rect 161566 2320 161572 2372
rect 161624 2360 161630 2372
rect 164620 2360 164648 2388
rect 161624 2332 164648 2360
rect 165433 2363 165491 2369
rect 161624 2320 161630 2332
rect 165433 2329 165445 2363
rect 165479 2360 165491 2363
rect 165798 2360 165804 2372
rect 165479 2332 165804 2360
rect 165479 2329 165491 2332
rect 165433 2323 165491 2329
rect 165798 2320 165804 2332
rect 165856 2320 165862 2372
rect 150437 2295 150495 2301
rect 150437 2261 150449 2295
rect 150483 2292 150495 2295
rect 150710 2292 150716 2304
rect 150483 2264 150716 2292
rect 150483 2261 150495 2264
rect 150437 2255 150495 2261
rect 150710 2252 150716 2264
rect 150768 2252 150774 2304
rect 154301 2295 154359 2301
rect 154301 2261 154313 2295
rect 154347 2292 154359 2295
rect 154390 2292 154396 2304
rect 154347 2264 154396 2292
rect 154347 2261 154359 2264
rect 154301 2255 154359 2261
rect 154390 2252 154396 2264
rect 154448 2252 154454 2304
rect 154758 2252 154764 2304
rect 154816 2292 154822 2304
rect 155218 2292 155224 2304
rect 154816 2264 155224 2292
rect 154816 2252 154822 2264
rect 155218 2252 155224 2264
rect 155276 2252 155282 2304
rect 157702 2292 157708 2304
rect 157663 2264 157708 2292
rect 157702 2252 157708 2264
rect 157760 2252 157766 2304
rect 160278 2252 160284 2304
rect 160336 2292 160342 2304
rect 160646 2292 160652 2304
rect 160336 2264 160652 2292
rect 160336 2252 160342 2264
rect 160646 2252 160652 2264
rect 160704 2252 160710 2304
rect 164053 2295 164111 2301
rect 164053 2261 164065 2295
rect 164099 2292 164111 2295
rect 164142 2292 164148 2304
rect 164099 2264 164148 2292
rect 164099 2261 164111 2264
rect 164053 2255 164111 2261
rect 164142 2252 164148 2264
rect 164200 2252 164206 2304
rect 368 2202 93012 2224
rect 368 2150 56667 2202
rect 56719 2150 56731 2202
rect 56783 2150 56795 2202
rect 56847 2150 56859 2202
rect 56911 2150 93012 2202
rect 368 2128 93012 2150
rect 102028 2202 169556 2224
rect 102028 2150 113088 2202
rect 113140 2150 113152 2202
rect 113204 2150 113216 2202
rect 113268 2150 113280 2202
rect 113332 2150 169556 2202
rect 102028 2128 169556 2150
rect 6270 2088 6276 2100
rect 6231 2060 6276 2088
rect 6270 2048 6276 2060
rect 6328 2048 6334 2100
rect 7282 2048 7288 2100
rect 7340 2088 7346 2100
rect 12158 2088 12164 2100
rect 7340 2060 12164 2088
rect 7340 2048 7346 2060
rect 12158 2048 12164 2060
rect 12216 2048 12222 2100
rect 17313 2091 17371 2097
rect 17313 2057 17325 2091
rect 17359 2088 17371 2091
rect 18506 2088 18512 2100
rect 17359 2060 18512 2088
rect 17359 2057 17371 2060
rect 17313 2051 17371 2057
rect 18506 2048 18512 2060
rect 18564 2048 18570 2100
rect 19610 2048 19616 2100
rect 19668 2088 19674 2100
rect 42610 2088 42616 2100
rect 19668 2060 42616 2088
rect 19668 2048 19674 2060
rect 42610 2048 42616 2060
rect 42668 2048 42674 2100
rect 42794 2088 42800 2100
rect 42755 2060 42800 2088
rect 42794 2048 42800 2060
rect 42852 2048 42858 2100
rect 43530 2088 43536 2100
rect 42904 2060 43536 2088
rect 2958 1980 2964 2032
rect 3016 2020 3022 2032
rect 3016 1992 10272 2020
rect 3016 1980 3022 1992
rect 3050 1912 3056 1964
rect 3108 1952 3114 1964
rect 4801 1955 4859 1961
rect 3108 1924 4384 1952
rect 3108 1912 3114 1924
rect 2225 1887 2283 1893
rect 2225 1853 2237 1887
rect 2271 1884 2283 1887
rect 3234 1884 3240 1896
rect 2271 1856 3240 1884
rect 2271 1853 2283 1856
rect 2225 1847 2283 1853
rect 3234 1844 3240 1856
rect 3292 1844 3298 1896
rect 4249 1887 4307 1893
rect 4249 1853 4261 1887
rect 4295 1853 4307 1887
rect 4356 1884 4384 1924
rect 4801 1921 4813 1955
rect 4847 1952 4859 1955
rect 5166 1952 5172 1964
rect 4847 1924 5172 1952
rect 4847 1921 4859 1924
rect 4801 1915 4859 1921
rect 5166 1912 5172 1924
rect 5224 1912 5230 1964
rect 8205 1955 8263 1961
rect 5276 1924 7788 1952
rect 5276 1884 5304 1924
rect 4356 1856 5304 1884
rect 6641 1887 6699 1893
rect 4249 1847 4307 1853
rect 6641 1853 6653 1887
rect 6687 1884 6699 1887
rect 7190 1884 7196 1896
rect 6687 1856 7196 1884
rect 6687 1853 6699 1856
rect 6641 1847 6699 1853
rect 2774 1776 2780 1828
rect 2832 1816 2838 1828
rect 4264 1816 4292 1847
rect 7190 1844 7196 1856
rect 7248 1844 7254 1896
rect 7653 1887 7711 1893
rect 7653 1853 7665 1887
rect 7699 1853 7711 1887
rect 7653 1847 7711 1853
rect 7668 1816 7696 1847
rect 2832 1788 4292 1816
rect 4632 1788 7696 1816
rect 7760 1816 7788 1924
rect 8205 1921 8217 1955
rect 8251 1952 8263 1955
rect 8386 1952 8392 1964
rect 8251 1924 8392 1952
rect 8251 1921 8263 1924
rect 8205 1915 8263 1921
rect 8386 1912 8392 1924
rect 8444 1912 8450 1964
rect 9214 1884 9220 1896
rect 9175 1856 9220 1884
rect 9214 1844 9220 1856
rect 9272 1844 9278 1896
rect 10244 1893 10272 1992
rect 10318 1980 10324 2032
rect 10376 2020 10382 2032
rect 32490 2020 32496 2032
rect 10376 1992 32496 2020
rect 10376 1980 10382 1992
rect 32490 1980 32496 1992
rect 32548 1980 32554 2032
rect 32674 1980 32680 2032
rect 32732 2020 32738 2032
rect 38470 2020 38476 2032
rect 32732 1992 38476 2020
rect 32732 1980 32738 1992
rect 38470 1980 38476 1992
rect 38528 1980 38534 2032
rect 38562 1980 38568 2032
rect 38620 2020 38626 2032
rect 41322 2020 41328 2032
rect 38620 1992 41328 2020
rect 38620 1980 38626 1992
rect 41322 1980 41328 1992
rect 41380 1980 41386 2032
rect 41414 1980 41420 2032
rect 41472 2020 41478 2032
rect 42061 2023 42119 2029
rect 41472 1992 41828 2020
rect 41472 1980 41478 1992
rect 10778 1952 10784 1964
rect 10739 1924 10784 1952
rect 10778 1912 10784 1924
rect 10836 1912 10842 1964
rect 15378 1912 15384 1964
rect 15436 1952 15442 1964
rect 20901 1955 20959 1961
rect 15436 1924 20392 1952
rect 15436 1912 15442 1924
rect 10229 1887 10287 1893
rect 10229 1853 10241 1887
rect 10275 1853 10287 1887
rect 11146 1884 11152 1896
rect 11059 1856 11152 1884
rect 10229 1847 10287 1853
rect 11146 1844 11152 1856
rect 11204 1884 11210 1896
rect 11701 1887 11759 1893
rect 11701 1884 11713 1887
rect 11204 1856 11713 1884
rect 11204 1844 11210 1856
rect 11701 1853 11713 1856
rect 11747 1853 11759 1887
rect 15102 1884 15108 1896
rect 15063 1856 15108 1884
rect 11701 1847 11759 1853
rect 15102 1844 15108 1856
rect 15160 1844 15166 1896
rect 18325 1887 18383 1893
rect 18325 1853 18337 1887
rect 18371 1884 18383 1887
rect 19337 1887 19395 1893
rect 19337 1884 19349 1887
rect 18371 1856 19349 1884
rect 18371 1853 18383 1856
rect 18325 1847 18383 1853
rect 19337 1853 19349 1856
rect 19383 1884 19395 1887
rect 19794 1884 19800 1896
rect 19383 1856 19800 1884
rect 19383 1853 19395 1856
rect 19337 1847 19395 1853
rect 19794 1844 19800 1856
rect 19852 1844 19858 1896
rect 20364 1893 20392 1924
rect 20901 1921 20913 1955
rect 20947 1952 20959 1955
rect 20993 1955 21051 1961
rect 20993 1952 21005 1955
rect 20947 1924 21005 1952
rect 20947 1921 20959 1924
rect 20901 1915 20959 1921
rect 20993 1921 21005 1924
rect 21039 1921 21051 1955
rect 20993 1915 21051 1921
rect 21266 1912 21272 1964
rect 21324 1952 21330 1964
rect 21324 1924 24716 1952
rect 21324 1912 21330 1924
rect 20349 1887 20407 1893
rect 20349 1853 20361 1887
rect 20395 1853 20407 1887
rect 20349 1847 20407 1853
rect 21729 1887 21787 1893
rect 21729 1853 21741 1887
rect 21775 1884 21787 1887
rect 22554 1884 22560 1896
rect 21775 1856 22560 1884
rect 21775 1853 21787 1856
rect 21729 1847 21787 1853
rect 22554 1844 22560 1856
rect 22612 1844 22618 1896
rect 23658 1884 23664 1896
rect 23619 1856 23664 1884
rect 23658 1844 23664 1856
rect 23716 1844 23722 1896
rect 24688 1893 24716 1924
rect 25038 1912 25044 1964
rect 25096 1952 25102 1964
rect 25225 1955 25283 1961
rect 25225 1952 25237 1955
rect 25096 1924 25237 1952
rect 25096 1912 25102 1924
rect 25225 1921 25237 1924
rect 25271 1952 25283 1955
rect 25271 1924 26188 1952
rect 25271 1921 25283 1924
rect 25225 1915 25283 1921
rect 24673 1887 24731 1893
rect 24673 1853 24685 1887
rect 24719 1853 24731 1887
rect 24673 1847 24731 1853
rect 26053 1887 26111 1893
rect 26053 1853 26065 1887
rect 26099 1853 26111 1887
rect 26160 1884 26188 1924
rect 26234 1912 26240 1964
rect 26292 1952 26298 1964
rect 26697 1955 26755 1961
rect 26697 1952 26709 1955
rect 26292 1924 26709 1952
rect 26292 1912 26298 1924
rect 26697 1921 26709 1924
rect 26743 1952 26755 1955
rect 26786 1952 26792 1964
rect 26743 1924 26792 1952
rect 26743 1921 26755 1924
rect 26697 1915 26755 1921
rect 26786 1912 26792 1924
rect 26844 1912 26850 1964
rect 28810 1952 28816 1964
rect 26896 1924 28816 1952
rect 26326 1884 26332 1896
rect 26160 1856 26332 1884
rect 26053 1847 26111 1853
rect 11790 1816 11796 1828
rect 7760 1788 11796 1816
rect 2832 1776 2838 1788
rect 4062 1708 4068 1760
rect 4120 1748 4126 1760
rect 4632 1748 4660 1788
rect 11790 1776 11796 1788
rect 11848 1776 11854 1828
rect 13814 1776 13820 1828
rect 13872 1816 13878 1828
rect 13872 1788 22692 1816
rect 13872 1776 13878 1788
rect 5166 1748 5172 1760
rect 4120 1720 4660 1748
rect 5127 1720 5172 1748
rect 4120 1708 4126 1720
rect 5166 1708 5172 1720
rect 5224 1708 5230 1760
rect 7558 1708 7564 1760
rect 7616 1748 7622 1760
rect 8662 1748 8668 1760
rect 7616 1720 8668 1748
rect 7616 1708 7622 1720
rect 8662 1708 8668 1720
rect 8720 1708 8726 1760
rect 20993 1751 21051 1757
rect 20993 1717 21005 1751
rect 21039 1748 21051 1751
rect 21266 1748 21272 1760
rect 21039 1720 21272 1748
rect 21039 1717 21051 1720
rect 20993 1711 21051 1717
rect 21266 1708 21272 1720
rect 21324 1708 21330 1760
rect 22554 1748 22560 1760
rect 22515 1720 22560 1748
rect 22554 1708 22560 1720
rect 22612 1708 22618 1760
rect 22664 1748 22692 1788
rect 22738 1776 22744 1828
rect 22796 1816 22802 1828
rect 26068 1816 26096 1847
rect 26326 1844 26332 1856
rect 26384 1844 26390 1896
rect 26602 1844 26608 1896
rect 26660 1884 26666 1896
rect 26896 1884 26924 1924
rect 28810 1912 28816 1924
rect 28868 1912 28874 1964
rect 30009 1955 30067 1961
rect 30009 1921 30021 1955
rect 30055 1921 30067 1955
rect 30009 1915 30067 1921
rect 26660 1856 26924 1884
rect 26660 1844 26666 1856
rect 28258 1844 28264 1896
rect 28316 1884 28322 1896
rect 28537 1887 28595 1893
rect 28537 1884 28549 1887
rect 28316 1856 28549 1884
rect 28316 1844 28322 1856
rect 28537 1853 28549 1856
rect 28583 1853 28595 1887
rect 30024 1884 30052 1915
rect 30098 1912 30104 1964
rect 30156 1952 30162 1964
rect 30466 1952 30472 1964
rect 30156 1924 30201 1952
rect 30379 1924 30472 1952
rect 30156 1912 30162 1924
rect 30466 1912 30472 1924
rect 30524 1952 30530 1964
rect 36630 1952 36636 1964
rect 30524 1924 36636 1952
rect 30524 1912 30530 1924
rect 36630 1912 36636 1924
rect 36688 1912 36694 1964
rect 36722 1912 36728 1964
rect 36780 1952 36786 1964
rect 41598 1952 41604 1964
rect 36780 1924 41604 1952
rect 36780 1912 36786 1924
rect 41598 1912 41604 1924
rect 41656 1912 41662 1964
rect 41800 1952 41828 1992
rect 42061 1989 42073 2023
rect 42107 2020 42119 2023
rect 42904 2020 42932 2060
rect 43530 2048 43536 2060
rect 43588 2048 43594 2100
rect 44174 2088 44180 2100
rect 44135 2060 44180 2088
rect 44174 2048 44180 2060
rect 44232 2048 44238 2100
rect 44266 2048 44272 2100
rect 44324 2088 44330 2100
rect 47302 2088 47308 2100
rect 44324 2060 47308 2088
rect 44324 2048 44330 2060
rect 47302 2048 47308 2060
rect 47360 2048 47366 2100
rect 47578 2048 47584 2100
rect 47636 2088 47642 2100
rect 48961 2091 49019 2097
rect 48961 2088 48973 2091
rect 47636 2060 48973 2088
rect 47636 2048 47642 2060
rect 48961 2057 48973 2060
rect 49007 2057 49019 2091
rect 48961 2051 49019 2057
rect 49050 2048 49056 2100
rect 49108 2088 49114 2100
rect 51074 2088 51080 2100
rect 49108 2060 51080 2088
rect 49108 2048 49114 2060
rect 51074 2048 51080 2060
rect 51132 2048 51138 2100
rect 51258 2048 51264 2100
rect 51316 2088 51322 2100
rect 52454 2088 52460 2100
rect 51316 2060 52460 2088
rect 51316 2048 51322 2060
rect 52454 2048 52460 2060
rect 52512 2048 52518 2100
rect 53098 2048 53104 2100
rect 53156 2088 53162 2100
rect 55490 2088 55496 2100
rect 53156 2060 55496 2088
rect 53156 2048 53162 2060
rect 55490 2048 55496 2060
rect 55548 2048 55554 2100
rect 59998 2088 60004 2100
rect 55784 2060 60004 2088
rect 42107 1992 42932 2020
rect 42981 2023 43039 2029
rect 42107 1989 42119 1992
rect 42061 1983 42119 1989
rect 42981 1989 42993 2023
rect 43027 2020 43039 2023
rect 47210 2020 47216 2032
rect 43027 1992 47216 2020
rect 43027 1989 43039 1992
rect 42981 1983 43039 1989
rect 47210 1980 47216 1992
rect 47268 1980 47274 2032
rect 47670 1980 47676 2032
rect 47728 2020 47734 2032
rect 47728 1992 49188 2020
rect 47728 1980 47734 1992
rect 43622 1952 43628 1964
rect 41800 1924 43628 1952
rect 43622 1912 43628 1924
rect 43680 1912 43686 1964
rect 43717 1955 43775 1961
rect 43717 1921 43729 1955
rect 43763 1952 43775 1955
rect 44174 1952 44180 1964
rect 43763 1924 44180 1952
rect 43763 1921 43775 1924
rect 43717 1915 43775 1921
rect 44174 1912 44180 1924
rect 44232 1912 44238 1964
rect 45094 1912 45100 1964
rect 45152 1952 45158 1964
rect 45557 1955 45615 1961
rect 45557 1952 45569 1955
rect 45152 1924 45569 1952
rect 45152 1912 45158 1924
rect 45557 1921 45569 1924
rect 45603 1921 45615 1955
rect 46106 1952 46112 1964
rect 46067 1924 46112 1952
rect 45557 1915 45615 1921
rect 46106 1912 46112 1924
rect 46164 1952 46170 1964
rect 46474 1952 46480 1964
rect 46164 1924 46480 1952
rect 46164 1912 46170 1924
rect 46474 1912 46480 1924
rect 46532 1912 46538 1964
rect 46842 1912 46848 1964
rect 46900 1952 46906 1964
rect 47578 1952 47584 1964
rect 46900 1924 47584 1952
rect 46900 1912 46906 1924
rect 47578 1912 47584 1924
rect 47636 1912 47642 1964
rect 47765 1955 47823 1961
rect 47765 1921 47777 1955
rect 47811 1952 47823 1955
rect 48130 1952 48136 1964
rect 47811 1924 48136 1952
rect 47811 1921 47823 1924
rect 47765 1915 47823 1921
rect 48130 1912 48136 1924
rect 48188 1912 48194 1964
rect 48682 1912 48688 1964
rect 48740 1952 48746 1964
rect 48777 1955 48835 1961
rect 48777 1952 48789 1955
rect 48740 1924 48789 1952
rect 48740 1912 48746 1924
rect 48777 1921 48789 1924
rect 48823 1921 48835 1955
rect 49160 1952 49188 1992
rect 49418 1980 49424 2032
rect 49476 2020 49482 2032
rect 50246 2020 50252 2032
rect 49476 1992 50252 2020
rect 49476 1980 49482 1992
rect 50246 1980 50252 1992
rect 50304 1980 50310 2032
rect 51169 2023 51227 2029
rect 50724 1992 51120 2020
rect 50724 1952 50752 1992
rect 49160 1924 50752 1952
rect 51092 1952 51120 1992
rect 51169 1989 51181 2023
rect 51215 2020 51227 2023
rect 53834 2020 53840 2032
rect 51215 1992 53840 2020
rect 51215 1989 51227 1992
rect 51169 1983 51227 1989
rect 53834 1980 53840 1992
rect 53892 2020 53898 2032
rect 54021 2023 54079 2029
rect 54021 2020 54033 2023
rect 53892 1992 54033 2020
rect 53892 1980 53898 1992
rect 54021 1989 54033 1992
rect 54067 1989 54079 2023
rect 54021 1983 54079 1989
rect 54110 1980 54116 2032
rect 54168 2020 54174 2032
rect 55784 2020 55812 2060
rect 59998 2048 60004 2060
rect 60056 2048 60062 2100
rect 60366 2088 60372 2100
rect 60327 2060 60372 2088
rect 60366 2048 60372 2060
rect 60424 2048 60430 2100
rect 60826 2088 60832 2100
rect 60568 2060 60832 2088
rect 54168 1992 55812 2020
rect 54168 1980 54174 1992
rect 55858 1980 55864 2032
rect 55916 2020 55922 2032
rect 55916 1992 56088 2020
rect 55916 1980 55922 1992
rect 51902 1952 51908 1964
rect 51092 1924 51908 1952
rect 48777 1915 48835 1921
rect 51902 1912 51908 1924
rect 51960 1912 51966 1964
rect 53650 1952 53656 1964
rect 52012 1924 53328 1952
rect 53611 1924 53656 1952
rect 30745 1887 30803 1893
rect 30745 1884 30757 1887
rect 30024 1856 30757 1884
rect 28537 1847 28595 1853
rect 30745 1853 30757 1856
rect 30791 1884 30803 1887
rect 31297 1887 31355 1893
rect 31297 1884 31309 1887
rect 30791 1856 31309 1884
rect 30791 1853 30803 1856
rect 30745 1847 30803 1853
rect 31297 1853 31309 1856
rect 31343 1853 31355 1887
rect 31297 1847 31355 1853
rect 32309 1887 32367 1893
rect 32309 1853 32321 1887
rect 32355 1884 32367 1887
rect 33594 1884 33600 1896
rect 32355 1856 33600 1884
rect 32355 1853 32367 1856
rect 32309 1847 32367 1853
rect 33594 1844 33600 1856
rect 33652 1844 33658 1896
rect 34517 1887 34575 1893
rect 34517 1853 34529 1887
rect 34563 1884 34575 1887
rect 35342 1884 35348 1896
rect 34563 1856 35348 1884
rect 34563 1853 34575 1856
rect 34517 1847 34575 1853
rect 35342 1844 35348 1856
rect 35400 1884 35406 1896
rect 35529 1887 35587 1893
rect 35529 1884 35541 1887
rect 35400 1856 35541 1884
rect 35400 1844 35406 1856
rect 35529 1853 35541 1856
rect 35575 1853 35587 1887
rect 35529 1847 35587 1853
rect 35897 1887 35955 1893
rect 35897 1853 35909 1887
rect 35943 1884 35955 1887
rect 36998 1884 37004 1896
rect 35943 1856 37004 1884
rect 35943 1853 35955 1856
rect 35897 1847 35955 1853
rect 36998 1844 37004 1856
rect 37056 1884 37062 1896
rect 37185 1887 37243 1893
rect 37185 1884 37197 1887
rect 37056 1856 37197 1884
rect 37056 1844 37062 1856
rect 37185 1853 37197 1856
rect 37231 1853 37243 1887
rect 37185 1847 37243 1853
rect 37274 1844 37280 1896
rect 37332 1884 37338 1896
rect 41046 1884 41052 1896
rect 37332 1856 41052 1884
rect 37332 1844 37338 1856
rect 41046 1844 41052 1856
rect 41104 1844 41110 1896
rect 41138 1844 41144 1896
rect 41196 1884 41202 1896
rect 50706 1884 50712 1896
rect 41196 1856 50712 1884
rect 41196 1844 41202 1856
rect 50706 1844 50712 1856
rect 50764 1844 50770 1896
rect 51442 1884 51448 1896
rect 50816 1856 51448 1884
rect 22796 1788 26096 1816
rect 26160 1788 30972 1816
rect 22796 1776 22802 1788
rect 26160 1748 26188 1788
rect 22664 1720 26188 1748
rect 26234 1708 26240 1760
rect 26292 1748 26298 1760
rect 28994 1748 29000 1760
rect 26292 1720 29000 1748
rect 26292 1708 26298 1720
rect 28994 1708 29000 1720
rect 29052 1708 29058 1760
rect 30944 1748 30972 1788
rect 33502 1776 33508 1828
rect 33560 1816 33566 1828
rect 36446 1816 36452 1828
rect 33560 1788 36452 1816
rect 33560 1776 33566 1788
rect 36446 1776 36452 1788
rect 36504 1776 36510 1828
rect 50816 1816 50844 1856
rect 51442 1844 51448 1856
rect 51500 1844 51506 1896
rect 52012 1884 52040 1924
rect 52178 1884 52184 1896
rect 51552 1856 52040 1884
rect 52139 1856 52184 1884
rect 51552 1816 51580 1856
rect 52178 1844 52184 1856
rect 52236 1844 52242 1896
rect 53193 1887 53251 1893
rect 53193 1853 53205 1887
rect 53239 1853 53251 1887
rect 53300 1884 53328 1924
rect 53650 1912 53656 1924
rect 53708 1912 53714 1964
rect 55214 1952 55220 1964
rect 55127 1924 55220 1952
rect 55214 1912 55220 1924
rect 55272 1952 55278 1964
rect 55950 1952 55956 1964
rect 55272 1924 55956 1952
rect 55272 1912 55278 1924
rect 55950 1912 55956 1924
rect 56008 1912 56014 1964
rect 56060 1952 56088 1992
rect 56318 1980 56324 2032
rect 56376 2020 56382 2032
rect 60568 2020 60596 2060
rect 60826 2048 60832 2060
rect 60884 2048 60890 2100
rect 63770 2088 63776 2100
rect 61396 2060 63776 2088
rect 61396 2020 61424 2060
rect 63770 2048 63776 2060
rect 63828 2048 63834 2100
rect 63865 2091 63923 2097
rect 63865 2057 63877 2091
rect 63911 2088 63923 2091
rect 64690 2088 64696 2100
rect 63911 2060 64696 2088
rect 63911 2057 63923 2060
rect 63865 2051 63923 2057
rect 64690 2048 64696 2060
rect 64748 2048 64754 2100
rect 65058 2048 65064 2100
rect 65116 2088 65122 2100
rect 65153 2091 65211 2097
rect 65153 2088 65165 2091
rect 65116 2060 65165 2088
rect 65116 2048 65122 2060
rect 65153 2057 65165 2060
rect 65199 2057 65211 2091
rect 66806 2088 66812 2100
rect 66767 2060 66812 2088
rect 65153 2051 65211 2057
rect 66806 2048 66812 2060
rect 66864 2048 66870 2100
rect 66898 2048 66904 2100
rect 66956 2088 66962 2100
rect 67726 2088 67732 2100
rect 66956 2060 67732 2088
rect 66956 2048 66962 2060
rect 67726 2048 67732 2060
rect 67784 2048 67790 2100
rect 67836 2060 69244 2088
rect 56376 1992 60596 2020
rect 60660 1992 61424 2020
rect 61657 2023 61715 2029
rect 56376 1980 56382 1992
rect 57698 1952 57704 1964
rect 56060 1924 57704 1952
rect 57698 1912 57704 1924
rect 57756 1912 57762 1964
rect 57882 1952 57888 1964
rect 57843 1924 57888 1952
rect 57882 1912 57888 1924
rect 57940 1912 57946 1964
rect 58434 1912 58440 1964
rect 58492 1952 58498 1964
rect 58802 1952 58808 1964
rect 58492 1924 58808 1952
rect 58492 1912 58498 1924
rect 58802 1912 58808 1924
rect 58860 1952 58866 1964
rect 58989 1955 59047 1961
rect 58989 1952 59001 1955
rect 58860 1924 59001 1952
rect 58860 1912 58866 1924
rect 58989 1921 59001 1924
rect 59035 1921 59047 1955
rect 58989 1915 59047 1921
rect 59541 1955 59599 1961
rect 59541 1921 59553 1955
rect 59587 1952 59599 1955
rect 60001 1955 60059 1961
rect 60001 1952 60013 1955
rect 59587 1924 60013 1952
rect 59587 1921 59599 1924
rect 59541 1915 59599 1921
rect 60001 1921 60013 1924
rect 60047 1921 60059 1955
rect 60001 1915 60059 1921
rect 54573 1887 54631 1893
rect 54573 1884 54585 1887
rect 53300 1856 54585 1884
rect 53193 1847 53251 1853
rect 54573 1853 54585 1856
rect 54619 1853 54631 1887
rect 54573 1847 54631 1853
rect 36556 1788 37228 1816
rect 36556 1748 36584 1788
rect 30944 1720 36584 1748
rect 36814 1708 36820 1760
rect 36872 1748 36878 1760
rect 37090 1748 37096 1760
rect 36872 1720 37096 1748
rect 36872 1708 36878 1720
rect 37090 1708 37096 1720
rect 37148 1708 37154 1760
rect 37200 1748 37228 1788
rect 37384 1788 50844 1816
rect 50908 1788 51580 1816
rect 37384 1748 37412 1788
rect 37200 1720 37412 1748
rect 38102 1708 38108 1760
rect 38160 1748 38166 1760
rect 38562 1748 38568 1760
rect 38160 1720 38568 1748
rect 38160 1708 38166 1720
rect 38562 1708 38568 1720
rect 38620 1708 38626 1760
rect 38654 1708 38660 1760
rect 38712 1748 38718 1760
rect 39022 1748 39028 1760
rect 38712 1720 39028 1748
rect 38712 1708 38718 1720
rect 39022 1708 39028 1720
rect 39080 1708 39086 1760
rect 41322 1708 41328 1760
rect 41380 1748 41386 1760
rect 42981 1751 43039 1757
rect 42981 1748 42993 1751
rect 41380 1720 42993 1748
rect 41380 1708 41386 1720
rect 42981 1717 42993 1720
rect 43027 1717 43039 1751
rect 42981 1711 43039 1717
rect 43533 1751 43591 1757
rect 43533 1717 43545 1751
rect 43579 1748 43591 1751
rect 43622 1748 43628 1760
rect 43579 1720 43628 1748
rect 43579 1717 43591 1720
rect 43533 1711 43591 1717
rect 43622 1708 43628 1720
rect 43680 1708 43686 1760
rect 43714 1708 43720 1760
rect 43772 1748 43778 1760
rect 44453 1751 44511 1757
rect 44453 1748 44465 1751
rect 43772 1720 44465 1748
rect 43772 1708 43778 1720
rect 44453 1717 44465 1720
rect 44499 1717 44511 1751
rect 44453 1711 44511 1717
rect 45462 1708 45468 1760
rect 45520 1748 45526 1760
rect 47397 1751 47455 1757
rect 47397 1748 47409 1751
rect 45520 1720 47409 1748
rect 45520 1708 45526 1720
rect 47397 1717 47409 1720
rect 47443 1717 47455 1751
rect 47397 1711 47455 1717
rect 47486 1708 47492 1760
rect 47544 1748 47550 1760
rect 49050 1748 49056 1760
rect 47544 1720 49056 1748
rect 47544 1708 47550 1720
rect 49050 1708 49056 1720
rect 49108 1708 49114 1760
rect 49142 1708 49148 1760
rect 49200 1748 49206 1760
rect 50614 1748 50620 1760
rect 49200 1720 50620 1748
rect 49200 1708 49206 1720
rect 50614 1708 50620 1720
rect 50672 1708 50678 1760
rect 50706 1708 50712 1760
rect 50764 1748 50770 1760
rect 50908 1748 50936 1788
rect 51810 1776 51816 1828
rect 51868 1816 51874 1828
rect 53208 1816 53236 1847
rect 54938 1844 54944 1896
rect 54996 1884 55002 1896
rect 57330 1884 57336 1896
rect 54996 1856 57336 1884
rect 54996 1844 55002 1856
rect 57330 1844 57336 1856
rect 57388 1844 57394 1896
rect 57425 1887 57483 1893
rect 57425 1853 57437 1887
rect 57471 1853 57483 1887
rect 57425 1847 57483 1853
rect 57440 1816 57468 1847
rect 57974 1844 57980 1896
rect 58032 1884 58038 1896
rect 59556 1884 59584 1915
rect 60366 1912 60372 1964
rect 60424 1952 60430 1964
rect 60553 1955 60611 1961
rect 60553 1952 60565 1955
rect 60424 1924 60565 1952
rect 60424 1912 60430 1924
rect 60553 1921 60565 1924
rect 60599 1921 60611 1955
rect 60553 1915 60611 1921
rect 58032 1856 59584 1884
rect 58032 1844 58038 1856
rect 59906 1844 59912 1896
rect 59964 1884 59970 1896
rect 60660 1884 60688 1992
rect 61657 1989 61669 2023
rect 61703 2020 61715 2023
rect 61746 2020 61752 2032
rect 61703 1992 61752 2020
rect 61703 1989 61715 1992
rect 61657 1983 61715 1989
rect 60734 1912 60740 1964
rect 60792 1952 60798 1964
rect 61289 1955 61347 1961
rect 60792 1924 61148 1952
rect 60792 1912 60798 1924
rect 59964 1856 60688 1884
rect 60921 1887 60979 1893
rect 59964 1844 59970 1856
rect 60921 1853 60933 1887
rect 60967 1884 60979 1887
rect 61010 1884 61016 1896
rect 60967 1856 61016 1884
rect 60967 1853 60979 1856
rect 60921 1847 60979 1853
rect 61010 1844 61016 1856
rect 61068 1844 61074 1896
rect 61120 1884 61148 1924
rect 61289 1921 61301 1955
rect 61335 1952 61347 1955
rect 61562 1952 61568 1964
rect 61335 1924 61568 1952
rect 61335 1921 61347 1924
rect 61289 1915 61347 1921
rect 61562 1912 61568 1924
rect 61620 1912 61626 1964
rect 61672 1884 61700 1983
rect 61746 1980 61752 1992
rect 61804 1980 61810 2032
rect 63678 2020 63684 2032
rect 63591 1992 63684 2020
rect 63678 1980 63684 1992
rect 63736 2020 63742 2032
rect 65334 2020 65340 2032
rect 63736 1992 65340 2020
rect 63736 1980 63742 1992
rect 65334 1980 65340 1992
rect 65392 1980 65398 2032
rect 65426 1980 65432 2032
rect 65484 2020 65490 2032
rect 67836 2020 67864 2060
rect 69216 2020 69244 2060
rect 69290 2048 69296 2100
rect 69348 2088 69354 2100
rect 70029 2091 70087 2097
rect 70029 2088 70041 2091
rect 69348 2060 70041 2088
rect 69348 2048 69354 2060
rect 70029 2057 70041 2060
rect 70075 2057 70087 2091
rect 71038 2088 71044 2100
rect 70999 2060 71044 2088
rect 70029 2051 70087 2057
rect 71038 2048 71044 2060
rect 71096 2048 71102 2100
rect 73246 2048 73252 2100
rect 73304 2088 73310 2100
rect 73525 2091 73583 2097
rect 73525 2088 73537 2091
rect 73304 2060 73537 2088
rect 73304 2048 73310 2060
rect 73525 2057 73537 2060
rect 73571 2057 73583 2091
rect 73525 2051 73583 2057
rect 73706 2048 73712 2100
rect 73764 2048 73770 2100
rect 77570 2088 77576 2100
rect 77531 2060 77576 2088
rect 77570 2048 77576 2060
rect 77628 2048 77634 2100
rect 78030 2088 78036 2100
rect 77991 2060 78036 2088
rect 78030 2048 78036 2060
rect 78088 2048 78094 2100
rect 79134 2088 79140 2100
rect 79095 2060 79140 2088
rect 79134 2048 79140 2060
rect 79192 2048 79198 2100
rect 79318 2048 79324 2100
rect 79376 2088 79382 2100
rect 79505 2091 79563 2097
rect 79505 2088 79517 2091
rect 79376 2060 79517 2088
rect 79376 2048 79382 2060
rect 79505 2057 79517 2060
rect 79551 2057 79563 2091
rect 79505 2051 79563 2057
rect 80882 2048 80888 2100
rect 80940 2088 80946 2100
rect 81342 2088 81348 2100
rect 80940 2060 81348 2088
rect 80940 2048 80946 2060
rect 81342 2048 81348 2060
rect 81400 2048 81406 2100
rect 82265 2091 82323 2097
rect 82265 2057 82277 2091
rect 82311 2088 82323 2091
rect 82814 2088 82820 2100
rect 82311 2060 82820 2088
rect 82311 2057 82323 2060
rect 82265 2051 82323 2057
rect 82814 2048 82820 2060
rect 82872 2048 82878 2100
rect 83090 2088 83096 2100
rect 83051 2060 83096 2088
rect 83090 2048 83096 2060
rect 83148 2048 83154 2100
rect 84746 2088 84752 2100
rect 84707 2060 84752 2088
rect 84746 2048 84752 2060
rect 84804 2048 84810 2100
rect 85758 2088 85764 2100
rect 85719 2060 85764 2088
rect 85758 2048 85764 2060
rect 85816 2048 85822 2100
rect 88886 2088 88892 2100
rect 88847 2060 88892 2088
rect 88886 2048 88892 2060
rect 88944 2048 88950 2100
rect 102318 2048 102324 2100
rect 102376 2088 102382 2100
rect 103241 2091 103299 2097
rect 103241 2088 103253 2091
rect 102376 2060 103253 2088
rect 102376 2048 102382 2060
rect 103241 2057 103253 2060
rect 103287 2088 103299 2091
rect 103330 2088 103336 2100
rect 103287 2060 103336 2088
rect 103287 2057 103299 2060
rect 103241 2051 103299 2057
rect 103330 2048 103336 2060
rect 103388 2048 103394 2100
rect 106550 2088 106556 2100
rect 106511 2060 106556 2088
rect 106550 2048 106556 2060
rect 106608 2048 106614 2100
rect 107010 2048 107016 2100
rect 107068 2088 107074 2100
rect 107841 2091 107899 2097
rect 107841 2088 107853 2091
rect 107068 2060 107853 2088
rect 107068 2048 107074 2060
rect 107841 2057 107853 2060
rect 107887 2057 107899 2091
rect 107841 2051 107899 2057
rect 108114 2048 108120 2100
rect 108172 2088 108178 2100
rect 130841 2091 130899 2097
rect 108172 2060 130792 2088
rect 108172 2048 108178 2060
rect 72878 2020 72884 2032
rect 65484 1992 67864 2020
rect 67928 1992 68600 2020
rect 69216 1992 72884 2020
rect 65484 1980 65490 1992
rect 62482 1912 62488 1964
rect 62540 1952 62546 1964
rect 62850 1952 62856 1964
rect 62540 1924 62585 1952
rect 62811 1924 62856 1952
rect 62540 1912 62546 1924
rect 62850 1912 62856 1924
rect 62908 1912 62914 1964
rect 63494 1912 63500 1964
rect 63552 1952 63558 1964
rect 63773 1955 63831 1961
rect 63773 1952 63785 1955
rect 63552 1924 63785 1952
rect 63552 1912 63558 1924
rect 63773 1921 63785 1924
rect 63819 1952 63831 1955
rect 64233 1955 64291 1961
rect 64233 1952 64245 1955
rect 63819 1924 64245 1952
rect 63819 1921 63831 1924
rect 63773 1915 63831 1921
rect 64233 1921 64245 1924
rect 64279 1921 64291 1955
rect 64233 1915 64291 1921
rect 65061 1955 65119 1961
rect 65061 1921 65073 1955
rect 65107 1952 65119 1955
rect 65610 1952 65616 1964
rect 65107 1924 65616 1952
rect 65107 1921 65119 1924
rect 65061 1915 65119 1921
rect 65610 1912 65616 1924
rect 65668 1912 65674 1964
rect 66717 1955 66775 1961
rect 66717 1921 66729 1955
rect 66763 1952 66775 1955
rect 67358 1952 67364 1964
rect 66763 1924 67364 1952
rect 66763 1921 66775 1924
rect 66717 1915 66775 1921
rect 67358 1912 67364 1924
rect 67416 1912 67422 1964
rect 62577 1887 62635 1893
rect 61120 1856 61700 1884
rect 61856 1856 62436 1884
rect 51868 1788 53236 1816
rect 53392 1788 57468 1816
rect 51868 1776 51874 1788
rect 50764 1720 50936 1748
rect 50764 1708 50770 1720
rect 51258 1708 51264 1760
rect 51316 1748 51322 1760
rect 53392 1748 53420 1788
rect 57698 1776 57704 1828
rect 57756 1816 57762 1828
rect 61856 1816 61884 1856
rect 57756 1788 61884 1816
rect 57756 1776 57762 1788
rect 62206 1776 62212 1828
rect 62264 1816 62270 1828
rect 62408 1816 62436 1856
rect 62577 1853 62589 1887
rect 62623 1884 62635 1887
rect 62666 1884 62672 1896
rect 62623 1856 62672 1884
rect 62623 1853 62635 1856
rect 62577 1847 62635 1853
rect 62666 1844 62672 1856
rect 62724 1844 62730 1896
rect 63034 1844 63040 1896
rect 63092 1884 63098 1896
rect 64598 1884 64604 1896
rect 63092 1856 64604 1884
rect 63092 1844 63098 1856
rect 64598 1844 64604 1856
rect 64656 1844 64662 1896
rect 66806 1844 66812 1896
rect 66864 1884 66870 1896
rect 67928 1884 67956 1992
rect 68094 1952 68100 1964
rect 68055 1924 68100 1952
rect 68094 1912 68100 1924
rect 68152 1912 68158 1964
rect 68572 1961 68600 1992
rect 72878 1980 72884 1992
rect 72936 1980 72942 2032
rect 72970 1980 72976 2032
rect 73028 2020 73034 2032
rect 73065 2023 73123 2029
rect 73065 2020 73077 2023
rect 73028 1992 73077 2020
rect 73028 1980 73034 1992
rect 73065 1989 73077 1992
rect 73111 2020 73123 2023
rect 73724 2020 73752 2048
rect 73111 1992 73752 2020
rect 73111 1989 73123 1992
rect 73065 1983 73123 1989
rect 73890 1980 73896 2032
rect 73948 2020 73954 2032
rect 88610 2020 88616 2032
rect 73948 1992 88616 2020
rect 73948 1980 73954 1992
rect 88610 1980 88616 1992
rect 88668 1980 88674 2032
rect 100662 1980 100668 2032
rect 100720 2020 100726 2032
rect 100720 1992 104756 2020
rect 100720 1980 100726 1992
rect 68557 1955 68615 1961
rect 68557 1921 68569 1955
rect 68603 1952 68615 1955
rect 68833 1955 68891 1961
rect 68833 1952 68845 1955
rect 68603 1924 68845 1952
rect 68603 1921 68615 1924
rect 68557 1915 68615 1921
rect 68833 1921 68845 1924
rect 68879 1921 68891 1955
rect 68833 1915 68891 1921
rect 69937 1955 69995 1961
rect 69937 1921 69949 1955
rect 69983 1952 69995 1955
rect 70302 1952 70308 1964
rect 69983 1924 70308 1952
rect 69983 1921 69995 1924
rect 69937 1915 69995 1921
rect 70302 1912 70308 1924
rect 70360 1912 70366 1964
rect 70946 1952 70952 1964
rect 70907 1924 70952 1952
rect 70946 1912 70952 1924
rect 71004 1912 71010 1964
rect 72329 1955 72387 1961
rect 72329 1921 72341 1955
rect 72375 1952 72387 1955
rect 72510 1952 72516 1964
rect 72375 1924 72516 1952
rect 72375 1921 72387 1924
rect 72329 1915 72387 1921
rect 72510 1912 72516 1924
rect 72568 1912 72574 1964
rect 73433 1955 73491 1961
rect 73433 1921 73445 1955
rect 73479 1952 73491 1955
rect 73709 1955 73767 1961
rect 73709 1952 73721 1955
rect 73479 1924 73721 1952
rect 73479 1921 73491 1924
rect 73433 1915 73491 1921
rect 73709 1921 73721 1924
rect 73755 1921 73767 1955
rect 73709 1915 73767 1921
rect 73801 1955 73859 1961
rect 73801 1921 73813 1955
rect 73847 1952 73859 1955
rect 73847 1924 74396 1952
rect 73847 1921 73859 1924
rect 73801 1915 73859 1921
rect 66864 1856 67956 1884
rect 68189 1887 68247 1893
rect 66864 1844 66870 1856
rect 68189 1853 68201 1887
rect 68235 1884 68247 1887
rect 69198 1884 69204 1896
rect 68235 1856 69204 1884
rect 68235 1853 68247 1856
rect 68189 1847 68247 1853
rect 69198 1844 69204 1856
rect 69256 1844 69262 1896
rect 72418 1884 72424 1896
rect 71332 1856 71728 1884
rect 72379 1856 72424 1884
rect 71332 1816 71360 1856
rect 62264 1788 62344 1816
rect 62408 1788 71360 1816
rect 71700 1816 71728 1856
rect 72418 1844 72424 1856
rect 72476 1844 72482 1896
rect 73801 1819 73859 1825
rect 73801 1816 73813 1819
rect 71700 1788 73813 1816
rect 62264 1776 62270 1788
rect 51316 1720 53420 1748
rect 51316 1708 51322 1720
rect 53650 1708 53656 1760
rect 53708 1748 53714 1760
rect 55398 1748 55404 1760
rect 53708 1720 55404 1748
rect 53708 1708 53714 1720
rect 55398 1708 55404 1720
rect 55456 1708 55462 1760
rect 55582 1748 55588 1760
rect 55543 1720 55588 1748
rect 55582 1708 55588 1720
rect 55640 1708 55646 1760
rect 56134 1708 56140 1760
rect 56192 1748 56198 1760
rect 56502 1748 56508 1760
rect 56192 1720 56508 1748
rect 56192 1708 56198 1720
rect 56502 1708 56508 1720
rect 56560 1708 56566 1760
rect 56962 1708 56968 1760
rect 57020 1748 57026 1760
rect 57149 1751 57207 1757
rect 57149 1748 57161 1751
rect 57020 1720 57161 1748
rect 57020 1708 57026 1720
rect 57149 1717 57161 1720
rect 57195 1717 57207 1751
rect 57149 1711 57207 1717
rect 57790 1708 57796 1760
rect 57848 1748 57854 1760
rect 59081 1751 59139 1757
rect 59081 1748 59093 1751
rect 57848 1720 59093 1748
rect 57848 1708 57854 1720
rect 59081 1717 59093 1720
rect 59127 1717 59139 1751
rect 59081 1711 59139 1717
rect 60090 1708 60096 1760
rect 60148 1748 60154 1760
rect 62114 1748 62120 1760
rect 60148 1720 62120 1748
rect 60148 1708 60154 1720
rect 62114 1708 62120 1720
rect 62172 1708 62178 1760
rect 62316 1748 62344 1788
rect 73801 1785 73813 1788
rect 73847 1785 73859 1819
rect 74368 1816 74396 1924
rect 74626 1912 74632 1964
rect 74684 1952 74690 1964
rect 75638 1952 75644 1964
rect 74684 1924 75644 1952
rect 74684 1912 74690 1924
rect 75638 1912 75644 1924
rect 75696 1912 75702 1964
rect 76653 1955 76711 1961
rect 76653 1921 76665 1955
rect 76699 1921 76711 1955
rect 76653 1915 76711 1921
rect 77481 1955 77539 1961
rect 77481 1921 77493 1955
rect 77527 1952 77539 1955
rect 78582 1952 78588 1964
rect 77527 1924 78588 1952
rect 77527 1921 77539 1924
rect 77481 1915 77539 1921
rect 75086 1884 75092 1896
rect 75047 1856 75092 1884
rect 75086 1844 75092 1856
rect 75144 1844 75150 1896
rect 75914 1844 75920 1896
rect 75972 1884 75978 1896
rect 76101 1887 76159 1893
rect 76101 1884 76113 1887
rect 75972 1856 76113 1884
rect 75972 1844 75978 1856
rect 76101 1853 76113 1856
rect 76147 1853 76159 1887
rect 76668 1884 76696 1915
rect 78582 1912 78588 1924
rect 78640 1912 78646 1964
rect 79042 1952 79048 1964
rect 79003 1924 79048 1952
rect 79042 1912 79048 1924
rect 79100 1912 79106 1964
rect 80425 1955 80483 1961
rect 80425 1921 80437 1955
rect 80471 1952 80483 1955
rect 80885 1955 80943 1961
rect 80471 1924 80836 1952
rect 80471 1921 80483 1924
rect 80425 1915 80483 1921
rect 77021 1887 77079 1893
rect 77021 1884 77033 1887
rect 76668 1856 77033 1884
rect 76101 1847 76159 1853
rect 77021 1853 77033 1856
rect 77067 1884 77079 1887
rect 80808 1884 80836 1924
rect 80885 1921 80897 1955
rect 80931 1952 80943 1955
rect 81342 1952 81348 1964
rect 80931 1924 81204 1952
rect 81303 1924 81348 1952
rect 80931 1921 80943 1924
rect 80885 1915 80943 1921
rect 80977 1887 81035 1893
rect 77067 1856 80560 1884
rect 80808 1856 80928 1884
rect 77067 1853 77079 1856
rect 77021 1847 77079 1853
rect 80425 1819 80483 1825
rect 80425 1816 80437 1819
rect 74368 1788 80437 1816
rect 73801 1779 73859 1785
rect 80425 1785 80437 1788
rect 80471 1785 80483 1819
rect 80532 1816 80560 1856
rect 80900 1816 80928 1856
rect 80977 1853 80989 1887
rect 81023 1884 81035 1887
rect 81066 1884 81072 1896
rect 81023 1856 81072 1884
rect 81023 1853 81035 1856
rect 80977 1847 81035 1853
rect 81066 1844 81072 1856
rect 81124 1844 81130 1896
rect 81176 1884 81204 1924
rect 81342 1912 81348 1924
rect 81400 1912 81406 1964
rect 82170 1952 82176 1964
rect 82131 1924 82176 1952
rect 82170 1912 82176 1924
rect 82228 1912 82234 1964
rect 83369 1955 83427 1961
rect 83369 1921 83381 1955
rect 83415 1952 83427 1955
rect 83645 1955 83703 1961
rect 83645 1952 83657 1955
rect 83415 1924 83657 1952
rect 83415 1921 83427 1924
rect 83369 1915 83427 1921
rect 83645 1921 83657 1924
rect 83691 1921 83703 1955
rect 84654 1952 84660 1964
rect 84615 1924 84660 1952
rect 83645 1915 83703 1921
rect 84654 1912 84660 1924
rect 84712 1912 84718 1964
rect 85666 1952 85672 1964
rect 85627 1924 85672 1952
rect 85666 1912 85672 1924
rect 85724 1912 85730 1964
rect 86310 1912 86316 1964
rect 86368 1952 86374 1964
rect 86865 1955 86923 1961
rect 86865 1952 86877 1955
rect 86368 1924 86877 1952
rect 86368 1912 86374 1924
rect 86865 1921 86877 1924
rect 86911 1952 86923 1955
rect 87230 1952 87236 1964
rect 86911 1924 87236 1952
rect 86911 1921 86923 1924
rect 86865 1915 86923 1921
rect 87230 1912 87236 1924
rect 87288 1912 87294 1964
rect 88245 1955 88303 1961
rect 88245 1921 88257 1955
rect 88291 1952 88303 1955
rect 88426 1952 88432 1964
rect 88291 1924 88432 1952
rect 88291 1921 88303 1924
rect 88245 1915 88303 1921
rect 88426 1912 88432 1924
rect 88484 1952 88490 1964
rect 89254 1952 89260 1964
rect 88484 1924 89260 1952
rect 88484 1912 88490 1924
rect 89254 1912 89260 1924
rect 89312 1912 89318 1964
rect 91922 1952 91928 1964
rect 91883 1924 91928 1952
rect 91922 1912 91928 1924
rect 91980 1912 91986 1964
rect 102321 1955 102379 1961
rect 102321 1921 102333 1955
rect 102367 1952 102379 1955
rect 103701 1955 103759 1961
rect 102367 1924 102456 1952
rect 102367 1921 102379 1924
rect 102321 1915 102379 1921
rect 81250 1884 81256 1896
rect 81176 1856 81256 1884
rect 81250 1844 81256 1856
rect 81308 1844 81314 1896
rect 83458 1884 83464 1896
rect 83419 1856 83464 1884
rect 83458 1844 83464 1856
rect 83516 1844 83522 1896
rect 84381 1887 84439 1893
rect 84381 1853 84393 1887
rect 84427 1884 84439 1887
rect 84562 1884 84568 1896
rect 84427 1856 84568 1884
rect 84427 1853 84439 1856
rect 84381 1847 84439 1853
rect 84562 1844 84568 1856
rect 84620 1884 84626 1896
rect 86681 1887 86739 1893
rect 86681 1884 86693 1887
rect 84620 1856 86693 1884
rect 84620 1844 84626 1856
rect 86681 1853 86693 1856
rect 86727 1853 86739 1887
rect 90361 1887 90419 1893
rect 86681 1847 86739 1853
rect 86880 1856 88288 1884
rect 86880 1816 86908 1856
rect 88150 1816 88156 1828
rect 80532 1788 80652 1816
rect 80900 1788 86908 1816
rect 88111 1788 88156 1816
rect 80425 1779 80483 1785
rect 66622 1748 66628 1760
rect 62316 1720 66628 1748
rect 66622 1708 66628 1720
rect 66680 1708 66686 1760
rect 66714 1708 66720 1760
rect 66772 1748 66778 1760
rect 67266 1748 67272 1760
rect 66772 1720 67272 1748
rect 66772 1708 66778 1720
rect 67266 1708 67272 1720
rect 67324 1748 67330 1760
rect 67637 1751 67695 1757
rect 67637 1748 67649 1751
rect 67324 1720 67649 1748
rect 67324 1708 67330 1720
rect 67637 1717 67649 1720
rect 67683 1717 67695 1751
rect 67637 1711 67695 1717
rect 67726 1708 67732 1760
rect 67784 1748 67790 1760
rect 70026 1748 70032 1760
rect 67784 1720 70032 1748
rect 67784 1708 67790 1720
rect 70026 1708 70032 1720
rect 70084 1708 70090 1760
rect 71498 1708 71504 1760
rect 71556 1748 71562 1760
rect 71685 1751 71743 1757
rect 71685 1748 71697 1751
rect 71556 1720 71697 1748
rect 71556 1708 71562 1720
rect 71685 1717 71697 1720
rect 71731 1748 71743 1751
rect 73614 1748 73620 1760
rect 71731 1720 73620 1748
rect 71731 1717 71743 1720
rect 71685 1711 71743 1717
rect 73614 1708 73620 1720
rect 73672 1708 73678 1760
rect 73709 1751 73767 1757
rect 73709 1717 73721 1751
rect 73755 1748 73767 1751
rect 73985 1751 74043 1757
rect 73985 1748 73997 1751
rect 73755 1720 73997 1748
rect 73755 1717 73767 1720
rect 73709 1711 73767 1717
rect 73985 1717 73997 1720
rect 74031 1748 74043 1751
rect 74166 1748 74172 1760
rect 74031 1720 74172 1748
rect 74031 1717 74043 1720
rect 73985 1711 74043 1717
rect 74166 1708 74172 1720
rect 74224 1708 74230 1760
rect 74258 1708 74264 1760
rect 74316 1748 74322 1760
rect 80514 1748 80520 1760
rect 74316 1720 80520 1748
rect 74316 1708 74322 1720
rect 80514 1708 80520 1720
rect 80572 1708 80578 1760
rect 80624 1748 80652 1788
rect 88150 1776 88156 1788
rect 88208 1776 88214 1828
rect 88260 1816 88288 1856
rect 90361 1853 90373 1887
rect 90407 1884 90419 1887
rect 91278 1884 91284 1896
rect 90407 1856 91284 1884
rect 90407 1853 90419 1856
rect 90361 1847 90419 1853
rect 91278 1844 91284 1856
rect 91336 1844 91342 1896
rect 91373 1887 91431 1893
rect 91373 1853 91385 1887
rect 91419 1853 91431 1887
rect 91373 1847 91431 1853
rect 91388 1816 91416 1847
rect 88260 1788 91416 1816
rect 95142 1776 95148 1828
rect 95200 1816 95206 1828
rect 96614 1816 96620 1828
rect 95200 1788 96620 1816
rect 95200 1776 95206 1788
rect 96614 1776 96620 1788
rect 96672 1776 96678 1828
rect 97718 1776 97724 1828
rect 97776 1816 97782 1828
rect 102428 1816 102456 1924
rect 103701 1921 103713 1955
rect 103747 1952 103759 1955
rect 104342 1952 104348 1964
rect 103747 1924 104348 1952
rect 103747 1921 103759 1924
rect 103701 1915 103759 1921
rect 104342 1912 104348 1924
rect 104400 1912 104406 1964
rect 104728 1893 104756 1992
rect 104894 1980 104900 2032
rect 104952 2020 104958 2032
rect 117774 2020 117780 2032
rect 104952 1992 114876 2020
rect 117735 1992 117780 2020
rect 104952 1980 104958 1992
rect 105262 1952 105268 1964
rect 105223 1924 105268 1952
rect 105262 1912 105268 1924
rect 105320 1912 105326 1964
rect 106461 1955 106519 1961
rect 106461 1921 106473 1955
rect 106507 1952 106519 1955
rect 106918 1952 106924 1964
rect 106507 1924 106924 1952
rect 106507 1921 106519 1924
rect 106461 1915 106519 1921
rect 106918 1912 106924 1924
rect 106976 1912 106982 1964
rect 107746 1952 107752 1964
rect 107707 1924 107752 1952
rect 107746 1912 107752 1924
rect 107804 1912 107810 1964
rect 108761 1955 108819 1961
rect 108761 1921 108773 1955
rect 108807 1952 108819 1955
rect 109034 1952 109040 1964
rect 108807 1924 109040 1952
rect 108807 1921 108819 1924
rect 108761 1915 108819 1921
rect 109034 1912 109040 1924
rect 109092 1912 109098 1964
rect 109586 1912 109592 1964
rect 109644 1952 109650 1964
rect 111058 1952 111064 1964
rect 109644 1924 111064 1952
rect 109644 1912 109650 1924
rect 111058 1912 111064 1924
rect 111116 1912 111122 1964
rect 111334 1952 111340 1964
rect 111295 1924 111340 1952
rect 111334 1912 111340 1924
rect 111392 1912 111398 1964
rect 112162 1952 112168 1964
rect 112123 1924 112168 1952
rect 112162 1912 112168 1924
rect 112220 1952 112226 1964
rect 112625 1955 112683 1961
rect 112625 1952 112637 1955
rect 112220 1924 112637 1952
rect 112220 1912 112226 1924
rect 112625 1921 112637 1924
rect 112671 1921 112683 1955
rect 112625 1915 112683 1921
rect 112898 1912 112904 1964
rect 112956 1952 112962 1964
rect 112956 1924 114692 1952
rect 112956 1912 112962 1924
rect 104713 1887 104771 1893
rect 104713 1853 104725 1887
rect 104759 1853 104771 1887
rect 104713 1847 104771 1853
rect 104802 1844 104808 1896
rect 104860 1884 104866 1896
rect 108574 1884 108580 1896
rect 104860 1856 108580 1884
rect 104860 1844 104866 1856
rect 108574 1844 108580 1856
rect 108632 1844 108638 1896
rect 108666 1844 108672 1896
rect 108724 1884 108730 1896
rect 108853 1887 108911 1893
rect 108853 1884 108865 1887
rect 108724 1856 108865 1884
rect 108724 1844 108730 1856
rect 108853 1853 108865 1856
rect 108899 1853 108911 1887
rect 109770 1884 109776 1896
rect 109731 1856 109776 1884
rect 108853 1847 108911 1853
rect 109770 1844 109776 1856
rect 109828 1844 109834 1896
rect 110690 1844 110696 1896
rect 110748 1884 110754 1896
rect 110785 1887 110843 1893
rect 110785 1884 110797 1887
rect 110748 1856 110797 1884
rect 110748 1844 110754 1856
rect 110785 1853 110797 1856
rect 110831 1853 110843 1887
rect 110785 1847 110843 1853
rect 111242 1844 111248 1896
rect 111300 1884 111306 1896
rect 112070 1884 112076 1896
rect 111300 1856 112076 1884
rect 111300 1844 111306 1856
rect 112070 1844 112076 1856
rect 112128 1844 112134 1896
rect 112254 1844 112260 1896
rect 112312 1884 112318 1896
rect 113450 1884 113456 1896
rect 112312 1856 113456 1884
rect 112312 1844 112318 1856
rect 113450 1844 113456 1856
rect 113508 1844 113514 1896
rect 113818 1884 113824 1896
rect 113779 1856 113824 1884
rect 113818 1844 113824 1856
rect 113876 1844 113882 1896
rect 102781 1819 102839 1825
rect 102781 1816 102793 1819
rect 97776 1788 102793 1816
rect 97776 1776 97782 1788
rect 102781 1785 102793 1788
rect 102827 1785 102839 1819
rect 114664 1816 114692 1924
rect 114848 1893 114876 1992
rect 117774 1980 117780 1992
rect 117832 1980 117838 2032
rect 117866 1980 117872 2032
rect 117924 2020 117930 2032
rect 118329 2023 118387 2029
rect 118329 2020 118341 2023
rect 117924 1992 118341 2020
rect 117924 1980 117930 1992
rect 118329 1989 118341 1992
rect 118375 1989 118387 2023
rect 118329 1983 118387 1989
rect 118786 1980 118792 2032
rect 118844 2020 118850 2032
rect 119065 2023 119123 2029
rect 119065 2020 119077 2023
rect 118844 1992 119077 2020
rect 118844 1980 118850 1992
rect 119065 1989 119077 1992
rect 119111 1989 119123 2023
rect 119065 1983 119123 1989
rect 119154 1980 119160 2032
rect 119212 2020 119218 2032
rect 120534 2020 120540 2032
rect 119212 1992 120540 2020
rect 119212 1980 119218 1992
rect 120534 1980 120540 1992
rect 120592 1980 120598 2032
rect 120626 1980 120632 2032
rect 120684 2020 120690 2032
rect 121089 2023 121147 2029
rect 121089 2020 121101 2023
rect 120684 1992 121101 2020
rect 120684 1980 120690 1992
rect 121089 1989 121101 1992
rect 121135 1989 121147 2023
rect 121089 1983 121147 1989
rect 121178 1980 121184 2032
rect 121236 2020 121242 2032
rect 122926 2020 122932 2032
rect 121236 1992 122512 2020
rect 122887 1992 122932 2020
rect 121236 1980 121242 1992
rect 115385 1955 115443 1961
rect 115385 1921 115397 1955
rect 115431 1952 115443 1955
rect 115566 1952 115572 1964
rect 115431 1924 115572 1952
rect 115431 1921 115443 1924
rect 115385 1915 115443 1921
rect 115566 1912 115572 1924
rect 115624 1912 115630 1964
rect 116210 1952 116216 1964
rect 116171 1924 116216 1952
rect 116210 1912 116216 1924
rect 116268 1912 116274 1964
rect 117682 1952 117688 1964
rect 117643 1924 117688 1952
rect 117682 1912 117688 1924
rect 117740 1912 117746 1964
rect 118602 1952 118608 1964
rect 117792 1924 118608 1952
rect 114833 1887 114891 1893
rect 114833 1853 114845 1887
rect 114879 1853 114891 1887
rect 116305 1887 116363 1893
rect 116305 1884 116317 1887
rect 114833 1847 114891 1853
rect 114940 1856 116317 1884
rect 114940 1816 114968 1856
rect 116305 1853 116317 1856
rect 116351 1853 116363 1887
rect 116305 1847 116363 1853
rect 116762 1844 116768 1896
rect 116820 1884 116826 1896
rect 117792 1884 117820 1924
rect 118602 1912 118608 1924
rect 118660 1912 118666 1964
rect 118973 1955 119031 1961
rect 118973 1921 118985 1955
rect 119019 1952 119031 1955
rect 119985 1955 120043 1961
rect 119019 1924 119568 1952
rect 119019 1921 119031 1924
rect 118973 1915 119031 1921
rect 119540 1893 119568 1924
rect 119985 1921 119997 1955
rect 120031 1952 120043 1955
rect 120166 1952 120172 1964
rect 120031 1924 120172 1952
rect 120031 1921 120043 1924
rect 119985 1915 120043 1921
rect 120166 1912 120172 1924
rect 120224 1912 120230 1964
rect 120994 1952 121000 1964
rect 120907 1924 121000 1952
rect 120994 1912 121000 1924
rect 121052 1952 121058 1964
rect 122374 1952 122380 1964
rect 121052 1924 122380 1952
rect 121052 1912 121058 1924
rect 122374 1912 122380 1924
rect 122432 1912 122438 1964
rect 116820 1856 117820 1884
rect 119525 1887 119583 1893
rect 116820 1844 116826 1856
rect 119525 1853 119537 1887
rect 119571 1884 119583 1887
rect 122006 1884 122012 1896
rect 119571 1856 122012 1884
rect 119571 1853 119583 1856
rect 119525 1847 119583 1853
rect 122006 1844 122012 1856
rect 122064 1844 122070 1896
rect 122484 1884 122512 1992
rect 122926 1980 122932 1992
rect 122984 1980 122990 2032
rect 124674 2020 124680 2032
rect 124635 1992 124680 2020
rect 124674 1980 124680 1992
rect 124732 1980 124738 2032
rect 125594 1980 125600 2032
rect 125652 2020 125658 2032
rect 126790 2020 126796 2032
rect 125652 1992 126796 2020
rect 125652 1980 125658 1992
rect 126790 1980 126796 1992
rect 126848 1980 126854 2032
rect 130654 2020 130660 2032
rect 126900 1992 130660 2020
rect 122834 1952 122840 1964
rect 122795 1924 122840 1952
rect 122834 1912 122840 1924
rect 122892 1912 122898 1964
rect 124585 1955 124643 1961
rect 124585 1921 124597 1955
rect 124631 1952 124643 1955
rect 124861 1955 124919 1961
rect 124861 1952 124873 1955
rect 124631 1924 124873 1952
rect 124631 1921 124643 1924
rect 124585 1915 124643 1921
rect 124861 1921 124873 1924
rect 124907 1921 124919 1955
rect 126900 1952 126928 1992
rect 130654 1980 130660 1992
rect 130712 1980 130718 2032
rect 130764 2020 130792 2060
rect 130841 2057 130853 2091
rect 130887 2088 130899 2091
rect 130930 2088 130936 2100
rect 130887 2060 130936 2088
rect 130887 2057 130899 2060
rect 130841 2051 130899 2057
rect 130930 2048 130936 2060
rect 130988 2048 130994 2100
rect 138658 2048 138664 2100
rect 138716 2088 138722 2100
rect 139029 2091 139087 2097
rect 139029 2088 139041 2091
rect 138716 2060 139041 2088
rect 138716 2048 138722 2060
rect 139029 2057 139041 2060
rect 139075 2088 139087 2091
rect 139394 2088 139400 2100
rect 139075 2060 139400 2088
rect 139075 2057 139087 2060
rect 139029 2051 139087 2057
rect 139394 2048 139400 2060
rect 139452 2048 139458 2100
rect 139578 2088 139584 2100
rect 139539 2060 139584 2088
rect 139578 2048 139584 2060
rect 139636 2048 139642 2100
rect 141142 2088 141148 2100
rect 141103 2060 141148 2088
rect 141142 2048 141148 2060
rect 141200 2048 141206 2100
rect 146021 2091 146079 2097
rect 146021 2057 146033 2091
rect 146067 2088 146079 2091
rect 146386 2088 146392 2100
rect 146067 2060 146392 2088
rect 146067 2057 146079 2060
rect 146021 2051 146079 2057
rect 146386 2048 146392 2060
rect 146444 2048 146450 2100
rect 150345 2091 150403 2097
rect 150345 2057 150357 2091
rect 150391 2088 150403 2091
rect 150986 2088 150992 2100
rect 150391 2060 150992 2088
rect 150391 2057 150403 2060
rect 150345 2051 150403 2057
rect 150986 2048 150992 2060
rect 151044 2048 151050 2100
rect 153746 2088 153752 2100
rect 153707 2060 153752 2088
rect 153746 2048 153752 2060
rect 153804 2048 153810 2100
rect 154761 2091 154819 2097
rect 154761 2057 154773 2091
rect 154807 2088 154819 2091
rect 154850 2088 154856 2100
rect 154807 2060 154856 2088
rect 154807 2057 154819 2060
rect 154761 2051 154819 2057
rect 154850 2048 154856 2060
rect 154908 2048 154914 2100
rect 155770 2088 155776 2100
rect 155731 2060 155776 2088
rect 155770 2048 155776 2060
rect 155828 2048 155834 2100
rect 160922 2088 160928 2100
rect 160883 2060 160928 2088
rect 160922 2048 160928 2060
rect 160980 2048 160986 2100
rect 162029 2091 162087 2097
rect 162029 2057 162041 2091
rect 162075 2088 162087 2091
rect 162394 2088 162400 2100
rect 162075 2060 162400 2088
rect 162075 2057 162087 2060
rect 162029 2051 162087 2057
rect 162394 2048 162400 2060
rect 162452 2048 162458 2100
rect 163961 2091 164019 2097
rect 163961 2057 163973 2091
rect 164007 2088 164019 2091
rect 164970 2088 164976 2100
rect 164007 2060 164976 2088
rect 164007 2057 164019 2060
rect 163961 2051 164019 2057
rect 164970 2048 164976 2060
rect 165028 2048 165034 2100
rect 136361 2023 136419 2029
rect 130764 1992 135484 2020
rect 127066 1952 127072 1964
rect 124861 1915 124919 1921
rect 124968 1924 126928 1952
rect 127027 1924 127072 1952
rect 124968 1884 124996 1924
rect 127066 1912 127072 1924
rect 127124 1912 127130 1964
rect 128173 1955 128231 1961
rect 128173 1921 128185 1955
rect 128219 1952 128231 1955
rect 128262 1952 128268 1964
rect 128219 1924 128268 1952
rect 128219 1921 128231 1924
rect 128173 1915 128231 1921
rect 128262 1912 128268 1924
rect 128320 1912 128326 1964
rect 130749 1955 130807 1961
rect 130749 1921 130761 1955
rect 130795 1952 130807 1955
rect 131206 1952 131212 1964
rect 130795 1924 131212 1952
rect 130795 1921 130807 1924
rect 130749 1915 130807 1921
rect 131206 1912 131212 1924
rect 131264 1912 131270 1964
rect 122484 1856 124996 1884
rect 125597 1887 125655 1893
rect 125597 1853 125609 1887
rect 125643 1884 125655 1887
rect 126146 1884 126152 1896
rect 125643 1856 126152 1884
rect 125643 1853 125655 1856
rect 125597 1847 125655 1853
rect 126146 1844 126152 1856
rect 126204 1844 126210 1896
rect 126606 1884 126612 1896
rect 126567 1856 126612 1884
rect 126606 1844 126612 1856
rect 126664 1844 126670 1896
rect 130565 1887 130623 1893
rect 126716 1856 130240 1884
rect 117774 1816 117780 1828
rect 102781 1779 102839 1785
rect 105004 1788 113864 1816
rect 114664 1788 114968 1816
rect 115032 1788 117780 1816
rect 83550 1748 83556 1760
rect 80624 1720 83556 1748
rect 83550 1708 83556 1720
rect 83608 1708 83614 1760
rect 83645 1751 83703 1757
rect 83645 1717 83657 1751
rect 83691 1748 83703 1751
rect 83921 1751 83979 1757
rect 83921 1748 83933 1751
rect 83691 1720 83933 1748
rect 83691 1717 83703 1720
rect 83645 1711 83703 1717
rect 83921 1717 83933 1720
rect 83967 1748 83979 1751
rect 85574 1748 85580 1760
rect 83967 1720 85580 1748
rect 83967 1717 83979 1720
rect 83921 1711 83979 1717
rect 85574 1708 85580 1720
rect 85632 1708 85638 1760
rect 86681 1751 86739 1757
rect 86681 1717 86693 1751
rect 86727 1748 86739 1751
rect 100018 1748 100024 1760
rect 86727 1720 100024 1748
rect 86727 1717 86739 1720
rect 86681 1711 86739 1717
rect 100018 1708 100024 1720
rect 100076 1708 100082 1760
rect 102410 1748 102416 1760
rect 102371 1720 102416 1748
rect 102410 1708 102416 1720
rect 102468 1708 102474 1760
rect 102502 1708 102508 1760
rect 102560 1748 102566 1760
rect 105004 1748 105032 1788
rect 102560 1720 105032 1748
rect 102560 1708 102566 1720
rect 106918 1708 106924 1760
rect 106976 1748 106982 1760
rect 110598 1748 110604 1760
rect 106976 1720 110604 1748
rect 106976 1708 106982 1720
rect 110598 1708 110604 1720
rect 110656 1708 110662 1760
rect 111610 1748 111616 1760
rect 111571 1720 111616 1748
rect 111610 1708 111616 1720
rect 111668 1708 111674 1760
rect 112254 1748 112260 1760
rect 112215 1720 112260 1748
rect 112254 1708 112260 1720
rect 112312 1708 112318 1760
rect 113836 1748 113864 1788
rect 115032 1748 115060 1788
rect 117774 1776 117780 1788
rect 117832 1776 117838 1828
rect 118329 1819 118387 1825
rect 118329 1785 118341 1819
rect 118375 1816 118387 1819
rect 126716 1816 126744 1856
rect 118375 1788 126744 1816
rect 128265 1819 128323 1825
rect 118375 1785 118387 1788
rect 118329 1779 118387 1785
rect 128265 1785 128277 1819
rect 128311 1816 128323 1819
rect 128538 1816 128544 1828
rect 128311 1788 128544 1816
rect 128311 1785 128323 1788
rect 128265 1779 128323 1785
rect 128538 1776 128544 1788
rect 128596 1776 128602 1828
rect 130212 1816 130240 1856
rect 130565 1853 130577 1887
rect 130611 1884 130623 1887
rect 131022 1884 131028 1896
rect 130611 1856 131028 1884
rect 130611 1853 130623 1856
rect 130565 1847 130623 1853
rect 131022 1844 131028 1856
rect 131080 1844 131086 1896
rect 133690 1884 133696 1896
rect 133651 1856 133696 1884
rect 133690 1844 133696 1856
rect 133748 1844 133754 1896
rect 134705 1887 134763 1893
rect 134705 1853 134717 1887
rect 134751 1884 134763 1887
rect 135346 1884 135352 1896
rect 134751 1856 135352 1884
rect 134751 1853 134763 1856
rect 134705 1847 134763 1853
rect 135346 1844 135352 1856
rect 135404 1844 135410 1896
rect 135456 1884 135484 1992
rect 136361 1989 136373 2023
rect 136407 2020 136419 2023
rect 138934 2020 138940 2032
rect 136407 1992 138940 2020
rect 136407 1989 136419 1992
rect 136361 1983 136419 1989
rect 135809 1955 135867 1961
rect 135809 1921 135821 1955
rect 135855 1952 135867 1955
rect 136376 1952 136404 1983
rect 138934 1980 138940 1992
rect 138992 1980 138998 2032
rect 139302 2020 139308 2032
rect 139263 1992 139308 2020
rect 139302 1980 139308 1992
rect 139360 1980 139366 2032
rect 144822 1980 144828 2032
rect 144880 2020 144886 2032
rect 152737 2023 152795 2029
rect 144880 1992 148916 2020
rect 144880 1980 144886 1992
rect 138661 1955 138719 1961
rect 135855 1924 136404 1952
rect 136468 1924 137692 1952
rect 135855 1921 135867 1924
rect 135809 1915 135867 1921
rect 136468 1884 136496 1924
rect 135456 1856 136496 1884
rect 137097 1887 137155 1893
rect 137097 1853 137109 1887
rect 137143 1884 137155 1887
rect 137278 1884 137284 1896
rect 137143 1856 137284 1884
rect 137143 1853 137155 1856
rect 137097 1847 137155 1853
rect 137278 1844 137284 1856
rect 137336 1884 137342 1896
rect 137554 1884 137560 1896
rect 137336 1856 137560 1884
rect 137336 1844 137342 1856
rect 137554 1844 137560 1856
rect 137612 1844 137618 1896
rect 137664 1884 137692 1924
rect 138661 1921 138673 1955
rect 138707 1952 138719 1955
rect 138750 1952 138756 1964
rect 138707 1924 138756 1952
rect 138707 1921 138719 1924
rect 138661 1915 138719 1921
rect 138750 1912 138756 1924
rect 138808 1912 138814 1964
rect 139486 1952 139492 1964
rect 139447 1924 139492 1952
rect 139486 1912 139492 1924
rect 139544 1912 139550 1964
rect 141421 1955 141479 1961
rect 141421 1921 141433 1955
rect 141467 1952 141479 1955
rect 141602 1952 141608 1964
rect 141467 1924 141608 1952
rect 141467 1921 141479 1924
rect 141421 1915 141479 1921
rect 141602 1912 141608 1924
rect 141660 1952 141666 1964
rect 141881 1955 141939 1961
rect 141881 1952 141893 1955
rect 141660 1924 141893 1952
rect 141660 1912 141666 1924
rect 141881 1921 141893 1924
rect 141927 1921 141939 1955
rect 144270 1952 144276 1964
rect 141881 1915 141939 1921
rect 143000 1924 143304 1952
rect 144231 1924 144276 1952
rect 138109 1887 138167 1893
rect 138109 1884 138121 1887
rect 137664 1856 138121 1884
rect 138109 1853 138121 1856
rect 138155 1853 138167 1887
rect 143000 1884 143028 1924
rect 143166 1884 143172 1896
rect 138109 1847 138167 1853
rect 138216 1856 143028 1884
rect 143127 1856 143172 1884
rect 138216 1816 138244 1856
rect 143166 1844 143172 1856
rect 143224 1844 143230 1896
rect 143276 1884 143304 1924
rect 144270 1912 144276 1924
rect 144328 1912 144334 1964
rect 145929 1955 145987 1961
rect 145929 1921 145941 1955
rect 145975 1952 145987 1955
rect 146662 1952 146668 1964
rect 145975 1924 146668 1952
rect 145975 1921 145987 1924
rect 145929 1915 145987 1921
rect 146662 1912 146668 1924
rect 146720 1912 146726 1964
rect 144181 1887 144239 1893
rect 144181 1884 144193 1887
rect 143276 1856 144193 1884
rect 144181 1853 144193 1856
rect 144227 1853 144239 1887
rect 147858 1884 147864 1896
rect 147819 1856 147864 1884
rect 144181 1847 144239 1853
rect 147858 1844 147864 1856
rect 147916 1844 147922 1896
rect 148888 1893 148916 1992
rect 152737 1989 152749 2023
rect 152783 2020 152795 2023
rect 154574 2020 154580 2032
rect 152783 1992 154580 2020
rect 152783 1989 152795 1992
rect 152737 1983 152795 1989
rect 154574 1980 154580 1992
rect 154632 1980 154638 2032
rect 149146 1952 149152 1964
rect 149107 1924 149152 1952
rect 149146 1912 149152 1924
rect 149204 1912 149210 1964
rect 150250 1952 150256 1964
rect 150211 1924 150256 1952
rect 150250 1912 150256 1924
rect 150308 1912 150314 1964
rect 152642 1952 152648 1964
rect 152603 1924 152648 1952
rect 152642 1912 152648 1924
rect 152700 1912 152706 1964
rect 153654 1952 153660 1964
rect 153615 1924 153660 1952
rect 153654 1912 153660 1924
rect 153712 1912 153718 1964
rect 154666 1952 154672 1964
rect 154627 1924 154672 1952
rect 154666 1912 154672 1924
rect 154724 1912 154730 1964
rect 155681 1955 155739 1961
rect 155681 1921 155693 1955
rect 155727 1952 155739 1955
rect 155862 1952 155868 1964
rect 155727 1924 155868 1952
rect 155727 1921 155739 1924
rect 155681 1915 155739 1921
rect 155862 1912 155868 1924
rect 155920 1912 155926 1964
rect 156690 1952 156696 1964
rect 156651 1924 156696 1952
rect 156690 1912 156696 1924
rect 156748 1952 156754 1964
rect 157153 1955 157211 1961
rect 157153 1952 157165 1955
rect 156748 1924 157165 1952
rect 156748 1912 156754 1924
rect 157153 1921 157165 1924
rect 157199 1921 157211 1955
rect 157153 1915 157211 1921
rect 158162 1912 158168 1964
rect 158220 1952 158226 1964
rect 158257 1955 158315 1961
rect 158257 1952 158269 1955
rect 158220 1924 158269 1952
rect 158220 1912 158226 1924
rect 158257 1921 158269 1924
rect 158303 1921 158315 1955
rect 159818 1952 159824 1964
rect 159779 1924 159824 1952
rect 158257 1915 158315 1921
rect 159818 1912 159824 1924
rect 159876 1912 159882 1964
rect 160830 1952 160836 1964
rect 160791 1924 160836 1952
rect 160830 1912 160836 1924
rect 160888 1912 160894 1964
rect 161934 1952 161940 1964
rect 161895 1924 161940 1952
rect 161934 1912 161940 1924
rect 161992 1912 161998 1964
rect 163869 1955 163927 1961
rect 163869 1921 163881 1955
rect 163915 1952 163927 1955
rect 163958 1952 163964 1964
rect 163915 1924 163964 1952
rect 163915 1921 163927 1924
rect 163869 1915 163927 1921
rect 163958 1912 163964 1924
rect 164016 1912 164022 1964
rect 164878 1952 164884 1964
rect 164839 1924 164884 1952
rect 164878 1912 164884 1924
rect 164936 1912 164942 1964
rect 166074 1912 166080 1964
rect 166132 1952 166138 1964
rect 166721 1955 166779 1961
rect 166721 1952 166733 1955
rect 166132 1924 166733 1952
rect 166132 1912 166138 1924
rect 166721 1921 166733 1924
rect 166767 1952 166779 1955
rect 166902 1952 166908 1964
rect 166767 1924 166908 1952
rect 166767 1921 166779 1924
rect 166721 1915 166779 1921
rect 166902 1912 166908 1924
rect 166960 1912 166966 1964
rect 148873 1887 148931 1893
rect 148873 1853 148885 1887
rect 148919 1853 148931 1887
rect 148873 1847 148931 1853
rect 165709 1887 165767 1893
rect 165709 1853 165721 1887
rect 165755 1884 165767 1887
rect 166166 1884 166172 1896
rect 165755 1856 166172 1884
rect 165755 1853 165767 1856
rect 165709 1847 165767 1853
rect 166166 1844 166172 1856
rect 166224 1844 166230 1896
rect 166534 1844 166540 1896
rect 166592 1884 166598 1896
rect 167089 1887 167147 1893
rect 167089 1884 167101 1887
rect 166592 1856 167101 1884
rect 166592 1844 166598 1856
rect 167089 1853 167101 1856
rect 167135 1853 167147 1887
rect 167089 1847 167147 1853
rect 129016 1788 129320 1816
rect 130212 1788 138244 1816
rect 113836 1720 115060 1748
rect 115106 1708 115112 1760
rect 115164 1748 115170 1760
rect 118234 1748 118240 1760
rect 115164 1720 118240 1748
rect 115164 1708 115170 1720
rect 118234 1708 118240 1720
rect 118292 1708 118298 1760
rect 118418 1748 118424 1760
rect 118379 1720 118424 1748
rect 118418 1708 118424 1720
rect 118476 1708 118482 1760
rect 118970 1708 118976 1760
rect 119028 1748 119034 1760
rect 119706 1748 119712 1760
rect 119028 1720 119712 1748
rect 119028 1708 119034 1720
rect 119706 1708 119712 1720
rect 119764 1708 119770 1760
rect 119890 1748 119896 1760
rect 119803 1720 119896 1748
rect 119890 1708 119896 1720
rect 119948 1748 119954 1760
rect 120077 1751 120135 1757
rect 120077 1748 120089 1751
rect 119948 1720 120089 1748
rect 119948 1708 119954 1720
rect 120077 1717 120089 1720
rect 120123 1717 120135 1751
rect 120077 1711 120135 1717
rect 120166 1708 120172 1760
rect 120224 1748 120230 1760
rect 120350 1748 120356 1760
rect 120224 1720 120356 1748
rect 120224 1708 120230 1720
rect 120350 1708 120356 1720
rect 120408 1748 120414 1760
rect 121178 1748 121184 1760
rect 120408 1720 121184 1748
rect 120408 1708 120414 1720
rect 121178 1708 121184 1720
rect 121236 1708 121242 1760
rect 123938 1748 123944 1760
rect 123899 1720 123944 1748
rect 123938 1708 123944 1720
rect 123996 1708 124002 1760
rect 124861 1751 124919 1757
rect 124861 1717 124873 1751
rect 124907 1748 124919 1751
rect 125137 1751 125195 1757
rect 125137 1748 125149 1751
rect 124907 1720 125149 1748
rect 124907 1717 124919 1720
rect 124861 1711 124919 1717
rect 125137 1717 125149 1720
rect 125183 1748 125195 1751
rect 126054 1748 126060 1760
rect 125183 1720 126060 1748
rect 125183 1717 125195 1720
rect 125137 1711 125195 1717
rect 126054 1708 126060 1720
rect 126112 1708 126118 1760
rect 126238 1708 126244 1760
rect 126296 1748 126302 1760
rect 129016 1748 129044 1788
rect 129182 1748 129188 1760
rect 126296 1720 129044 1748
rect 129143 1720 129188 1748
rect 126296 1708 126302 1720
rect 129182 1708 129188 1720
rect 129240 1708 129246 1760
rect 129292 1748 129320 1788
rect 132494 1748 132500 1760
rect 129292 1720 132500 1748
rect 132494 1708 132500 1720
rect 132552 1708 132558 1760
rect 133414 1708 133420 1760
rect 133472 1748 133478 1760
rect 134150 1748 134156 1760
rect 133472 1720 134156 1748
rect 133472 1708 133478 1720
rect 134150 1708 134156 1720
rect 134208 1708 134214 1760
rect 135898 1748 135904 1760
rect 135859 1720 135904 1748
rect 135898 1708 135904 1720
rect 135956 1708 135962 1760
rect 137830 1708 137836 1760
rect 137888 1748 137894 1760
rect 139486 1748 139492 1760
rect 137888 1720 139492 1748
rect 137888 1708 137894 1720
rect 139486 1708 139492 1720
rect 139544 1748 139550 1760
rect 139949 1751 140007 1757
rect 139949 1748 139961 1751
rect 139544 1720 139961 1748
rect 139544 1708 139550 1720
rect 139949 1717 139961 1720
rect 139995 1717 140007 1751
rect 139949 1711 140007 1717
rect 141050 1708 141056 1760
rect 141108 1748 141114 1760
rect 141513 1751 141571 1757
rect 141513 1748 141525 1751
rect 141108 1720 141525 1748
rect 141108 1708 141114 1720
rect 141513 1717 141525 1720
rect 141559 1717 141571 1751
rect 141513 1711 141571 1717
rect 155862 1708 155868 1760
rect 155920 1748 155926 1760
rect 156141 1751 156199 1757
rect 156141 1748 156153 1751
rect 155920 1720 156153 1748
rect 155920 1708 155926 1720
rect 156141 1717 156153 1720
rect 156187 1717 156199 1751
rect 156141 1711 156199 1717
rect 156785 1751 156843 1757
rect 156785 1717 156797 1751
rect 156831 1748 156843 1751
rect 156874 1748 156880 1760
rect 156831 1720 156880 1748
rect 156831 1717 156843 1720
rect 156785 1711 156843 1717
rect 156874 1708 156880 1720
rect 156932 1708 156938 1760
rect 158346 1748 158352 1760
rect 158307 1720 158352 1748
rect 158346 1708 158352 1720
rect 158404 1708 158410 1760
rect 158714 1748 158720 1760
rect 158675 1720 158720 1748
rect 158714 1708 158720 1720
rect 158772 1708 158778 1760
rect 159634 1748 159640 1760
rect 159547 1720 159640 1748
rect 159634 1708 159640 1720
rect 159692 1748 159698 1760
rect 159913 1751 159971 1757
rect 159913 1748 159925 1751
rect 159692 1720 159925 1748
rect 159692 1708 159698 1720
rect 159913 1717 159925 1720
rect 159959 1717 159971 1751
rect 159913 1711 159971 1717
rect 368 1658 93012 1680
rect 368 1606 28456 1658
rect 28508 1606 28520 1658
rect 28572 1606 28584 1658
rect 28636 1606 28648 1658
rect 28700 1606 84878 1658
rect 84930 1606 84942 1658
rect 84994 1606 85006 1658
rect 85058 1606 85070 1658
rect 85122 1606 93012 1658
rect 95050 1640 95056 1692
rect 95108 1680 95114 1692
rect 96982 1680 96988 1692
rect 95108 1652 96988 1680
rect 95108 1640 95114 1652
rect 96982 1640 96988 1652
rect 97040 1640 97046 1692
rect 98641 1683 98699 1689
rect 98641 1649 98653 1683
rect 98687 1680 98699 1683
rect 100294 1680 100300 1692
rect 98687 1652 100300 1680
rect 98687 1649 98699 1652
rect 98641 1643 98699 1649
rect 100294 1640 100300 1652
rect 100352 1640 100358 1692
rect 102028 1658 169556 1680
rect 368 1584 93012 1606
rect 95970 1572 95976 1624
rect 96028 1612 96034 1624
rect 99377 1615 99435 1621
rect 99377 1612 99389 1615
rect 96028 1584 99389 1612
rect 96028 1572 96034 1584
rect 99377 1581 99389 1584
rect 99423 1581 99435 1615
rect 99377 1575 99435 1581
rect 99466 1572 99472 1624
rect 99524 1612 99530 1624
rect 100110 1612 100116 1624
rect 99524 1584 100116 1612
rect 99524 1572 99530 1584
rect 100110 1572 100116 1584
rect 100168 1572 100174 1624
rect 102028 1606 141299 1658
rect 141351 1606 141363 1658
rect 141415 1606 141427 1658
rect 141479 1606 141491 1658
rect 141543 1606 169556 1658
rect 102028 1584 169556 1606
rect 2038 1504 2044 1556
rect 2096 1544 2102 1556
rect 3050 1544 3056 1556
rect 2096 1516 3056 1544
rect 2096 1504 2102 1516
rect 3050 1504 3056 1516
rect 3108 1504 3114 1556
rect 3234 1504 3240 1556
rect 3292 1544 3298 1556
rect 3789 1547 3847 1553
rect 3789 1544 3801 1547
rect 3292 1516 3801 1544
rect 3292 1504 3298 1516
rect 3789 1513 3801 1516
rect 3835 1513 3847 1547
rect 7190 1544 7196 1556
rect 7151 1516 7196 1544
rect 3789 1507 3847 1513
rect 7190 1504 7196 1516
rect 7248 1504 7254 1556
rect 9214 1544 9220 1556
rect 9175 1516 9220 1544
rect 9214 1504 9220 1516
rect 9272 1544 9278 1556
rect 10505 1547 10563 1553
rect 9272 1516 9536 1544
rect 9272 1504 9278 1516
rect 1670 1436 1676 1488
rect 1728 1476 1734 1488
rect 7466 1476 7472 1488
rect 1728 1448 7472 1476
rect 1728 1436 1734 1448
rect 7466 1436 7472 1448
rect 7524 1436 7530 1488
rect 2406 1368 2412 1420
rect 2464 1408 2470 1420
rect 9508 1417 9536 1516
rect 10505 1513 10517 1547
rect 10551 1544 10563 1547
rect 10778 1544 10784 1556
rect 10551 1516 10784 1544
rect 10551 1513 10563 1516
rect 10505 1507 10563 1513
rect 10778 1504 10784 1516
rect 10836 1504 10842 1556
rect 15102 1544 15108 1556
rect 15063 1516 15108 1544
rect 15102 1504 15108 1516
rect 15160 1504 15166 1556
rect 22186 1544 22192 1556
rect 21284 1516 22192 1544
rect 18598 1436 18604 1488
rect 18656 1476 18662 1488
rect 21284 1476 21312 1516
rect 22186 1504 22192 1516
rect 22244 1504 22250 1556
rect 25038 1544 25044 1556
rect 24999 1516 25044 1544
rect 25038 1504 25044 1516
rect 25096 1504 25102 1556
rect 26786 1544 26792 1556
rect 26747 1516 26792 1544
rect 26786 1504 26792 1516
rect 26844 1504 26850 1556
rect 28258 1544 28264 1556
rect 28219 1516 28264 1544
rect 28258 1504 28264 1516
rect 28316 1504 28322 1556
rect 30466 1544 30472 1556
rect 28368 1516 29500 1544
rect 30427 1516 30472 1544
rect 18656 1448 21312 1476
rect 18656 1436 18662 1448
rect 22094 1436 22100 1488
rect 22152 1476 22158 1488
rect 23845 1479 23903 1485
rect 23845 1476 23857 1479
rect 22152 1448 23857 1476
rect 22152 1436 22158 1448
rect 23845 1445 23857 1448
rect 23891 1445 23903 1479
rect 23845 1439 23903 1445
rect 24026 1436 24032 1488
rect 24084 1476 24090 1488
rect 28368 1476 28396 1516
rect 24084 1448 28396 1476
rect 24084 1436 24090 1448
rect 5353 1411 5411 1417
rect 5353 1408 5365 1411
rect 2464 1380 5365 1408
rect 2464 1368 2470 1380
rect 5353 1377 5365 1380
rect 5399 1377 5411 1411
rect 5353 1371 5411 1377
rect 9493 1411 9551 1417
rect 9493 1377 9505 1411
rect 9539 1377 9551 1411
rect 11606 1408 11612 1420
rect 11567 1380 11612 1408
rect 9493 1371 9551 1377
rect 11606 1368 11612 1380
rect 11664 1368 11670 1420
rect 11790 1368 11796 1420
rect 11848 1408 11854 1420
rect 16209 1411 16267 1417
rect 16209 1408 16221 1411
rect 11848 1380 16221 1408
rect 11848 1368 11854 1380
rect 16209 1377 16221 1380
rect 16255 1377 16267 1411
rect 16209 1371 16267 1377
rect 20714 1368 20720 1420
rect 20772 1408 20778 1420
rect 21177 1411 21235 1417
rect 21177 1408 21189 1411
rect 20772 1380 21189 1408
rect 20772 1368 20778 1380
rect 21177 1377 21189 1380
rect 21223 1377 21235 1411
rect 22554 1408 22560 1420
rect 22515 1380 22560 1408
rect 21177 1371 21235 1377
rect 22554 1368 22560 1380
rect 22612 1368 22618 1420
rect 28074 1408 28080 1420
rect 24136 1380 28080 1408
rect 4341 1343 4399 1349
rect 4341 1340 4353 1343
rect 4172 1312 4353 1340
rect 4172 1281 4200 1312
rect 4341 1309 4353 1312
rect 4387 1309 4399 1343
rect 4341 1303 4399 1309
rect 5905 1343 5963 1349
rect 5905 1309 5917 1343
rect 5951 1340 5963 1343
rect 7742 1340 7748 1352
rect 5951 1312 6316 1340
rect 7703 1312 7748 1340
rect 5951 1309 5963 1312
rect 5905 1303 5963 1309
rect 3329 1275 3387 1281
rect 3329 1241 3341 1275
rect 3375 1272 3387 1275
rect 4157 1275 4215 1281
rect 4157 1272 4169 1275
rect 3375 1244 4169 1272
rect 3375 1241 3387 1244
rect 3329 1235 3387 1241
rect 4157 1241 4169 1244
rect 4203 1241 4215 1275
rect 4157 1235 4215 1241
rect 6288 1216 6316 1312
rect 7742 1300 7748 1312
rect 7800 1300 7806 1352
rect 10597 1343 10655 1349
rect 10597 1309 10609 1343
rect 10643 1340 10655 1343
rect 11146 1340 11152 1352
rect 10643 1312 11152 1340
rect 10643 1309 10655 1312
rect 10597 1303 10655 1309
rect 11146 1300 11152 1312
rect 11204 1300 11210 1352
rect 12161 1343 12219 1349
rect 12161 1309 12173 1343
rect 12207 1309 12219 1343
rect 12161 1303 12219 1309
rect 2225 1207 2283 1213
rect 2225 1173 2237 1207
rect 2271 1204 2283 1207
rect 5994 1204 6000 1216
rect 2271 1176 6000 1204
rect 2271 1173 2283 1176
rect 2225 1167 2283 1173
rect 5994 1164 6000 1176
rect 6052 1164 6058 1216
rect 6270 1204 6276 1216
rect 6231 1176 6276 1204
rect 6270 1164 6276 1176
rect 6328 1164 6334 1216
rect 6730 1204 6736 1216
rect 6691 1176 6736 1204
rect 6730 1164 6736 1176
rect 6788 1164 6794 1216
rect 8297 1207 8355 1213
rect 8297 1173 8309 1207
rect 8343 1204 8355 1207
rect 8386 1204 8392 1216
rect 8343 1176 8392 1204
rect 8343 1173 8355 1176
rect 8297 1167 8355 1173
rect 8386 1164 8392 1176
rect 8444 1164 8450 1216
rect 12176 1204 12204 1303
rect 15102 1300 15108 1352
rect 15160 1340 15166 1352
rect 15197 1343 15255 1349
rect 15197 1340 15209 1343
rect 15160 1312 15209 1340
rect 15160 1300 15166 1312
rect 15197 1309 15209 1312
rect 15243 1309 15255 1343
rect 15197 1303 15255 1309
rect 16761 1343 16819 1349
rect 16761 1309 16773 1343
rect 16807 1309 16819 1343
rect 18874 1340 18880 1352
rect 18835 1312 18880 1340
rect 16761 1303 16819 1309
rect 12529 1207 12587 1213
rect 12529 1204 12541 1207
rect 12176 1176 12541 1204
rect 12529 1173 12541 1176
rect 12575 1204 12587 1207
rect 12802 1204 12808 1216
rect 12575 1176 12808 1204
rect 12575 1173 12587 1176
rect 12529 1167 12587 1173
rect 12802 1164 12808 1176
rect 12860 1164 12866 1216
rect 12986 1204 12992 1216
rect 12947 1176 12992 1204
rect 12986 1164 12992 1176
rect 13044 1164 13050 1216
rect 16776 1204 16804 1303
rect 18874 1300 18880 1312
rect 18932 1340 18938 1352
rect 19521 1343 19579 1349
rect 19521 1340 19533 1343
rect 18932 1312 19533 1340
rect 18932 1300 18938 1312
rect 19521 1309 19533 1312
rect 19567 1309 19579 1343
rect 19521 1303 19579 1309
rect 19797 1343 19855 1349
rect 19797 1309 19809 1343
rect 19843 1340 19855 1343
rect 20165 1343 20223 1349
rect 20165 1340 20177 1343
rect 19843 1312 20177 1340
rect 19843 1309 19855 1312
rect 19797 1303 19855 1309
rect 20165 1309 20177 1312
rect 20211 1309 20223 1343
rect 20165 1303 20223 1309
rect 21729 1343 21787 1349
rect 21729 1309 21741 1343
rect 21775 1340 21787 1343
rect 22097 1343 22155 1349
rect 22097 1340 22109 1343
rect 21775 1312 22109 1340
rect 21775 1309 21787 1312
rect 21729 1303 21787 1309
rect 22097 1309 22109 1312
rect 22143 1340 22155 1343
rect 23474 1340 23480 1352
rect 22143 1312 23480 1340
rect 22143 1309 22155 1312
rect 22097 1303 22155 1309
rect 23474 1300 23480 1312
rect 23532 1300 23538 1352
rect 23566 1300 23572 1352
rect 23624 1340 23630 1352
rect 23661 1343 23719 1349
rect 23661 1340 23673 1343
rect 23624 1312 23673 1340
rect 23624 1300 23630 1312
rect 23661 1309 23673 1312
rect 23707 1309 23719 1343
rect 23661 1303 23719 1309
rect 17494 1232 17500 1284
rect 17552 1272 17558 1284
rect 18690 1272 18696 1284
rect 17552 1244 18696 1272
rect 17552 1232 17558 1244
rect 18690 1232 18696 1244
rect 18748 1232 18754 1284
rect 19245 1275 19303 1281
rect 19245 1241 19257 1275
rect 19291 1272 19303 1275
rect 24136 1272 24164 1380
rect 28074 1368 28080 1380
rect 28132 1368 28138 1420
rect 28184 1380 28580 1408
rect 26142 1340 26148 1352
rect 26103 1312 26148 1340
rect 26142 1300 26148 1312
rect 26200 1300 26206 1352
rect 26510 1340 26516 1352
rect 26471 1312 26516 1340
rect 26510 1300 26516 1312
rect 26568 1300 26574 1352
rect 27338 1300 27344 1352
rect 27396 1340 27402 1352
rect 27396 1312 27441 1340
rect 27396 1300 27402 1312
rect 27706 1300 27712 1352
rect 27764 1340 27770 1352
rect 28184 1340 28212 1380
rect 27764 1312 28212 1340
rect 27764 1300 27770 1312
rect 28350 1300 28356 1352
rect 28408 1340 28414 1352
rect 28552 1340 28580 1380
rect 28626 1368 28632 1420
rect 28684 1408 28690 1420
rect 29365 1411 29423 1417
rect 29365 1408 29377 1411
rect 28684 1380 29377 1408
rect 28684 1368 28690 1380
rect 29365 1377 29377 1380
rect 29411 1377 29423 1411
rect 29472 1408 29500 1516
rect 30466 1504 30472 1516
rect 30524 1504 30530 1556
rect 30742 1504 30748 1556
rect 30800 1544 30806 1556
rect 32766 1544 32772 1556
rect 30800 1516 32772 1544
rect 30800 1504 30806 1516
rect 32766 1504 32772 1516
rect 32824 1504 32830 1556
rect 33410 1504 33416 1556
rect 33468 1544 33474 1556
rect 40494 1544 40500 1556
rect 33468 1516 40500 1544
rect 33468 1504 33474 1516
rect 40494 1504 40500 1516
rect 40552 1504 40558 1556
rect 40678 1504 40684 1556
rect 40736 1544 40742 1556
rect 41966 1544 41972 1556
rect 40736 1516 41972 1544
rect 40736 1504 40742 1516
rect 41966 1504 41972 1516
rect 42024 1504 42030 1556
rect 42242 1504 42248 1556
rect 42300 1544 42306 1556
rect 46293 1547 46351 1553
rect 46293 1544 46305 1547
rect 42300 1516 46305 1544
rect 42300 1504 42306 1516
rect 46293 1513 46305 1516
rect 46339 1513 46351 1547
rect 46474 1544 46480 1556
rect 46435 1516 46480 1544
rect 46293 1507 46351 1513
rect 46474 1504 46480 1516
rect 46532 1504 46538 1556
rect 48590 1544 48596 1556
rect 46584 1516 48596 1544
rect 30282 1436 30288 1488
rect 30340 1476 30346 1488
rect 33502 1476 33508 1488
rect 30340 1448 33508 1476
rect 30340 1436 30346 1448
rect 33502 1436 33508 1448
rect 33560 1436 33566 1488
rect 33870 1476 33876 1488
rect 33831 1448 33876 1476
rect 33870 1436 33876 1448
rect 33928 1436 33934 1488
rect 34330 1436 34336 1488
rect 34388 1476 34394 1488
rect 40126 1476 40132 1488
rect 34388 1448 40132 1476
rect 34388 1436 34394 1448
rect 40126 1436 40132 1448
rect 40184 1436 40190 1488
rect 43990 1476 43996 1488
rect 40236 1448 43996 1476
rect 32401 1411 32459 1417
rect 32401 1408 32413 1411
rect 29472 1380 32413 1408
rect 29365 1371 29423 1377
rect 32401 1377 32413 1380
rect 32447 1377 32459 1411
rect 32401 1371 32459 1377
rect 32490 1368 32496 1420
rect 32548 1408 32554 1420
rect 32548 1380 36400 1408
rect 32548 1368 32554 1380
rect 29917 1343 29975 1349
rect 28408 1312 28453 1340
rect 28552 1312 28764 1340
rect 28408 1300 28414 1312
rect 19291 1244 24164 1272
rect 19291 1241 19303 1244
rect 19245 1235 19303 1241
rect 24670 1232 24676 1284
rect 24728 1272 24734 1284
rect 25317 1275 25375 1281
rect 25317 1272 25329 1275
rect 24728 1244 25329 1272
rect 24728 1232 24734 1244
rect 25317 1241 25329 1244
rect 25363 1241 25375 1275
rect 25317 1235 25375 1241
rect 26050 1232 26056 1284
rect 26108 1272 26114 1284
rect 28626 1272 28632 1284
rect 26108 1244 28632 1272
rect 26108 1232 26114 1244
rect 28626 1232 28632 1244
rect 28684 1232 28690 1284
rect 28736 1272 28764 1312
rect 29917 1309 29929 1343
rect 29963 1340 29975 1343
rect 30561 1343 30619 1349
rect 30561 1340 30573 1343
rect 29963 1312 30573 1340
rect 29963 1309 29975 1312
rect 29917 1303 29975 1309
rect 30561 1309 30573 1312
rect 30607 1309 30619 1343
rect 30561 1303 30619 1309
rect 30834 1300 30840 1352
rect 30892 1340 30898 1352
rect 31113 1343 31171 1349
rect 31113 1340 31125 1343
rect 30892 1312 31125 1340
rect 30892 1300 30898 1312
rect 31113 1309 31125 1312
rect 31159 1340 31171 1343
rect 31389 1343 31447 1349
rect 31389 1340 31401 1343
rect 31159 1312 31401 1340
rect 31159 1309 31171 1312
rect 31113 1303 31171 1309
rect 31389 1309 31401 1312
rect 31435 1309 31447 1343
rect 31389 1303 31447 1309
rect 32953 1343 33011 1349
rect 32953 1309 32965 1343
rect 32999 1340 33011 1343
rect 33045 1343 33103 1349
rect 33045 1340 33057 1343
rect 32999 1312 33057 1340
rect 32999 1309 33011 1312
rect 32953 1303 33011 1309
rect 33045 1309 33057 1312
rect 33091 1309 33103 1343
rect 33594 1340 33600 1352
rect 33555 1312 33600 1340
rect 33045 1303 33103 1309
rect 33594 1300 33600 1312
rect 33652 1340 33658 1352
rect 33781 1343 33839 1349
rect 33781 1340 33793 1343
rect 33652 1312 33793 1340
rect 33652 1300 33658 1312
rect 33781 1309 33793 1312
rect 33827 1309 33839 1343
rect 33781 1303 33839 1309
rect 34517 1343 34575 1349
rect 34517 1309 34529 1343
rect 34563 1309 34575 1343
rect 35342 1340 35348 1352
rect 35303 1312 35348 1340
rect 34517 1303 34575 1309
rect 33134 1272 33140 1284
rect 28736 1244 33140 1272
rect 33134 1232 33140 1244
rect 33192 1232 33198 1284
rect 34532 1272 34560 1303
rect 35342 1300 35348 1312
rect 35400 1300 35406 1352
rect 35434 1300 35440 1352
rect 35492 1340 35498 1352
rect 35713 1343 35771 1349
rect 35713 1340 35725 1343
rect 35492 1312 35725 1340
rect 35492 1300 35498 1312
rect 35713 1309 35725 1312
rect 35759 1340 35771 1343
rect 35894 1340 35900 1352
rect 35759 1312 35900 1340
rect 35759 1309 35771 1312
rect 35713 1303 35771 1309
rect 35894 1300 35900 1312
rect 35952 1300 35958 1352
rect 36081 1343 36139 1349
rect 36081 1309 36093 1343
rect 36127 1309 36139 1343
rect 36372 1340 36400 1380
rect 36446 1368 36452 1420
rect 36504 1408 36510 1420
rect 39574 1408 39580 1420
rect 36504 1380 39580 1408
rect 36504 1368 36510 1380
rect 39574 1368 39580 1380
rect 39632 1368 39638 1420
rect 39666 1368 39672 1420
rect 39724 1408 39730 1420
rect 40236 1408 40264 1448
rect 43990 1436 43996 1448
rect 44048 1436 44054 1488
rect 44100 1448 45324 1476
rect 40862 1408 40868 1420
rect 39724 1380 40264 1408
rect 40328 1380 40868 1408
rect 39724 1368 39730 1380
rect 36814 1340 36820 1352
rect 36372 1312 36820 1340
rect 36081 1303 36139 1309
rect 34882 1272 34888 1284
rect 34532 1244 34888 1272
rect 34882 1232 34888 1244
rect 34940 1232 34946 1284
rect 35066 1232 35072 1284
rect 35124 1272 35130 1284
rect 35986 1272 35992 1284
rect 35124 1244 35992 1272
rect 35124 1232 35130 1244
rect 35986 1232 35992 1244
rect 36044 1232 36050 1284
rect 36096 1272 36124 1303
rect 36814 1300 36820 1312
rect 36872 1300 36878 1352
rect 36998 1340 37004 1352
rect 36959 1312 37004 1340
rect 36998 1300 37004 1312
rect 37056 1300 37062 1352
rect 37369 1343 37427 1349
rect 37369 1309 37381 1343
rect 37415 1340 37427 1343
rect 37550 1340 37556 1352
rect 37415 1312 37556 1340
rect 37415 1309 37427 1312
rect 37369 1303 37427 1309
rect 37550 1300 37556 1312
rect 37608 1300 37614 1352
rect 37737 1343 37795 1349
rect 37737 1309 37749 1343
rect 37783 1340 37795 1343
rect 38105 1343 38163 1349
rect 38105 1340 38117 1343
rect 37783 1312 38117 1340
rect 37783 1309 37795 1312
rect 37737 1303 37795 1309
rect 38105 1309 38117 1312
rect 38151 1340 38163 1343
rect 39022 1340 39028 1352
rect 38151 1312 39028 1340
rect 38151 1309 38163 1312
rect 38105 1303 38163 1309
rect 39022 1300 39028 1312
rect 39080 1300 39086 1352
rect 39114 1300 39120 1352
rect 39172 1340 39178 1352
rect 39209 1343 39267 1349
rect 39209 1340 39221 1343
rect 39172 1312 39221 1340
rect 39172 1300 39178 1312
rect 39209 1309 39221 1312
rect 39255 1340 39267 1343
rect 40129 1343 40187 1349
rect 40129 1340 40141 1343
rect 39255 1312 40141 1340
rect 39255 1309 39267 1312
rect 39209 1303 39267 1309
rect 40129 1309 40141 1312
rect 40175 1309 40187 1343
rect 40129 1303 40187 1309
rect 40218 1300 40224 1352
rect 40276 1340 40282 1352
rect 40328 1340 40356 1380
rect 40862 1368 40868 1380
rect 40920 1368 40926 1420
rect 40954 1368 40960 1420
rect 41012 1408 41018 1420
rect 41322 1408 41328 1420
rect 41012 1380 41328 1408
rect 41012 1368 41018 1380
rect 41322 1368 41328 1380
rect 41380 1368 41386 1420
rect 41506 1408 41512 1420
rect 41467 1380 41512 1408
rect 41506 1368 41512 1380
rect 41564 1368 41570 1420
rect 43717 1411 43775 1417
rect 43717 1408 43729 1411
rect 41616 1380 43729 1408
rect 40276 1312 40356 1340
rect 40276 1300 40282 1312
rect 40402 1300 40408 1352
rect 40460 1340 40466 1352
rect 41616 1340 41644 1380
rect 43717 1377 43729 1380
rect 43763 1377 43775 1411
rect 43717 1371 43775 1377
rect 43806 1368 43812 1420
rect 43864 1408 43870 1420
rect 44100 1408 44128 1448
rect 44910 1408 44916 1420
rect 43864 1380 44128 1408
rect 44192 1380 44916 1408
rect 43864 1368 43870 1380
rect 40460 1312 41644 1340
rect 40460 1300 40466 1312
rect 41690 1300 41696 1352
rect 41748 1340 41754 1352
rect 42518 1340 42524 1352
rect 41748 1312 42524 1340
rect 41748 1300 41754 1312
rect 42518 1300 42524 1312
rect 42576 1300 42582 1352
rect 42610 1300 42616 1352
rect 42668 1340 42674 1352
rect 42705 1343 42763 1349
rect 42705 1340 42717 1343
rect 42668 1312 42717 1340
rect 42668 1300 42674 1312
rect 42705 1309 42717 1312
rect 42751 1309 42763 1343
rect 42705 1303 42763 1309
rect 36449 1275 36507 1281
rect 36449 1272 36461 1275
rect 36096 1244 36461 1272
rect 36449 1241 36461 1244
rect 36495 1272 36507 1275
rect 39482 1272 39488 1284
rect 36495 1244 39488 1272
rect 36495 1241 36507 1244
rect 36449 1235 36507 1241
rect 39482 1232 39488 1244
rect 39540 1232 39546 1284
rect 39853 1275 39911 1281
rect 39853 1241 39865 1275
rect 39899 1272 39911 1275
rect 39899 1244 40540 1272
rect 39899 1241 39911 1244
rect 39853 1235 39911 1241
rect 17129 1207 17187 1213
rect 17129 1204 17141 1207
rect 16776 1176 17141 1204
rect 17129 1173 17141 1176
rect 17175 1204 17187 1207
rect 17218 1204 17224 1216
rect 17175 1176 17224 1204
rect 17175 1173 17187 1176
rect 17129 1167 17187 1173
rect 17218 1164 17224 1176
rect 17276 1164 17282 1216
rect 19610 1164 19616 1216
rect 19668 1204 19674 1216
rect 19797 1207 19855 1213
rect 19797 1204 19809 1207
rect 19668 1176 19809 1204
rect 19668 1164 19674 1176
rect 19797 1173 19809 1176
rect 19843 1204 19855 1207
rect 19889 1207 19947 1213
rect 19889 1204 19901 1207
rect 19843 1176 19901 1204
rect 19843 1173 19855 1176
rect 19797 1167 19855 1173
rect 19889 1173 19901 1176
rect 19935 1173 19947 1207
rect 19889 1167 19947 1173
rect 20806 1164 20812 1216
rect 20864 1204 20870 1216
rect 22738 1204 22744 1216
rect 20864 1176 22744 1204
rect 20864 1164 20870 1176
rect 22738 1164 22744 1176
rect 22796 1164 22802 1216
rect 23566 1164 23572 1216
rect 23624 1204 23630 1216
rect 24489 1207 24547 1213
rect 24489 1204 24501 1207
rect 23624 1176 24501 1204
rect 23624 1164 23630 1176
rect 24489 1173 24501 1176
rect 24535 1204 24547 1207
rect 24578 1204 24584 1216
rect 24535 1176 24584 1204
rect 24535 1173 24547 1176
rect 24489 1167 24547 1173
rect 24578 1164 24584 1176
rect 24636 1164 24642 1216
rect 25774 1164 25780 1216
rect 25832 1204 25838 1216
rect 30282 1204 30288 1216
rect 25832 1176 30288 1204
rect 25832 1164 25838 1176
rect 30282 1164 30288 1176
rect 30340 1164 30346 1216
rect 30561 1207 30619 1213
rect 30561 1173 30573 1207
rect 30607 1204 30619 1207
rect 30834 1204 30840 1216
rect 30607 1176 30840 1204
rect 30607 1173 30619 1176
rect 30561 1167 30619 1173
rect 30834 1164 30840 1176
rect 30892 1164 30898 1216
rect 33045 1207 33103 1213
rect 33045 1173 33057 1207
rect 33091 1204 33103 1207
rect 33321 1207 33379 1213
rect 33321 1204 33333 1207
rect 33091 1176 33333 1204
rect 33091 1173 33103 1176
rect 33045 1167 33103 1173
rect 33321 1173 33333 1176
rect 33367 1204 33379 1207
rect 40402 1204 40408 1216
rect 33367 1176 40408 1204
rect 33367 1173 33379 1176
rect 33321 1167 33379 1173
rect 40402 1164 40408 1176
rect 40460 1164 40466 1216
rect 40512 1204 40540 1244
rect 40586 1232 40592 1284
rect 40644 1272 40650 1284
rect 44192 1272 44220 1380
rect 44910 1368 44916 1380
rect 44968 1368 44974 1420
rect 44269 1343 44327 1349
rect 44269 1309 44281 1343
rect 44315 1309 44327 1343
rect 44269 1303 44327 1309
rect 40644 1244 44220 1272
rect 40644 1232 40650 1244
rect 43254 1204 43260 1216
rect 40512 1176 43260 1204
rect 43254 1164 43260 1176
rect 43312 1164 43318 1216
rect 44284 1204 44312 1303
rect 44358 1300 44364 1352
rect 44416 1340 44422 1352
rect 45296 1349 45324 1448
rect 45646 1436 45652 1488
rect 45704 1476 45710 1488
rect 46584 1476 46612 1516
rect 48590 1504 48596 1516
rect 48648 1504 48654 1556
rect 48682 1504 48688 1556
rect 48740 1544 48746 1556
rect 49605 1547 49663 1553
rect 49605 1544 49617 1547
rect 48740 1516 49617 1544
rect 48740 1504 48746 1516
rect 49605 1513 49617 1516
rect 49651 1544 49663 1547
rect 50982 1544 50988 1556
rect 49651 1516 50988 1544
rect 49651 1513 49663 1516
rect 49605 1507 49663 1513
rect 50982 1504 50988 1516
rect 51040 1504 51046 1556
rect 51074 1504 51080 1556
rect 51132 1544 51138 1556
rect 57057 1547 57115 1553
rect 57057 1544 57069 1547
rect 51132 1516 57069 1544
rect 51132 1504 51138 1516
rect 57057 1513 57069 1516
rect 57103 1513 57115 1547
rect 58802 1544 58808 1556
rect 58763 1516 58808 1544
rect 57057 1507 57115 1513
rect 58802 1504 58808 1516
rect 58860 1504 58866 1556
rect 59078 1504 59084 1556
rect 59136 1544 59142 1556
rect 61105 1547 61163 1553
rect 61105 1544 61117 1547
rect 59136 1516 61117 1544
rect 59136 1504 59142 1516
rect 61105 1513 61117 1516
rect 61151 1513 61163 1547
rect 61105 1507 61163 1513
rect 61381 1547 61439 1553
rect 61381 1513 61393 1547
rect 61427 1544 61439 1547
rect 61562 1544 61568 1556
rect 61427 1516 61568 1544
rect 61427 1513 61439 1516
rect 61381 1507 61439 1513
rect 61562 1504 61568 1516
rect 61620 1504 61626 1556
rect 62114 1544 62120 1556
rect 62075 1516 62120 1544
rect 62114 1504 62120 1516
rect 62172 1504 62178 1556
rect 62482 1504 62488 1556
rect 62540 1544 62546 1556
rect 63310 1544 63316 1556
rect 62540 1516 63316 1544
rect 62540 1504 62546 1516
rect 63310 1504 63316 1516
rect 63368 1504 63374 1556
rect 63770 1504 63776 1556
rect 63828 1544 63834 1556
rect 69842 1544 69848 1556
rect 63828 1516 69848 1544
rect 63828 1504 63834 1516
rect 69842 1504 69848 1516
rect 69900 1504 69906 1556
rect 70029 1547 70087 1553
rect 70029 1513 70041 1547
rect 70075 1544 70087 1547
rect 70302 1544 70308 1556
rect 70075 1516 70308 1544
rect 70075 1513 70087 1516
rect 70029 1507 70087 1513
rect 70302 1504 70308 1516
rect 70360 1504 70366 1556
rect 70394 1504 70400 1556
rect 70452 1544 70458 1556
rect 72602 1544 72608 1556
rect 70452 1516 72608 1544
rect 70452 1504 70458 1516
rect 72602 1504 72608 1516
rect 72660 1504 72666 1556
rect 72697 1547 72755 1553
rect 72697 1513 72709 1547
rect 72743 1544 72755 1547
rect 74994 1544 75000 1556
rect 72743 1516 75000 1544
rect 72743 1513 72755 1516
rect 72697 1507 72755 1513
rect 74994 1504 75000 1516
rect 75052 1504 75058 1556
rect 75086 1504 75092 1556
rect 75144 1544 75150 1556
rect 75181 1547 75239 1553
rect 75181 1544 75193 1547
rect 75144 1516 75193 1544
rect 75144 1504 75150 1516
rect 75181 1513 75193 1516
rect 75227 1513 75239 1547
rect 75181 1507 75239 1513
rect 80974 1504 80980 1556
rect 81032 1544 81038 1556
rect 81250 1544 81256 1556
rect 81032 1516 81256 1544
rect 81032 1504 81038 1516
rect 81250 1504 81256 1516
rect 81308 1544 81314 1556
rect 81621 1547 81679 1553
rect 81621 1544 81633 1547
rect 81308 1516 81633 1544
rect 81308 1504 81314 1516
rect 81621 1513 81633 1516
rect 81667 1513 81679 1547
rect 81621 1507 81679 1513
rect 84654 1504 84660 1556
rect 84712 1544 84718 1556
rect 84841 1547 84899 1553
rect 84841 1544 84853 1547
rect 84712 1516 84853 1544
rect 84712 1504 84718 1516
rect 84841 1513 84853 1516
rect 84887 1513 84899 1547
rect 87414 1544 87420 1556
rect 84841 1507 84899 1513
rect 85040 1516 87420 1544
rect 45704 1448 46612 1476
rect 45704 1436 45710 1448
rect 46750 1436 46756 1488
rect 46808 1476 46814 1488
rect 50338 1476 50344 1488
rect 46808 1448 50344 1476
rect 46808 1436 46814 1448
rect 50338 1436 50344 1448
rect 50396 1436 50402 1488
rect 55214 1476 55220 1488
rect 50448 1448 55076 1476
rect 55175 1448 55220 1476
rect 45370 1368 45376 1420
rect 45428 1408 45434 1420
rect 46474 1408 46480 1420
rect 45428 1380 46480 1408
rect 45428 1368 45434 1380
rect 46474 1368 46480 1380
rect 46532 1368 46538 1420
rect 46566 1368 46572 1420
rect 46624 1408 46630 1420
rect 46661 1411 46719 1417
rect 46661 1408 46673 1411
rect 46624 1380 46673 1408
rect 46624 1368 46630 1380
rect 46661 1377 46673 1380
rect 46707 1377 46719 1411
rect 50448 1408 50476 1448
rect 46661 1371 46719 1377
rect 46768 1380 50476 1408
rect 45097 1343 45155 1349
rect 45097 1340 45109 1343
rect 44416 1312 45109 1340
rect 44416 1300 44422 1312
rect 45097 1309 45109 1312
rect 45143 1309 45155 1343
rect 45097 1303 45155 1309
rect 45281 1343 45339 1349
rect 45281 1309 45293 1343
rect 45327 1340 45339 1343
rect 46109 1343 46167 1349
rect 46109 1340 46121 1343
rect 45327 1312 46121 1340
rect 45327 1309 45339 1312
rect 45281 1303 45339 1309
rect 46109 1309 46121 1312
rect 46155 1309 46167 1343
rect 46109 1303 46167 1309
rect 46293 1343 46351 1349
rect 46293 1309 46305 1343
rect 46339 1340 46351 1343
rect 46768 1340 46796 1380
rect 50522 1368 50528 1420
rect 50580 1408 50586 1420
rect 53190 1408 53196 1420
rect 50580 1380 53196 1408
rect 50580 1368 50586 1380
rect 53190 1368 53196 1380
rect 53248 1368 53254 1420
rect 53466 1368 53472 1420
rect 53524 1408 53530 1420
rect 54294 1408 54300 1420
rect 53524 1380 54300 1408
rect 53524 1368 53530 1380
rect 54294 1368 54300 1380
rect 54352 1368 54358 1420
rect 55048 1408 55076 1448
rect 55214 1436 55220 1448
rect 55272 1436 55278 1488
rect 55490 1436 55496 1488
rect 55548 1476 55554 1488
rect 84749 1479 84807 1485
rect 84749 1476 84761 1479
rect 55548 1448 84761 1476
rect 55548 1436 55554 1448
rect 84749 1445 84761 1448
rect 84795 1445 84807 1479
rect 84749 1439 84807 1445
rect 57698 1408 57704 1420
rect 55048 1380 57704 1408
rect 57698 1368 57704 1380
rect 57756 1368 57762 1420
rect 59906 1368 59912 1420
rect 59964 1408 59970 1420
rect 59964 1380 60688 1408
rect 59964 1368 59970 1380
rect 46339 1312 46796 1340
rect 46339 1309 46351 1312
rect 46293 1303 46351 1309
rect 46934 1300 46940 1352
rect 46992 1340 46998 1352
rect 48774 1340 48780 1352
rect 46992 1312 48780 1340
rect 46992 1300 46998 1312
rect 48774 1300 48780 1312
rect 48832 1300 48838 1352
rect 48869 1343 48927 1349
rect 48869 1309 48881 1343
rect 48915 1309 48927 1343
rect 48869 1303 48927 1309
rect 44726 1232 44732 1284
rect 44784 1272 44790 1284
rect 45646 1272 45652 1284
rect 44784 1244 45652 1272
rect 44784 1232 44790 1244
rect 45646 1232 45652 1244
rect 45704 1232 45710 1284
rect 45830 1232 45836 1284
rect 45888 1272 45894 1284
rect 47302 1272 47308 1284
rect 45888 1244 47308 1272
rect 45888 1232 45894 1244
rect 47302 1232 47308 1244
rect 47360 1232 47366 1284
rect 47412 1244 47716 1272
rect 44634 1204 44640 1216
rect 44284 1176 44640 1204
rect 44634 1164 44640 1176
rect 44692 1164 44698 1216
rect 44910 1164 44916 1216
rect 44968 1204 44974 1216
rect 47412 1204 47440 1244
rect 47578 1204 47584 1216
rect 44968 1176 47440 1204
rect 47539 1176 47584 1204
rect 44968 1164 44974 1176
rect 47578 1164 47584 1176
rect 47636 1164 47642 1216
rect 47688 1204 47716 1244
rect 47762 1232 47768 1284
rect 47820 1272 47826 1284
rect 48225 1275 48283 1281
rect 48225 1272 48237 1275
rect 47820 1244 48237 1272
rect 47820 1232 47826 1244
rect 48225 1241 48237 1244
rect 48271 1241 48283 1275
rect 48884 1272 48912 1303
rect 49050 1300 49056 1352
rect 49108 1340 49114 1352
rect 49789 1343 49847 1349
rect 49789 1340 49801 1343
rect 49108 1312 49801 1340
rect 49108 1300 49114 1312
rect 49789 1309 49801 1312
rect 49835 1309 49847 1343
rect 49789 1303 49847 1309
rect 50062 1300 50068 1352
rect 50120 1340 50126 1352
rect 50338 1340 50344 1352
rect 50120 1312 50344 1340
rect 50120 1300 50126 1312
rect 50338 1300 50344 1312
rect 50396 1300 50402 1352
rect 50433 1343 50491 1349
rect 50433 1309 50445 1343
rect 50479 1340 50491 1343
rect 50893 1343 50951 1349
rect 50893 1340 50905 1343
rect 50479 1312 50905 1340
rect 50479 1309 50491 1312
rect 50433 1303 50491 1309
rect 50893 1309 50905 1312
rect 50939 1340 50951 1343
rect 51902 1340 51908 1352
rect 50939 1312 51908 1340
rect 50939 1309 50951 1312
rect 50893 1303 50951 1309
rect 51902 1300 51908 1312
rect 51960 1300 51966 1352
rect 51997 1343 52055 1349
rect 51997 1309 52009 1343
rect 52043 1340 52055 1343
rect 52178 1340 52184 1352
rect 52043 1312 52184 1340
rect 52043 1309 52055 1312
rect 51997 1303 52055 1309
rect 52178 1300 52184 1312
rect 52236 1340 52242 1352
rect 52457 1343 52515 1349
rect 52457 1340 52469 1343
rect 52236 1312 52469 1340
rect 52236 1300 52242 1312
rect 52457 1309 52469 1312
rect 52503 1309 52515 1343
rect 52457 1303 52515 1309
rect 53561 1343 53619 1349
rect 53561 1309 53573 1343
rect 53607 1340 53619 1343
rect 53650 1340 53656 1352
rect 53607 1312 53656 1340
rect 53607 1309 53619 1312
rect 53561 1303 53619 1309
rect 53650 1300 53656 1312
rect 53708 1300 53714 1352
rect 53834 1340 53840 1352
rect 53795 1312 53840 1340
rect 53834 1300 53840 1312
rect 53892 1300 53898 1352
rect 54205 1343 54263 1349
rect 54205 1309 54217 1343
rect 54251 1309 54263 1343
rect 54205 1303 54263 1309
rect 54573 1343 54631 1349
rect 54573 1309 54585 1343
rect 54619 1340 54631 1343
rect 54941 1343 54999 1349
rect 54941 1340 54953 1343
rect 54619 1312 54953 1340
rect 54619 1309 54631 1312
rect 54573 1303 54631 1309
rect 54941 1309 54953 1312
rect 54987 1340 54999 1343
rect 55214 1340 55220 1352
rect 54987 1312 55220 1340
rect 54987 1309 54999 1312
rect 54941 1303 54999 1309
rect 49329 1275 49387 1281
rect 49329 1272 49341 1275
rect 48884 1244 49341 1272
rect 48225 1235 48283 1241
rect 49329 1241 49341 1244
rect 49375 1272 49387 1275
rect 54220 1272 54248 1303
rect 55214 1300 55220 1312
rect 55272 1300 55278 1352
rect 55582 1340 55588 1352
rect 55543 1312 55588 1340
rect 55582 1300 55588 1312
rect 55640 1300 55646 1352
rect 55769 1343 55827 1349
rect 55769 1309 55781 1343
rect 55815 1309 55827 1343
rect 55769 1303 55827 1309
rect 56137 1343 56195 1349
rect 56137 1309 56149 1343
rect 56183 1309 56195 1343
rect 56137 1303 56195 1309
rect 55784 1272 55812 1303
rect 49375 1244 54248 1272
rect 54312 1244 55812 1272
rect 49375 1241 49387 1244
rect 49329 1235 49387 1241
rect 50062 1204 50068 1216
rect 47688 1176 50068 1204
rect 50062 1164 50068 1176
rect 50120 1164 50126 1216
rect 50154 1164 50160 1216
rect 50212 1204 50218 1216
rect 54312 1204 54340 1244
rect 50212 1176 54340 1204
rect 50212 1164 50218 1176
rect 55306 1164 55312 1216
rect 55364 1204 55370 1216
rect 56042 1204 56048 1216
rect 55364 1176 56048 1204
rect 55364 1164 55370 1176
rect 56042 1164 56048 1176
rect 56100 1164 56106 1216
rect 56152 1204 56180 1303
rect 56226 1300 56232 1352
rect 56284 1340 56290 1352
rect 56962 1340 56968 1352
rect 56284 1312 56640 1340
rect 56923 1312 56968 1340
rect 56284 1300 56290 1312
rect 56502 1204 56508 1216
rect 56152 1176 56508 1204
rect 56502 1164 56508 1176
rect 56560 1164 56566 1216
rect 56612 1204 56640 1312
rect 56962 1300 56968 1312
rect 57020 1300 57026 1352
rect 57517 1343 57575 1349
rect 57517 1309 57529 1343
rect 57563 1309 57575 1343
rect 57517 1303 57575 1309
rect 57238 1232 57244 1284
rect 57296 1272 57302 1284
rect 57532 1272 57560 1303
rect 57882 1300 57888 1352
rect 57940 1340 57946 1352
rect 58345 1343 58403 1349
rect 58345 1340 58357 1343
rect 57940 1312 58357 1340
rect 57940 1300 57946 1312
rect 58345 1309 58357 1312
rect 58391 1309 58403 1343
rect 58345 1303 58403 1309
rect 59081 1343 59139 1349
rect 59081 1309 59093 1343
rect 59127 1340 59139 1343
rect 59449 1343 59507 1349
rect 59449 1340 59461 1343
rect 59127 1312 59461 1340
rect 59127 1309 59139 1312
rect 59081 1303 59139 1309
rect 59449 1309 59461 1312
rect 59495 1309 59507 1343
rect 59449 1303 59507 1309
rect 60553 1343 60611 1349
rect 60553 1309 60565 1343
rect 60599 1309 60611 1343
rect 60660 1340 60688 1380
rect 60826 1368 60832 1420
rect 60884 1408 60890 1420
rect 61105 1411 61163 1417
rect 60884 1380 60929 1408
rect 60884 1368 60890 1380
rect 61105 1377 61117 1411
rect 61151 1408 61163 1411
rect 62850 1408 62856 1420
rect 61151 1380 62856 1408
rect 61151 1377 61163 1380
rect 61105 1371 61163 1377
rect 62850 1368 62856 1380
rect 62908 1368 62914 1420
rect 63678 1408 63684 1420
rect 63604 1380 63684 1408
rect 61010 1340 61016 1352
rect 60660 1312 61016 1340
rect 60553 1303 60611 1309
rect 57977 1275 58035 1281
rect 57977 1272 57989 1275
rect 57296 1244 57989 1272
rect 57296 1232 57302 1244
rect 57977 1241 57989 1244
rect 58023 1241 58035 1275
rect 60274 1272 60280 1284
rect 57977 1235 58035 1241
rect 58084 1244 60280 1272
rect 58084 1204 58112 1244
rect 60274 1232 60280 1244
rect 60332 1232 60338 1284
rect 56612 1176 58112 1204
rect 58986 1164 58992 1216
rect 59044 1204 59050 1216
rect 59081 1207 59139 1213
rect 59081 1204 59093 1207
rect 59044 1176 59093 1204
rect 59044 1164 59050 1176
rect 59081 1173 59093 1176
rect 59127 1204 59139 1207
rect 59173 1207 59231 1213
rect 59173 1204 59185 1207
rect 59127 1176 59185 1204
rect 59127 1173 59139 1176
rect 59081 1167 59139 1173
rect 59173 1173 59185 1176
rect 59219 1173 59231 1207
rect 60568 1204 60596 1303
rect 61010 1300 61016 1312
rect 61068 1300 61074 1352
rect 61749 1343 61807 1349
rect 61749 1309 61761 1343
rect 61795 1340 61807 1343
rect 62298 1340 62304 1352
rect 61795 1312 62304 1340
rect 61795 1309 61807 1312
rect 61749 1303 61807 1309
rect 62298 1300 62304 1312
rect 62356 1300 62362 1352
rect 63604 1349 63632 1380
rect 63678 1368 63684 1380
rect 63736 1368 63742 1420
rect 65610 1408 65616 1420
rect 65523 1380 65616 1408
rect 65610 1368 65616 1380
rect 65668 1408 65674 1420
rect 66806 1408 66812 1420
rect 65668 1380 66812 1408
rect 65668 1368 65674 1380
rect 66806 1368 66812 1380
rect 66864 1368 66870 1420
rect 67358 1408 67364 1420
rect 67319 1380 67364 1408
rect 67358 1368 67364 1380
rect 67416 1368 67422 1420
rect 68554 1408 68560 1420
rect 68515 1380 68560 1408
rect 68554 1368 68560 1380
rect 68612 1368 68618 1420
rect 68738 1368 68744 1420
rect 68796 1408 68802 1420
rect 72697 1411 72755 1417
rect 72697 1408 72709 1411
rect 68796 1380 72709 1408
rect 68796 1368 68802 1380
rect 72697 1377 72709 1380
rect 72743 1377 72755 1411
rect 72970 1408 72976 1420
rect 72931 1380 72976 1408
rect 72697 1371 72755 1377
rect 72970 1368 72976 1380
rect 73028 1368 73034 1420
rect 74350 1408 74356 1420
rect 74311 1380 74356 1408
rect 74350 1368 74356 1380
rect 74408 1368 74414 1420
rect 76742 1408 76748 1420
rect 74460 1380 76748 1408
rect 63589 1343 63647 1349
rect 63589 1309 63601 1343
rect 63635 1309 63647 1343
rect 63770 1340 63776 1352
rect 63731 1312 63776 1340
rect 63589 1303 63647 1309
rect 63770 1300 63776 1312
rect 63828 1300 63834 1352
rect 63954 1340 63960 1352
rect 63915 1312 63960 1340
rect 63954 1300 63960 1312
rect 64012 1340 64018 1352
rect 64417 1343 64475 1349
rect 64417 1340 64429 1343
rect 64012 1312 64429 1340
rect 64012 1300 64018 1312
rect 64417 1309 64429 1312
rect 64463 1309 64475 1343
rect 64417 1303 64475 1309
rect 65061 1343 65119 1349
rect 65061 1309 65073 1343
rect 65107 1340 65119 1343
rect 65978 1340 65984 1352
rect 65107 1312 65984 1340
rect 65107 1309 65119 1312
rect 65061 1303 65119 1309
rect 65978 1300 65984 1312
rect 66036 1300 66042 1352
rect 66533 1343 66591 1349
rect 66533 1309 66545 1343
rect 66579 1309 66591 1343
rect 66533 1303 66591 1309
rect 66625 1343 66683 1349
rect 66625 1309 66637 1343
rect 66671 1340 66683 1343
rect 67082 1340 67088 1352
rect 66671 1312 67088 1340
rect 66671 1309 66683 1312
rect 66625 1303 66683 1309
rect 60642 1232 60648 1284
rect 60700 1272 60706 1284
rect 60700 1244 60872 1272
rect 60700 1232 60706 1244
rect 60734 1204 60740 1216
rect 60568 1176 60740 1204
rect 59173 1167 59231 1173
rect 60734 1164 60740 1176
rect 60792 1164 60798 1216
rect 60844 1204 60872 1244
rect 61194 1232 61200 1284
rect 61252 1272 61258 1284
rect 66548 1272 66576 1303
rect 67082 1300 67088 1312
rect 67140 1300 67146 1352
rect 67266 1300 67272 1352
rect 67324 1340 67330 1352
rect 67545 1343 67603 1349
rect 67545 1340 67557 1343
rect 67324 1312 67557 1340
rect 67324 1300 67330 1312
rect 67545 1309 67557 1312
rect 67591 1309 67603 1343
rect 67545 1303 67603 1309
rect 69017 1343 69075 1349
rect 69017 1309 69029 1343
rect 69063 1309 69075 1343
rect 70946 1340 70952 1352
rect 70907 1312 70952 1340
rect 69017 1303 69075 1309
rect 66898 1272 66904 1284
rect 61252 1244 65288 1272
rect 66548 1244 66904 1272
rect 61252 1232 61258 1244
rect 61470 1204 61476 1216
rect 60844 1176 61476 1204
rect 61470 1164 61476 1176
rect 61528 1164 61534 1216
rect 62298 1164 62304 1216
rect 62356 1204 62362 1216
rect 62666 1204 62672 1216
rect 62356 1176 62672 1204
rect 62356 1164 62362 1176
rect 62666 1164 62672 1176
rect 62724 1164 62730 1216
rect 65150 1204 65156 1216
rect 65111 1176 65156 1204
rect 65150 1164 65156 1176
rect 65208 1164 65214 1216
rect 65260 1204 65288 1244
rect 66898 1232 66904 1244
rect 66956 1232 66962 1284
rect 69032 1272 69060 1303
rect 70946 1300 70952 1312
rect 71004 1300 71010 1352
rect 71498 1340 71504 1352
rect 71459 1312 71504 1340
rect 71498 1300 71504 1312
rect 71556 1300 71562 1352
rect 71774 1340 71780 1352
rect 71735 1312 71780 1340
rect 71774 1300 71780 1312
rect 71832 1300 71838 1352
rect 72050 1340 72056 1352
rect 72011 1312 72056 1340
rect 72050 1300 72056 1312
rect 72108 1340 72114 1352
rect 72421 1343 72479 1349
rect 72421 1340 72433 1343
rect 72108 1312 72433 1340
rect 72108 1300 72114 1312
rect 72421 1309 72433 1312
rect 72467 1309 72479 1343
rect 72421 1303 72479 1309
rect 72510 1300 72516 1352
rect 72568 1340 72574 1352
rect 72881 1343 72939 1349
rect 72881 1340 72893 1343
rect 72568 1312 72893 1340
rect 72568 1300 72574 1312
rect 72881 1309 72893 1312
rect 72927 1340 72939 1343
rect 74460 1340 74488 1380
rect 76742 1368 76748 1380
rect 76800 1368 76806 1420
rect 77294 1408 77300 1420
rect 77255 1380 77300 1408
rect 77294 1368 77300 1380
rect 77352 1368 77358 1420
rect 78030 1408 78036 1420
rect 77864 1380 78036 1408
rect 72927 1312 74488 1340
rect 74537 1343 74595 1349
rect 72927 1309 72939 1312
rect 72881 1303 72939 1309
rect 74537 1309 74549 1343
rect 74583 1340 74595 1343
rect 76098 1340 76104 1352
rect 74583 1312 74948 1340
rect 76059 1312 76104 1340
rect 74583 1309 74595 1312
rect 74537 1303 74595 1309
rect 69477 1275 69535 1281
rect 69477 1272 69489 1275
rect 67008 1244 68784 1272
rect 69032 1244 69489 1272
rect 67008 1204 67036 1244
rect 65260 1176 67036 1204
rect 67082 1164 67088 1216
rect 67140 1204 67146 1216
rect 68646 1204 68652 1216
rect 67140 1176 68652 1204
rect 67140 1164 67146 1176
rect 68646 1164 68652 1176
rect 68704 1164 68710 1216
rect 68756 1204 68784 1244
rect 69477 1241 69489 1244
rect 69523 1272 69535 1275
rect 73890 1272 73896 1284
rect 69523 1244 73896 1272
rect 69523 1241 69535 1244
rect 69477 1235 69535 1241
rect 73890 1232 73896 1244
rect 73948 1232 73954 1284
rect 71866 1204 71872 1216
rect 68756 1176 71872 1204
rect 71866 1164 71872 1176
rect 71924 1164 71930 1216
rect 72602 1164 72608 1216
rect 72660 1204 72666 1216
rect 73062 1204 73068 1216
rect 72660 1176 73068 1204
rect 72660 1164 72666 1176
rect 73062 1164 73068 1176
rect 73120 1164 73126 1216
rect 74920 1213 74948 1312
rect 76098 1300 76104 1312
rect 76156 1340 76162 1352
rect 77864 1349 77892 1380
rect 78030 1368 78036 1380
rect 78088 1408 78094 1420
rect 83001 1411 83059 1417
rect 78088 1380 82768 1408
rect 78088 1368 78094 1380
rect 76285 1343 76343 1349
rect 76285 1340 76297 1343
rect 76156 1312 76297 1340
rect 76156 1300 76162 1312
rect 76285 1309 76297 1312
rect 76331 1309 76343 1343
rect 76285 1303 76343 1309
rect 77849 1343 77907 1349
rect 77849 1309 77861 1343
rect 77895 1309 77907 1343
rect 79318 1340 79324 1352
rect 79279 1312 79324 1340
rect 77849 1303 77907 1309
rect 79318 1300 79324 1312
rect 79376 1300 79382 1352
rect 79410 1300 79416 1352
rect 79468 1340 79474 1352
rect 79594 1340 79600 1352
rect 79468 1312 79513 1340
rect 79555 1312 79600 1340
rect 79468 1300 79474 1312
rect 79594 1300 79600 1312
rect 79652 1340 79658 1352
rect 80057 1343 80115 1349
rect 80057 1340 80069 1343
rect 79652 1312 80069 1340
rect 79652 1300 79658 1312
rect 80057 1309 80069 1312
rect 80103 1309 80115 1343
rect 80057 1303 80115 1309
rect 80609 1343 80667 1349
rect 80609 1309 80621 1343
rect 80655 1340 80667 1343
rect 81897 1343 81955 1349
rect 80655 1312 80836 1340
rect 80655 1309 80667 1312
rect 80609 1303 80667 1309
rect 80146 1232 80152 1284
rect 80204 1272 80210 1284
rect 80701 1275 80759 1281
rect 80701 1272 80713 1275
rect 80204 1244 80713 1272
rect 80204 1232 80210 1244
rect 80701 1241 80713 1244
rect 80747 1241 80759 1275
rect 80701 1235 80759 1241
rect 74905 1207 74963 1213
rect 74905 1173 74917 1207
rect 74951 1204 74963 1207
rect 75178 1204 75184 1216
rect 74951 1176 75184 1204
rect 74951 1173 74963 1176
rect 74905 1167 74963 1173
rect 75178 1164 75184 1176
rect 75236 1164 75242 1216
rect 78217 1207 78275 1213
rect 78217 1173 78229 1207
rect 78263 1204 78275 1207
rect 78582 1204 78588 1216
rect 78263 1176 78588 1204
rect 78263 1173 78275 1176
rect 78217 1167 78275 1173
rect 78582 1164 78588 1176
rect 78640 1164 78646 1216
rect 78953 1207 79011 1213
rect 78953 1173 78965 1207
rect 78999 1204 79011 1207
rect 79042 1204 79048 1216
rect 78999 1176 79048 1204
rect 78999 1173 79011 1176
rect 78953 1167 79011 1173
rect 79042 1164 79048 1176
rect 79100 1204 79106 1216
rect 79962 1204 79968 1216
rect 79100 1176 79968 1204
rect 79100 1164 79106 1176
rect 79962 1164 79968 1176
rect 80020 1164 80026 1216
rect 80517 1207 80575 1213
rect 80517 1173 80529 1207
rect 80563 1204 80575 1207
rect 80808 1204 80836 1312
rect 81897 1309 81909 1343
rect 81943 1340 81955 1343
rect 82740 1340 82768 1380
rect 83001 1377 83013 1411
rect 83047 1408 83059 1411
rect 83090 1408 83096 1420
rect 83047 1380 83096 1408
rect 83047 1377 83059 1380
rect 83001 1371 83059 1377
rect 83090 1368 83096 1380
rect 83148 1368 83154 1420
rect 84194 1408 84200 1420
rect 84155 1380 84200 1408
rect 84194 1368 84200 1380
rect 84252 1368 84258 1420
rect 85040 1408 85068 1516
rect 87414 1504 87420 1516
rect 87472 1504 87478 1556
rect 91189 1547 91247 1553
rect 91189 1513 91201 1547
rect 91235 1544 91247 1547
rect 91278 1544 91284 1556
rect 91235 1516 91284 1544
rect 91235 1513 91247 1516
rect 91189 1507 91247 1513
rect 91278 1504 91284 1516
rect 91336 1504 91342 1556
rect 92290 1504 92296 1556
rect 92348 1544 92354 1556
rect 98641 1547 98699 1553
rect 98641 1544 98653 1547
rect 92348 1516 98653 1544
rect 92348 1504 92354 1516
rect 98641 1513 98653 1516
rect 98687 1513 98699 1547
rect 98641 1507 98699 1513
rect 99190 1504 99196 1556
rect 99248 1544 99254 1556
rect 99248 1516 101720 1544
rect 99248 1504 99254 1516
rect 100202 1476 100208 1488
rect 84304 1380 85068 1408
rect 85132 1448 100208 1476
rect 84304 1340 84332 1380
rect 84562 1340 84568 1352
rect 81943 1312 82676 1340
rect 82740 1312 84332 1340
rect 84523 1312 84568 1340
rect 81943 1309 81955 1312
rect 81897 1303 81955 1309
rect 81342 1272 81348 1284
rect 81303 1244 81348 1272
rect 81342 1232 81348 1244
rect 81400 1232 81406 1284
rect 81526 1232 81532 1284
rect 81584 1272 81590 1284
rect 82170 1272 82176 1284
rect 81584 1244 82176 1272
rect 81584 1232 81590 1244
rect 82170 1232 82176 1244
rect 82228 1272 82234 1284
rect 82357 1275 82415 1281
rect 82357 1272 82369 1275
rect 82228 1244 82369 1272
rect 82228 1232 82234 1244
rect 82357 1241 82369 1244
rect 82403 1241 82415 1275
rect 82357 1235 82415 1241
rect 82648 1216 82676 1312
rect 84562 1300 84568 1312
rect 84620 1300 84626 1352
rect 84749 1343 84807 1349
rect 84749 1309 84761 1343
rect 84795 1340 84807 1343
rect 85132 1340 85160 1448
rect 100202 1436 100208 1448
rect 100260 1436 100266 1488
rect 101692 1476 101720 1516
rect 101766 1504 101772 1556
rect 101824 1544 101830 1556
rect 102502 1544 102508 1556
rect 101824 1516 102508 1544
rect 101824 1504 101830 1516
rect 102502 1504 102508 1516
rect 102560 1504 102566 1556
rect 104342 1504 104348 1556
rect 104400 1544 104406 1556
rect 104529 1547 104587 1553
rect 104529 1544 104541 1547
rect 104400 1516 104541 1544
rect 104400 1504 104406 1516
rect 104529 1513 104541 1516
rect 104575 1513 104587 1547
rect 104529 1507 104587 1513
rect 105262 1504 105268 1556
rect 105320 1544 105326 1556
rect 105817 1547 105875 1553
rect 105817 1544 105829 1547
rect 105320 1516 105829 1544
rect 105320 1504 105326 1516
rect 105817 1513 105829 1516
rect 105863 1513 105875 1547
rect 105817 1507 105875 1513
rect 107930 1504 107936 1556
rect 107988 1544 107994 1556
rect 110966 1544 110972 1556
rect 107988 1516 110972 1544
rect 107988 1504 107994 1516
rect 110966 1504 110972 1516
rect 111024 1504 111030 1556
rect 112530 1504 112536 1556
rect 112588 1544 112594 1556
rect 117406 1544 117412 1556
rect 112588 1516 117412 1544
rect 112588 1504 112594 1516
rect 117406 1504 117412 1516
rect 117464 1504 117470 1556
rect 117682 1504 117688 1556
rect 117740 1544 117746 1556
rect 117961 1547 118019 1553
rect 117961 1544 117973 1547
rect 117740 1516 117973 1544
rect 117740 1504 117746 1516
rect 117961 1513 117973 1516
rect 118007 1544 118019 1547
rect 118050 1544 118056 1556
rect 118007 1516 118056 1544
rect 118007 1513 118019 1516
rect 117961 1507 118019 1513
rect 118050 1504 118056 1516
rect 118108 1504 118114 1556
rect 118786 1504 118792 1556
rect 118844 1544 118850 1556
rect 135898 1544 135904 1556
rect 118844 1516 135904 1544
rect 118844 1504 118850 1516
rect 135898 1504 135904 1516
rect 135956 1504 135962 1556
rect 137554 1544 137560 1556
rect 137515 1516 137560 1544
rect 137554 1504 137560 1516
rect 137612 1504 137618 1556
rect 138477 1547 138535 1553
rect 138477 1513 138489 1547
rect 138523 1544 138535 1547
rect 138750 1544 138756 1556
rect 138523 1516 138756 1544
rect 138523 1513 138535 1516
rect 138477 1507 138535 1513
rect 138750 1504 138756 1516
rect 138808 1504 138814 1556
rect 143166 1504 143172 1556
rect 143224 1544 143230 1556
rect 143353 1547 143411 1553
rect 143353 1544 143365 1547
rect 143224 1516 143365 1544
rect 143224 1504 143230 1516
rect 143353 1513 143365 1516
rect 143399 1513 143411 1547
rect 158162 1544 158168 1556
rect 158123 1516 158168 1544
rect 143353 1507 143411 1513
rect 158162 1504 158168 1516
rect 158220 1504 158226 1556
rect 159818 1504 159824 1556
rect 159876 1544 159882 1556
rect 160097 1547 160155 1553
rect 160097 1544 160109 1547
rect 159876 1516 160109 1544
rect 159876 1504 159882 1516
rect 160097 1513 160109 1516
rect 160143 1513 160155 1547
rect 160097 1507 160155 1513
rect 164878 1504 164884 1556
rect 164936 1544 164942 1556
rect 166074 1544 166080 1556
rect 164936 1516 166080 1544
rect 164936 1504 164942 1516
rect 166074 1504 166080 1516
rect 166132 1504 166138 1556
rect 126146 1476 126152 1488
rect 101692 1448 118556 1476
rect 85666 1368 85672 1420
rect 85724 1408 85730 1420
rect 86313 1411 86371 1417
rect 86313 1408 86325 1411
rect 85724 1380 86325 1408
rect 85724 1368 85730 1380
rect 86313 1377 86325 1380
rect 86359 1408 86371 1411
rect 87414 1408 87420 1420
rect 86359 1380 87420 1408
rect 86359 1377 86371 1380
rect 86313 1371 86371 1377
rect 87414 1368 87420 1380
rect 87472 1368 87478 1420
rect 88886 1408 88892 1420
rect 88847 1380 88892 1408
rect 88886 1368 88892 1380
rect 88944 1368 88950 1420
rect 89714 1368 89720 1420
rect 89772 1408 89778 1420
rect 89901 1411 89959 1417
rect 89901 1408 89913 1411
rect 89772 1380 89913 1408
rect 89772 1368 89778 1380
rect 89901 1377 89913 1380
rect 89947 1377 89959 1411
rect 89901 1371 89959 1377
rect 91922 1368 91928 1420
rect 91980 1408 91986 1420
rect 92201 1411 92259 1417
rect 92201 1408 92213 1411
rect 91980 1380 92213 1408
rect 91980 1368 91986 1380
rect 92201 1377 92213 1380
rect 92247 1408 92259 1411
rect 99466 1408 99472 1420
rect 92247 1380 99472 1408
rect 92247 1377 92259 1380
rect 92201 1371 92259 1377
rect 99466 1368 99472 1380
rect 99524 1368 99530 1420
rect 99558 1368 99564 1420
rect 99616 1408 99622 1420
rect 100570 1408 100576 1420
rect 99616 1380 100576 1408
rect 99616 1368 99622 1380
rect 100570 1368 100576 1380
rect 100628 1368 100634 1420
rect 102318 1408 102324 1420
rect 100680 1380 102180 1408
rect 102279 1380 102324 1408
rect 84795 1312 85160 1340
rect 85393 1343 85451 1349
rect 84795 1309 84807 1312
rect 84749 1303 84807 1309
rect 85393 1309 85405 1343
rect 85439 1309 85451 1343
rect 85393 1303 85451 1309
rect 86405 1343 86463 1349
rect 86405 1309 86417 1343
rect 86451 1340 86463 1343
rect 87230 1340 87236 1352
rect 86451 1312 87000 1340
rect 87191 1312 87236 1340
rect 86451 1309 86463 1312
rect 86405 1303 86463 1309
rect 85408 1272 85436 1303
rect 86972 1281 87000 1312
rect 87230 1300 87236 1312
rect 87288 1300 87294 1352
rect 87509 1343 87567 1349
rect 87509 1309 87521 1343
rect 87555 1340 87567 1343
rect 88426 1340 88432 1352
rect 87555 1312 88104 1340
rect 88387 1312 88432 1340
rect 87555 1309 87567 1312
rect 87509 1303 87567 1309
rect 85945 1275 86003 1281
rect 85945 1272 85957 1275
rect 85408 1244 85957 1272
rect 85945 1241 85957 1244
rect 85991 1272 86003 1275
rect 86957 1275 87015 1281
rect 85991 1244 86632 1272
rect 85991 1241 86003 1244
rect 85945 1235 86003 1241
rect 81158 1204 81164 1216
rect 80563 1176 81164 1204
rect 80563 1173 80575 1176
rect 80517 1167 80575 1173
rect 81158 1164 81164 1176
rect 81216 1164 81222 1216
rect 81986 1204 81992 1216
rect 81947 1176 81992 1204
rect 81986 1164 81992 1176
rect 82044 1164 82050 1216
rect 82630 1164 82636 1216
rect 82688 1204 82694 1216
rect 82725 1207 82783 1213
rect 82725 1204 82737 1207
rect 82688 1176 82737 1204
rect 82688 1164 82694 1176
rect 82725 1173 82737 1176
rect 82771 1173 82783 1207
rect 85482 1204 85488 1216
rect 85443 1176 85488 1204
rect 82725 1167 82783 1173
rect 85482 1164 85488 1176
rect 85540 1164 85546 1216
rect 86494 1204 86500 1216
rect 86455 1176 86500 1204
rect 86494 1164 86500 1176
rect 86552 1164 86558 1216
rect 86604 1204 86632 1244
rect 86957 1241 86969 1275
rect 87003 1272 87015 1275
rect 87782 1272 87788 1284
rect 87003 1244 87788 1272
rect 87003 1241 87015 1244
rect 86957 1235 87015 1241
rect 87782 1232 87788 1244
rect 87840 1232 87846 1284
rect 87046 1204 87052 1216
rect 86604 1176 87052 1204
rect 87046 1164 87052 1176
rect 87104 1164 87110 1216
rect 87598 1204 87604 1216
rect 87559 1176 87604 1204
rect 87598 1164 87604 1176
rect 87656 1164 87662 1216
rect 88076 1213 88104 1312
rect 88426 1300 88432 1312
rect 88484 1300 88490 1352
rect 90174 1300 90180 1352
rect 90232 1340 90238 1352
rect 90453 1343 90511 1349
rect 90453 1340 90465 1343
rect 90232 1312 90465 1340
rect 90232 1300 90238 1312
rect 90453 1309 90465 1312
rect 90499 1340 90511 1343
rect 90729 1343 90787 1349
rect 90729 1340 90741 1343
rect 90499 1312 90741 1340
rect 90499 1309 90511 1312
rect 90453 1303 90511 1309
rect 90729 1309 90741 1312
rect 90775 1309 90787 1343
rect 90729 1303 90787 1309
rect 91094 1300 91100 1352
rect 91152 1340 91158 1352
rect 91281 1343 91339 1349
rect 91281 1340 91293 1343
rect 91152 1312 91293 1340
rect 91152 1300 91158 1312
rect 91281 1309 91293 1312
rect 91327 1340 91339 1343
rect 91741 1343 91799 1349
rect 91741 1340 91753 1343
rect 91327 1312 91753 1340
rect 91327 1309 91339 1312
rect 91281 1303 91339 1309
rect 91741 1309 91753 1312
rect 91787 1309 91799 1343
rect 91741 1303 91799 1309
rect 94774 1300 94780 1352
rect 94832 1340 94838 1352
rect 100680 1340 100708 1380
rect 94832 1312 100708 1340
rect 102152 1340 102180 1380
rect 102318 1368 102324 1380
rect 102376 1368 102382 1420
rect 103514 1408 103520 1420
rect 102428 1380 103376 1408
rect 103475 1380 103520 1408
rect 102428 1340 102456 1380
rect 102152 1312 102456 1340
rect 103348 1340 103376 1380
rect 103514 1368 103520 1380
rect 103572 1368 103578 1420
rect 106366 1408 106372 1420
rect 103624 1380 106372 1408
rect 103624 1340 103652 1380
rect 106366 1368 106372 1380
rect 106424 1368 106430 1420
rect 106918 1408 106924 1420
rect 106879 1380 106924 1408
rect 106918 1368 106924 1380
rect 106976 1368 106982 1420
rect 107746 1368 107752 1420
rect 107804 1408 107810 1420
rect 107841 1411 107899 1417
rect 107841 1408 107853 1411
rect 107804 1380 107853 1408
rect 107804 1368 107810 1380
rect 107841 1377 107853 1380
rect 107887 1408 107899 1411
rect 109218 1408 109224 1420
rect 107887 1380 109224 1408
rect 107887 1377 107899 1380
rect 107841 1371 107899 1377
rect 109218 1368 109224 1380
rect 109276 1368 109282 1420
rect 110693 1411 110751 1417
rect 110693 1377 110705 1411
rect 110739 1408 110751 1411
rect 110782 1408 110788 1420
rect 110739 1380 110788 1408
rect 110739 1377 110751 1380
rect 110693 1371 110751 1377
rect 110782 1368 110788 1380
rect 110840 1368 110846 1420
rect 111794 1368 111800 1420
rect 111852 1408 111858 1420
rect 112438 1408 112444 1420
rect 111852 1380 112444 1408
rect 111852 1368 111858 1380
rect 112438 1368 112444 1380
rect 112496 1368 112502 1420
rect 112622 1408 112628 1420
rect 112583 1380 112628 1408
rect 112622 1368 112628 1380
rect 112680 1368 112686 1420
rect 113818 1408 113824 1420
rect 113779 1380 113824 1408
rect 113818 1368 113824 1380
rect 113876 1408 113882 1420
rect 114005 1411 114063 1417
rect 114005 1408 114017 1411
rect 113876 1380 114017 1408
rect 113876 1368 113882 1380
rect 114005 1377 114017 1380
rect 114051 1377 114063 1411
rect 114005 1371 114063 1377
rect 115014 1368 115020 1420
rect 115072 1408 115078 1420
rect 116210 1408 116216 1420
rect 115072 1380 116216 1408
rect 115072 1368 115078 1380
rect 116210 1368 116216 1380
rect 116268 1408 116274 1420
rect 116673 1411 116731 1417
rect 116673 1408 116685 1411
rect 116268 1380 116685 1408
rect 116268 1368 116274 1380
rect 116673 1377 116685 1380
rect 116719 1377 116731 1411
rect 116673 1371 116731 1377
rect 117409 1411 117467 1417
rect 117409 1377 117421 1411
rect 117455 1408 117467 1411
rect 118418 1408 118424 1420
rect 117455 1380 118424 1408
rect 117455 1377 117467 1380
rect 117409 1371 117467 1377
rect 118418 1368 118424 1380
rect 118476 1368 118482 1420
rect 103348 1312 103652 1340
rect 103885 1343 103943 1349
rect 94832 1300 94838 1312
rect 103885 1309 103897 1343
rect 103931 1309 103943 1343
rect 103885 1303 103943 1309
rect 104989 1343 105047 1349
rect 104989 1309 105001 1343
rect 105035 1340 105047 1343
rect 105035 1312 105216 1340
rect 105035 1309 105047 1312
rect 104989 1303 105047 1309
rect 96246 1232 96252 1284
rect 96304 1272 96310 1284
rect 102226 1272 102232 1284
rect 96304 1244 102232 1272
rect 96304 1232 96310 1244
rect 102226 1232 102232 1244
rect 102284 1232 102290 1284
rect 103900 1272 103928 1303
rect 104253 1275 104311 1281
rect 104253 1272 104265 1275
rect 103900 1244 104265 1272
rect 104253 1241 104265 1244
rect 104299 1272 104311 1275
rect 105081 1275 105139 1281
rect 105081 1272 105093 1275
rect 104299 1244 105093 1272
rect 104299 1241 104311 1244
rect 104253 1235 104311 1241
rect 105081 1241 105093 1244
rect 105127 1241 105139 1275
rect 105081 1235 105139 1241
rect 105188 1272 105216 1312
rect 105262 1300 105268 1352
rect 105320 1340 105326 1352
rect 106001 1343 106059 1349
rect 106001 1340 106013 1343
rect 105320 1312 106013 1340
rect 105320 1300 105326 1312
rect 106001 1309 106013 1312
rect 106047 1340 106059 1343
rect 106461 1343 106519 1349
rect 106461 1340 106473 1343
rect 106047 1312 106473 1340
rect 106047 1309 106059 1312
rect 106001 1303 106059 1309
rect 106461 1309 106473 1312
rect 106507 1309 106519 1343
rect 109034 1340 109040 1352
rect 108995 1312 109040 1340
rect 106461 1303 106519 1309
rect 109034 1300 109040 1312
rect 109092 1300 109098 1352
rect 109770 1340 109776 1352
rect 109144 1312 109776 1340
rect 105449 1275 105507 1281
rect 105449 1272 105461 1275
rect 105188 1244 105461 1272
rect 88061 1207 88119 1213
rect 88061 1173 88073 1207
rect 88107 1204 88119 1207
rect 88150 1204 88156 1216
rect 88107 1176 88156 1204
rect 88107 1173 88119 1176
rect 88061 1167 88119 1173
rect 88150 1164 88156 1176
rect 88208 1164 88214 1216
rect 89990 1164 89996 1216
rect 90048 1204 90054 1216
rect 91094 1204 91100 1216
rect 90048 1176 91100 1204
rect 90048 1164 90054 1176
rect 91094 1164 91100 1176
rect 91152 1164 91158 1216
rect 91370 1204 91376 1216
rect 91331 1176 91376 1204
rect 91370 1164 91376 1176
rect 91428 1164 91434 1216
rect 94038 1164 94044 1216
rect 94096 1204 94102 1216
rect 105188 1204 105216 1244
rect 105449 1241 105461 1244
rect 105495 1241 105507 1275
rect 105449 1235 105507 1241
rect 105814 1232 105820 1284
rect 105872 1272 105878 1284
rect 108485 1275 108543 1281
rect 105872 1244 107148 1272
rect 105872 1232 105878 1244
rect 106090 1204 106096 1216
rect 94096 1176 105216 1204
rect 106051 1176 106096 1204
rect 94096 1164 94102 1176
rect 106090 1164 106096 1176
rect 106148 1164 106154 1216
rect 107010 1204 107016 1216
rect 106971 1176 107016 1204
rect 107010 1164 107016 1176
rect 107068 1164 107074 1216
rect 107120 1204 107148 1244
rect 108485 1241 108497 1275
rect 108531 1272 108543 1275
rect 109144 1272 109172 1312
rect 109770 1300 109776 1312
rect 109828 1340 109834 1352
rect 109957 1343 110015 1349
rect 109957 1340 109969 1343
rect 109828 1312 109969 1340
rect 109828 1300 109834 1312
rect 109957 1309 109969 1312
rect 110003 1309 110015 1343
rect 109957 1303 110015 1309
rect 110601 1343 110659 1349
rect 110601 1309 110613 1343
rect 110647 1309 110659 1343
rect 110601 1303 110659 1309
rect 108531 1244 109172 1272
rect 108531 1241 108543 1244
rect 108485 1235 108543 1241
rect 109218 1232 109224 1284
rect 109276 1272 109282 1284
rect 109276 1244 109356 1272
rect 109276 1232 109282 1244
rect 109034 1204 109040 1216
rect 107120 1176 109040 1204
rect 109034 1164 109040 1176
rect 109092 1164 109098 1216
rect 109328 1204 109356 1244
rect 109402 1232 109408 1284
rect 109460 1272 109466 1284
rect 110608 1272 110636 1303
rect 111242 1300 111248 1352
rect 111300 1340 111306 1352
rect 111610 1340 111616 1352
rect 111300 1312 111616 1340
rect 111300 1300 111306 1312
rect 111610 1300 111616 1312
rect 111668 1300 111674 1352
rect 112254 1300 112260 1352
rect 112312 1340 112318 1352
rect 112717 1343 112775 1349
rect 112717 1340 112729 1343
rect 112312 1312 112729 1340
rect 112312 1300 112318 1312
rect 112717 1309 112729 1312
rect 112763 1340 112775 1343
rect 113453 1343 113511 1349
rect 113453 1340 113465 1343
rect 112763 1312 113465 1340
rect 112763 1309 112775 1312
rect 112717 1303 112775 1309
rect 113453 1309 113465 1312
rect 113499 1309 113511 1343
rect 118528 1340 118556 1448
rect 119540 1448 124996 1476
rect 126107 1448 126152 1476
rect 118878 1368 118884 1420
rect 118936 1408 118942 1420
rect 119433 1411 119491 1417
rect 119433 1408 119445 1411
rect 118936 1380 119445 1408
rect 118936 1368 118942 1380
rect 119433 1377 119445 1380
rect 119479 1377 119491 1411
rect 119433 1371 119491 1377
rect 119540 1340 119568 1448
rect 119706 1368 119712 1420
rect 119764 1408 119770 1420
rect 120994 1408 121000 1420
rect 119764 1380 120856 1408
rect 120955 1380 121000 1408
rect 119764 1368 119770 1380
rect 119890 1340 119896 1352
rect 113453 1303 113511 1309
rect 113560 1312 118280 1340
rect 118528 1312 119568 1340
rect 119851 1312 119896 1340
rect 111061 1275 111119 1281
rect 111061 1272 111073 1275
rect 109460 1244 111073 1272
rect 109460 1232 109466 1244
rect 111061 1241 111073 1244
rect 111107 1241 111119 1275
rect 111061 1235 111119 1241
rect 111334 1232 111340 1284
rect 111392 1272 111398 1284
rect 111521 1275 111579 1281
rect 111521 1272 111533 1275
rect 111392 1244 111533 1272
rect 111392 1232 111398 1244
rect 111521 1241 111533 1244
rect 111567 1272 111579 1275
rect 113560 1272 113588 1312
rect 111567 1244 113588 1272
rect 111567 1241 111579 1244
rect 111521 1235 111579 1241
rect 114094 1232 114100 1284
rect 114152 1272 114158 1284
rect 118142 1272 118148 1284
rect 114152 1244 118148 1272
rect 114152 1232 114158 1244
rect 118142 1232 118148 1244
rect 118200 1232 118206 1284
rect 118252 1272 118280 1312
rect 119890 1300 119896 1312
rect 119948 1300 119954 1352
rect 120350 1340 120356 1352
rect 120311 1312 120356 1340
rect 120350 1300 120356 1312
rect 120408 1300 120414 1352
rect 120828 1340 120856 1380
rect 120994 1368 121000 1380
rect 121052 1368 121058 1420
rect 123938 1408 123944 1420
rect 121104 1380 123800 1408
rect 123899 1380 123944 1408
rect 121104 1340 121132 1380
rect 120828 1312 121132 1340
rect 121825 1343 121883 1349
rect 121825 1309 121837 1343
rect 121871 1340 121883 1343
rect 122282 1340 122288 1352
rect 121871 1312 122288 1340
rect 121871 1309 121883 1312
rect 121825 1303 121883 1309
rect 122282 1300 122288 1312
rect 122340 1300 122346 1352
rect 123772 1340 123800 1380
rect 123938 1368 123944 1380
rect 123996 1368 124002 1420
rect 124968 1417 124996 1448
rect 126146 1436 126152 1448
rect 126204 1476 126210 1488
rect 126204 1448 126376 1476
rect 126204 1436 126210 1448
rect 124953 1411 125011 1417
rect 124048 1380 124904 1408
rect 124048 1340 124076 1380
rect 123772 1312 124076 1340
rect 124876 1340 124904 1380
rect 124953 1377 124965 1411
rect 124999 1377 125011 1411
rect 126238 1408 126244 1420
rect 124953 1371 125011 1377
rect 125060 1380 126244 1408
rect 125060 1340 125088 1380
rect 126238 1368 126244 1380
rect 126296 1368 126302 1420
rect 126348 1417 126376 1448
rect 130654 1436 130660 1488
rect 130712 1476 130718 1488
rect 135254 1476 135260 1488
rect 130712 1448 135260 1476
rect 130712 1436 130718 1448
rect 135254 1436 135260 1448
rect 135312 1436 135318 1488
rect 139854 1436 139860 1488
rect 139912 1476 139918 1488
rect 139912 1448 142200 1476
rect 139912 1436 139918 1448
rect 126333 1411 126391 1417
rect 126333 1377 126345 1411
rect 126379 1377 126391 1411
rect 129182 1408 129188 1420
rect 129143 1380 129188 1408
rect 126333 1371 126391 1377
rect 129182 1368 129188 1380
rect 129240 1368 129246 1420
rect 129826 1368 129832 1420
rect 129884 1408 129890 1420
rect 130197 1411 130255 1417
rect 130197 1408 130209 1411
rect 129884 1380 130209 1408
rect 129884 1368 129890 1380
rect 130197 1377 130209 1380
rect 130243 1377 130255 1411
rect 133693 1411 133751 1417
rect 133693 1408 133705 1411
rect 130197 1371 130255 1377
rect 133156 1380 133705 1408
rect 124876 1312 125088 1340
rect 125505 1343 125563 1349
rect 125505 1309 125517 1343
rect 125551 1340 125563 1343
rect 125778 1340 125784 1352
rect 125551 1312 125784 1340
rect 125551 1309 125563 1312
rect 125505 1303 125563 1309
rect 125778 1300 125784 1312
rect 125836 1300 125842 1352
rect 130749 1343 130807 1349
rect 130749 1309 130761 1343
rect 130795 1340 130807 1343
rect 131022 1340 131028 1352
rect 130795 1312 131028 1340
rect 130795 1309 130807 1312
rect 130749 1303 130807 1309
rect 131022 1300 131028 1312
rect 131080 1300 131086 1352
rect 133156 1349 133184 1380
rect 133693 1377 133705 1380
rect 133739 1408 133751 1411
rect 134610 1408 134616 1420
rect 133739 1380 134616 1408
rect 133739 1377 133751 1380
rect 133693 1371 133751 1377
rect 134610 1368 134616 1380
rect 134668 1368 134674 1420
rect 135346 1408 135352 1420
rect 135307 1380 135352 1408
rect 135346 1368 135352 1380
rect 135404 1368 135410 1420
rect 135438 1368 135444 1420
rect 135496 1408 135502 1420
rect 136361 1411 136419 1417
rect 136361 1408 136373 1411
rect 135496 1380 136373 1408
rect 135496 1368 135502 1380
rect 136361 1377 136373 1380
rect 136407 1377 136419 1411
rect 138658 1408 138664 1420
rect 136361 1371 136419 1377
rect 136468 1380 137324 1408
rect 138619 1380 138664 1408
rect 131945 1343 132003 1349
rect 131945 1309 131957 1343
rect 131991 1340 132003 1343
rect 132221 1343 132279 1349
rect 132221 1340 132233 1343
rect 131991 1312 132233 1340
rect 131991 1309 132003 1312
rect 131945 1303 132003 1309
rect 132221 1309 132233 1312
rect 132267 1309 132279 1343
rect 132221 1303 132279 1309
rect 133141 1343 133199 1349
rect 133141 1309 133153 1343
rect 133187 1309 133199 1343
rect 136468 1340 136496 1380
rect 136634 1340 136640 1352
rect 133141 1303 133199 1309
rect 133340 1312 136496 1340
rect 136595 1312 136640 1340
rect 133233 1275 133291 1281
rect 133233 1272 133245 1275
rect 118252 1244 133245 1272
rect 133233 1241 133245 1244
rect 133279 1241 133291 1275
rect 133233 1235 133291 1241
rect 109497 1207 109555 1213
rect 109497 1204 109509 1207
rect 109328 1176 109509 1204
rect 109497 1173 109509 1176
rect 109543 1173 109555 1207
rect 109497 1167 109555 1173
rect 109678 1164 109684 1216
rect 109736 1204 109742 1216
rect 111150 1204 111156 1216
rect 109736 1176 111156 1204
rect 109736 1164 109742 1176
rect 111150 1164 111156 1176
rect 111208 1164 111214 1216
rect 114002 1164 114008 1216
rect 114060 1204 114066 1216
rect 115017 1207 115075 1213
rect 115017 1204 115029 1207
rect 114060 1176 115029 1204
rect 114060 1164 114066 1176
rect 115017 1173 115029 1176
rect 115063 1173 115075 1207
rect 115566 1204 115572 1216
rect 115527 1176 115572 1204
rect 115017 1167 115075 1173
rect 115566 1164 115572 1176
rect 115624 1164 115630 1216
rect 116210 1204 116216 1216
rect 116171 1176 116216 1204
rect 116210 1164 116216 1176
rect 116268 1164 116274 1216
rect 116302 1164 116308 1216
rect 116360 1204 116366 1216
rect 121917 1207 121975 1213
rect 121917 1204 121929 1207
rect 116360 1176 121929 1204
rect 116360 1164 116366 1176
rect 121917 1173 121929 1176
rect 121963 1173 121975 1207
rect 121917 1167 121975 1173
rect 122834 1164 122840 1216
rect 122892 1204 122898 1216
rect 122929 1207 122987 1213
rect 122929 1204 122941 1207
rect 122892 1176 122941 1204
rect 122892 1164 122898 1176
rect 122929 1173 122941 1176
rect 122975 1204 122987 1207
rect 124122 1204 124128 1216
rect 122975 1176 124128 1204
rect 122975 1173 122987 1176
rect 122929 1167 122987 1173
rect 124122 1164 124128 1176
rect 124180 1164 124186 1216
rect 126974 1204 126980 1216
rect 126935 1176 126980 1204
rect 126974 1164 126980 1176
rect 127032 1164 127038 1216
rect 128262 1204 128268 1216
rect 128223 1176 128268 1204
rect 128262 1164 128268 1176
rect 128320 1164 128326 1216
rect 131117 1207 131175 1213
rect 131117 1173 131129 1207
rect 131163 1204 131175 1207
rect 131206 1204 131212 1216
rect 131163 1176 131212 1204
rect 131163 1173 131175 1176
rect 131117 1167 131175 1173
rect 131206 1164 131212 1176
rect 131264 1164 131270 1216
rect 132034 1204 132040 1216
rect 131995 1176 132040 1204
rect 132034 1164 132040 1176
rect 132092 1164 132098 1216
rect 132221 1207 132279 1213
rect 132221 1173 132233 1207
rect 132267 1204 132279 1207
rect 132497 1207 132555 1213
rect 132497 1204 132509 1207
rect 132267 1176 132509 1204
rect 132267 1173 132279 1176
rect 132221 1167 132279 1173
rect 132497 1173 132509 1176
rect 132543 1204 132555 1207
rect 133340 1204 133368 1312
rect 136634 1300 136640 1312
rect 136692 1340 136698 1352
rect 137189 1343 137247 1349
rect 137189 1340 137201 1343
rect 136692 1312 137201 1340
rect 136692 1300 136698 1312
rect 137189 1309 137201 1312
rect 137235 1309 137247 1343
rect 137296 1340 137324 1380
rect 138658 1368 138664 1380
rect 138716 1368 138722 1420
rect 139946 1408 139952 1420
rect 139907 1380 139952 1408
rect 139946 1368 139952 1380
rect 140004 1368 140010 1420
rect 141142 1408 141148 1420
rect 141103 1380 141148 1408
rect 141142 1368 141148 1380
rect 141200 1368 141206 1420
rect 142172 1417 142200 1448
rect 151906 1436 151912 1488
rect 151964 1476 151970 1488
rect 151964 1448 159312 1476
rect 151964 1436 151970 1448
rect 142157 1411 142215 1417
rect 142157 1377 142169 1411
rect 142203 1377 142215 1411
rect 147858 1408 147864 1420
rect 147819 1380 147864 1408
rect 142157 1371 142215 1377
rect 147858 1368 147864 1380
rect 147916 1408 147922 1420
rect 148321 1411 148379 1417
rect 148321 1408 148333 1411
rect 147916 1380 148333 1408
rect 147916 1368 147922 1380
rect 148321 1377 148333 1380
rect 148367 1377 148379 1411
rect 148321 1371 148379 1377
rect 148502 1368 148508 1420
rect 148560 1408 148566 1420
rect 150250 1408 150256 1420
rect 148560 1380 150256 1408
rect 148560 1368 148566 1380
rect 150250 1368 150256 1380
rect 150308 1408 150314 1420
rect 150345 1411 150403 1417
rect 150345 1408 150357 1411
rect 150308 1380 150357 1408
rect 150308 1368 150314 1380
rect 150345 1377 150357 1380
rect 150391 1377 150403 1411
rect 156782 1408 156788 1420
rect 156743 1380 156788 1408
rect 150345 1371 150403 1377
rect 156782 1368 156788 1380
rect 156840 1368 156846 1420
rect 159284 1417 159312 1448
rect 159269 1411 159327 1417
rect 159269 1377 159281 1411
rect 159315 1377 159327 1411
rect 159269 1371 159327 1377
rect 163958 1368 163964 1420
rect 164016 1408 164022 1420
rect 165430 1408 165436 1420
rect 164016 1380 164464 1408
rect 165391 1380 165436 1408
rect 164016 1368 164022 1380
rect 137296 1312 138980 1340
rect 137189 1303 137247 1309
rect 134610 1232 134616 1284
rect 134668 1272 134674 1284
rect 138952 1272 138980 1312
rect 139670 1300 139676 1352
rect 139728 1340 139734 1352
rect 139765 1343 139823 1349
rect 139765 1340 139777 1343
rect 139728 1312 139777 1340
rect 139728 1300 139734 1312
rect 139765 1309 139777 1312
rect 139811 1340 139823 1343
rect 140501 1343 140559 1349
rect 140501 1340 140513 1343
rect 139811 1312 140513 1340
rect 139811 1309 139823 1312
rect 139765 1303 139823 1309
rect 140501 1309 140513 1312
rect 140547 1309 140559 1343
rect 140501 1303 140559 1309
rect 142709 1343 142767 1349
rect 142709 1309 142721 1343
rect 142755 1340 142767 1343
rect 142985 1343 143043 1349
rect 142985 1340 142997 1343
rect 142755 1312 142997 1340
rect 142755 1309 142767 1312
rect 142709 1303 142767 1309
rect 142985 1309 142997 1312
rect 143031 1340 143043 1343
rect 143166 1340 143172 1352
rect 143031 1312 143172 1340
rect 143031 1309 143043 1312
rect 142985 1303 143043 1309
rect 143166 1300 143172 1312
rect 143224 1300 143230 1352
rect 144914 1340 144920 1352
rect 144875 1312 144920 1340
rect 144914 1300 144920 1312
rect 144972 1340 144978 1352
rect 145377 1343 145435 1349
rect 145377 1340 145389 1343
rect 144972 1312 145389 1340
rect 144972 1300 144978 1312
rect 145377 1309 145389 1312
rect 145423 1309 145435 1343
rect 145377 1303 145435 1309
rect 145742 1300 145748 1352
rect 145800 1340 145806 1352
rect 145929 1343 145987 1349
rect 145929 1340 145941 1343
rect 145800 1312 145941 1340
rect 145800 1300 145806 1312
rect 145929 1309 145941 1312
rect 145975 1340 145987 1343
rect 146389 1343 146447 1349
rect 146389 1340 146401 1343
rect 145975 1312 146401 1340
rect 145975 1309 145987 1312
rect 145929 1303 145987 1309
rect 146389 1309 146401 1312
rect 146435 1309 146447 1343
rect 146389 1303 146447 1309
rect 149054 1300 149060 1352
rect 149112 1340 149118 1352
rect 149885 1343 149943 1349
rect 149885 1340 149897 1343
rect 149112 1312 149897 1340
rect 149112 1300 149118 1312
rect 149885 1309 149897 1312
rect 149931 1309 149943 1343
rect 149885 1303 149943 1309
rect 149977 1343 150035 1349
rect 149977 1309 149989 1343
rect 150023 1340 150035 1343
rect 150066 1340 150072 1352
rect 150023 1312 150072 1340
rect 150023 1309 150035 1312
rect 149977 1303 150035 1309
rect 140038 1272 140044 1284
rect 134668 1244 136220 1272
rect 138952 1244 140044 1272
rect 134668 1232 134674 1244
rect 134334 1204 134340 1216
rect 132543 1176 133368 1204
rect 134295 1176 134340 1204
rect 132543 1173 132555 1176
rect 132497 1167 132555 1173
rect 134334 1164 134340 1176
rect 134392 1164 134398 1216
rect 134426 1164 134432 1216
rect 134484 1204 134490 1216
rect 136082 1204 136088 1216
rect 134484 1176 136088 1204
rect 134484 1164 134490 1176
rect 136082 1164 136088 1176
rect 136140 1164 136146 1216
rect 136192 1204 136220 1244
rect 140038 1232 140044 1244
rect 140096 1232 140102 1284
rect 140958 1232 140964 1284
rect 141016 1272 141022 1284
rect 141142 1272 141148 1284
rect 141016 1244 141148 1272
rect 141016 1232 141022 1244
rect 141142 1232 141148 1244
rect 141200 1232 141206 1284
rect 145009 1275 145067 1281
rect 145009 1241 145021 1275
rect 145055 1272 145067 1275
rect 149146 1272 149152 1284
rect 145055 1244 149152 1272
rect 145055 1241 145067 1244
rect 145009 1235 145067 1241
rect 149146 1232 149152 1244
rect 149204 1232 149210 1284
rect 149900 1272 149928 1303
rect 150066 1300 150072 1312
rect 150124 1300 150130 1352
rect 151354 1340 151360 1352
rect 151315 1312 151360 1340
rect 151354 1300 151360 1312
rect 151412 1300 151418 1352
rect 151446 1300 151452 1352
rect 151504 1340 151510 1352
rect 152642 1340 152648 1352
rect 151504 1312 152648 1340
rect 151504 1300 151510 1312
rect 152642 1300 152648 1312
rect 152700 1300 152706 1352
rect 154393 1343 154451 1349
rect 154393 1309 154405 1343
rect 154439 1340 154451 1343
rect 155770 1340 155776 1352
rect 154439 1312 155776 1340
rect 154439 1309 154451 1312
rect 154393 1303 154451 1309
rect 155770 1300 155776 1312
rect 155828 1300 155834 1352
rect 156874 1340 156880 1352
rect 156835 1312 156880 1340
rect 156874 1300 156880 1312
rect 156932 1340 156938 1352
rect 157613 1343 157671 1349
rect 157613 1340 157625 1343
rect 156932 1312 157625 1340
rect 156932 1300 156938 1312
rect 157613 1309 157625 1312
rect 157659 1309 157671 1343
rect 157613 1303 157671 1309
rect 158257 1343 158315 1349
rect 158257 1309 158269 1343
rect 158303 1340 158315 1343
rect 158714 1340 158720 1352
rect 158303 1312 158720 1340
rect 158303 1309 158315 1312
rect 158257 1303 158315 1309
rect 150713 1275 150771 1281
rect 150713 1272 150725 1275
rect 149900 1244 150725 1272
rect 150713 1241 150725 1244
rect 150759 1241 150771 1275
rect 151372 1272 151400 1300
rect 151817 1275 151875 1281
rect 151817 1272 151829 1275
rect 151372 1244 151829 1272
rect 150713 1235 150771 1241
rect 151817 1241 151829 1244
rect 151863 1241 151875 1275
rect 151817 1235 151875 1241
rect 155218 1232 155224 1284
rect 155276 1272 155282 1284
rect 158272 1272 158300 1303
rect 158714 1300 158720 1312
rect 158772 1300 158778 1352
rect 159634 1340 159640 1352
rect 159595 1312 159640 1340
rect 159634 1300 159640 1312
rect 159692 1300 159698 1352
rect 161106 1340 161112 1352
rect 161067 1312 161112 1340
rect 161106 1300 161112 1312
rect 161164 1340 161170 1352
rect 161569 1343 161627 1349
rect 161569 1340 161581 1343
rect 161164 1312 161581 1340
rect 161164 1300 161170 1312
rect 161569 1309 161581 1312
rect 161615 1309 161627 1343
rect 161569 1303 161627 1309
rect 162302 1300 162308 1352
rect 162360 1340 162366 1352
rect 162397 1343 162455 1349
rect 162397 1340 162409 1343
rect 162360 1312 162409 1340
rect 162360 1300 162366 1312
rect 162397 1309 162409 1312
rect 162443 1309 162455 1343
rect 162397 1303 162455 1309
rect 155276 1244 158300 1272
rect 155276 1232 155282 1244
rect 159542 1232 159548 1284
rect 159600 1272 159606 1284
rect 160830 1272 160836 1284
rect 159600 1244 160836 1272
rect 159600 1232 159606 1244
rect 160830 1232 160836 1244
rect 160888 1232 160894 1284
rect 162412 1272 162440 1303
rect 162854 1300 162860 1352
rect 162912 1340 162918 1352
rect 164436 1349 164464 1380
rect 165430 1368 165436 1380
rect 165488 1368 165494 1420
rect 163593 1343 163651 1349
rect 163593 1340 163605 1343
rect 162912 1312 163605 1340
rect 162912 1300 162918 1312
rect 163593 1309 163605 1312
rect 163639 1340 163651 1343
rect 164053 1343 164111 1349
rect 164053 1340 164065 1343
rect 163639 1312 164065 1340
rect 163639 1309 163651 1312
rect 163593 1303 163651 1309
rect 164053 1309 164065 1312
rect 164099 1309 164111 1343
rect 164053 1303 164111 1309
rect 164421 1343 164479 1349
rect 164421 1309 164433 1343
rect 164467 1309 164479 1343
rect 164421 1303 164479 1309
rect 164973 1343 165031 1349
rect 164973 1309 164985 1343
rect 165019 1340 165031 1343
rect 166445 1343 166503 1349
rect 166445 1340 166457 1343
rect 165019 1312 166457 1340
rect 165019 1309 165031 1312
rect 164973 1303 165031 1309
rect 166445 1309 166457 1312
rect 166491 1309 166503 1343
rect 166718 1340 166724 1352
rect 166679 1312 166724 1340
rect 166445 1303 166503 1309
rect 162949 1275 163007 1281
rect 162949 1272 162961 1275
rect 162412 1244 162961 1272
rect 162949 1241 162961 1244
rect 162995 1241 163007 1275
rect 166460 1272 166488 1303
rect 166718 1300 166724 1312
rect 166776 1340 166782 1352
rect 167181 1343 167239 1349
rect 167181 1340 167193 1343
rect 166776 1312 167193 1340
rect 166776 1300 166782 1312
rect 167181 1309 167193 1312
rect 167227 1309 167239 1343
rect 167181 1303 167239 1309
rect 167733 1275 167791 1281
rect 167733 1272 167745 1275
rect 166460 1244 167745 1272
rect 162949 1235 163007 1241
rect 167733 1241 167745 1244
rect 167779 1241 167791 1275
rect 167733 1235 167791 1241
rect 139670 1204 139676 1216
rect 136192 1176 139676 1204
rect 139670 1164 139676 1176
rect 139728 1164 139734 1216
rect 143994 1164 144000 1216
rect 144052 1204 144058 1216
rect 144270 1204 144276 1216
rect 144052 1176 144276 1204
rect 144052 1164 144058 1176
rect 144270 1164 144276 1176
rect 144328 1204 144334 1216
rect 144457 1207 144515 1213
rect 144457 1204 144469 1207
rect 144328 1176 144469 1204
rect 144328 1164 144334 1176
rect 144457 1173 144469 1176
rect 144503 1173 144515 1207
rect 146018 1204 146024 1216
rect 145979 1176 146024 1204
rect 144457 1167 144515 1173
rect 146018 1164 146024 1176
rect 146076 1164 146082 1216
rect 146662 1164 146668 1216
rect 146720 1204 146726 1216
rect 146757 1207 146815 1213
rect 146757 1204 146769 1207
rect 146720 1176 146769 1204
rect 146720 1164 146726 1176
rect 146757 1173 146769 1176
rect 146803 1173 146815 1207
rect 146757 1167 146815 1173
rect 151449 1207 151507 1213
rect 151449 1173 151461 1207
rect 151495 1204 151507 1207
rect 151722 1204 151728 1216
rect 151495 1176 151728 1204
rect 151495 1173 151507 1176
rect 151449 1167 151507 1173
rect 151722 1164 151728 1176
rect 151780 1164 151786 1216
rect 152918 1164 152924 1216
rect 152976 1204 152982 1216
rect 153654 1204 153660 1216
rect 152976 1176 153660 1204
rect 152976 1164 152982 1176
rect 153654 1164 153660 1176
rect 153712 1164 153718 1216
rect 154022 1164 154028 1216
rect 154080 1204 154086 1216
rect 154666 1204 154672 1216
rect 154080 1176 154672 1204
rect 154080 1164 154086 1176
rect 154666 1164 154672 1176
rect 154724 1204 154730 1216
rect 154853 1207 154911 1213
rect 154853 1204 154865 1207
rect 154724 1176 154865 1204
rect 154724 1164 154730 1176
rect 154853 1173 154865 1176
rect 154899 1173 154911 1207
rect 154853 1167 154911 1173
rect 161201 1207 161259 1213
rect 161201 1173 161213 1207
rect 161247 1204 161259 1207
rect 161290 1204 161296 1216
rect 161247 1176 161296 1204
rect 161247 1173 161259 1176
rect 161201 1167 161259 1173
rect 161290 1164 161296 1176
rect 161348 1164 161354 1216
rect 161474 1164 161480 1216
rect 161532 1204 161538 1216
rect 161934 1204 161940 1216
rect 161532 1176 161940 1204
rect 161532 1164 161538 1176
rect 161934 1164 161940 1176
rect 161992 1164 161998 1216
rect 162489 1207 162547 1213
rect 162489 1173 162501 1207
rect 162535 1204 162547 1207
rect 162762 1204 162768 1216
rect 162535 1176 162768 1204
rect 162535 1173 162547 1176
rect 162489 1167 162547 1173
rect 162762 1164 162768 1176
rect 162820 1164 162826 1216
rect 163685 1207 163743 1213
rect 163685 1173 163697 1207
rect 163731 1204 163743 1207
rect 164418 1204 164424 1216
rect 163731 1176 164424 1204
rect 163731 1173 163743 1176
rect 163685 1167 163743 1173
rect 164418 1164 164424 1176
rect 164476 1164 164482 1216
rect 166810 1204 166816 1216
rect 166771 1176 166816 1204
rect 166810 1164 166816 1176
rect 166868 1164 166874 1216
rect 166902 1164 166908 1216
rect 166960 1204 166966 1216
rect 167549 1207 167607 1213
rect 167549 1204 167561 1207
rect 166960 1176 167561 1204
rect 166960 1164 166966 1176
rect 167549 1173 167561 1176
rect 167595 1173 167607 1207
rect 167549 1167 167607 1173
rect 368 1114 93012 1136
rect 368 1062 56667 1114
rect 56719 1062 56731 1114
rect 56783 1062 56795 1114
rect 56847 1062 56859 1114
rect 56911 1062 93012 1114
rect 102028 1114 169556 1136
rect 368 1040 93012 1062
rect 97350 1028 97356 1080
rect 97408 1068 97414 1080
rect 100849 1071 100907 1077
rect 100849 1068 100861 1071
rect 97408 1040 100861 1068
rect 97408 1028 97414 1040
rect 100849 1037 100861 1040
rect 100895 1037 100907 1071
rect 102028 1062 113088 1114
rect 113140 1062 113152 1114
rect 113204 1062 113216 1114
rect 113268 1062 113280 1114
rect 113332 1062 169556 1114
rect 102028 1040 169556 1062
rect 100849 1031 100907 1037
rect 3421 1003 3479 1009
rect 3421 969 3433 1003
rect 3467 1000 3479 1003
rect 3605 1003 3663 1009
rect 3605 1000 3617 1003
rect 3467 972 3617 1000
rect 3467 969 3479 972
rect 3421 963 3479 969
rect 3605 969 3617 972
rect 3651 1000 3663 1003
rect 6730 1000 6736 1012
rect 3651 972 6736 1000
rect 3651 969 3663 972
rect 3605 963 3663 969
rect 6730 960 6736 972
rect 6788 960 6794 1012
rect 12161 1003 12219 1009
rect 12161 969 12173 1003
rect 12207 1000 12219 1003
rect 12986 1000 12992 1012
rect 12207 972 12992 1000
rect 12207 969 12219 972
rect 12161 963 12219 969
rect 2225 935 2283 941
rect 2225 901 2237 935
rect 2271 932 2283 935
rect 5905 935 5963 941
rect 5905 932 5917 935
rect 2271 904 5917 932
rect 2271 901 2283 904
rect 2225 895 2283 901
rect 5905 901 5917 904
rect 5951 901 5963 935
rect 5905 895 5963 901
rect 3421 867 3479 873
rect 3421 833 3433 867
rect 3467 864 3479 867
rect 3697 867 3755 873
rect 3697 864 3709 867
rect 3467 836 3709 864
rect 3467 833 3479 836
rect 3421 827 3479 833
rect 3697 833 3709 836
rect 3743 833 3755 867
rect 3697 827 3755 833
rect 5261 867 5319 873
rect 5261 833 5273 867
rect 5307 864 5319 867
rect 5626 864 5632 876
rect 5307 836 5632 864
rect 5307 833 5319 836
rect 5261 827 5319 833
rect 5626 824 5632 836
rect 5684 824 5690 876
rect 5920 864 5948 895
rect 5994 892 6000 944
rect 6052 932 6058 944
rect 8757 935 8815 941
rect 8757 932 8769 935
rect 6052 904 8769 932
rect 6052 892 6058 904
rect 8757 901 8769 904
rect 8803 932 8815 935
rect 8803 904 9076 932
rect 8803 901 8815 904
rect 8757 895 8815 901
rect 6181 867 6239 873
rect 6181 864 6193 867
rect 5920 836 6193 864
rect 6181 833 6193 836
rect 6227 833 6239 867
rect 6181 827 6239 833
rect 7745 867 7803 873
rect 7745 833 7757 867
rect 7791 864 7803 867
rect 8110 864 8116 876
rect 7791 836 8116 864
rect 7791 833 7803 836
rect 7745 827 7803 833
rect 8110 824 8116 836
rect 8168 824 8174 876
rect 9048 873 9076 904
rect 9033 867 9091 873
rect 9033 833 9045 867
rect 9079 833 9091 867
rect 9033 827 9091 833
rect 10597 867 10655 873
rect 10597 833 10609 867
rect 10643 864 10655 867
rect 10962 864 10968 876
rect 10643 836 10968 864
rect 10643 833 10655 836
rect 10597 827 10655 833
rect 10962 824 10968 836
rect 11020 824 11026 876
rect 12268 873 12296 972
rect 12986 960 12992 972
rect 13044 960 13050 1012
rect 19337 1003 19395 1009
rect 19337 969 19349 1003
rect 19383 1000 19395 1003
rect 19610 1000 19616 1012
rect 19383 972 19616 1000
rect 19383 969 19395 972
rect 19337 963 19395 969
rect 19610 960 19616 972
rect 19668 960 19674 1012
rect 19794 960 19800 1012
rect 19852 1000 19858 1012
rect 22189 1003 22247 1009
rect 19852 972 19897 1000
rect 19852 960 19858 972
rect 22189 969 22201 1003
rect 22235 1000 22247 1003
rect 23658 1000 23664 1012
rect 22235 972 23664 1000
rect 22235 969 22247 972
rect 22189 963 22247 969
rect 23658 960 23664 972
rect 23716 1000 23722 1012
rect 24670 1000 24676 1012
rect 23716 972 24676 1000
rect 23716 960 23722 972
rect 24670 960 24676 972
rect 24728 960 24734 1012
rect 24946 1000 24952 1012
rect 24907 972 24952 1000
rect 24946 960 24952 972
rect 25004 960 25010 1012
rect 25866 1000 25872 1012
rect 25827 972 25872 1000
rect 25866 960 25872 972
rect 25924 960 25930 1012
rect 26142 960 26148 1012
rect 26200 1000 26206 1012
rect 26329 1003 26387 1009
rect 26329 1000 26341 1003
rect 26200 972 26341 1000
rect 26200 960 26206 972
rect 26329 969 26341 972
rect 26375 969 26387 1003
rect 26329 963 26387 969
rect 27982 960 27988 1012
rect 28040 1000 28046 1012
rect 30190 1000 30196 1012
rect 28040 972 30196 1000
rect 28040 960 28046 972
rect 30190 960 30196 972
rect 30248 960 30254 1012
rect 30282 960 30288 1012
rect 30340 1000 30346 1012
rect 31849 1003 31907 1009
rect 31849 1000 31861 1003
rect 30340 972 31861 1000
rect 30340 960 30346 972
rect 31849 969 31861 972
rect 31895 969 31907 1003
rect 31849 963 31907 969
rect 31938 960 31944 1012
rect 31996 1000 32002 1012
rect 35710 1000 35716 1012
rect 31996 972 35716 1000
rect 31996 960 32002 972
rect 35710 960 35716 972
rect 35768 960 35774 1012
rect 36354 1000 36360 1012
rect 36315 972 36360 1000
rect 36354 960 36360 972
rect 36412 960 36418 1012
rect 36446 960 36452 1012
rect 36504 1000 36510 1012
rect 38473 1003 38531 1009
rect 38473 1000 38485 1003
rect 36504 972 38485 1000
rect 36504 960 36510 972
rect 38473 969 38485 972
rect 38519 969 38531 1003
rect 40770 1000 40776 1012
rect 38473 963 38531 969
rect 38672 972 40776 1000
rect 35066 932 35072 944
rect 12360 904 35072 932
rect 12253 867 12311 873
rect 12253 833 12265 867
rect 12299 833 12311 867
rect 12253 827 12311 833
rect 4338 756 4344 808
rect 4396 796 4402 808
rect 4709 799 4767 805
rect 4709 796 4721 799
rect 4396 768 4721 796
rect 4396 756 4402 768
rect 4709 765 4721 768
rect 4755 765 4767 799
rect 4709 759 4767 765
rect 4890 756 4896 808
rect 4948 796 4954 808
rect 7193 799 7251 805
rect 7193 796 7205 799
rect 4948 768 7205 796
rect 4948 756 4954 768
rect 7193 765 7205 768
rect 7239 765 7251 799
rect 7193 759 7251 765
rect 9674 756 9680 808
rect 9732 796 9738 808
rect 10045 799 10103 805
rect 10045 796 10057 799
rect 9732 768 10057 796
rect 9732 756 9738 768
rect 10045 765 10057 768
rect 10091 765 10103 799
rect 10045 759 10103 765
rect 5626 728 5632 740
rect 5587 700 5632 728
rect 5626 688 5632 700
rect 5684 688 5690 740
rect 7834 688 7840 740
rect 7892 728 7898 740
rect 12360 728 12388 904
rect 35066 892 35072 904
rect 35124 892 35130 944
rect 37458 932 37464 944
rect 35268 904 37464 932
rect 13817 867 13875 873
rect 13817 833 13829 867
rect 13863 864 13875 867
rect 15933 867 15991 873
rect 13863 836 14228 864
rect 13863 833 13875 836
rect 13817 827 13875 833
rect 12434 756 12440 808
rect 12492 796 12498 808
rect 13265 799 13323 805
rect 13265 796 13277 799
rect 12492 768 13277 796
rect 12492 756 12498 768
rect 13265 765 13277 768
rect 13311 765 13323 799
rect 13265 759 13323 765
rect 7892 700 12388 728
rect 7892 688 7898 700
rect 10962 660 10968 672
rect 10923 632 10968 660
rect 10962 620 10968 632
rect 11020 620 11026 672
rect 14200 669 14228 836
rect 15933 833 15945 867
rect 15979 833 15991 867
rect 15933 827 15991 833
rect 16669 867 16727 873
rect 16669 833 16681 867
rect 16715 864 16727 867
rect 16761 867 16819 873
rect 16761 864 16773 867
rect 16715 836 16773 864
rect 16715 833 16727 836
rect 16669 827 16727 833
rect 16761 833 16773 836
rect 16807 833 16819 867
rect 16761 827 16819 833
rect 18233 867 18291 873
rect 18233 833 18245 867
rect 18279 864 18291 867
rect 18601 867 18659 873
rect 18601 864 18613 867
rect 18279 836 18613 864
rect 18279 833 18291 836
rect 18233 827 18291 833
rect 18601 833 18613 836
rect 18647 833 18659 867
rect 18601 827 18659 833
rect 14921 799 14979 805
rect 14921 765 14933 799
rect 14967 796 14979 799
rect 15749 799 15807 805
rect 15749 796 15761 799
rect 14967 768 15761 796
rect 14967 765 14979 768
rect 14921 759 14979 765
rect 15749 765 15761 768
rect 15795 796 15807 799
rect 15948 796 15976 827
rect 15795 768 15976 796
rect 16301 799 16359 805
rect 15795 765 15807 768
rect 15749 759 15807 765
rect 16301 765 16313 799
rect 16347 796 16359 799
rect 18248 796 18276 827
rect 20622 824 20628 876
rect 20680 864 20686 876
rect 20717 867 20775 873
rect 20717 864 20729 867
rect 20680 836 20729 864
rect 20680 824 20686 836
rect 20717 833 20729 836
rect 20763 864 20775 867
rect 21453 867 21511 873
rect 21453 864 21465 867
rect 20763 836 21465 864
rect 20763 833 20775 836
rect 20717 827 20775 833
rect 21453 833 21465 836
rect 21499 833 21511 867
rect 21453 827 21511 833
rect 22002 824 22008 876
rect 22060 864 22066 876
rect 23477 867 23535 873
rect 23477 864 23489 867
rect 22060 836 23489 864
rect 22060 824 22066 836
rect 23477 833 23489 836
rect 23523 864 23535 867
rect 24305 867 24363 873
rect 24305 864 24317 867
rect 23523 836 24317 864
rect 23523 833 23535 836
rect 23477 827 23535 833
rect 24305 833 24317 836
rect 24351 833 24363 867
rect 24305 827 24363 833
rect 24857 867 24915 873
rect 24857 833 24869 867
rect 24903 833 24915 867
rect 24857 827 24915 833
rect 16347 768 18276 796
rect 16347 765 16359 768
rect 16301 759 16359 765
rect 18322 756 18328 808
rect 18380 796 18386 808
rect 20441 799 20499 805
rect 20441 796 20453 799
rect 18380 768 20453 796
rect 18380 756 18386 768
rect 20441 765 20453 768
rect 20487 765 20499 799
rect 24026 796 24032 808
rect 23987 768 24032 796
rect 20441 759 20499 765
rect 24026 756 24032 768
rect 24084 756 24090 808
rect 24872 796 24900 827
rect 25866 824 25872 876
rect 25924 864 25930 876
rect 26513 867 26571 873
rect 26513 864 26525 867
rect 25924 836 26525 864
rect 25924 824 25930 836
rect 26513 833 26525 836
rect 26559 833 26571 867
rect 27890 864 27896 876
rect 26513 827 26571 833
rect 26620 836 27660 864
rect 27851 836 27896 864
rect 25409 799 25467 805
rect 25409 796 25421 799
rect 24872 768 25421 796
rect 25409 765 25421 768
rect 25455 796 25467 799
rect 26620 796 26648 836
rect 27522 796 27528 808
rect 25455 768 26648 796
rect 27483 768 27528 796
rect 25455 765 25467 768
rect 25409 759 25467 765
rect 27522 756 27528 768
rect 27580 756 27586 808
rect 27632 796 27660 836
rect 27890 824 27896 836
rect 27948 864 27954 876
rect 28353 867 28411 873
rect 28353 864 28365 867
rect 27948 836 28365 864
rect 27948 824 27954 836
rect 28353 833 28365 836
rect 28399 833 28411 867
rect 28353 827 28411 833
rect 30098 824 30104 876
rect 30156 864 30162 876
rect 30377 867 30435 873
rect 30377 864 30389 867
rect 30156 836 30389 864
rect 30156 824 30162 836
rect 30377 833 30389 836
rect 30423 864 30435 867
rect 30745 867 30803 873
rect 30745 864 30757 867
rect 30423 836 30757 864
rect 30423 833 30435 836
rect 30377 827 30435 833
rect 30745 833 30757 836
rect 30791 833 30803 867
rect 33410 864 33416 876
rect 30745 827 30803 833
rect 31680 836 33416 864
rect 28994 796 29000 808
rect 27632 768 29000 796
rect 28994 756 29000 768
rect 29052 756 29058 808
rect 30469 799 30527 805
rect 30469 765 30481 799
rect 30515 796 30527 799
rect 31680 796 31708 836
rect 33410 824 33416 836
rect 33468 824 33474 876
rect 33505 867 33563 873
rect 33505 833 33517 867
rect 33551 864 33563 867
rect 33870 864 33876 876
rect 33551 836 33876 864
rect 33551 833 33563 836
rect 33505 827 33563 833
rect 33870 824 33876 836
rect 33928 824 33934 876
rect 34698 824 34704 876
rect 34756 864 34762 876
rect 35268 864 35296 904
rect 37458 892 37464 904
rect 37516 892 37522 944
rect 38565 935 38623 941
rect 38565 932 38577 935
rect 37660 904 38577 932
rect 35434 864 35440 876
rect 34756 836 35296 864
rect 35395 836 35440 864
rect 34756 824 34762 836
rect 35434 824 35440 836
rect 35492 824 35498 876
rect 35989 867 36047 873
rect 35989 833 36001 867
rect 36035 864 36047 867
rect 36035 836 37504 864
rect 36035 833 36047 836
rect 35989 827 36047 833
rect 37476 796 37504 836
rect 37550 824 37556 876
rect 37608 864 37614 876
rect 37660 873 37688 904
rect 38565 901 38577 904
rect 38611 901 38623 935
rect 38565 895 38623 901
rect 37645 867 37703 873
rect 37645 864 37657 867
rect 37608 836 37657 864
rect 37608 824 37614 836
rect 37645 833 37657 836
rect 37691 833 37703 867
rect 37645 827 37703 833
rect 37826 824 37832 876
rect 37884 864 37890 876
rect 38672 864 38700 972
rect 40770 960 40776 972
rect 40828 960 40834 1012
rect 40954 960 40960 1012
rect 41012 1000 41018 1012
rect 42242 1000 42248 1012
rect 41012 972 42248 1000
rect 41012 960 41018 972
rect 42242 960 42248 972
rect 42300 960 42306 1012
rect 42334 960 42340 1012
rect 42392 1000 42398 1012
rect 44542 1000 44548 1012
rect 42392 972 44548 1000
rect 42392 960 42398 972
rect 44542 960 44548 972
rect 44600 960 44606 1012
rect 44818 1000 44824 1012
rect 44779 972 44824 1000
rect 44818 960 44824 972
rect 44876 960 44882 1012
rect 44910 960 44916 1012
rect 44968 1000 44974 1012
rect 47210 1000 47216 1012
rect 44968 972 47216 1000
rect 44968 960 44974 972
rect 47210 960 47216 972
rect 47268 960 47274 1012
rect 47673 1003 47731 1009
rect 47673 969 47685 1003
rect 47719 1000 47731 1003
rect 47854 1000 47860 1012
rect 47719 972 47860 1000
rect 47719 969 47731 972
rect 47673 963 47731 969
rect 47854 960 47860 972
rect 47912 960 47918 1012
rect 48777 1003 48835 1009
rect 48777 969 48789 1003
rect 48823 1000 48835 1003
rect 49602 1000 49608 1012
rect 48823 972 49608 1000
rect 48823 969 48835 972
rect 48777 963 48835 969
rect 49602 960 49608 972
rect 49660 960 49666 1012
rect 50065 1003 50123 1009
rect 50065 969 50077 1003
rect 50111 1000 50123 1003
rect 50154 1000 50160 1012
rect 50111 972 50160 1000
rect 50111 969 50123 972
rect 50065 963 50123 969
rect 50154 960 50160 972
rect 50212 960 50218 1012
rect 50430 960 50436 1012
rect 50488 1000 50494 1012
rect 102410 1000 102416 1012
rect 50488 972 102416 1000
rect 50488 960 50494 972
rect 102410 960 102416 972
rect 102468 960 102474 1012
rect 103977 1003 104035 1009
rect 103716 972 103928 1000
rect 40678 932 40684 944
rect 37884 836 38700 864
rect 38764 904 40684 932
rect 37884 824 37890 836
rect 38286 796 38292 808
rect 30515 768 31708 796
rect 31772 768 36952 796
rect 37476 768 38292 796
rect 30515 765 30527 768
rect 30469 759 30527 765
rect 16761 731 16819 737
rect 16761 697 16773 731
rect 16807 728 16819 731
rect 17037 731 17095 737
rect 17037 728 17049 731
rect 16807 700 17049 728
rect 16807 697 16819 700
rect 16761 691 16819 697
rect 17037 697 17049 700
rect 17083 728 17095 731
rect 27982 728 27988 740
rect 17083 700 27988 728
rect 17083 697 17095 700
rect 17037 691 17095 697
rect 27982 688 27988 700
rect 28040 688 28046 740
rect 28074 688 28080 740
rect 28132 728 28138 740
rect 31772 728 31800 768
rect 33321 731 33379 737
rect 28132 700 31800 728
rect 31864 700 33272 728
rect 28132 688 28138 700
rect 14185 663 14243 669
rect 14185 629 14197 663
rect 14231 660 14243 663
rect 14274 660 14280 672
rect 14231 632 14280 660
rect 14231 629 14243 632
rect 14185 623 14243 629
rect 14274 620 14280 632
rect 14332 620 14338 672
rect 18046 660 18052 672
rect 18007 632 18052 660
rect 18046 620 18052 632
rect 18104 620 18110 672
rect 26510 620 26516 672
rect 26568 660 26574 672
rect 28810 660 28816 672
rect 26568 632 28816 660
rect 26568 620 26574 632
rect 28810 620 28816 632
rect 28868 620 28874 672
rect 30190 620 30196 672
rect 30248 660 30254 672
rect 31864 660 31892 700
rect 30248 632 31892 660
rect 33244 660 33272 700
rect 33321 697 33333 731
rect 33367 728 33379 731
rect 34698 728 34704 740
rect 33367 700 34704 728
rect 33367 697 33379 700
rect 33321 691 33379 697
rect 34698 688 34704 700
rect 34756 688 34762 740
rect 34882 688 34888 740
rect 34940 728 34946 740
rect 36538 728 36544 740
rect 34940 700 36544 728
rect 34940 688 34946 700
rect 36538 688 36544 700
rect 36596 688 36602 740
rect 36924 728 36952 768
rect 38286 756 38292 768
rect 38344 756 38350 808
rect 38764 796 38792 904
rect 40678 892 40684 904
rect 40736 892 40742 944
rect 40862 892 40868 944
rect 40920 932 40926 944
rect 40920 904 41920 932
rect 40920 892 40926 904
rect 38930 824 38936 876
rect 38988 864 38994 876
rect 39117 867 39175 873
rect 39117 864 39129 867
rect 38988 836 39129 864
rect 38988 824 38994 836
rect 39117 833 39129 836
rect 39163 833 39175 867
rect 41506 864 41512 876
rect 39117 827 39175 833
rect 39224 836 41092 864
rect 41467 836 41512 864
rect 38396 768 38792 796
rect 38396 728 38424 768
rect 39022 756 39028 808
rect 39080 796 39086 808
rect 39224 796 39252 836
rect 39080 768 39252 796
rect 39080 756 39086 768
rect 39298 756 39304 808
rect 39356 796 39362 808
rect 40494 796 40500 808
rect 39356 768 40500 796
rect 39356 756 39362 768
rect 40494 756 40500 768
rect 40552 756 40558 808
rect 40586 756 40592 808
rect 40644 796 40650 808
rect 41064 796 41092 836
rect 41506 824 41512 836
rect 41564 864 41570 876
rect 41601 867 41659 873
rect 41601 864 41613 867
rect 41564 836 41613 864
rect 41564 824 41570 836
rect 41601 833 41613 836
rect 41647 833 41659 867
rect 41601 827 41659 833
rect 40644 768 41000 796
rect 41064 768 41828 796
rect 40644 756 40650 768
rect 36924 700 38424 728
rect 38473 731 38531 737
rect 38473 697 38485 731
rect 38519 728 38531 731
rect 38519 700 39620 728
rect 38519 697 38531 700
rect 38473 691 38531 697
rect 36446 660 36452 672
rect 33244 632 36452 660
rect 30248 620 30254 632
rect 36446 620 36452 632
rect 36504 620 36510 672
rect 38013 663 38071 669
rect 38013 629 38025 663
rect 38059 660 38071 663
rect 39298 660 39304 672
rect 38059 632 39304 660
rect 38059 629 38071 632
rect 38013 623 38071 629
rect 39298 620 39304 632
rect 39356 620 39362 672
rect 39592 660 39620 700
rect 40402 688 40408 740
rect 40460 728 40466 740
rect 40862 728 40868 740
rect 40460 700 40868 728
rect 40460 688 40466 700
rect 40862 688 40868 700
rect 40920 688 40926 740
rect 40972 728 41000 768
rect 41690 728 41696 740
rect 40972 700 41696 728
rect 41690 688 41696 700
rect 41748 688 41754 740
rect 41598 660 41604 672
rect 39592 632 41604 660
rect 41598 620 41604 632
rect 41656 620 41662 672
rect 41800 660 41828 768
rect 41892 728 41920 904
rect 41966 892 41972 944
rect 42024 932 42030 944
rect 42518 932 42524 944
rect 42024 904 42524 932
rect 42024 892 42030 904
rect 42518 892 42524 904
rect 42576 892 42582 944
rect 43070 892 43076 944
rect 43128 932 43134 944
rect 65150 932 65156 944
rect 43128 904 65156 932
rect 43128 892 43134 904
rect 65150 892 65156 904
rect 65208 892 65214 944
rect 66346 932 66352 944
rect 66307 904 66352 932
rect 66346 892 66352 904
rect 66404 932 66410 944
rect 68373 935 68431 941
rect 68373 932 68385 935
rect 66404 904 66484 932
rect 66404 892 66410 904
rect 42337 867 42395 873
rect 42337 833 42349 867
rect 42383 864 42395 867
rect 42705 867 42763 873
rect 42705 864 42717 867
rect 42383 836 42717 864
rect 42383 833 42395 836
rect 42337 827 42395 833
rect 42705 833 42717 836
rect 42751 864 42763 867
rect 42978 864 42984 876
rect 42751 836 42984 864
rect 42751 833 42763 836
rect 42705 827 42763 833
rect 42978 824 42984 836
rect 43036 824 43042 876
rect 43809 867 43867 873
rect 43809 833 43821 867
rect 43855 833 43867 867
rect 43809 827 43867 833
rect 41969 799 42027 805
rect 41969 765 41981 799
rect 42015 796 42027 799
rect 43824 796 43852 827
rect 43898 824 43904 876
rect 43956 864 43962 876
rect 43993 867 44051 873
rect 43993 864 44005 867
rect 43956 836 44005 864
rect 43956 824 43962 836
rect 43993 833 44005 836
rect 44039 833 44051 867
rect 43993 827 44051 833
rect 44082 824 44088 876
rect 44140 864 44146 876
rect 44910 864 44916 876
rect 44140 836 44916 864
rect 44140 824 44146 836
rect 44910 824 44916 836
rect 44968 824 44974 876
rect 45646 824 45652 876
rect 45704 864 45710 876
rect 46109 867 46167 873
rect 46109 864 46121 867
rect 45704 836 46121 864
rect 45704 824 45710 836
rect 46109 833 46121 836
rect 46155 833 46167 867
rect 46290 864 46296 876
rect 46251 836 46296 864
rect 46109 827 46167 833
rect 46290 824 46296 836
rect 46348 864 46354 876
rect 47121 867 47179 873
rect 47121 864 47133 867
rect 46348 836 47133 864
rect 46348 824 46354 836
rect 47121 833 47133 836
rect 47167 833 47179 867
rect 49418 864 49424 876
rect 47121 827 47179 833
rect 47228 836 49424 864
rect 44269 799 44327 805
rect 44269 796 44281 799
rect 42015 768 44281 796
rect 42015 765 42027 768
rect 41969 759 42027 765
rect 44269 765 44281 768
rect 44315 765 44327 799
rect 44269 759 44327 765
rect 44634 756 44640 808
rect 44692 796 44698 808
rect 47228 796 47256 836
rect 49418 824 49424 836
rect 49476 824 49482 876
rect 49605 867 49663 873
rect 49605 833 49617 867
rect 49651 864 49663 867
rect 50154 864 50160 876
rect 49651 836 50160 864
rect 49651 833 49663 836
rect 49605 827 49663 833
rect 50154 824 50160 836
rect 50212 824 50218 876
rect 50525 867 50583 873
rect 50525 833 50537 867
rect 50571 864 50583 867
rect 51629 867 51687 873
rect 51629 864 51641 867
rect 50571 836 51641 864
rect 50571 833 50583 836
rect 50525 827 50583 833
rect 51629 833 51641 836
rect 51675 864 51687 867
rect 51813 867 51871 873
rect 51813 864 51825 867
rect 51675 836 51825 864
rect 51675 833 51687 836
rect 51629 827 51687 833
rect 51813 833 51825 836
rect 51859 833 51871 867
rect 52546 864 52552 876
rect 52507 836 52552 864
rect 51813 827 51871 833
rect 52546 824 52552 836
rect 52604 824 52610 876
rect 52641 867 52699 873
rect 52641 833 52653 867
rect 52687 864 52699 867
rect 53006 864 53012 876
rect 52687 836 53012 864
rect 52687 833 52699 836
rect 52641 827 52699 833
rect 53006 824 53012 836
rect 53064 824 53070 876
rect 53469 867 53527 873
rect 53469 833 53481 867
rect 53515 864 53527 867
rect 54021 867 54079 873
rect 54021 864 54033 867
rect 53515 836 54033 864
rect 53515 833 53527 836
rect 53469 827 53527 833
rect 54021 833 54033 836
rect 54067 864 54079 867
rect 55306 864 55312 876
rect 54067 836 55312 864
rect 54067 833 54079 836
rect 54021 827 54079 833
rect 55306 824 55312 836
rect 55364 824 55370 876
rect 55490 824 55496 876
rect 55548 864 55554 876
rect 55861 867 55919 873
rect 55861 864 55873 867
rect 55548 836 55873 864
rect 55548 824 55554 836
rect 55861 833 55873 836
rect 55907 833 55919 867
rect 55861 827 55919 833
rect 56505 867 56563 873
rect 56505 833 56517 867
rect 56551 864 56563 867
rect 56873 867 56931 873
rect 56873 864 56885 867
rect 56551 836 56885 864
rect 56551 833 56563 836
rect 56505 827 56563 833
rect 56873 833 56885 836
rect 56919 864 56931 867
rect 57790 864 57796 876
rect 56919 836 57796 864
rect 56919 833 56931 836
rect 56873 827 56931 833
rect 57790 824 57796 836
rect 57848 824 57854 876
rect 58526 864 58532 876
rect 58487 836 58532 864
rect 58526 824 58532 836
rect 58584 824 58590 876
rect 59173 867 59231 873
rect 59173 833 59185 867
rect 59219 833 59231 867
rect 59173 827 59231 833
rect 44692 768 47256 796
rect 44692 756 44698 768
rect 47394 756 47400 808
rect 47452 796 47458 808
rect 48777 799 48835 805
rect 48777 796 48789 799
rect 47452 768 48789 796
rect 47452 756 47458 768
rect 48777 765 48789 768
rect 48823 765 48835 799
rect 48777 759 48835 765
rect 48961 799 49019 805
rect 48961 765 48973 799
rect 49007 765 49019 799
rect 50798 796 50804 808
rect 48961 759 49019 765
rect 49988 768 50804 796
rect 45370 728 45376 740
rect 41892 700 45376 728
rect 45370 688 45376 700
rect 45428 688 45434 740
rect 46106 688 46112 740
rect 46164 728 46170 740
rect 48976 728 49004 759
rect 46164 700 49004 728
rect 46164 688 46170 700
rect 49050 688 49056 740
rect 49108 728 49114 740
rect 49694 728 49700 740
rect 49108 700 49700 728
rect 49108 688 49114 700
rect 49694 688 49700 700
rect 49752 688 49758 740
rect 49786 688 49792 740
rect 49844 728 49850 740
rect 49988 728 50016 768
rect 50798 756 50804 768
rect 50856 756 50862 808
rect 50890 756 50896 808
rect 50948 796 50954 808
rect 54478 796 54484 808
rect 50948 768 54484 796
rect 50948 756 50954 768
rect 54478 756 54484 768
rect 54536 756 54542 808
rect 54849 799 54907 805
rect 54849 765 54861 799
rect 54895 796 54907 799
rect 56962 796 56968 808
rect 54895 768 56968 796
rect 54895 765 54907 768
rect 54849 759 54907 765
rect 56962 756 56968 768
rect 57020 756 57026 808
rect 57517 799 57575 805
rect 57517 765 57529 799
rect 57563 796 57575 799
rect 58986 796 58992 808
rect 57563 768 58992 796
rect 57563 765 57575 768
rect 57517 759 57575 765
rect 58986 756 58992 768
rect 59044 756 59050 808
rect 59188 796 59216 827
rect 59722 824 59728 876
rect 59780 864 59786 876
rect 60369 867 60427 873
rect 60369 864 60381 867
rect 59780 836 60381 864
rect 59780 824 59786 836
rect 60369 833 60381 836
rect 60415 833 60427 867
rect 60369 827 60427 833
rect 60458 824 60464 876
rect 60516 864 60522 876
rect 61381 867 61439 873
rect 61381 864 61393 867
rect 60516 836 61393 864
rect 60516 824 60522 836
rect 61381 833 61393 836
rect 61427 833 61439 867
rect 61381 827 61439 833
rect 61470 824 61476 876
rect 61528 864 61534 876
rect 63770 864 63776 876
rect 61528 836 63632 864
rect 63731 836 63776 864
rect 61528 824 61534 836
rect 59633 799 59691 805
rect 59633 796 59645 799
rect 59188 768 59645 796
rect 59633 765 59645 768
rect 59679 796 59691 799
rect 59906 796 59912 808
rect 59679 768 59912 796
rect 59679 765 59691 768
rect 59633 759 59691 765
rect 59906 756 59912 768
rect 59964 756 59970 808
rect 61933 799 61991 805
rect 61933 796 61945 799
rect 61120 768 61945 796
rect 49844 700 50016 728
rect 49844 688 49850 700
rect 50154 688 50160 740
rect 50212 728 50218 740
rect 51905 731 51963 737
rect 51905 728 51917 731
rect 50212 700 51917 728
rect 50212 688 50218 700
rect 51905 697 51917 700
rect 51951 697 51963 731
rect 51905 691 51963 697
rect 51994 688 52000 740
rect 52052 728 52058 740
rect 52641 731 52699 737
rect 52641 728 52653 731
rect 52052 700 52653 728
rect 52052 688 52058 700
rect 52641 697 52653 700
rect 52687 697 52699 731
rect 52914 728 52920 740
rect 52827 700 52920 728
rect 52641 691 52699 697
rect 52914 688 52920 700
rect 52972 728 52978 740
rect 52972 700 53788 728
rect 52972 688 52978 700
rect 53466 660 53472 672
rect 41800 632 53472 660
rect 53466 620 53472 632
rect 53524 620 53530 672
rect 53561 663 53619 669
rect 53561 629 53573 663
rect 53607 660 53619 663
rect 53650 660 53656 672
rect 53607 632 53656 660
rect 53607 629 53619 632
rect 53561 623 53619 629
rect 53650 620 53656 632
rect 53708 620 53714 672
rect 53760 660 53788 700
rect 55214 688 55220 740
rect 55272 728 55278 740
rect 56410 728 56416 740
rect 55272 700 56416 728
rect 55272 688 55278 700
rect 56410 688 56416 700
rect 56468 688 56474 740
rect 60366 688 60372 740
rect 60424 728 60430 740
rect 61120 728 61148 768
rect 61933 765 61945 768
rect 61979 765 61991 799
rect 61933 759 61991 765
rect 63497 799 63555 805
rect 63497 765 63509 799
rect 63543 765 63555 799
rect 63604 796 63632 836
rect 63770 824 63776 836
rect 63828 864 63834 876
rect 66456 873 66484 904
rect 68020 904 68385 932
rect 68020 873 68048 904
rect 68373 901 68385 904
rect 68419 932 68431 935
rect 68738 932 68744 944
rect 68419 904 68744 932
rect 68419 901 68431 904
rect 68373 895 68431 901
rect 68738 892 68744 904
rect 68796 892 68802 944
rect 68830 892 68836 944
rect 68888 932 68894 944
rect 70118 932 70124 944
rect 68888 904 70124 932
rect 68888 892 68894 904
rect 70118 892 70124 904
rect 70176 892 70182 944
rect 70581 935 70639 941
rect 70581 901 70593 935
rect 70627 932 70639 935
rect 70670 932 70676 944
rect 70627 904 70676 932
rect 70627 901 70639 904
rect 70581 895 70639 901
rect 70670 892 70676 904
rect 70728 892 70734 944
rect 70854 892 70860 944
rect 70912 932 70918 944
rect 70949 935 71007 941
rect 70949 932 70961 935
rect 70912 904 70961 932
rect 70912 892 70918 904
rect 70949 901 70961 904
rect 70995 901 71007 935
rect 71866 932 71872 944
rect 71827 904 71872 932
rect 70949 895 71007 901
rect 71866 892 71872 904
rect 71924 892 71930 944
rect 74813 935 74871 941
rect 74813 901 74825 935
rect 74859 932 74871 935
rect 75086 932 75092 944
rect 74859 904 75092 932
rect 74859 901 74871 904
rect 74813 895 74871 901
rect 75086 892 75092 904
rect 75144 892 75150 944
rect 75178 892 75184 944
rect 75236 932 75242 944
rect 80514 932 80520 944
rect 75236 904 80284 932
rect 80475 904 80520 932
rect 75236 892 75242 904
rect 64509 867 64567 873
rect 64509 864 64521 867
rect 63828 836 64521 864
rect 63828 824 63834 836
rect 64509 833 64521 836
rect 64555 833 64567 867
rect 64509 827 64567 833
rect 66441 867 66499 873
rect 66441 833 66453 867
rect 66487 833 66499 867
rect 66441 827 66499 833
rect 68005 867 68063 873
rect 68005 833 68017 867
rect 68051 833 68063 867
rect 69198 864 69204 876
rect 69159 836 69204 864
rect 68005 827 68063 833
rect 69198 824 69204 836
rect 69256 864 69262 876
rect 69937 867 69995 873
rect 69937 864 69949 867
rect 69256 836 69949 864
rect 69256 824 69262 836
rect 69937 833 69949 836
rect 69983 833 69995 867
rect 69937 827 69995 833
rect 70489 867 70547 873
rect 70489 833 70501 867
rect 70535 864 70547 867
rect 70872 864 70900 892
rect 70535 836 70900 864
rect 70535 833 70547 836
rect 70489 827 70547 833
rect 71774 824 71780 876
rect 71832 864 71838 876
rect 71961 867 72019 873
rect 71961 864 71973 867
rect 71832 836 71973 864
rect 71832 824 71838 836
rect 71961 833 71973 836
rect 72007 864 72019 867
rect 72881 867 72939 873
rect 72881 864 72893 867
rect 72007 836 72893 864
rect 72007 833 72019 836
rect 71961 827 72019 833
rect 72881 833 72893 836
rect 72927 833 72939 867
rect 72881 827 72939 833
rect 72970 824 72976 876
rect 73028 864 73034 876
rect 73433 867 73491 873
rect 73433 864 73445 867
rect 73028 836 73445 864
rect 73028 824 73034 836
rect 73433 833 73445 836
rect 73479 833 73491 867
rect 73433 827 73491 833
rect 76469 867 76527 873
rect 76469 833 76481 867
rect 76515 864 76527 867
rect 76650 864 76656 876
rect 76515 836 76656 864
rect 76515 833 76527 836
rect 76469 827 76527 833
rect 76650 824 76656 836
rect 76708 864 76714 876
rect 76837 867 76895 873
rect 76837 864 76849 867
rect 76708 836 76849 864
rect 76708 824 76714 836
rect 76837 833 76849 836
rect 76883 833 76895 867
rect 76837 827 76895 833
rect 77481 867 77539 873
rect 77481 833 77493 867
rect 77527 864 77539 867
rect 78033 867 78091 873
rect 78033 864 78045 867
rect 77527 836 78045 864
rect 77527 833 77539 836
rect 77481 827 77539 833
rect 78033 833 78045 836
rect 78079 864 78091 867
rect 79226 864 79232 876
rect 78079 836 79232 864
rect 78079 833 78091 836
rect 78033 827 78091 833
rect 79226 824 79232 836
rect 79284 824 79290 876
rect 79321 867 79379 873
rect 79321 833 79333 867
rect 79367 864 79379 867
rect 79410 864 79416 876
rect 79367 836 79416 864
rect 79367 833 79379 836
rect 79321 827 79379 833
rect 79410 824 79416 836
rect 79468 864 79474 876
rect 79689 867 79747 873
rect 79689 864 79701 867
rect 79468 836 79701 864
rect 79468 824 79474 836
rect 79689 833 79701 836
rect 79735 833 79747 867
rect 79689 827 79747 833
rect 67453 799 67511 805
rect 67453 796 67465 799
rect 63604 768 67465 796
rect 63497 759 63555 765
rect 67453 765 67465 768
rect 67499 765 67511 799
rect 68922 796 68928 808
rect 68883 768 68928 796
rect 67453 759 67511 765
rect 60424 700 61148 728
rect 60424 688 60430 700
rect 61194 688 61200 740
rect 61252 728 61258 740
rect 63512 728 63540 759
rect 68922 756 68928 768
rect 68980 756 68986 808
rect 69842 756 69848 808
rect 69900 796 69906 808
rect 74258 796 74264 808
rect 69900 768 74264 796
rect 69900 756 69906 768
rect 74258 756 74264 768
rect 74316 756 74322 808
rect 75822 796 75828 808
rect 75783 768 75828 796
rect 75822 756 75828 768
rect 75880 756 75886 808
rect 77570 796 77576 808
rect 77531 768 77576 796
rect 77570 756 77576 768
rect 77628 756 77634 808
rect 78674 796 78680 808
rect 78635 768 78680 796
rect 78674 756 78680 768
rect 78732 756 78738 808
rect 61252 700 63540 728
rect 61252 688 61258 700
rect 65058 688 65064 740
rect 65116 728 65122 740
rect 65610 728 65616 740
rect 65116 700 65616 728
rect 65116 688 65122 700
rect 65610 688 65616 700
rect 65668 688 65674 740
rect 68094 688 68100 740
rect 68152 728 68158 740
rect 68741 731 68799 737
rect 68741 728 68753 731
rect 68152 700 68753 728
rect 68152 688 68158 700
rect 68741 697 68753 700
rect 68787 728 68799 731
rect 69106 728 69112 740
rect 68787 700 69112 728
rect 68787 697 68799 700
rect 68741 691 68799 697
rect 69106 688 69112 700
rect 69164 688 69170 740
rect 70210 688 70216 740
rect 70268 728 70274 740
rect 75730 728 75736 740
rect 70268 700 75736 728
rect 70268 688 70274 700
rect 75730 688 75736 700
rect 75788 688 75794 740
rect 79594 728 79600 740
rect 75840 700 79600 728
rect 56042 660 56048 672
rect 53760 632 56048 660
rect 56042 620 56048 632
rect 56100 620 56106 672
rect 56226 620 56232 672
rect 56284 660 56290 672
rect 57422 660 57428 672
rect 56284 632 57428 660
rect 56284 620 56290 632
rect 57422 620 57428 632
rect 57480 620 57486 672
rect 59630 620 59636 672
rect 59688 660 59694 672
rect 60458 660 60464 672
rect 59688 632 60464 660
rect 59688 620 59694 632
rect 60458 620 60464 632
rect 60516 620 60522 672
rect 60642 620 60648 672
rect 60700 660 60706 672
rect 65426 660 65432 672
rect 60700 632 65432 660
rect 60700 620 60706 632
rect 65426 620 65432 632
rect 65484 620 65490 672
rect 65518 620 65524 672
rect 65576 660 65582 672
rect 75840 660 75868 700
rect 79594 688 79600 700
rect 79652 688 79658 740
rect 65576 632 75868 660
rect 80256 660 80284 904
rect 80514 892 80520 904
rect 80572 892 80578 944
rect 84749 935 84807 941
rect 84749 932 84761 935
rect 84212 904 84761 932
rect 81066 824 81072 876
rect 81124 864 81130 876
rect 81161 867 81219 873
rect 81161 864 81173 867
rect 81124 836 81173 864
rect 81124 824 81130 836
rect 81161 833 81173 836
rect 81207 864 81219 867
rect 81529 867 81587 873
rect 81529 864 81541 867
rect 81207 836 81541 864
rect 81207 833 81219 836
rect 81161 827 81219 833
rect 81529 833 81541 836
rect 81575 833 81587 867
rect 81529 827 81587 833
rect 82081 867 82139 873
rect 82081 833 82093 867
rect 82127 833 82139 867
rect 82081 827 82139 833
rect 83185 867 83243 873
rect 83185 833 83197 867
rect 83231 864 83243 867
rect 83458 864 83464 876
rect 83231 836 83464 864
rect 83231 833 83243 836
rect 83185 827 83243 833
rect 82096 796 82124 827
rect 83458 824 83464 836
rect 83516 864 83522 876
rect 84212 873 84240 904
rect 84749 901 84761 904
rect 84795 932 84807 935
rect 84838 932 84844 944
rect 84795 904 84844 932
rect 84795 901 84807 904
rect 84749 895 84807 901
rect 84838 892 84844 904
rect 84896 892 84902 944
rect 86310 892 86316 944
rect 86368 892 86374 944
rect 87969 935 88027 941
rect 87969 932 87981 935
rect 87432 904 87981 932
rect 83645 867 83703 873
rect 83645 864 83657 867
rect 83516 836 83657 864
rect 83516 824 83522 836
rect 83645 833 83657 836
rect 83691 833 83703 867
rect 83645 827 83703 833
rect 84197 867 84255 873
rect 84197 833 84209 867
rect 84243 833 84255 867
rect 84197 827 84255 833
rect 86037 867 86095 873
rect 86037 833 86049 867
rect 86083 864 86095 867
rect 86328 864 86356 892
rect 87432 873 87460 904
rect 87969 901 87981 904
rect 88015 932 88027 935
rect 89622 932 89628 944
rect 88015 904 89628 932
rect 88015 901 88027 904
rect 87969 895 88027 901
rect 89622 892 89628 904
rect 89680 892 89686 944
rect 89993 935 90051 941
rect 89993 901 90005 935
rect 90039 932 90051 935
rect 90174 932 90180 944
rect 90039 904 90180 932
rect 90039 901 90051 904
rect 89993 895 90051 901
rect 90174 892 90180 904
rect 90232 892 90238 944
rect 91833 935 91891 941
rect 91833 901 91845 935
rect 91879 932 91891 935
rect 92014 932 92020 944
rect 91879 904 92020 932
rect 91879 901 91891 904
rect 91833 895 91891 901
rect 92014 892 92020 904
rect 92072 892 92078 944
rect 92293 935 92351 941
rect 92293 901 92305 935
rect 92339 932 92351 935
rect 93670 932 93676 944
rect 92339 904 93676 932
rect 92339 901 92351 904
rect 92293 895 92351 901
rect 86497 867 86555 873
rect 86497 864 86509 867
rect 86083 836 86509 864
rect 86083 833 86095 836
rect 86037 827 86095 833
rect 86497 833 86509 836
rect 86543 833 86555 867
rect 86497 827 86555 833
rect 87417 867 87475 873
rect 87417 833 87429 867
rect 87463 833 87475 867
rect 87417 827 87475 833
rect 88610 824 88616 876
rect 88668 864 88674 876
rect 88889 867 88947 873
rect 88889 864 88901 867
rect 88668 836 88901 864
rect 88668 824 88674 836
rect 88889 833 88901 836
rect 88935 833 88947 867
rect 88889 827 88947 833
rect 82633 799 82691 805
rect 82633 796 82645 799
rect 82096 768 82645 796
rect 82633 765 82645 768
rect 82679 796 82691 799
rect 84010 796 84016 808
rect 82679 768 84016 796
rect 82679 765 82691 768
rect 82633 759 82691 765
rect 84010 756 84016 768
rect 84068 756 84074 808
rect 88904 796 88932 827
rect 89346 824 89352 876
rect 89404 864 89410 876
rect 89901 867 89959 873
rect 89901 864 89913 867
rect 89404 836 89913 864
rect 89404 824 89410 836
rect 89901 833 89913 836
rect 89947 864 89959 867
rect 90361 867 90419 873
rect 90361 864 90373 867
rect 89947 836 90373 864
rect 89947 833 89959 836
rect 89901 827 89959 833
rect 90361 833 90373 836
rect 90407 833 90419 867
rect 90361 827 90419 833
rect 91741 867 91799 873
rect 91741 833 91753 867
rect 91787 864 91799 867
rect 92308 864 92336 895
rect 93670 892 93676 904
rect 93728 892 93734 944
rect 94406 892 94412 944
rect 94464 932 94470 944
rect 103716 932 103744 972
rect 94464 904 103744 932
rect 103900 932 103928 972
rect 103977 969 103989 1003
rect 104023 1000 104035 1003
rect 104621 1003 104679 1009
rect 104621 1000 104633 1003
rect 104023 972 104633 1000
rect 104023 969 104035 972
rect 103977 963 104035 969
rect 104621 969 104633 972
rect 104667 1000 104679 1003
rect 104986 1000 104992 1012
rect 104667 972 104992 1000
rect 104667 969 104679 972
rect 104621 963 104679 969
rect 104986 960 104992 972
rect 105044 960 105050 1012
rect 105265 1003 105323 1009
rect 105265 969 105277 1003
rect 105311 1000 105323 1003
rect 107010 1000 107016 1012
rect 105311 972 107016 1000
rect 105311 969 105323 972
rect 105265 963 105323 969
rect 105170 932 105176 944
rect 103900 904 105176 932
rect 94464 892 94470 904
rect 105170 892 105176 904
rect 105228 892 105234 944
rect 91787 836 92336 864
rect 102321 867 102379 873
rect 91787 833 91799 836
rect 91741 827 91799 833
rect 102321 833 102333 867
rect 102367 864 102379 867
rect 103885 867 103943 873
rect 102367 836 103836 864
rect 102367 833 102379 836
rect 102321 827 102379 833
rect 89441 799 89499 805
rect 89441 796 89453 799
rect 88904 768 89453 796
rect 89441 765 89453 768
rect 89487 765 89499 799
rect 89441 759 89499 765
rect 102594 756 102600 808
rect 102652 796 102658 808
rect 103333 799 103391 805
rect 103333 796 103345 799
rect 102652 768 103345 796
rect 102652 756 102658 768
rect 103333 765 103345 768
rect 103379 765 103391 799
rect 103808 796 103836 836
rect 103885 833 103897 867
rect 103931 864 103943 867
rect 104250 864 104256 876
rect 103931 836 104256 864
rect 103931 833 103943 836
rect 103885 827 103943 833
rect 104250 824 104256 836
rect 104308 824 104314 876
rect 105372 873 105400 972
rect 107010 960 107016 972
rect 107068 960 107074 1012
rect 107838 1000 107844 1012
rect 107799 972 107844 1000
rect 107838 960 107844 972
rect 107896 960 107902 1012
rect 133509 1003 133567 1009
rect 133509 1000 133521 1003
rect 109144 972 133521 1000
rect 109144 932 109172 972
rect 133509 969 133521 972
rect 133555 969 133567 1003
rect 133690 1000 133696 1012
rect 133651 972 133696 1000
rect 133509 963 133567 969
rect 133690 960 133696 972
rect 133748 960 133754 1012
rect 133874 960 133880 1012
rect 133932 1000 133938 1012
rect 135622 1000 135628 1012
rect 133932 972 135628 1000
rect 133932 960 133938 972
rect 135622 960 135628 972
rect 135680 960 135686 1012
rect 136082 1000 136088 1012
rect 136043 972 136088 1000
rect 136082 960 136088 972
rect 136140 1000 136146 1012
rect 136361 1003 136419 1009
rect 136361 1000 136373 1003
rect 136140 972 136373 1000
rect 136140 960 136146 972
rect 136361 969 136373 972
rect 136407 969 136419 1003
rect 136361 963 136419 969
rect 139029 1003 139087 1009
rect 139029 969 139041 1003
rect 139075 1000 139087 1003
rect 139210 1000 139216 1012
rect 139075 972 139216 1000
rect 139075 969 139087 972
rect 139029 963 139087 969
rect 139210 960 139216 972
rect 139268 1000 139274 1012
rect 140774 1000 140780 1012
rect 139268 972 140780 1000
rect 139268 960 139274 972
rect 140774 960 140780 972
rect 140832 960 140838 1012
rect 141050 1000 141056 1012
rect 141011 972 141056 1000
rect 141050 960 141056 972
rect 141108 960 141114 1012
rect 143166 1000 143172 1012
rect 143127 972 143172 1000
rect 143166 960 143172 972
rect 143224 960 143230 1012
rect 155218 1000 155224 1012
rect 155179 972 155224 1000
rect 155218 960 155224 972
rect 155276 960 155282 1012
rect 155770 1000 155776 1012
rect 155731 972 155776 1000
rect 155770 960 155776 972
rect 155828 960 155834 1012
rect 156601 1003 156659 1009
rect 156601 969 156613 1003
rect 156647 1000 156659 1003
rect 158254 1000 158260 1012
rect 156647 972 158260 1000
rect 156647 969 156659 972
rect 156601 963 156659 969
rect 105464 904 109172 932
rect 105357 867 105415 873
rect 105357 833 105369 867
rect 105403 833 105415 867
rect 105357 827 105415 833
rect 103977 799 104035 805
rect 103977 796 103989 799
rect 103808 768 103989 796
rect 103333 759 103391 765
rect 103977 765 103989 768
rect 104023 765 104035 799
rect 103977 759 104035 765
rect 104986 756 104992 808
rect 105044 796 105050 808
rect 105464 796 105492 904
rect 109218 892 109224 944
rect 109276 932 109282 944
rect 110417 935 110475 941
rect 110417 932 110429 935
rect 109276 904 110429 932
rect 109276 892 109282 904
rect 110417 901 110429 904
rect 110463 901 110475 935
rect 110417 895 110475 901
rect 106090 824 106096 876
rect 106148 864 106154 876
rect 106461 867 106519 873
rect 106461 864 106473 867
rect 106148 836 106473 864
rect 106148 824 106154 836
rect 106461 833 106473 836
rect 106507 864 106519 867
rect 107197 867 107255 873
rect 107197 864 107209 867
rect 106507 836 107209 864
rect 106507 833 106519 836
rect 106461 827 106519 833
rect 107197 833 107209 836
rect 107243 833 107255 867
rect 110432 864 110460 895
rect 110782 892 110788 944
rect 110840 932 110846 944
rect 112717 935 112775 941
rect 112717 932 112729 935
rect 110840 904 112729 932
rect 110840 892 110846 904
rect 110877 867 110935 873
rect 110877 864 110889 867
rect 107197 827 107255 833
rect 107304 836 110368 864
rect 110432 836 110889 864
rect 106366 796 106372 808
rect 105044 768 105492 796
rect 106327 768 106372 796
rect 105044 756 105050 768
rect 106366 756 106372 768
rect 106424 756 106430 808
rect 82170 728 82176 740
rect 82131 700 82176 728
rect 82170 688 82176 700
rect 82228 688 82234 740
rect 87509 731 87567 737
rect 87509 728 87521 731
rect 82372 700 87521 728
rect 82372 660 82400 700
rect 87509 697 87521 700
rect 87555 697 87567 731
rect 88978 728 88984 740
rect 88939 700 88984 728
rect 87509 691 87567 697
rect 88978 688 88984 700
rect 89036 688 89042 740
rect 89070 688 89076 740
rect 89128 728 89134 740
rect 107304 728 107332 836
rect 107930 756 107936 808
rect 107988 796 107994 808
rect 109402 796 109408 808
rect 107988 768 109408 796
rect 107988 756 107994 768
rect 109402 756 109408 768
rect 109460 756 109466 808
rect 109589 799 109647 805
rect 109589 765 109601 799
rect 109635 765 109647 799
rect 110340 796 110368 836
rect 110877 833 110889 836
rect 110923 833 110935 867
rect 110877 827 110935 833
rect 111150 824 111156 876
rect 111208 864 111214 876
rect 111996 873 112024 904
rect 112717 901 112729 904
rect 112763 901 112775 935
rect 112717 895 112775 901
rect 113821 935 113879 941
rect 113821 901 113833 935
rect 113867 932 113879 935
rect 114002 932 114008 944
rect 113867 904 114008 932
rect 113867 901 113879 904
rect 113821 895 113879 901
rect 113928 873 113956 904
rect 114002 892 114008 904
rect 114060 892 114066 944
rect 116210 932 116216 944
rect 116171 904 116216 932
rect 116210 892 116216 904
rect 116268 932 116274 944
rect 116268 904 116440 932
rect 116268 892 116274 904
rect 111981 867 112039 873
rect 111208 836 111472 864
rect 111208 824 111214 836
rect 111444 796 111472 836
rect 111981 833 111993 867
rect 112027 833 112039 867
rect 111981 827 112039 833
rect 113913 867 113971 873
rect 113913 833 113925 867
rect 113959 833 113971 867
rect 115477 867 115535 873
rect 113913 827 113971 833
rect 114020 836 115060 864
rect 114020 796 114048 836
rect 114922 796 114928 808
rect 110340 768 111380 796
rect 111444 768 114048 796
rect 114883 768 114928 796
rect 109589 759 109647 765
rect 89128 700 107332 728
rect 109604 728 109632 759
rect 111242 728 111248 740
rect 109604 700 111248 728
rect 89128 688 89134 700
rect 111242 688 111248 700
rect 111300 688 111306 740
rect 111352 728 111380 768
rect 114922 756 114928 768
rect 114980 756 114986 808
rect 115032 796 115060 836
rect 115477 833 115489 867
rect 115523 864 115535 867
rect 115845 867 115903 873
rect 115845 864 115857 867
rect 115523 836 115857 864
rect 115523 833 115535 836
rect 115477 827 115535 833
rect 115845 833 115857 836
rect 115891 864 115903 867
rect 116302 864 116308 876
rect 115891 836 116308 864
rect 115891 833 115903 836
rect 115845 827 115903 833
rect 116302 824 116308 836
rect 116360 824 116366 876
rect 116412 873 116440 904
rect 116504 904 144224 932
rect 116397 867 116455 873
rect 116397 833 116409 867
rect 116443 833 116455 867
rect 116397 827 116455 833
rect 116504 796 116532 904
rect 117961 867 118019 873
rect 117961 833 117973 867
rect 118007 833 118019 867
rect 117961 827 118019 833
rect 115032 768 116532 796
rect 117409 799 117467 805
rect 117409 765 117421 799
rect 117455 765 117467 799
rect 117976 796 118004 827
rect 118142 824 118148 876
rect 118200 864 118206 876
rect 119065 867 119123 873
rect 118200 836 118556 864
rect 118200 824 118206 836
rect 118329 799 118387 805
rect 118329 796 118341 799
rect 117976 768 118341 796
rect 117409 759 117467 765
rect 118329 765 118341 768
rect 118375 796 118387 799
rect 118418 796 118424 808
rect 118375 768 118424 796
rect 118375 765 118387 768
rect 118329 759 118387 765
rect 112165 731 112223 737
rect 112165 728 112177 731
rect 111352 700 112177 728
rect 112165 697 112177 700
rect 112211 697 112223 731
rect 117424 728 117452 759
rect 118418 756 118424 768
rect 118476 756 118482 808
rect 118528 796 118556 836
rect 119065 833 119077 867
rect 119111 864 119123 867
rect 119249 867 119307 873
rect 119249 864 119261 867
rect 119111 836 119261 864
rect 119111 833 119123 836
rect 119065 827 119123 833
rect 119249 833 119261 836
rect 119295 864 119307 867
rect 119338 864 119344 876
rect 119295 836 119344 864
rect 119295 833 119307 836
rect 119249 827 119307 833
rect 119338 824 119344 836
rect 119396 824 119402 876
rect 120813 867 120871 873
rect 120813 833 120825 867
rect 120859 864 120871 867
rect 120905 867 120963 873
rect 120905 864 120917 867
rect 120859 836 120917 864
rect 120859 833 120871 836
rect 120813 827 120871 833
rect 120905 833 120917 836
rect 120951 833 120963 867
rect 120905 827 120963 833
rect 122101 867 122159 873
rect 122101 833 122113 867
rect 122147 864 122159 867
rect 122650 864 122656 876
rect 122147 836 122656 864
rect 122147 833 122159 836
rect 122101 827 122159 833
rect 122650 824 122656 836
rect 122708 824 122714 876
rect 123757 867 123815 873
rect 123757 833 123769 867
rect 123803 864 123815 867
rect 123938 864 123944 876
rect 123803 836 123944 864
rect 123803 833 123815 836
rect 123757 827 123815 833
rect 123938 824 123944 836
rect 123996 824 124002 876
rect 125594 824 125600 876
rect 125652 873 125658 876
rect 125652 864 125663 873
rect 126146 864 126152 876
rect 125652 836 125697 864
rect 126107 836 126152 864
rect 125652 827 125663 836
rect 125652 824 125658 827
rect 126146 824 126152 836
rect 126204 824 126210 876
rect 128265 867 128323 873
rect 128265 833 128277 867
rect 128311 864 128323 867
rect 128633 867 128691 873
rect 128633 864 128645 867
rect 128311 836 128645 864
rect 128311 833 128323 836
rect 128265 827 128323 833
rect 128633 833 128645 836
rect 128679 833 128691 867
rect 128633 827 128691 833
rect 129182 824 129188 876
rect 129240 864 129246 876
rect 129277 867 129335 873
rect 129277 864 129289 867
rect 129240 836 129289 864
rect 129240 824 129246 836
rect 129277 833 129289 836
rect 129323 833 129335 867
rect 129277 827 129335 833
rect 131117 867 131175 873
rect 131117 833 131129 867
rect 131163 864 131175 867
rect 131393 867 131451 873
rect 131393 864 131405 867
rect 131163 836 131405 864
rect 131163 833 131175 836
rect 131117 827 131175 833
rect 131393 833 131405 836
rect 131439 833 131451 867
rect 131393 827 131451 833
rect 132405 867 132463 873
rect 132405 833 132417 867
rect 132451 864 132463 867
rect 132954 864 132960 876
rect 132451 836 132960 864
rect 132451 833 132463 836
rect 132405 827 132463 833
rect 132954 824 132960 836
rect 133012 824 133018 876
rect 133690 824 133696 876
rect 133748 864 133754 876
rect 133877 867 133935 873
rect 133877 864 133889 867
rect 133748 836 133889 864
rect 133748 824 133754 836
rect 133877 833 133889 836
rect 133923 833 133935 867
rect 133877 827 133935 833
rect 135441 867 135499 873
rect 135441 833 135453 867
rect 135487 864 135499 867
rect 135809 867 135867 873
rect 135809 864 135821 867
rect 135487 836 135821 864
rect 135487 833 135499 836
rect 135441 827 135499 833
rect 135809 833 135821 836
rect 135855 864 135867 867
rect 136910 864 136916 876
rect 135855 836 136916 864
rect 135855 833 135867 836
rect 135809 827 135867 833
rect 136910 824 136916 836
rect 136968 824 136974 876
rect 137646 864 137652 876
rect 137607 836 137652 864
rect 137646 824 137652 836
rect 137704 864 137710 876
rect 138293 867 138351 873
rect 138293 864 138305 867
rect 137704 836 138305 864
rect 137704 824 137710 836
rect 138293 833 138305 836
rect 138339 833 138351 867
rect 138293 827 138351 833
rect 138845 867 138903 873
rect 138845 833 138857 867
rect 138891 864 138903 867
rect 140777 867 140835 873
rect 138891 836 140268 864
rect 138891 833 138903 836
rect 138845 827 138903 833
rect 133966 796 133972 808
rect 118528 768 133972 796
rect 133966 756 133972 768
rect 134024 756 134030 808
rect 134058 756 134064 808
rect 134116 796 134122 808
rect 134889 799 134947 805
rect 134889 796 134901 799
rect 134116 768 134901 796
rect 134116 756 134122 768
rect 134889 765 134901 768
rect 134935 765 134947 799
rect 134889 759 134947 765
rect 136361 799 136419 805
rect 136361 765 136373 799
rect 136407 796 136419 799
rect 136453 799 136511 805
rect 136453 796 136465 799
rect 136407 768 136465 796
rect 136407 765 136419 768
rect 136361 759 136419 765
rect 136453 765 136465 768
rect 136499 765 136511 799
rect 139210 796 139216 808
rect 139171 768 139216 796
rect 136453 759 136511 765
rect 139210 756 139216 768
rect 139268 756 139274 808
rect 140240 805 140268 836
rect 140777 833 140789 867
rect 140823 864 140835 867
rect 141050 864 141056 876
rect 140823 836 141056 864
rect 140823 833 140835 836
rect 140777 827 140835 833
rect 141050 824 141056 836
rect 141108 824 141114 876
rect 142057 867 142115 873
rect 142057 833 142069 867
rect 142103 833 142115 867
rect 142057 827 142115 833
rect 140225 799 140283 805
rect 140225 765 140237 799
rect 140271 765 140283 799
rect 140225 759 140283 765
rect 140866 756 140872 808
rect 140924 796 140930 808
rect 142080 796 142108 827
rect 142154 824 142160 876
rect 142212 864 142218 876
rect 143077 867 143135 873
rect 143077 864 143089 867
rect 142212 836 143089 864
rect 142212 824 142218 836
rect 143077 833 143089 836
rect 143123 864 143135 867
rect 143537 867 143595 873
rect 143537 864 143549 867
rect 143123 836 143549 864
rect 143123 833 143135 836
rect 143077 827 143135 833
rect 143537 833 143549 836
rect 143583 833 143595 867
rect 143537 827 143595 833
rect 142525 799 142583 805
rect 142525 796 142537 799
rect 140924 768 142537 796
rect 140924 756 140930 768
rect 142525 765 142537 768
rect 142571 765 142583 799
rect 142525 759 142583 765
rect 112165 691 112223 697
rect 113284 700 117452 728
rect 83274 660 83280 672
rect 80256 632 82400 660
rect 83235 632 83280 660
rect 65576 620 65582 632
rect 83274 620 83280 632
rect 83332 620 83338 672
rect 84286 660 84292 672
rect 84247 632 84292 660
rect 84286 620 84292 632
rect 84344 620 84350 672
rect 86126 660 86132 672
rect 86087 632 86132 660
rect 86126 620 86132 632
rect 86184 620 86190 672
rect 95602 620 95608 672
rect 95660 660 95666 672
rect 103054 660 103060 672
rect 95660 632 103060 660
rect 95660 620 95666 632
rect 103054 620 103060 632
rect 103112 620 103118 672
rect 104250 660 104256 672
rect 104211 632 104256 660
rect 104250 620 104256 632
rect 104308 620 104314 672
rect 106366 620 106372 672
rect 106424 660 106430 672
rect 113284 660 113312 700
rect 120074 688 120080 740
rect 120132 728 120138 740
rect 120537 731 120595 737
rect 120537 728 120549 731
rect 120132 700 120549 728
rect 120132 688 120138 700
rect 120537 697 120549 700
rect 120583 697 120595 731
rect 122193 731 122251 737
rect 122193 728 122205 731
rect 120537 691 120595 697
rect 120644 700 122205 728
rect 106424 632 113312 660
rect 106424 620 106430 632
rect 115566 620 115572 672
rect 115624 660 115630 672
rect 120644 660 120672 700
rect 122193 697 122205 700
rect 122239 697 122251 731
rect 122193 691 122251 697
rect 125689 731 125747 737
rect 125689 697 125701 731
rect 125735 728 125747 731
rect 125778 728 125784 740
rect 125735 700 125784 728
rect 125735 697 125747 700
rect 125689 691 125747 697
rect 125778 688 125784 700
rect 125836 688 125842 740
rect 131209 731 131267 737
rect 131209 728 131221 731
rect 126164 700 131221 728
rect 115624 632 120672 660
rect 120905 663 120963 669
rect 115624 620 115630 632
rect 120905 629 120917 663
rect 120951 660 120963 663
rect 121181 663 121239 669
rect 121181 660 121193 663
rect 120951 632 121193 660
rect 120951 629 120963 632
rect 120905 623 120963 629
rect 121181 629 121193 632
rect 121227 660 121239 663
rect 126164 660 126192 700
rect 131209 697 131221 700
rect 131255 697 131267 731
rect 131758 728 131764 740
rect 131209 691 131267 697
rect 131316 700 131764 728
rect 121227 632 126192 660
rect 121227 629 121239 632
rect 121181 623 121239 629
rect 126974 620 126980 672
rect 127032 660 127038 672
rect 128357 663 128415 669
rect 128357 660 128369 663
rect 127032 632 128369 660
rect 127032 620 127038 632
rect 128357 629 128369 632
rect 128403 629 128415 663
rect 128357 623 128415 629
rect 128633 663 128691 669
rect 128633 629 128645 663
rect 128679 660 128691 663
rect 128817 663 128875 669
rect 128817 660 128829 663
rect 128679 632 128829 660
rect 128679 629 128691 632
rect 128633 623 128691 629
rect 128817 629 128829 632
rect 128863 660 128875 663
rect 131316 660 131344 700
rect 131758 688 131764 700
rect 131816 688 131822 740
rect 137738 728 137744 740
rect 137699 700 137744 728
rect 137738 688 137744 700
rect 137796 688 137802 740
rect 137922 688 137928 740
rect 137980 728 137986 740
rect 144196 728 144224 904
rect 146018 824 146024 876
rect 146076 864 146082 876
rect 146297 867 146355 873
rect 146297 864 146309 867
rect 146076 836 146309 864
rect 146076 824 146082 836
rect 146297 833 146309 836
rect 146343 864 146355 867
rect 147033 867 147091 873
rect 147033 864 147045 867
rect 146343 836 147045 864
rect 146343 833 146355 836
rect 146297 827 146355 833
rect 147033 833 147045 836
rect 147079 833 147091 867
rect 151722 864 151728 876
rect 151683 836 151728 864
rect 147033 827 147091 833
rect 151722 824 151728 836
rect 151780 864 151786 876
rect 152461 867 152519 873
rect 152461 864 152473 867
rect 151780 836 152473 864
rect 151780 824 151786 836
rect 152461 833 152473 836
rect 152507 833 152519 867
rect 152461 827 152519 833
rect 156708 805 156736 972
rect 158254 960 158260 972
rect 158312 960 158318 1012
rect 158346 960 158352 1012
rect 158404 1000 158410 1012
rect 158533 1003 158591 1009
rect 158533 1000 158545 1003
rect 158404 972 158545 1000
rect 158404 960 158410 972
rect 158533 969 158545 972
rect 158579 969 158591 1003
rect 161290 1000 161296 1012
rect 158533 963 158591 969
rect 161032 972 161296 1000
rect 158257 867 158315 873
rect 158257 833 158269 867
rect 158303 864 158315 867
rect 158364 864 158392 960
rect 158303 836 158392 864
rect 158993 867 159051 873
rect 158303 833 158315 836
rect 158257 827 158315 833
rect 158993 833 159005 867
rect 159039 864 159051 867
rect 159450 864 159456 876
rect 159039 836 159456 864
rect 159039 833 159051 836
rect 158993 827 159051 833
rect 159450 824 159456 836
rect 159508 824 159514 876
rect 161032 873 161060 972
rect 161290 960 161296 972
rect 161348 960 161354 1012
rect 166629 1003 166687 1009
rect 166629 969 166641 1003
rect 166675 1000 166687 1003
rect 166810 1000 166816 1012
rect 166675 972 166816 1000
rect 166675 969 166687 972
rect 166629 963 166687 969
rect 166810 960 166816 972
rect 166868 960 166874 1012
rect 167733 935 167791 941
rect 167733 932 167745 935
rect 164988 904 167745 932
rect 161017 867 161075 873
rect 161017 833 161029 867
rect 161063 833 161075 867
rect 161017 827 161075 833
rect 161845 867 161903 873
rect 161845 833 161857 867
rect 161891 864 161903 867
rect 162026 864 162032 876
rect 161891 836 162032 864
rect 161891 833 161903 836
rect 161845 827 161903 833
rect 162026 824 162032 836
rect 162084 824 162090 876
rect 162762 824 162768 876
rect 162820 864 162826 876
rect 164988 873 165016 904
rect 167733 901 167745 904
rect 167779 901 167791 935
rect 167733 895 167791 901
rect 163133 867 163191 873
rect 163133 864 163145 867
rect 162820 836 163145 864
rect 162820 824 162826 836
rect 163133 833 163145 836
rect 163179 864 163191 867
rect 163869 867 163927 873
rect 163869 864 163881 867
rect 163179 836 163881 864
rect 163179 833 163191 836
rect 163133 827 163191 833
rect 163869 833 163881 836
rect 163915 833 163927 867
rect 163869 827 163927 833
rect 164697 867 164755 873
rect 164697 833 164709 867
rect 164743 864 164755 867
rect 164973 867 165031 873
rect 164973 864 164985 867
rect 164743 836 164985 864
rect 164743 833 164755 836
rect 164697 827 164755 833
rect 164973 833 164985 836
rect 165019 833 165031 867
rect 164973 827 165031 833
rect 166537 867 166595 873
rect 166537 833 166549 867
rect 166583 864 166595 867
rect 166629 867 166687 873
rect 166629 864 166641 867
rect 166583 836 166641 864
rect 166583 833 166595 836
rect 166537 827 166595 833
rect 166629 833 166641 836
rect 166675 833 166687 867
rect 166629 827 166687 833
rect 144733 799 144791 805
rect 144733 765 144745 799
rect 144779 796 144791 799
rect 145193 799 145251 805
rect 145193 796 145205 799
rect 144779 768 145205 796
rect 144779 765 144791 768
rect 144733 759 144791 765
rect 145193 765 145205 768
rect 145239 796 145251 799
rect 147769 799 147827 805
rect 147769 796 147781 799
rect 145239 768 147781 796
rect 145239 765 145251 768
rect 145193 759 145251 765
rect 147769 765 147781 768
rect 147815 765 147827 799
rect 147769 759 147827 765
rect 149517 799 149575 805
rect 149517 765 149529 799
rect 149563 796 149575 799
rect 150345 799 150403 805
rect 150345 796 150357 799
rect 149563 768 150357 796
rect 149563 765 149575 768
rect 149517 759 149575 765
rect 150345 765 150357 768
rect 150391 796 150403 799
rect 150621 799 150679 805
rect 150621 796 150633 799
rect 150391 768 150633 796
rect 150391 765 150403 768
rect 150345 759 150403 765
rect 150621 765 150633 768
rect 150667 765 150679 799
rect 156693 799 156751 805
rect 150621 759 150679 765
rect 150728 768 156644 796
rect 146481 731 146539 737
rect 146481 728 146493 731
rect 137980 700 144132 728
rect 144196 700 146493 728
rect 137980 688 137986 700
rect 128863 632 131344 660
rect 131393 663 131451 669
rect 128863 629 128875 632
rect 128817 623 128875 629
rect 131393 629 131405 663
rect 131439 660 131451 663
rect 131669 663 131727 669
rect 131669 660 131681 663
rect 131439 632 131681 660
rect 131439 629 131451 632
rect 131393 623 131451 629
rect 131669 629 131681 632
rect 131715 660 131727 663
rect 132126 660 132132 672
rect 131715 632 132132 660
rect 131715 629 131727 632
rect 131669 623 131727 629
rect 132126 620 132132 632
rect 132184 620 132190 672
rect 132494 660 132500 672
rect 132455 632 132500 660
rect 132494 620 132500 632
rect 132552 620 132558 672
rect 132954 660 132960 672
rect 132915 632 132960 660
rect 132954 620 132960 632
rect 133012 620 133018 672
rect 133601 663 133659 669
rect 133601 629 133613 663
rect 133647 660 133659 663
rect 138845 663 138903 669
rect 138845 660 138857 663
rect 133647 632 138857 660
rect 133647 629 133659 632
rect 133601 623 133659 629
rect 138845 629 138857 632
rect 138891 629 138903 663
rect 138845 623 138903 629
rect 142157 663 142215 669
rect 142157 629 142169 663
rect 142203 660 142215 663
rect 143994 660 144000 672
rect 142203 632 144000 660
rect 142203 629 142215 632
rect 142157 623 142215 629
rect 143994 620 144000 632
rect 144052 620 144058 672
rect 144104 660 144132 700
rect 146481 697 146493 700
rect 146527 697 146539 731
rect 146481 691 146539 697
rect 150728 660 150756 768
rect 151906 728 151912 740
rect 151867 700 151912 728
rect 151906 688 151912 700
rect 151964 688 151970 740
rect 156616 728 156644 768
rect 156693 765 156705 799
rect 156739 765 156751 799
rect 156693 759 156751 765
rect 156782 756 156788 808
rect 156840 796 156846 808
rect 157705 799 157763 805
rect 157705 796 157717 799
rect 156840 768 157717 796
rect 156840 756 156846 768
rect 157705 765 157717 768
rect 157751 765 157763 799
rect 160462 796 160468 808
rect 160423 768 160468 796
rect 157705 759 157763 765
rect 160462 756 160468 768
rect 160520 756 160526 808
rect 163041 799 163099 805
rect 163041 765 163053 799
rect 163087 765 163099 799
rect 165982 796 165988 808
rect 165943 768 165988 796
rect 163041 759 163099 765
rect 163056 728 163084 759
rect 165982 756 165988 768
rect 166040 756 166046 808
rect 156616 700 163084 728
rect 144104 632 150756 660
rect 368 570 93012 592
rect 368 518 28456 570
rect 28508 518 28520 570
rect 28572 518 28584 570
rect 28636 518 28648 570
rect 28700 518 84878 570
rect 84930 518 84942 570
rect 84994 518 85006 570
rect 85058 518 85070 570
rect 85122 518 93012 570
rect 368 496 93012 518
rect 102028 570 169556 592
rect 102028 518 141299 570
rect 141351 518 141363 570
rect 141415 518 141427 570
rect 141479 518 141491 570
rect 141543 518 169556 570
rect 102028 496 169556 518
rect 8754 416 8760 468
rect 8812 456 8818 468
rect 27522 456 27528 468
rect 8812 428 27528 456
rect 8812 416 8818 428
rect 27522 416 27528 428
rect 27580 416 27586 468
rect 28810 416 28816 468
rect 28868 456 28874 468
rect 32766 456 32772 468
rect 28868 428 32772 456
rect 28868 416 28874 428
rect 32766 416 32772 428
rect 32824 416 32830 468
rect 32858 416 32864 468
rect 32916 456 32922 468
rect 42334 456 42340 468
rect 32916 428 42340 456
rect 32916 416 32922 428
rect 42334 416 42340 428
rect 42392 416 42398 468
rect 42429 459 42487 465
rect 42429 425 42441 459
rect 42475 456 42487 459
rect 42794 456 42800 468
rect 42475 428 42800 456
rect 42475 425 42487 428
rect 42429 419 42487 425
rect 42794 416 42800 428
rect 42852 416 42858 468
rect 42978 416 42984 468
rect 43036 456 43042 468
rect 50890 456 50896 468
rect 43036 428 50896 456
rect 43036 416 43042 428
rect 50890 416 50896 428
rect 50948 416 50954 468
rect 50985 459 51043 465
rect 50985 425 50997 459
rect 51031 456 51043 459
rect 52730 456 52736 468
rect 51031 428 52736 456
rect 51031 425 51043 428
rect 50985 419 51043 425
rect 52730 416 52736 428
rect 52788 416 52794 468
rect 53006 416 53012 468
rect 53064 456 53070 468
rect 57146 456 57152 468
rect 53064 428 57152 456
rect 53064 416 53070 428
rect 57146 416 57152 428
rect 57204 416 57210 468
rect 57422 416 57428 468
rect 57480 456 57486 468
rect 68922 456 68928 468
rect 57480 428 68928 456
rect 57480 416 57486 428
rect 68922 416 68928 428
rect 68980 416 68986 468
rect 69106 416 69112 468
rect 69164 456 69170 468
rect 72970 456 72976 468
rect 69164 428 72976 456
rect 69164 416 69170 428
rect 72970 416 72976 428
rect 73028 416 73034 468
rect 81618 416 81624 468
rect 81676 456 81682 468
rect 89070 456 89076 468
rect 81676 428 89076 456
rect 81676 416 81682 428
rect 89070 416 89076 428
rect 89128 416 89134 468
rect 101122 416 101128 468
rect 101180 456 101186 468
rect 137738 456 137744 468
rect 101180 428 137744 456
rect 101180 416 101186 428
rect 137738 416 137744 428
rect 137796 416 137802 468
rect 138290 416 138296 468
rect 138348 456 138354 468
rect 140866 456 140872 468
rect 138348 428 140872 456
rect 138348 416 138354 428
rect 140866 416 140872 428
rect 140924 416 140930 468
rect 10962 348 10968 400
rect 11020 388 11026 400
rect 19242 388 19248 400
rect 11020 360 19248 388
rect 11020 348 11026 360
rect 19242 348 19248 360
rect 19300 348 19306 400
rect 23474 348 23480 400
rect 23532 388 23538 400
rect 81986 388 81992 400
rect 23532 360 81992 388
rect 23532 348 23538 360
rect 81986 348 81992 360
rect 82044 348 82050 400
rect 98546 348 98552 400
rect 98604 388 98610 400
rect 114922 388 114928 400
rect 98604 360 114928 388
rect 98604 348 98610 360
rect 114922 348 114928 360
rect 114980 348 114986 400
rect 132126 348 132132 400
rect 132184 388 132190 400
rect 140314 388 140320 400
rect 132184 360 140320 388
rect 132184 348 132190 360
rect 140314 348 140320 360
rect 140372 348 140378 400
rect 17218 280 17224 332
rect 17276 320 17282 332
rect 82170 320 82176 332
rect 17276 292 82176 320
rect 17276 280 17282 292
rect 82170 280 82176 292
rect 82228 280 82234 332
rect 95050 280 95056 332
rect 95108 320 95114 332
rect 95108 292 96660 320
rect 95108 280 95114 292
rect 21266 212 21272 264
rect 21324 252 21330 264
rect 83274 252 83280 264
rect 21324 224 83280 252
rect 21324 212 21330 224
rect 83274 212 83280 224
rect 83332 212 83338 264
rect 96632 252 96660 292
rect 104802 280 104808 332
rect 104860 320 104866 332
rect 111337 323 111395 329
rect 111337 320 111349 323
rect 104860 292 111349 320
rect 104860 280 104866 292
rect 111337 289 111349 292
rect 111383 289 111395 323
rect 111337 283 111395 289
rect 111429 323 111487 329
rect 111429 289 111441 323
rect 111475 320 111487 323
rect 114462 320 114468 332
rect 111475 292 114468 320
rect 111475 289 111487 292
rect 111429 283 111487 289
rect 114462 280 114468 292
rect 114520 280 114526 332
rect 118418 280 118424 332
rect 118476 320 118482 332
rect 132034 320 132040 332
rect 118476 292 132040 320
rect 118476 280 118482 292
rect 132034 280 132040 292
rect 132092 280 132098 332
rect 132954 280 132960 332
rect 133012 320 133018 332
rect 134153 323 134211 329
rect 134153 320 134165 323
rect 133012 292 134165 320
rect 133012 280 133018 292
rect 134153 289 134165 292
rect 134199 289 134211 323
rect 134153 283 134211 289
rect 107930 252 107936 264
rect 96632 224 107936 252
rect 107930 212 107936 224
rect 107988 212 107994 264
rect 108114 212 108120 264
rect 108172 252 108178 264
rect 160462 252 160468 264
rect 108172 224 160468 252
rect 108172 212 108178 224
rect 160462 212 160468 224
rect 160520 212 160526 264
rect 30834 144 30840 196
rect 30892 184 30898 196
rect 91370 184 91376 196
rect 30892 156 91376 184
rect 30892 144 30898 156
rect 91370 144 91376 156
rect 91428 144 91434 196
rect 106274 144 106280 196
rect 106332 184 106338 196
rect 151906 184 151912 196
rect 106332 156 151912 184
rect 106332 144 106338 156
rect 151906 144 151912 156
rect 151964 144 151970 196
rect 24026 76 24032 128
rect 24084 116 24090 128
rect 36446 116 36452 128
rect 24084 88 36308 116
rect 36407 88 36452 116
rect 24084 76 24090 88
rect 18046 8 18052 60
rect 18104 48 18110 60
rect 34330 48 34336 60
rect 18104 20 34336 48
rect 18104 8 18110 20
rect 34330 8 34336 20
rect 34388 8 34394 60
rect 34514 8 34520 60
rect 34572 48 34578 60
rect 35802 48 35808 60
rect 34572 20 35808 48
rect 34572 8 34578 20
rect 35802 8 35808 20
rect 35860 8 35866 60
rect 36280 48 36308 88
rect 36446 76 36452 88
rect 36504 76 36510 128
rect 36538 76 36544 128
rect 36596 116 36602 128
rect 36633 119 36691 125
rect 36633 116 36645 119
rect 36596 88 36645 116
rect 36596 76 36602 88
rect 36633 85 36645 88
rect 36679 85 36691 119
rect 36633 79 36691 85
rect 36722 76 36728 128
rect 36780 116 36786 128
rect 40954 116 40960 128
rect 36780 88 40960 116
rect 36780 76 36786 88
rect 40954 76 40960 88
rect 41012 76 41018 128
rect 41049 119 41107 125
rect 41049 85 41061 119
rect 41095 116 41107 119
rect 41095 88 41276 116
rect 41095 85 41107 88
rect 41049 79 41107 85
rect 41138 48 41144 60
rect 36280 20 41144 48
rect 41138 8 41144 20
rect 41196 8 41202 60
rect 41248 48 41276 88
rect 41322 76 41328 128
rect 41380 116 41386 128
rect 42153 119 42211 125
rect 42153 116 42165 119
rect 41380 88 42165 116
rect 41380 76 41386 88
rect 42153 85 42165 88
rect 42199 85 42211 119
rect 42153 79 42211 85
rect 42245 119 42303 125
rect 42245 85 42257 119
rect 42291 116 42303 119
rect 47394 116 47400 128
rect 42291 88 47400 116
rect 42291 85 42303 88
rect 42245 79 42303 85
rect 47394 76 47400 88
rect 47452 76 47458 128
rect 47578 76 47584 128
rect 47636 116 47642 128
rect 48130 116 48136 128
rect 47636 88 48136 116
rect 47636 76 47642 88
rect 48130 76 48136 88
rect 48188 116 48194 128
rect 50154 116 50160 128
rect 48188 88 50160 116
rect 48188 76 48194 88
rect 50154 76 50160 88
rect 50212 76 50218 128
rect 50338 76 50344 128
rect 50396 116 50402 128
rect 78674 116 78680 128
rect 50396 88 78680 116
rect 50396 76 50402 88
rect 78674 76 78680 88
rect 78732 76 78738 128
rect 104250 76 104256 128
rect 104308 116 104314 128
rect 111245 119 111303 125
rect 111245 116 111257 119
rect 104308 88 111257 116
rect 104308 76 104314 88
rect 111245 85 111257 88
rect 111291 85 111303 119
rect 111245 79 111303 85
rect 111337 119 111395 125
rect 111337 85 111349 119
rect 111383 116 111395 119
rect 134058 116 134064 128
rect 111383 88 134064 116
rect 111383 85 111395 88
rect 111337 79 111395 85
rect 134058 76 134064 88
rect 134116 76 134122 128
rect 134153 119 134211 125
rect 134153 85 134165 119
rect 134199 116 134211 119
rect 139118 116 139124 128
rect 134199 88 139124 116
rect 134199 85 134211 88
rect 134153 79 134211 85
rect 139118 76 139124 88
rect 139176 76 139182 128
rect 49881 51 49939 57
rect 49881 48 49893 51
rect 41248 20 49893 48
rect 49881 17 49893 20
rect 49927 17 49939 51
rect 49881 11 49939 17
rect 49970 8 49976 60
rect 50028 48 50034 60
rect 75822 48 75828 60
rect 50028 20 75828 48
rect 50028 8 50034 20
rect 75822 8 75828 20
rect 75880 8 75886 60
rect 107746 8 107752 60
rect 107804 48 107810 60
rect 156782 48 156788 60
rect 107804 20 156788 48
rect 107804 8 107810 20
rect 156782 8 156788 20
rect 156840 8 156846 60
<< via1 >>
rect 50896 12928 50948 12980
rect 56508 12928 56560 12980
rect 66076 12928 66128 12980
rect 32220 12860 32272 12912
rect 35900 12860 35952 12912
rect 35992 12860 36044 12912
rect 41328 12792 41380 12844
rect 46296 12860 46348 12912
rect 70860 12860 70912 12912
rect 22376 12724 22428 12776
rect 40408 12724 40460 12776
rect 45928 12724 45980 12776
rect 46480 12724 46532 12776
rect 83280 12656 83332 12708
rect 26240 12588 26292 12640
rect 41696 12588 41748 12640
rect 41788 12588 41840 12640
rect 66352 12588 66404 12640
rect 98184 12588 98236 12640
rect 121644 12588 121696 12640
rect 23296 12520 23348 12572
rect 38016 12520 38068 12572
rect 38936 12520 38988 12572
rect 40960 12520 41012 12572
rect 41052 12520 41104 12572
rect 41512 12520 41564 12572
rect 55680 12520 55732 12572
rect 61292 12520 61344 12572
rect 109960 12520 110012 12572
rect 123208 12520 123260 12572
rect 50712 12452 50764 12504
rect 56140 12452 56192 12504
rect 56968 12452 57020 12504
rect 59452 12452 59504 12504
rect 96896 12452 96948 12504
rect 121368 12452 121420 12504
rect 136640 12452 136692 12504
rect 145104 12452 145156 12504
rect 29000 12384 29052 12436
rect 32496 12384 32548 12436
rect 34428 12384 34480 12436
rect 35624 12427 35676 12436
rect 35624 12393 35633 12427
rect 35633 12393 35667 12427
rect 35667 12393 35676 12427
rect 35624 12384 35676 12393
rect 83004 12384 83056 12436
rect 110512 12384 110564 12436
rect 123484 12384 123536 12436
rect 137008 12384 137060 12436
rect 152464 12384 152516 12436
rect 11520 12316 11572 12368
rect 75000 12316 75052 12368
rect 144736 12316 144788 12368
rect 163872 12316 163924 12368
rect 24584 12248 24636 12300
rect 32496 12248 32548 12300
rect 24492 12180 24544 12232
rect 28448 12180 28500 12232
rect 29184 12180 29236 12232
rect 38384 12248 38436 12300
rect 38568 12248 38620 12300
rect 58256 12248 58308 12300
rect 67824 12248 67876 12300
rect 72424 12248 72476 12300
rect 83096 12248 83148 12300
rect 108488 12248 108540 12300
rect 121276 12248 121328 12300
rect 121920 12248 121972 12300
rect 126888 12248 126940 12300
rect 137376 12248 137428 12300
rect 162952 12248 163004 12300
rect 53104 12180 53156 12232
rect 55404 12180 55456 12232
rect 65616 12180 65668 12232
rect 79048 12180 79100 12232
rect 108028 12180 108080 12232
rect 125600 12180 125652 12232
rect 137192 12180 137244 12232
rect 137836 12180 137888 12232
rect 165896 12180 165948 12232
rect 4528 12112 4580 12164
rect 27620 12112 27672 12164
rect 32496 12155 32548 12164
rect 32496 12121 32505 12155
rect 32505 12121 32539 12155
rect 32539 12121 32548 12155
rect 32496 12112 32548 12121
rect 34060 12112 34112 12164
rect 46204 12112 46256 12164
rect 61200 12112 61252 12164
rect 68008 12112 68060 12164
rect 80428 12112 80480 12164
rect 103152 12112 103204 12164
rect 111524 12112 111576 12164
rect 113364 12112 113416 12164
rect 119620 12112 119672 12164
rect 119988 12112 120040 12164
rect 23388 12087 23440 12096
rect 23388 12053 23397 12087
rect 23397 12053 23431 12087
rect 23431 12053 23440 12087
rect 23388 12044 23440 12053
rect 24216 12044 24268 12096
rect 26884 12044 26936 12096
rect 27528 12044 27580 12096
rect 27896 12044 27948 12096
rect 30656 12044 30708 12096
rect 30748 12044 30800 12096
rect 31944 12044 31996 12096
rect 37096 12044 37148 12096
rect 37188 12044 37240 12096
rect 39580 12044 39632 12096
rect 55864 12044 55916 12096
rect 64512 12044 64564 12096
rect 73620 12044 73672 12096
rect 76840 12044 76892 12096
rect 77944 12087 77996 12096
rect 77944 12053 77953 12087
rect 77953 12053 77987 12087
rect 77987 12053 77996 12087
rect 77944 12044 77996 12053
rect 80244 12044 80296 12096
rect 82912 12044 82964 12096
rect 101404 12044 101456 12096
rect 118332 12044 118384 12096
rect 118700 12044 118752 12096
rect 127900 12112 127952 12164
rect 132868 12112 132920 12164
rect 134340 12112 134392 12164
rect 146760 12112 146812 12164
rect 149060 12112 149112 12164
rect 153292 12112 153344 12164
rect 135260 12044 135312 12096
rect 135444 12044 135496 12096
rect 160376 12044 160428 12096
rect 56667 11942 56719 11994
rect 56731 11942 56783 11994
rect 56795 11942 56847 11994
rect 56859 11942 56911 11994
rect 113088 11942 113140 11994
rect 113152 11942 113204 11994
rect 113216 11942 113268 11994
rect 113280 11942 113332 11994
rect 9680 11772 9732 11824
rect 14464 11772 14516 11824
rect 4804 11747 4856 11756
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 8024 11704 8076 11756
rect 20720 11704 20772 11756
rect 22376 11747 22428 11756
rect 6276 11636 6328 11688
rect 9680 11636 9732 11688
rect 14464 11636 14516 11688
rect 20168 11636 20220 11688
rect 20812 11679 20864 11688
rect 20812 11645 20821 11679
rect 20821 11645 20855 11679
rect 20855 11645 20864 11679
rect 20812 11636 20864 11645
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 24584 11704 24636 11756
rect 29092 11840 29144 11892
rect 32036 11840 32088 11892
rect 26608 11704 26660 11756
rect 29000 11704 29052 11756
rect 30932 11772 30984 11824
rect 41144 11840 41196 11892
rect 41236 11840 41288 11892
rect 42248 11840 42300 11892
rect 42432 11840 42484 11892
rect 43812 11840 43864 11892
rect 46204 11840 46256 11892
rect 55864 11840 55916 11892
rect 60832 11840 60884 11892
rect 63224 11883 63276 11892
rect 63224 11849 63233 11883
rect 63233 11849 63267 11883
rect 63267 11849 63276 11883
rect 63224 11840 63276 11849
rect 33508 11772 33560 11824
rect 17684 11568 17736 11620
rect 27252 11636 27304 11688
rect 27344 11636 27396 11688
rect 32588 11704 32640 11756
rect 29368 11636 29420 11688
rect 31576 11636 31628 11688
rect 35256 11704 35308 11756
rect 37188 11772 37240 11824
rect 34244 11636 34296 11688
rect 37004 11679 37056 11688
rect 37004 11645 37013 11679
rect 37013 11645 37047 11679
rect 37047 11645 37056 11679
rect 37004 11636 37056 11645
rect 37188 11636 37240 11688
rect 38568 11747 38620 11756
rect 38568 11713 38577 11747
rect 38577 11713 38611 11747
rect 38611 11713 38620 11747
rect 38568 11704 38620 11713
rect 39212 11704 39264 11756
rect 39856 11704 39908 11756
rect 40776 11704 40828 11756
rect 41052 11747 41104 11756
rect 41052 11713 41061 11747
rect 41061 11713 41095 11747
rect 41095 11713 41104 11747
rect 41052 11704 41104 11713
rect 41144 11704 41196 11756
rect 41788 11704 41840 11756
rect 37648 11636 37700 11688
rect 47124 11704 47176 11756
rect 49148 11704 49200 11756
rect 49608 11747 49660 11756
rect 49608 11713 49617 11747
rect 49617 11713 49651 11747
rect 49651 11713 49660 11747
rect 49608 11704 49660 11713
rect 49792 11704 49844 11756
rect 52736 11704 52788 11756
rect 53472 11704 53524 11756
rect 54576 11704 54628 11756
rect 56324 11704 56376 11756
rect 56508 11747 56560 11756
rect 56508 11713 56517 11747
rect 56517 11713 56551 11747
rect 56551 11713 56560 11747
rect 56508 11704 56560 11713
rect 56876 11704 56928 11756
rect 57428 11704 57480 11756
rect 57796 11747 57848 11756
rect 57796 11713 57805 11747
rect 57805 11713 57839 11747
rect 57839 11713 57848 11747
rect 57796 11704 57848 11713
rect 58072 11747 58124 11756
rect 58072 11713 58081 11747
rect 58081 11713 58115 11747
rect 58115 11713 58124 11747
rect 58072 11704 58124 11713
rect 58256 11772 58308 11824
rect 65616 11772 65668 11824
rect 61384 11704 61436 11756
rect 61660 11704 61712 11756
rect 62488 11704 62540 11756
rect 64696 11747 64748 11756
rect 64696 11713 64705 11747
rect 64705 11713 64739 11747
rect 64739 11713 64748 11747
rect 64696 11704 64748 11713
rect 65156 11747 65208 11756
rect 65156 11713 65165 11747
rect 65165 11713 65199 11747
rect 65199 11713 65208 11747
rect 65156 11704 65208 11713
rect 42064 11636 42116 11688
rect 46296 11636 46348 11688
rect 46480 11636 46532 11688
rect 49240 11636 49292 11688
rect 49424 11636 49476 11688
rect 49700 11636 49752 11688
rect 50712 11636 50764 11688
rect 51172 11636 51224 11688
rect 51816 11679 51868 11688
rect 51816 11645 51825 11679
rect 51825 11645 51859 11679
rect 51859 11645 51868 11679
rect 51816 11636 51868 11645
rect 54944 11636 54996 11688
rect 55128 11636 55180 11688
rect 56784 11636 56836 11688
rect 60924 11636 60976 11688
rect 65892 11636 65944 11688
rect 67824 11679 67876 11688
rect 67824 11645 67833 11679
rect 67833 11645 67867 11679
rect 67867 11645 67876 11679
rect 67824 11636 67876 11645
rect 67916 11636 67968 11688
rect 70308 11704 70360 11756
rect 71688 11704 71740 11756
rect 71872 11704 71924 11756
rect 72332 11747 72384 11756
rect 72332 11713 72341 11747
rect 72341 11713 72375 11747
rect 72375 11713 72384 11747
rect 72332 11704 72384 11713
rect 74356 11840 74408 11892
rect 74448 11840 74500 11892
rect 79048 11883 79100 11892
rect 75828 11772 75880 11824
rect 79048 11849 79057 11883
rect 79057 11849 79091 11883
rect 79091 11849 79100 11883
rect 79048 11840 79100 11849
rect 83280 11883 83332 11892
rect 83280 11849 83289 11883
rect 83289 11849 83323 11883
rect 83323 11849 83332 11883
rect 83280 11840 83332 11849
rect 108212 11840 108264 11892
rect 108488 11840 108540 11892
rect 108948 11840 109000 11892
rect 118700 11840 118752 11892
rect 118792 11883 118844 11892
rect 118792 11849 118801 11883
rect 118801 11849 118835 11883
rect 118835 11849 118844 11883
rect 118792 11840 118844 11849
rect 124036 11840 124088 11892
rect 125600 11840 125652 11892
rect 132684 11840 132736 11892
rect 134708 11840 134760 11892
rect 152464 11840 152516 11892
rect 74816 11747 74868 11756
rect 74816 11713 74825 11747
rect 74825 11713 74859 11747
rect 74859 11713 74868 11747
rect 74816 11704 74868 11713
rect 70492 11679 70544 11688
rect 70492 11645 70501 11679
rect 70501 11645 70535 11679
rect 70535 11645 70544 11679
rect 70492 11636 70544 11645
rect 72884 11636 72936 11688
rect 75460 11704 75512 11756
rect 77668 11704 77720 11756
rect 78772 11704 78824 11756
rect 82176 11772 82228 11824
rect 96896 11815 96948 11824
rect 80980 11704 81032 11756
rect 75368 11636 75420 11688
rect 77576 11679 77628 11688
rect 77576 11645 77585 11679
rect 77585 11645 77619 11679
rect 77619 11645 77628 11679
rect 77576 11636 77628 11645
rect 80060 11636 80112 11688
rect 80152 11636 80204 11688
rect 28356 11568 28408 11620
rect 28448 11568 28500 11620
rect 81716 11636 81768 11688
rect 82544 11704 82596 11756
rect 83372 11704 83424 11756
rect 96896 11781 96905 11815
rect 96905 11781 96939 11815
rect 96939 11781 96948 11815
rect 96896 11772 96948 11781
rect 84752 11704 84804 11756
rect 87144 11747 87196 11756
rect 87144 11713 87153 11747
rect 87153 11713 87187 11747
rect 87187 11713 87196 11747
rect 87144 11704 87196 11713
rect 92664 11704 92716 11756
rect 93308 11747 93360 11756
rect 93308 11713 93317 11747
rect 93317 11713 93351 11747
rect 93351 11713 93360 11747
rect 93308 11704 93360 11713
rect 98184 11747 98236 11756
rect 98184 11713 98193 11747
rect 98193 11713 98227 11747
rect 98227 11713 98236 11747
rect 98184 11704 98236 11713
rect 104072 11704 104124 11756
rect 86960 11636 87012 11688
rect 91744 11679 91796 11688
rect 91744 11645 91753 11679
rect 91753 11645 91787 11679
rect 91787 11645 91796 11679
rect 91744 11636 91796 11645
rect 93124 11679 93176 11688
rect 93124 11645 93133 11679
rect 93133 11645 93167 11679
rect 93167 11645 93176 11679
rect 93124 11636 93176 11645
rect 93676 11679 93728 11688
rect 93676 11645 93685 11679
rect 93685 11645 93719 11679
rect 93719 11645 93728 11679
rect 93676 11636 93728 11645
rect 99472 11636 99524 11688
rect 101864 11636 101916 11688
rect 112260 11772 112312 11824
rect 107752 11747 107804 11756
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 6092 11500 6144 11552
rect 9680 11500 9732 11552
rect 9772 11500 9824 11552
rect 17316 11500 17368 11552
rect 20076 11500 20128 11552
rect 27068 11500 27120 11552
rect 27436 11500 27488 11552
rect 27528 11500 27580 11552
rect 35532 11500 35584 11552
rect 35624 11500 35676 11552
rect 41328 11500 41380 11552
rect 50160 11500 50212 11552
rect 50252 11500 50304 11552
rect 52184 11500 52236 11552
rect 52460 11543 52512 11552
rect 52460 11509 52469 11543
rect 52469 11509 52503 11543
rect 52503 11509 52512 11543
rect 52460 11500 52512 11509
rect 53104 11543 53156 11552
rect 53104 11509 53113 11543
rect 53113 11509 53147 11543
rect 53147 11509 53156 11543
rect 53104 11500 53156 11509
rect 53196 11500 53248 11552
rect 56140 11500 56192 11552
rect 59728 11543 59780 11552
rect 59728 11509 59737 11543
rect 59737 11509 59771 11543
rect 59771 11509 59780 11543
rect 59728 11500 59780 11509
rect 60648 11500 60700 11552
rect 61200 11500 61252 11552
rect 64512 11543 64564 11552
rect 64512 11509 64521 11543
rect 64521 11509 64555 11543
rect 64555 11509 64564 11543
rect 64512 11500 64564 11509
rect 69020 11543 69072 11552
rect 69020 11509 69029 11543
rect 69029 11509 69063 11543
rect 69063 11509 69072 11543
rect 69020 11500 69072 11509
rect 70584 11500 70636 11552
rect 72792 11543 72844 11552
rect 72792 11509 72801 11543
rect 72801 11509 72835 11543
rect 72835 11509 72844 11543
rect 72792 11500 72844 11509
rect 74632 11500 74684 11552
rect 76288 11543 76340 11552
rect 76288 11509 76297 11543
rect 76297 11509 76331 11543
rect 76331 11509 76340 11543
rect 76288 11500 76340 11509
rect 76748 11500 76800 11552
rect 80152 11543 80204 11552
rect 80152 11509 80161 11543
rect 80161 11509 80195 11543
rect 80195 11509 80204 11543
rect 80152 11500 80204 11509
rect 88340 11500 88392 11552
rect 95516 11543 95568 11552
rect 95516 11509 95525 11543
rect 95525 11509 95559 11543
rect 95559 11509 95568 11543
rect 95516 11500 95568 11509
rect 96620 11500 96672 11552
rect 98276 11543 98328 11552
rect 98276 11509 98285 11543
rect 98285 11509 98319 11543
rect 98319 11509 98328 11543
rect 98276 11500 98328 11509
rect 106556 11636 106608 11688
rect 107752 11713 107761 11747
rect 107761 11713 107795 11747
rect 107795 11713 107804 11747
rect 107752 11704 107804 11713
rect 109868 11704 109920 11756
rect 109960 11704 110012 11756
rect 122196 11772 122248 11824
rect 124772 11772 124824 11824
rect 128452 11772 128504 11824
rect 112996 11747 113048 11756
rect 109040 11636 109092 11688
rect 104900 11568 104952 11620
rect 112996 11713 113005 11747
rect 113005 11713 113039 11747
rect 113039 11713 113048 11747
rect 112996 11704 113048 11713
rect 111708 11679 111760 11688
rect 111708 11645 111717 11679
rect 111717 11645 111751 11679
rect 111751 11645 111760 11679
rect 111708 11636 111760 11645
rect 115572 11704 115624 11756
rect 116492 11704 116544 11756
rect 114652 11636 114704 11688
rect 116308 11636 116360 11688
rect 114100 11568 114152 11620
rect 118332 11747 118384 11756
rect 118332 11713 118341 11747
rect 118341 11713 118375 11747
rect 118375 11713 118384 11747
rect 118332 11704 118384 11713
rect 118884 11704 118936 11756
rect 120264 11679 120316 11688
rect 120264 11645 120273 11679
rect 120273 11645 120307 11679
rect 120307 11645 120316 11679
rect 120264 11636 120316 11645
rect 121920 11704 121972 11756
rect 123116 11747 123168 11756
rect 123116 11713 123125 11747
rect 123125 11713 123159 11747
rect 123159 11713 123168 11747
rect 123116 11704 123168 11713
rect 123208 11747 123260 11756
rect 123208 11713 123217 11747
rect 123217 11713 123251 11747
rect 123251 11713 123260 11747
rect 123208 11704 123260 11713
rect 124312 11704 124364 11756
rect 125140 11704 125192 11756
rect 105268 11500 105320 11552
rect 107108 11543 107160 11552
rect 107108 11509 107117 11543
rect 107117 11509 107151 11543
rect 107151 11509 107160 11543
rect 107108 11500 107160 11509
rect 107844 11543 107896 11552
rect 107844 11509 107853 11543
rect 107853 11509 107887 11543
rect 107887 11509 107896 11543
rect 107844 11500 107896 11509
rect 109960 11500 110012 11552
rect 110880 11500 110932 11552
rect 111248 11543 111300 11552
rect 111248 11509 111257 11543
rect 111257 11509 111291 11543
rect 111291 11509 111300 11543
rect 111248 11500 111300 11509
rect 116492 11543 116544 11552
rect 116492 11509 116501 11543
rect 116501 11509 116535 11543
rect 116535 11509 116544 11543
rect 116492 11500 116544 11509
rect 117964 11543 118016 11552
rect 117964 11509 117973 11543
rect 117973 11509 118007 11543
rect 118007 11509 118016 11543
rect 117964 11500 118016 11509
rect 118608 11568 118660 11620
rect 126980 11636 127032 11688
rect 121736 11568 121788 11620
rect 124404 11568 124456 11620
rect 127716 11636 127768 11688
rect 128084 11704 128136 11756
rect 130660 11772 130712 11824
rect 130476 11704 130528 11756
rect 131764 11704 131816 11756
rect 133236 11747 133288 11756
rect 129740 11636 129792 11688
rect 132500 11636 132552 11688
rect 132684 11679 132736 11688
rect 132684 11645 132693 11679
rect 132693 11645 132727 11679
rect 132727 11645 132736 11679
rect 132684 11636 132736 11645
rect 133236 11713 133245 11747
rect 133245 11713 133279 11747
rect 133279 11713 133288 11747
rect 133236 11704 133288 11713
rect 135076 11772 135128 11824
rect 137192 11704 137244 11756
rect 138388 11747 138440 11756
rect 138388 11713 138397 11747
rect 138397 11713 138431 11747
rect 138431 11713 138440 11747
rect 138388 11704 138440 11713
rect 143356 11704 143408 11756
rect 143908 11704 143960 11756
rect 144828 11704 144880 11756
rect 146760 11704 146812 11756
rect 150440 11704 150492 11756
rect 151452 11704 151504 11756
rect 154488 11747 154540 11756
rect 154488 11713 154497 11747
rect 154497 11713 154531 11747
rect 154531 11713 154540 11747
rect 154488 11704 154540 11713
rect 136088 11636 136140 11688
rect 160192 11747 160244 11756
rect 160192 11713 160201 11747
rect 160201 11713 160235 11747
rect 160235 11713 160244 11747
rect 160192 11704 160244 11713
rect 160376 11704 160428 11756
rect 162216 11704 162268 11756
rect 162952 11704 163004 11756
rect 165896 11747 165948 11756
rect 165896 11713 165905 11747
rect 165905 11713 165939 11747
rect 165939 11713 165948 11747
rect 165896 11704 165948 11713
rect 167184 11704 167236 11756
rect 140228 11679 140280 11688
rect 140228 11645 140237 11679
rect 140237 11645 140271 11679
rect 140271 11645 140280 11679
rect 140228 11636 140280 11645
rect 140320 11636 140372 11688
rect 144552 11679 144604 11688
rect 144552 11645 144561 11679
rect 144561 11645 144595 11679
rect 144595 11645 144604 11679
rect 144552 11636 144604 11645
rect 146484 11636 146536 11688
rect 118792 11500 118844 11552
rect 119252 11500 119304 11552
rect 130660 11568 130712 11620
rect 144920 11568 144972 11620
rect 145104 11568 145156 11620
rect 156144 11636 156196 11688
rect 156880 11636 156932 11688
rect 166080 11636 166132 11688
rect 151636 11568 151688 11620
rect 159548 11568 159600 11620
rect 164332 11568 164384 11620
rect 124680 11543 124732 11552
rect 124680 11509 124689 11543
rect 124689 11509 124723 11543
rect 124723 11509 124732 11543
rect 124680 11500 124732 11509
rect 126152 11500 126204 11552
rect 130200 11500 130252 11552
rect 131304 11500 131356 11552
rect 134340 11543 134392 11552
rect 134340 11509 134349 11543
rect 134349 11509 134383 11543
rect 134383 11509 134392 11543
rect 134340 11500 134392 11509
rect 135628 11543 135680 11552
rect 135628 11509 135637 11543
rect 135637 11509 135671 11543
rect 135671 11509 135680 11543
rect 135628 11500 135680 11509
rect 135996 11543 136048 11552
rect 135996 11509 136005 11543
rect 136005 11509 136039 11543
rect 136039 11509 136048 11543
rect 135996 11500 136048 11509
rect 137468 11543 137520 11552
rect 137468 11509 137477 11543
rect 137477 11509 137511 11543
rect 137511 11509 137520 11543
rect 137468 11500 137520 11509
rect 138112 11543 138164 11552
rect 138112 11509 138121 11543
rect 138121 11509 138155 11543
rect 138155 11509 138164 11543
rect 138112 11500 138164 11509
rect 144000 11543 144052 11552
rect 144000 11509 144009 11543
rect 144009 11509 144043 11543
rect 144043 11509 144052 11543
rect 144000 11500 144052 11509
rect 146944 11543 146996 11552
rect 146944 11509 146953 11543
rect 146953 11509 146987 11543
rect 146987 11509 146996 11543
rect 146944 11500 146996 11509
rect 150992 11543 151044 11552
rect 150992 11509 151001 11543
rect 151001 11509 151035 11543
rect 151035 11509 151044 11543
rect 150992 11500 151044 11509
rect 153200 11500 153252 11552
rect 155960 11500 156012 11552
rect 157432 11543 157484 11552
rect 157432 11509 157441 11543
rect 157441 11509 157475 11543
rect 157475 11509 157484 11543
rect 157432 11500 157484 11509
rect 163044 11500 163096 11552
rect 166724 11500 166776 11552
rect 28456 11398 28508 11450
rect 28520 11398 28572 11450
rect 28584 11398 28636 11450
rect 28648 11398 28700 11450
rect 84878 11398 84930 11450
rect 84942 11398 84994 11450
rect 85006 11398 85058 11450
rect 85070 11398 85122 11450
rect 141299 11398 141351 11450
rect 141363 11398 141415 11450
rect 141427 11398 141479 11450
rect 141491 11398 141543 11450
rect 4804 11339 4856 11348
rect 4804 11305 4813 11339
rect 4813 11305 4847 11339
rect 4847 11305 4856 11339
rect 4804 11296 4856 11305
rect 11520 11296 11572 11348
rect 16488 11339 16540 11348
rect 16488 11305 16497 11339
rect 16497 11305 16531 11339
rect 16531 11305 16540 11339
rect 16488 11296 16540 11305
rect 22376 11339 22428 11348
rect 22376 11305 22385 11339
rect 22385 11305 22419 11339
rect 22419 11305 22428 11339
rect 22376 11296 22428 11305
rect 27988 11296 28040 11348
rect 29184 11339 29236 11348
rect 29184 11305 29193 11339
rect 29193 11305 29227 11339
rect 29227 11305 29236 11339
rect 29184 11296 29236 11305
rect 29368 11296 29420 11348
rect 31300 11296 31352 11348
rect 33140 11296 33192 11348
rect 34060 11339 34112 11348
rect 34060 11305 34069 11339
rect 34069 11305 34103 11339
rect 34103 11305 34112 11339
rect 34060 11296 34112 11305
rect 34980 11296 35032 11348
rect 39764 11296 39816 11348
rect 43720 11339 43772 11348
rect 43720 11305 43729 11339
rect 43729 11305 43763 11339
rect 43763 11305 43772 11339
rect 43720 11296 43772 11305
rect 45836 11296 45888 11348
rect 46296 11296 46348 11348
rect 46572 11296 46624 11348
rect 70768 11339 70820 11348
rect 70768 11305 70777 11339
rect 70777 11305 70811 11339
rect 70811 11305 70820 11339
rect 70768 11296 70820 11305
rect 72332 11339 72384 11348
rect 72332 11305 72341 11339
rect 72341 11305 72375 11339
rect 72375 11305 72384 11339
rect 72332 11296 72384 11305
rect 74448 11339 74500 11348
rect 74448 11305 74457 11339
rect 74457 11305 74491 11339
rect 74491 11305 74500 11339
rect 74448 11296 74500 11305
rect 75000 11339 75052 11348
rect 75000 11305 75009 11339
rect 75009 11305 75043 11339
rect 75043 11305 75052 11339
rect 75000 11296 75052 11305
rect 75368 11339 75420 11348
rect 75368 11305 75377 11339
rect 75377 11305 75411 11339
rect 75411 11305 75420 11339
rect 75368 11296 75420 11305
rect 77668 11339 77720 11348
rect 77668 11305 77677 11339
rect 77677 11305 77711 11339
rect 77711 11305 77720 11339
rect 77668 11296 77720 11305
rect 77944 11339 77996 11348
rect 77944 11305 77953 11339
rect 77953 11305 77987 11339
rect 77987 11305 77996 11339
rect 77944 11296 77996 11305
rect 78772 11296 78824 11348
rect 80980 11296 81032 11348
rect 83004 11339 83056 11348
rect 83004 11305 83013 11339
rect 83013 11305 83047 11339
rect 83047 11305 83056 11339
rect 83004 11296 83056 11305
rect 83372 11339 83424 11348
rect 83372 11305 83381 11339
rect 83381 11305 83415 11339
rect 83415 11305 83424 11339
rect 83372 11296 83424 11305
rect 84752 11339 84804 11348
rect 84752 11305 84761 11339
rect 84761 11305 84795 11339
rect 84795 11305 84804 11339
rect 84752 11296 84804 11305
rect 87144 11339 87196 11348
rect 87144 11305 87153 11339
rect 87153 11305 87187 11339
rect 87187 11305 87196 11339
rect 87144 11296 87196 11305
rect 98184 11339 98236 11348
rect 98184 11305 98193 11339
rect 98193 11305 98227 11339
rect 98227 11305 98236 11339
rect 98184 11296 98236 11305
rect 101404 11339 101456 11348
rect 101404 11305 101413 11339
rect 101413 11305 101447 11339
rect 101447 11305 101456 11339
rect 101404 11296 101456 11305
rect 104072 11339 104124 11348
rect 104072 11305 104081 11339
rect 104081 11305 104115 11339
rect 104115 11305 104124 11339
rect 104072 11296 104124 11305
rect 104900 11339 104952 11348
rect 104900 11305 104909 11339
rect 104909 11305 104943 11339
rect 104943 11305 104952 11339
rect 104900 11296 104952 11305
rect 105268 11339 105320 11348
rect 105268 11305 105277 11339
rect 105277 11305 105311 11339
rect 105311 11305 105320 11339
rect 105268 11296 105320 11305
rect 106556 11339 106608 11348
rect 106556 11305 106565 11339
rect 106565 11305 106599 11339
rect 106599 11305 106608 11339
rect 106556 11296 106608 11305
rect 3700 11228 3752 11280
rect 5724 11228 5776 11280
rect 9772 11228 9824 11280
rect 19892 11228 19944 11280
rect 22100 11228 22152 11280
rect 24216 11271 24268 11280
rect 24216 11237 24225 11271
rect 24225 11237 24259 11271
rect 24259 11237 24268 11271
rect 24216 11228 24268 11237
rect 24584 11271 24636 11280
rect 24584 11237 24593 11271
rect 24593 11237 24627 11271
rect 24627 11237 24636 11271
rect 24584 11228 24636 11237
rect 26608 11271 26660 11280
rect 26608 11237 26617 11271
rect 26617 11237 26651 11271
rect 26651 11237 26660 11271
rect 26608 11228 26660 11237
rect 4344 11160 4396 11212
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 7656 11203 7708 11212
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 6092 11092 6144 11144
rect 7656 11169 7665 11203
rect 7665 11169 7699 11203
rect 7699 11169 7708 11203
rect 7656 11160 7708 11169
rect 9680 11160 9732 11212
rect 16948 11160 17000 11212
rect 19156 11160 19208 11212
rect 28724 11228 28776 11280
rect 30748 11271 30800 11280
rect 30748 11237 30757 11271
rect 30757 11237 30791 11271
rect 30791 11237 30800 11271
rect 30748 11228 30800 11237
rect 33416 11228 33468 11280
rect 37740 11228 37792 11280
rect 27068 11160 27120 11212
rect 28264 11203 28316 11212
rect 28264 11169 28273 11203
rect 28273 11169 28307 11203
rect 28307 11169 28316 11203
rect 28264 11160 28316 11169
rect 8024 11135 8076 11144
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 4068 11024 4120 11076
rect 8576 11024 8628 11076
rect 12624 11024 12676 11076
rect 16488 11092 16540 11144
rect 20076 11092 20128 11144
rect 23388 11092 23440 11144
rect 24216 11092 24268 11144
rect 31944 11160 31996 11212
rect 32404 11160 32456 11212
rect 32588 11160 32640 11212
rect 35532 11203 35584 11212
rect 19708 11024 19760 11076
rect 20812 11024 20864 11076
rect 24860 11024 24912 11076
rect 11428 10956 11480 11008
rect 24308 10956 24360 11008
rect 24676 10999 24728 11008
rect 24676 10965 24685 10999
rect 24685 10965 24719 10999
rect 24719 10965 24728 10999
rect 24676 10956 24728 10965
rect 24768 10956 24820 11008
rect 27436 11024 27488 11076
rect 29644 11092 29696 11144
rect 30748 11092 30800 11144
rect 32496 11092 32548 11144
rect 29092 11024 29144 11076
rect 32128 11024 32180 11076
rect 35532 11169 35541 11203
rect 35541 11169 35575 11203
rect 35575 11169 35584 11203
rect 35532 11160 35584 11169
rect 36728 11160 36780 11212
rect 37004 11203 37056 11212
rect 37004 11169 37013 11203
rect 37013 11169 37047 11203
rect 37047 11169 37056 11203
rect 37004 11160 37056 11169
rect 37096 11160 37148 11212
rect 48780 11228 48832 11280
rect 49148 11271 49200 11280
rect 49148 11237 49157 11271
rect 49157 11237 49191 11271
rect 49191 11237 49200 11271
rect 49148 11228 49200 11237
rect 49240 11228 49292 11280
rect 51080 11228 51132 11280
rect 56968 11228 57020 11280
rect 58900 11228 58952 11280
rect 59084 11228 59136 11280
rect 60924 11228 60976 11280
rect 61292 11228 61344 11280
rect 61384 11228 61436 11280
rect 69940 11228 69992 11280
rect 38016 11203 38068 11212
rect 38016 11169 38025 11203
rect 38025 11169 38059 11203
rect 38059 11169 38068 11203
rect 38016 11160 38068 11169
rect 34612 11024 34664 11076
rect 36176 11092 36228 11144
rect 37648 11092 37700 11144
rect 72424 11160 72476 11212
rect 72792 11160 72844 11212
rect 38936 11067 38988 11076
rect 38936 11033 38945 11067
rect 38945 11033 38979 11067
rect 38979 11033 38988 11067
rect 38936 11024 38988 11033
rect 27252 10956 27304 11008
rect 27528 10956 27580 11008
rect 27620 10956 27672 11008
rect 32312 10956 32364 11008
rect 32496 10956 32548 11008
rect 37556 10956 37608 11008
rect 37648 10956 37700 11008
rect 38752 10956 38804 11008
rect 39396 10956 39448 11008
rect 41052 11092 41104 11144
rect 40592 11024 40644 11076
rect 42800 11092 42852 11144
rect 45652 11092 45704 11144
rect 45836 11135 45888 11144
rect 45836 11101 45845 11135
rect 45845 11101 45879 11135
rect 45879 11101 45888 11135
rect 45836 11092 45888 11101
rect 45928 11092 45980 11144
rect 46664 11092 46716 11144
rect 47124 11135 47176 11144
rect 47124 11101 47133 11135
rect 47133 11101 47167 11135
rect 47167 11101 47176 11135
rect 47124 11092 47176 11101
rect 48688 11092 48740 11144
rect 48780 11092 48832 11144
rect 49424 11092 49476 11144
rect 49700 11135 49752 11144
rect 49700 11101 49709 11135
rect 49709 11101 49743 11135
rect 49743 11101 49752 11135
rect 49700 11092 49752 11101
rect 46388 11024 46440 11076
rect 49608 11067 49660 11076
rect 40776 10999 40828 11008
rect 40776 10965 40785 10999
rect 40785 10965 40819 10999
rect 40819 10965 40828 10999
rect 40776 10956 40828 10965
rect 40960 10956 41012 11008
rect 41788 10956 41840 11008
rect 42064 10956 42116 11008
rect 46664 10956 46716 11008
rect 47032 10956 47084 11008
rect 48228 10999 48280 11008
rect 48228 10965 48237 10999
rect 48237 10965 48271 10999
rect 48271 10965 48280 10999
rect 48228 10956 48280 10965
rect 49608 11033 49617 11067
rect 49617 11033 49651 11067
rect 49651 11033 49660 11067
rect 50252 11092 50304 11144
rect 50528 11092 50580 11144
rect 50712 11092 50764 11144
rect 50988 11135 51040 11144
rect 50988 11101 50997 11135
rect 50997 11101 51031 11135
rect 51031 11101 51040 11135
rect 50988 11092 51040 11101
rect 52460 11135 52512 11144
rect 52460 11101 52469 11135
rect 52469 11101 52503 11135
rect 52503 11101 52512 11135
rect 52460 11092 52512 11101
rect 55128 11135 55180 11144
rect 49608 11024 49660 11033
rect 50160 11024 50212 11076
rect 53564 11067 53616 11076
rect 53564 11033 53573 11067
rect 53573 11033 53607 11067
rect 53607 11033 53616 11067
rect 53564 11024 53616 11033
rect 54668 11024 54720 11076
rect 55128 11101 55137 11135
rect 55137 11101 55171 11135
rect 55171 11101 55180 11135
rect 55128 11092 55180 11101
rect 55312 11135 55364 11144
rect 55312 11101 55321 11135
rect 55321 11101 55355 11135
rect 55355 11101 55364 11135
rect 55312 11092 55364 11101
rect 55496 11135 55548 11144
rect 55496 11101 55505 11135
rect 55505 11101 55539 11135
rect 55539 11101 55548 11135
rect 55496 11092 55548 11101
rect 56048 11135 56100 11144
rect 56048 11101 56057 11135
rect 56057 11101 56091 11135
rect 56091 11101 56100 11135
rect 56048 11092 56100 11101
rect 56508 11092 56560 11144
rect 56784 11135 56836 11144
rect 56784 11101 56793 11135
rect 56793 11101 56827 11135
rect 56827 11101 56836 11135
rect 56784 11092 56836 11101
rect 57152 11092 57204 11144
rect 59544 11092 59596 11144
rect 59728 11135 59780 11144
rect 59728 11101 59737 11135
rect 59737 11101 59771 11135
rect 59771 11101 59780 11135
rect 59728 11092 59780 11101
rect 61292 11135 61344 11144
rect 61292 11101 61301 11135
rect 61301 11101 61335 11135
rect 61335 11101 61344 11135
rect 61292 11092 61344 11101
rect 63408 11092 63460 11144
rect 63592 11135 63644 11144
rect 63592 11101 63601 11135
rect 63601 11101 63635 11135
rect 63635 11101 63644 11135
rect 63592 11092 63644 11101
rect 64696 11135 64748 11144
rect 64696 11101 64705 11135
rect 64705 11101 64739 11135
rect 64739 11101 64748 11135
rect 64696 11092 64748 11101
rect 67916 11092 67968 11144
rect 68928 11135 68980 11144
rect 68928 11101 68937 11135
rect 68937 11101 68971 11135
rect 68971 11101 68980 11135
rect 68928 11092 68980 11101
rect 70308 11092 70360 11144
rect 70584 11092 70636 11144
rect 71136 11092 71188 11144
rect 57796 11024 57848 11076
rect 65156 11024 65208 11076
rect 69572 11024 69624 11076
rect 79140 11228 79192 11280
rect 73528 11203 73580 11212
rect 73528 11169 73537 11203
rect 73537 11169 73571 11203
rect 73571 11169 73580 11203
rect 73528 11160 73580 11169
rect 76196 11160 76248 11212
rect 74724 11092 74776 11144
rect 76012 11092 76064 11144
rect 76748 11092 76800 11144
rect 76840 11135 76892 11144
rect 76840 11101 76849 11135
rect 76849 11101 76883 11135
rect 76883 11101 76892 11135
rect 80428 11203 80480 11212
rect 80428 11169 80437 11203
rect 80437 11169 80471 11203
rect 80471 11169 80480 11203
rect 80428 11160 80480 11169
rect 81716 11203 81768 11212
rect 81716 11169 81725 11203
rect 81725 11169 81759 11203
rect 81759 11169 81768 11203
rect 81716 11160 81768 11169
rect 76840 11092 76892 11101
rect 80060 11092 80112 11144
rect 82452 11228 82504 11280
rect 81992 11160 82044 11212
rect 82912 11135 82964 11144
rect 74816 11067 74868 11076
rect 74816 11033 74825 11067
rect 74825 11033 74859 11067
rect 74859 11033 74868 11067
rect 74816 11024 74868 11033
rect 82912 11101 82921 11135
rect 82921 11101 82955 11135
rect 82955 11101 82964 11135
rect 93308 11228 93360 11280
rect 96804 11228 96856 11280
rect 93676 11160 93728 11212
rect 93860 11160 93912 11212
rect 95516 11203 95568 11212
rect 95516 11169 95525 11203
rect 95525 11169 95559 11203
rect 95559 11169 95568 11203
rect 95516 11160 95568 11169
rect 99472 11203 99524 11212
rect 99472 11169 99481 11203
rect 99481 11169 99515 11203
rect 99515 11169 99524 11203
rect 99472 11160 99524 11169
rect 82912 11092 82964 11101
rect 96620 11135 96672 11144
rect 51448 10956 51500 11008
rect 51540 10956 51592 11008
rect 53012 10956 53064 11008
rect 54576 10956 54628 11008
rect 55128 10956 55180 11008
rect 57152 10956 57204 11008
rect 58072 10999 58124 11008
rect 58072 10965 58081 10999
rect 58081 10965 58115 10999
rect 58115 10965 58124 10999
rect 58072 10956 58124 10965
rect 58440 10956 58492 11008
rect 60464 10956 60516 11008
rect 61936 10956 61988 11008
rect 62488 10999 62540 11008
rect 62488 10965 62497 10999
rect 62497 10965 62531 10999
rect 62531 10965 62540 10999
rect 62488 10956 62540 10965
rect 65248 10956 65300 11008
rect 65340 10956 65392 11008
rect 85764 11024 85816 11076
rect 87512 11067 87564 11076
rect 87512 11033 87521 11067
rect 87521 11033 87555 11067
rect 87555 11033 87564 11067
rect 87512 11024 87564 11033
rect 91744 11067 91796 11076
rect 91744 11033 91753 11067
rect 91753 11033 91787 11067
rect 91787 11033 91796 11067
rect 91744 11024 91796 11033
rect 92020 11067 92072 11076
rect 92020 11033 92029 11067
rect 92029 11033 92063 11067
rect 92063 11033 92072 11067
rect 92020 11024 92072 11033
rect 96620 11101 96629 11135
rect 96629 11101 96663 11135
rect 96663 11101 96672 11135
rect 96620 11092 96672 11101
rect 108028 11228 108080 11280
rect 101864 11203 101916 11212
rect 101864 11169 101873 11203
rect 101873 11169 101907 11203
rect 101907 11169 101916 11203
rect 101864 11160 101916 11169
rect 103152 11203 103204 11212
rect 103152 11169 103161 11203
rect 103161 11169 103195 11203
rect 103195 11169 103204 11203
rect 103152 11160 103204 11169
rect 100668 11024 100720 11076
rect 107108 11160 107160 11212
rect 110880 11203 110932 11212
rect 110880 11169 110889 11203
rect 110889 11169 110923 11203
rect 110923 11169 110932 11203
rect 111248 11203 111300 11212
rect 110880 11160 110932 11169
rect 111248 11169 111257 11203
rect 111257 11169 111291 11203
rect 111291 11169 111300 11203
rect 111248 11160 111300 11169
rect 108212 11135 108264 11144
rect 108212 11101 108221 11135
rect 108221 11101 108255 11135
rect 108255 11101 108264 11135
rect 108212 11092 108264 11101
rect 108580 11135 108632 11144
rect 108580 11101 108589 11135
rect 108589 11101 108623 11135
rect 108623 11101 108632 11135
rect 108580 11092 108632 11101
rect 110512 11135 110564 11144
rect 110512 11101 110521 11135
rect 110521 11101 110555 11135
rect 110555 11101 110564 11135
rect 110512 11092 110564 11101
rect 78312 10956 78364 11008
rect 85948 10999 86000 11008
rect 85948 10965 85957 10999
rect 85957 10965 85991 10999
rect 85991 10965 86000 10999
rect 85948 10956 86000 10965
rect 90364 10999 90416 11008
rect 90364 10965 90373 10999
rect 90373 10965 90407 10999
rect 90407 10965 90416 10999
rect 90364 10956 90416 10965
rect 107752 10956 107804 11008
rect 108580 10956 108632 11008
rect 109040 10999 109092 11008
rect 109040 10965 109049 10999
rect 109049 10965 109083 10999
rect 109083 10965 109092 10999
rect 110972 11024 111024 11076
rect 118608 11296 118660 11348
rect 121276 11339 121328 11348
rect 121276 11305 121285 11339
rect 121285 11305 121319 11339
rect 121319 11305 121328 11339
rect 121276 11296 121328 11305
rect 121736 11339 121788 11348
rect 121736 11305 121745 11339
rect 121745 11305 121779 11339
rect 121779 11305 121788 11339
rect 121736 11296 121788 11305
rect 121920 11296 121972 11348
rect 123116 11339 123168 11348
rect 123116 11305 123125 11339
rect 123125 11305 123159 11339
rect 123159 11305 123168 11339
rect 123116 11296 123168 11305
rect 124312 11296 124364 11348
rect 114468 11228 114520 11280
rect 112996 11160 113048 11212
rect 123392 11271 123444 11280
rect 123392 11237 123401 11271
rect 123401 11237 123435 11271
rect 123435 11237 123444 11271
rect 123392 11228 123444 11237
rect 125508 11228 125560 11280
rect 115020 11203 115072 11212
rect 115020 11169 115029 11203
rect 115029 11169 115063 11203
rect 115063 11169 115072 11203
rect 115020 11160 115072 11169
rect 115204 11160 115256 11212
rect 117964 11203 118016 11212
rect 117964 11169 117973 11203
rect 117973 11169 118007 11203
rect 118007 11169 118016 11203
rect 117964 11160 118016 11169
rect 118700 11160 118752 11212
rect 115572 11135 115624 11144
rect 115572 11101 115581 11135
rect 115581 11101 115615 11135
rect 115615 11101 115624 11135
rect 115572 11092 115624 11101
rect 113732 11024 113784 11076
rect 114652 11024 114704 11076
rect 116584 11024 116636 11076
rect 122932 11160 122984 11212
rect 125324 11203 125376 11212
rect 120264 11067 120316 11076
rect 120264 11033 120273 11067
rect 120273 11033 120307 11067
rect 120307 11033 120316 11067
rect 120264 11024 120316 11033
rect 124680 11092 124732 11144
rect 125324 11169 125333 11203
rect 125333 11169 125367 11203
rect 125367 11169 125376 11203
rect 125324 11160 125376 11169
rect 127164 11296 127216 11348
rect 127716 11339 127768 11348
rect 127716 11305 127725 11339
rect 127725 11305 127759 11339
rect 127759 11305 127768 11339
rect 127716 11296 127768 11305
rect 130476 11339 130528 11348
rect 130476 11305 130485 11339
rect 130485 11305 130519 11339
rect 130519 11305 130528 11339
rect 130476 11296 130528 11305
rect 133236 11339 133288 11348
rect 133236 11305 133245 11339
rect 133245 11305 133279 11339
rect 133279 11305 133288 11339
rect 133236 11296 133288 11305
rect 136088 11339 136140 11348
rect 136088 11305 136097 11339
rect 136097 11305 136131 11339
rect 136131 11305 136140 11339
rect 136088 11296 136140 11305
rect 137192 11296 137244 11348
rect 126152 11271 126204 11280
rect 126152 11237 126161 11271
rect 126161 11237 126195 11271
rect 126195 11237 126204 11271
rect 126152 11228 126204 11237
rect 126244 11092 126296 11144
rect 131948 11228 132000 11280
rect 135628 11228 135680 11280
rect 122196 11067 122248 11076
rect 122196 11033 122205 11067
rect 122205 11033 122239 11067
rect 122239 11033 122248 11067
rect 122196 11024 122248 11033
rect 126980 11024 127032 11076
rect 127808 11024 127860 11076
rect 127900 11024 127952 11076
rect 130292 11160 130344 11212
rect 130200 11135 130252 11144
rect 130200 11101 130209 11135
rect 130209 11101 130243 11135
rect 130243 11101 130252 11135
rect 130200 11092 130252 11101
rect 135260 11203 135312 11212
rect 135260 11169 135269 11203
rect 135269 11169 135303 11203
rect 135303 11169 135312 11203
rect 135260 11160 135312 11169
rect 137468 11160 137520 11212
rect 139492 11228 139544 11280
rect 128820 11024 128872 11076
rect 134340 11092 134392 11144
rect 135168 11092 135220 11144
rect 135996 11092 136048 11144
rect 136640 11135 136692 11144
rect 136640 11101 136649 11135
rect 136649 11101 136683 11135
rect 136683 11101 136692 11135
rect 136640 11092 136692 11101
rect 138112 11092 138164 11144
rect 140872 11160 140924 11212
rect 144552 11296 144604 11348
rect 144828 11296 144880 11348
rect 141240 11228 141292 11280
rect 150440 11271 150492 11280
rect 142344 11203 142396 11212
rect 142344 11169 142353 11203
rect 142353 11169 142387 11203
rect 142387 11169 142396 11203
rect 150440 11237 150449 11271
rect 150449 11237 150483 11271
rect 150483 11237 150492 11271
rect 150440 11228 150492 11237
rect 142344 11160 142396 11169
rect 146484 11203 146536 11212
rect 146484 11169 146493 11203
rect 146493 11169 146527 11203
rect 146527 11169 146536 11203
rect 146484 11160 146536 11169
rect 147496 11203 147548 11212
rect 147496 11169 147505 11203
rect 147505 11169 147539 11203
rect 147539 11169 147548 11203
rect 147496 11160 147548 11169
rect 150992 11160 151044 11212
rect 151544 11203 151596 11212
rect 151544 11169 151553 11203
rect 151553 11169 151587 11203
rect 151587 11169 151596 11203
rect 151544 11160 151596 11169
rect 156144 11296 156196 11348
rect 160192 11339 160244 11348
rect 160192 11305 160201 11339
rect 160201 11305 160235 11339
rect 160235 11305 160244 11339
rect 160192 11296 160244 11305
rect 162216 11296 162268 11348
rect 165896 11339 165948 11348
rect 165896 11305 165905 11339
rect 165905 11305 165939 11339
rect 165939 11305 165948 11339
rect 165896 11296 165948 11305
rect 153292 11228 153344 11280
rect 163872 11203 163924 11212
rect 163872 11169 163881 11203
rect 163881 11169 163915 11203
rect 163915 11169 163924 11203
rect 163872 11160 163924 11169
rect 166080 11203 166132 11212
rect 166080 11169 166089 11203
rect 166089 11169 166123 11203
rect 166123 11169 166132 11203
rect 166080 11160 166132 11169
rect 131120 11067 131172 11076
rect 131120 11033 131129 11067
rect 131129 11033 131163 11067
rect 131163 11033 131172 11067
rect 131120 11024 131172 11033
rect 132500 11024 132552 11076
rect 133144 11024 133196 11076
rect 143356 11135 143408 11144
rect 143356 11101 143365 11135
rect 143365 11101 143399 11135
rect 143399 11101 143408 11135
rect 143356 11092 143408 11101
rect 140228 11067 140280 11076
rect 140228 11033 140237 11067
rect 140237 11033 140271 11067
rect 140271 11033 140280 11067
rect 140228 11024 140280 11033
rect 140688 11024 140740 11076
rect 144000 11092 144052 11144
rect 145012 11135 145064 11144
rect 145012 11101 145021 11135
rect 145021 11101 145055 11135
rect 145055 11101 145064 11135
rect 145012 11092 145064 11101
rect 146944 11092 146996 11144
rect 151636 11135 151688 11144
rect 151636 11101 151645 11135
rect 151645 11101 151679 11135
rect 151679 11101 151688 11135
rect 151636 11092 151688 11101
rect 150716 11024 150768 11076
rect 151452 11024 151504 11076
rect 156880 11135 156932 11144
rect 156880 11101 156889 11135
rect 156889 11101 156923 11135
rect 156923 11101 156932 11135
rect 156880 11092 156932 11101
rect 157432 11092 157484 11144
rect 151820 11024 151872 11076
rect 154120 11024 154172 11076
rect 154488 11067 154540 11076
rect 154488 11033 154497 11067
rect 154497 11033 154531 11067
rect 154531 11033 154540 11067
rect 154488 11024 154540 11033
rect 163044 11092 163096 11144
rect 167184 11135 167236 11144
rect 167184 11101 167193 11135
rect 167193 11101 167227 11135
rect 167227 11101 167236 11135
rect 167184 11092 167236 11101
rect 109040 10956 109092 10965
rect 110788 10956 110840 11008
rect 110880 10956 110932 11008
rect 111892 10956 111944 11008
rect 114560 10999 114612 11008
rect 114560 10965 114569 10999
rect 114569 10965 114603 10999
rect 114603 10965 114612 10999
rect 114560 10956 114612 10965
rect 117780 10956 117832 11008
rect 119712 10956 119764 11008
rect 120448 10956 120500 11008
rect 128268 10956 128320 11008
rect 155316 10956 155368 11008
rect 159272 10999 159324 11008
rect 159272 10965 159281 10999
rect 159281 10965 159315 10999
rect 159315 10965 159324 10999
rect 159272 10956 159324 10965
rect 56667 10854 56719 10906
rect 56731 10854 56783 10906
rect 56795 10854 56847 10906
rect 56859 10854 56911 10906
rect 113088 10854 113140 10906
rect 113152 10854 113204 10906
rect 113216 10854 113268 10906
rect 113280 10854 113332 10906
rect 6276 10795 6328 10804
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 9680 10752 9732 10804
rect 23572 10795 23624 10804
rect 23572 10761 23581 10795
rect 23581 10761 23615 10795
rect 23615 10761 23624 10795
rect 23572 10752 23624 10761
rect 24676 10752 24728 10804
rect 3700 10616 3752 10668
rect 3976 10616 4028 10668
rect 4344 10659 4396 10668
rect 4344 10625 4353 10659
rect 4353 10625 4387 10659
rect 4387 10625 4396 10659
rect 4344 10616 4396 10625
rect 4804 10616 4856 10668
rect 5080 10659 5132 10668
rect 5080 10625 5089 10659
rect 5089 10625 5123 10659
rect 5123 10625 5132 10659
rect 5080 10616 5132 10625
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 14004 10616 14056 10668
rect 19708 10659 19760 10668
rect 8300 10548 8352 10600
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 18052 10480 18104 10532
rect 18420 10480 18472 10532
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 26056 10752 26108 10804
rect 51172 10752 51224 10804
rect 51264 10752 51316 10804
rect 60464 10752 60516 10804
rect 28816 10684 28868 10736
rect 18788 10548 18840 10600
rect 21640 10659 21692 10668
rect 21640 10625 21649 10659
rect 21649 10625 21683 10659
rect 21683 10625 21692 10659
rect 21640 10616 21692 10625
rect 24768 10616 24820 10668
rect 25872 10659 25924 10668
rect 25872 10625 25881 10659
rect 25881 10625 25915 10659
rect 25915 10625 25924 10659
rect 25872 10616 25924 10625
rect 27252 10616 27304 10668
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 29092 10684 29144 10736
rect 29000 10659 29052 10668
rect 29000 10625 29009 10659
rect 29009 10625 29043 10659
rect 29043 10625 29052 10659
rect 29000 10616 29052 10625
rect 30564 10684 30616 10736
rect 31668 10684 31720 10736
rect 32772 10684 32824 10736
rect 33876 10684 33928 10736
rect 30748 10659 30800 10668
rect 30748 10625 30757 10659
rect 30757 10625 30791 10659
rect 30791 10625 30800 10659
rect 30748 10616 30800 10625
rect 31392 10616 31444 10668
rect 32220 10659 32272 10668
rect 16580 10412 16632 10464
rect 18696 10412 18748 10464
rect 24124 10412 24176 10464
rect 27804 10548 27856 10600
rect 29460 10548 29512 10600
rect 29552 10548 29604 10600
rect 32220 10625 32229 10659
rect 32229 10625 32263 10659
rect 32263 10625 32272 10659
rect 32220 10616 32272 10625
rect 32312 10616 32364 10668
rect 41972 10684 42024 10736
rect 42064 10684 42116 10736
rect 42340 10684 42392 10736
rect 42432 10684 42484 10736
rect 45836 10684 45888 10736
rect 35164 10659 35216 10668
rect 35164 10625 35173 10659
rect 35173 10625 35207 10659
rect 35207 10625 35216 10659
rect 35164 10616 35216 10625
rect 35348 10616 35400 10668
rect 37464 10659 37516 10668
rect 24308 10480 24360 10532
rect 31576 10480 31628 10532
rect 35624 10548 35676 10600
rect 36084 10591 36136 10600
rect 36084 10557 36093 10591
rect 36093 10557 36127 10591
rect 36127 10557 36136 10591
rect 36084 10548 36136 10557
rect 36360 10548 36412 10600
rect 37004 10548 37056 10600
rect 37464 10625 37473 10659
rect 37473 10625 37507 10659
rect 37507 10625 37516 10659
rect 37464 10616 37516 10625
rect 37556 10616 37608 10668
rect 41052 10616 41104 10668
rect 41604 10616 41656 10668
rect 41696 10616 41748 10668
rect 37648 10548 37700 10600
rect 38660 10480 38712 10532
rect 41696 10480 41748 10532
rect 41788 10480 41840 10532
rect 41972 10480 42024 10532
rect 26148 10412 26200 10464
rect 27436 10412 27488 10464
rect 27528 10412 27580 10464
rect 27804 10412 27856 10464
rect 27988 10412 28040 10464
rect 31484 10412 31536 10464
rect 32588 10412 32640 10464
rect 35072 10412 35124 10464
rect 35624 10412 35676 10464
rect 42064 10412 42116 10464
rect 43352 10616 43404 10668
rect 46388 10659 46440 10668
rect 43168 10548 43220 10600
rect 45836 10548 45888 10600
rect 46388 10625 46397 10659
rect 46397 10625 46431 10659
rect 46431 10625 46440 10659
rect 46388 10616 46440 10625
rect 47124 10659 47176 10668
rect 47124 10625 47133 10659
rect 47133 10625 47167 10659
rect 47167 10625 47176 10659
rect 47124 10616 47176 10625
rect 48228 10616 48280 10668
rect 49700 10616 49752 10668
rect 50620 10616 50672 10668
rect 50712 10616 50764 10668
rect 51448 10684 51500 10736
rect 55312 10684 55364 10736
rect 51724 10659 51776 10668
rect 48964 10591 49016 10600
rect 48964 10557 48973 10591
rect 48973 10557 49007 10591
rect 49007 10557 49016 10591
rect 48964 10548 49016 10557
rect 49056 10548 49108 10600
rect 51724 10625 51733 10659
rect 51733 10625 51767 10659
rect 51767 10625 51776 10659
rect 51724 10616 51776 10625
rect 51816 10616 51868 10668
rect 52368 10616 52420 10668
rect 53472 10616 53524 10668
rect 54944 10659 54996 10668
rect 54944 10625 54953 10659
rect 54953 10625 54987 10659
rect 54987 10625 54996 10659
rect 54944 10616 54996 10625
rect 55864 10684 55916 10736
rect 58072 10684 58124 10736
rect 60740 10752 60792 10804
rect 60924 10752 60976 10804
rect 61752 10752 61804 10804
rect 63776 10752 63828 10804
rect 71688 10752 71740 10804
rect 71780 10752 71832 10804
rect 73252 10752 73304 10804
rect 74356 10752 74408 10804
rect 74540 10752 74592 10804
rect 78036 10752 78088 10804
rect 82912 10752 82964 10804
rect 83924 10752 83976 10804
rect 86960 10795 87012 10804
rect 86960 10761 86969 10795
rect 86969 10761 87003 10795
rect 87003 10761 87012 10795
rect 86960 10752 87012 10761
rect 56232 10616 56284 10668
rect 56416 10616 56468 10668
rect 56968 10548 57020 10600
rect 57888 10616 57940 10668
rect 59452 10616 59504 10668
rect 70676 10684 70728 10736
rect 72516 10684 72568 10736
rect 46572 10480 46624 10532
rect 43352 10412 43404 10464
rect 45560 10412 45612 10464
rect 49792 10412 49844 10464
rect 49976 10455 50028 10464
rect 49976 10421 49985 10455
rect 49985 10421 50019 10455
rect 50019 10421 50028 10455
rect 49976 10412 50028 10421
rect 50160 10412 50212 10464
rect 51448 10412 51500 10464
rect 51632 10412 51684 10464
rect 52828 10412 52880 10464
rect 55220 10412 55272 10464
rect 55496 10412 55548 10464
rect 56048 10412 56100 10464
rect 56324 10455 56376 10464
rect 56324 10421 56333 10455
rect 56333 10421 56367 10455
rect 56367 10421 56376 10455
rect 56324 10412 56376 10421
rect 56508 10480 56560 10532
rect 57428 10480 57480 10532
rect 57980 10548 58032 10600
rect 60648 10616 60700 10668
rect 62304 10616 62356 10668
rect 65340 10616 65392 10668
rect 66260 10659 66312 10668
rect 66260 10625 66269 10659
rect 66269 10625 66303 10659
rect 66303 10625 66312 10659
rect 66260 10616 66312 10625
rect 67824 10616 67876 10668
rect 68744 10616 68796 10668
rect 69388 10659 69440 10668
rect 69388 10625 69397 10659
rect 69397 10625 69431 10659
rect 69431 10625 69440 10659
rect 69388 10616 69440 10625
rect 70492 10616 70544 10668
rect 73620 10659 73672 10668
rect 73620 10625 73629 10659
rect 73629 10625 73663 10659
rect 73663 10625 73672 10659
rect 73620 10616 73672 10625
rect 74448 10616 74500 10668
rect 60740 10548 60792 10600
rect 60924 10548 60976 10600
rect 58624 10412 58676 10464
rect 60188 10412 60240 10464
rect 60372 10480 60424 10532
rect 61936 10548 61988 10600
rect 65248 10548 65300 10600
rect 80428 10684 80480 10736
rect 75092 10616 75144 10668
rect 66168 10523 66220 10532
rect 66168 10489 66177 10523
rect 66177 10489 66211 10523
rect 66211 10489 66220 10523
rect 66168 10480 66220 10489
rect 66352 10480 66404 10532
rect 71504 10523 71556 10532
rect 71504 10489 71513 10523
rect 71513 10489 71547 10523
rect 71547 10489 71556 10523
rect 71504 10480 71556 10489
rect 72056 10480 72108 10532
rect 61660 10455 61712 10464
rect 61660 10421 61669 10455
rect 61669 10421 61703 10455
rect 61703 10421 61712 10455
rect 61660 10412 61712 10421
rect 72424 10455 72476 10464
rect 72424 10421 72433 10455
rect 72433 10421 72467 10455
rect 72467 10421 72476 10455
rect 72424 10412 72476 10421
rect 76288 10548 76340 10600
rect 77392 10591 77444 10600
rect 77392 10557 77401 10591
rect 77401 10557 77435 10591
rect 77435 10557 77444 10591
rect 77392 10548 77444 10557
rect 77760 10616 77812 10668
rect 79048 10659 79100 10668
rect 79048 10625 79057 10659
rect 79057 10625 79091 10659
rect 79091 10625 79100 10659
rect 79048 10616 79100 10625
rect 81532 10616 81584 10668
rect 80244 10548 80296 10600
rect 81164 10591 81216 10600
rect 81164 10557 81173 10591
rect 81173 10557 81207 10591
rect 81207 10557 81216 10591
rect 81164 10548 81216 10557
rect 81440 10548 81492 10600
rect 83188 10616 83240 10668
rect 83556 10659 83608 10668
rect 83556 10625 83565 10659
rect 83565 10625 83599 10659
rect 83599 10625 83608 10659
rect 83556 10616 83608 10625
rect 85764 10659 85816 10668
rect 85764 10625 85773 10659
rect 85773 10625 85807 10659
rect 85807 10625 85816 10659
rect 90364 10752 90416 10804
rect 91744 10752 91796 10804
rect 95516 10752 95568 10804
rect 106188 10752 106240 10804
rect 111064 10752 111116 10804
rect 120264 10752 120316 10804
rect 120724 10752 120776 10804
rect 123760 10752 123812 10804
rect 124772 10795 124824 10804
rect 124772 10761 124781 10795
rect 124781 10761 124815 10795
rect 124815 10761 124824 10795
rect 124772 10752 124824 10761
rect 127164 10752 127216 10804
rect 128268 10752 128320 10804
rect 131948 10795 132000 10804
rect 85764 10616 85816 10625
rect 88340 10659 88392 10668
rect 88340 10625 88349 10659
rect 88349 10625 88383 10659
rect 88383 10625 88392 10659
rect 88340 10616 88392 10625
rect 90916 10616 90968 10668
rect 82728 10548 82780 10600
rect 84660 10591 84712 10600
rect 84660 10557 84669 10591
rect 84669 10557 84703 10591
rect 84703 10557 84712 10591
rect 84660 10548 84712 10557
rect 85672 10591 85724 10600
rect 85672 10557 85681 10591
rect 85681 10557 85715 10591
rect 85715 10557 85724 10591
rect 85672 10548 85724 10557
rect 88064 10591 88116 10600
rect 88064 10557 88073 10591
rect 88073 10557 88107 10591
rect 88107 10557 88116 10591
rect 88064 10548 88116 10557
rect 93124 10548 93176 10600
rect 73896 10480 73948 10532
rect 74080 10412 74132 10464
rect 78220 10480 78272 10532
rect 96068 10616 96120 10668
rect 98920 10659 98972 10668
rect 95884 10591 95936 10600
rect 95884 10557 95893 10591
rect 95893 10557 95927 10591
rect 95927 10557 95936 10591
rect 95884 10548 95936 10557
rect 98368 10548 98420 10600
rect 98920 10625 98929 10659
rect 98929 10625 98963 10659
rect 98963 10625 98972 10659
rect 98920 10616 98972 10625
rect 101772 10616 101824 10668
rect 104256 10616 104308 10668
rect 106188 10659 106240 10668
rect 106188 10625 106197 10659
rect 106197 10625 106231 10659
rect 106231 10625 106240 10659
rect 106188 10616 106240 10625
rect 99564 10548 99616 10600
rect 102232 10591 102284 10600
rect 102232 10557 102241 10591
rect 102241 10557 102275 10591
rect 102275 10557 102284 10591
rect 102232 10548 102284 10557
rect 103244 10591 103296 10600
rect 103244 10557 103253 10591
rect 103253 10557 103287 10591
rect 103287 10557 103296 10591
rect 103244 10548 103296 10557
rect 104624 10591 104676 10600
rect 104624 10557 104633 10591
rect 104633 10557 104667 10591
rect 104667 10557 104676 10591
rect 104624 10548 104676 10557
rect 110880 10684 110932 10736
rect 107844 10616 107896 10668
rect 108948 10616 109000 10668
rect 111340 10659 111392 10668
rect 111340 10625 111349 10659
rect 111349 10625 111383 10659
rect 111383 10625 111392 10659
rect 111340 10616 111392 10625
rect 107660 10591 107712 10600
rect 107660 10557 107669 10591
rect 107669 10557 107703 10591
rect 107703 10557 107712 10591
rect 107660 10548 107712 10557
rect 110052 10591 110104 10600
rect 110052 10557 110061 10591
rect 110061 10557 110095 10591
rect 110095 10557 110104 10591
rect 110052 10548 110104 10557
rect 112628 10616 112680 10668
rect 105636 10480 105688 10532
rect 108856 10480 108908 10532
rect 112904 10548 112956 10600
rect 113456 10548 113508 10600
rect 110972 10480 111024 10532
rect 111340 10480 111392 10532
rect 117136 10616 117188 10668
rect 119620 10684 119672 10736
rect 119712 10684 119764 10736
rect 121092 10659 121144 10668
rect 121092 10625 121101 10659
rect 121101 10625 121135 10659
rect 121135 10625 121144 10659
rect 121092 10616 121144 10625
rect 123116 10616 123168 10668
rect 114836 10548 114888 10600
rect 115848 10548 115900 10600
rect 116676 10591 116728 10600
rect 116676 10557 116685 10591
rect 116685 10557 116719 10591
rect 116719 10557 116728 10591
rect 116676 10548 116728 10557
rect 119528 10591 119580 10600
rect 119528 10557 119537 10591
rect 119537 10557 119571 10591
rect 119571 10557 119580 10591
rect 119528 10548 119580 10557
rect 120540 10591 120592 10600
rect 120540 10557 120549 10591
rect 120549 10557 120583 10591
rect 120583 10557 120592 10591
rect 120540 10548 120592 10557
rect 114652 10480 114704 10532
rect 123392 10548 123444 10600
rect 124956 10616 125008 10668
rect 127072 10616 127124 10668
rect 127624 10616 127676 10668
rect 128360 10616 128412 10668
rect 129188 10616 129240 10668
rect 125600 10548 125652 10600
rect 126244 10548 126296 10600
rect 129556 10591 129608 10600
rect 129556 10557 129565 10591
rect 129565 10557 129599 10591
rect 129599 10557 129608 10591
rect 129556 10548 129608 10557
rect 130660 10659 130712 10668
rect 130660 10625 130669 10659
rect 130669 10625 130703 10659
rect 130703 10625 130712 10659
rect 130660 10616 130712 10625
rect 131948 10761 131957 10795
rect 131957 10761 131991 10795
rect 131991 10761 132000 10795
rect 131948 10752 132000 10761
rect 148324 10752 148376 10804
rect 131580 10684 131632 10736
rect 135076 10684 135128 10736
rect 134064 10659 134116 10668
rect 134064 10625 134073 10659
rect 134073 10625 134107 10659
rect 134107 10625 134116 10659
rect 134064 10616 134116 10625
rect 139124 10684 139176 10736
rect 132960 10591 133012 10600
rect 132960 10557 132969 10591
rect 132969 10557 133003 10591
rect 133003 10557 133012 10591
rect 132960 10548 133012 10557
rect 137468 10616 137520 10668
rect 139032 10659 139084 10668
rect 139032 10625 139041 10659
rect 139041 10625 139075 10659
rect 139075 10625 139084 10659
rect 139032 10616 139084 10625
rect 145012 10684 145064 10736
rect 146852 10684 146904 10736
rect 142160 10659 142212 10668
rect 136272 10548 136324 10600
rect 142160 10625 142169 10659
rect 142169 10625 142203 10659
rect 142203 10625 142212 10659
rect 142160 10616 142212 10625
rect 144920 10659 144972 10668
rect 144920 10625 144929 10659
rect 144929 10625 144963 10659
rect 144963 10625 144972 10659
rect 144920 10616 144972 10625
rect 147864 10659 147916 10668
rect 147864 10625 147873 10659
rect 147873 10625 147907 10659
rect 147907 10625 147916 10659
rect 147864 10616 147916 10625
rect 151636 10616 151688 10668
rect 153200 10659 153252 10668
rect 153200 10625 153209 10659
rect 153209 10625 153243 10659
rect 153243 10625 153252 10659
rect 153200 10616 153252 10625
rect 155960 10659 156012 10668
rect 155960 10625 155969 10659
rect 155969 10625 156003 10659
rect 156003 10625 156012 10659
rect 155960 10616 156012 10625
rect 158720 10616 158772 10668
rect 159272 10616 159324 10668
rect 141056 10548 141108 10600
rect 144184 10548 144236 10600
rect 146944 10548 146996 10600
rect 148784 10548 148836 10600
rect 152096 10548 152148 10600
rect 155316 10548 155368 10600
rect 156144 10591 156196 10600
rect 156144 10557 156153 10591
rect 156153 10557 156187 10591
rect 156187 10557 156196 10591
rect 156144 10548 156196 10557
rect 157248 10548 157300 10600
rect 159548 10659 159600 10668
rect 159548 10625 159557 10659
rect 159557 10625 159591 10659
rect 159591 10625 159600 10659
rect 159548 10616 159600 10625
rect 162860 10659 162912 10668
rect 162860 10625 162869 10659
rect 162869 10625 162903 10659
rect 162903 10625 162912 10659
rect 162860 10616 162912 10625
rect 164332 10659 164384 10668
rect 164332 10625 164341 10659
rect 164341 10625 164375 10659
rect 164375 10625 164384 10659
rect 164332 10616 164384 10625
rect 142252 10523 142304 10532
rect 109684 10412 109736 10464
rect 111156 10412 111208 10464
rect 111708 10412 111760 10464
rect 112904 10455 112956 10464
rect 112904 10421 112913 10455
rect 112913 10421 112947 10455
rect 112947 10421 112956 10455
rect 112904 10412 112956 10421
rect 112996 10412 113048 10464
rect 142252 10489 142261 10523
rect 142261 10489 142295 10523
rect 142295 10489 142304 10523
rect 142252 10480 142304 10489
rect 145104 10523 145156 10532
rect 145104 10489 145113 10523
rect 145113 10489 145147 10523
rect 145147 10489 145156 10523
rect 145104 10480 145156 10489
rect 149796 10480 149848 10532
rect 152372 10480 152424 10532
rect 153292 10523 153344 10532
rect 153292 10489 153301 10523
rect 153301 10489 153335 10523
rect 153335 10489 153344 10523
rect 153292 10480 153344 10489
rect 162676 10548 162728 10600
rect 165620 10591 165672 10600
rect 165620 10557 165629 10591
rect 165629 10557 165663 10591
rect 165663 10557 165672 10591
rect 165620 10548 165672 10557
rect 166724 10659 166776 10668
rect 166724 10625 166733 10659
rect 166733 10625 166767 10659
rect 166767 10625 166776 10659
rect 166724 10616 166776 10625
rect 121184 10412 121236 10464
rect 122748 10412 122800 10464
rect 122932 10455 122984 10464
rect 122932 10421 122941 10455
rect 122941 10421 122975 10455
rect 122975 10421 122984 10455
rect 122932 10412 122984 10421
rect 123760 10412 123812 10464
rect 127440 10412 127492 10464
rect 127624 10455 127676 10464
rect 127624 10421 127633 10455
rect 127633 10421 127667 10455
rect 127667 10421 127676 10455
rect 127624 10412 127676 10421
rect 128084 10412 128136 10464
rect 132408 10455 132460 10464
rect 132408 10421 132417 10455
rect 132417 10421 132451 10455
rect 132451 10421 132460 10455
rect 132408 10412 132460 10421
rect 133512 10412 133564 10464
rect 138020 10455 138072 10464
rect 138020 10421 138029 10455
rect 138029 10421 138063 10455
rect 138063 10421 138072 10455
rect 140412 10455 140464 10464
rect 138020 10412 138072 10421
rect 140412 10421 140421 10455
rect 140421 10421 140455 10455
rect 140455 10421 140464 10455
rect 140412 10412 140464 10421
rect 147588 10412 147640 10464
rect 157248 10412 157300 10464
rect 157984 10455 158036 10464
rect 157984 10421 157993 10455
rect 157993 10421 158027 10455
rect 158027 10421 158036 10455
rect 157984 10412 158036 10421
rect 160468 10455 160520 10464
rect 160468 10421 160477 10455
rect 160477 10421 160511 10455
rect 160511 10421 160520 10455
rect 160468 10412 160520 10421
rect 28456 10310 28508 10362
rect 28520 10310 28572 10362
rect 28584 10310 28636 10362
rect 28648 10310 28700 10362
rect 84878 10310 84930 10362
rect 84942 10310 84994 10362
rect 85006 10310 85058 10362
rect 85070 10310 85122 10362
rect 141299 10310 141351 10362
rect 141363 10310 141415 10362
rect 141427 10310 141479 10362
rect 141491 10310 141543 10362
rect 4344 10208 4396 10260
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 9312 10208 9364 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 14004 10251 14056 10260
rect 14004 10217 14013 10251
rect 14013 10217 14047 10251
rect 14047 10217 14056 10251
rect 14004 10208 14056 10217
rect 17316 10251 17368 10260
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 19708 10251 19760 10260
rect 19708 10217 19717 10251
rect 19717 10217 19751 10251
rect 19751 10217 19760 10251
rect 19708 10208 19760 10217
rect 29092 10208 29144 10260
rect 30748 10208 30800 10260
rect 33876 10208 33928 10260
rect 35164 10208 35216 10260
rect 2872 10140 2924 10192
rect 9680 10140 9732 10192
rect 19524 10140 19576 10192
rect 4160 10115 4212 10124
rect 4160 10081 4169 10115
rect 4169 10081 4203 10115
rect 4203 10081 4212 10115
rect 4160 10072 4212 10081
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 4068 10004 4120 10056
rect 4712 10004 4764 10056
rect 7012 10072 7064 10124
rect 3608 9868 3660 9920
rect 4436 9868 4488 9920
rect 5080 9911 5132 9920
rect 5080 9877 5089 9911
rect 5089 9877 5123 9911
rect 5123 9877 5132 9911
rect 5080 9868 5132 9877
rect 20076 10072 20128 10124
rect 20168 10115 20220 10124
rect 20168 10081 20177 10115
rect 20177 10081 20211 10115
rect 20211 10081 20220 10115
rect 20168 10072 20220 10081
rect 20720 10072 20772 10124
rect 24032 10140 24084 10192
rect 25136 10140 25188 10192
rect 25872 10140 25924 10192
rect 24768 10115 24820 10124
rect 17316 10004 17368 10056
rect 23388 10004 23440 10056
rect 23572 10047 23624 10056
rect 23572 10013 23581 10047
rect 23581 10013 23615 10047
rect 23615 10013 23624 10047
rect 23572 10004 23624 10013
rect 23940 10004 23992 10056
rect 24768 10081 24777 10115
rect 24777 10081 24811 10115
rect 24811 10081 24820 10115
rect 24768 10072 24820 10081
rect 26976 10140 27028 10192
rect 27896 10140 27948 10192
rect 29000 10140 29052 10192
rect 34336 10140 34388 10192
rect 34520 10140 34572 10192
rect 35440 10140 35492 10192
rect 36820 10208 36872 10260
rect 41604 10208 41656 10260
rect 41880 10208 41932 10260
rect 42064 10208 42116 10260
rect 42432 10208 42484 10260
rect 42800 10208 42852 10260
rect 46572 10208 46624 10260
rect 48228 10208 48280 10260
rect 48596 10208 48648 10260
rect 50804 10208 50856 10260
rect 50988 10208 51040 10260
rect 51540 10208 51592 10260
rect 51724 10208 51776 10260
rect 52368 10208 52420 10260
rect 54944 10208 54996 10260
rect 55404 10251 55456 10260
rect 55404 10217 55413 10251
rect 55413 10217 55447 10251
rect 55447 10217 55456 10251
rect 55404 10208 55456 10217
rect 55496 10208 55548 10260
rect 60740 10208 60792 10260
rect 60924 10208 60976 10260
rect 64236 10208 64288 10260
rect 65248 10251 65300 10260
rect 65248 10217 65257 10251
rect 65257 10217 65291 10251
rect 65291 10217 65300 10251
rect 65248 10208 65300 10217
rect 68744 10251 68796 10260
rect 68744 10217 68753 10251
rect 68753 10217 68787 10251
rect 68787 10217 68796 10251
rect 68744 10208 68796 10217
rect 69388 10251 69440 10260
rect 69388 10217 69397 10251
rect 69397 10217 69431 10251
rect 69431 10217 69440 10251
rect 69388 10208 69440 10217
rect 70492 10208 70544 10260
rect 70860 10208 70912 10260
rect 74448 10208 74500 10260
rect 75092 10208 75144 10260
rect 76380 10251 76432 10260
rect 76380 10217 76389 10251
rect 76389 10217 76423 10251
rect 76423 10217 76432 10251
rect 76380 10208 76432 10217
rect 76564 10208 76616 10260
rect 78220 10251 78272 10260
rect 78220 10217 78229 10251
rect 78229 10217 78263 10251
rect 78263 10217 78272 10251
rect 78220 10208 78272 10217
rect 78312 10208 78364 10260
rect 79048 10251 79100 10260
rect 79048 10217 79057 10251
rect 79057 10217 79091 10251
rect 79091 10217 79100 10251
rect 79048 10208 79100 10217
rect 80244 10251 80296 10260
rect 80244 10217 80253 10251
rect 80253 10217 80287 10251
rect 80287 10217 80296 10251
rect 80244 10208 80296 10217
rect 80428 10251 80480 10260
rect 80428 10217 80437 10251
rect 80437 10217 80471 10251
rect 80471 10217 80480 10251
rect 80428 10208 80480 10217
rect 81532 10251 81584 10260
rect 81532 10217 81541 10251
rect 81541 10217 81575 10251
rect 81575 10217 81584 10251
rect 81532 10208 81584 10217
rect 82728 10251 82780 10260
rect 82728 10217 82737 10251
rect 82737 10217 82771 10251
rect 82771 10217 82780 10251
rect 82728 10208 82780 10217
rect 83556 10251 83608 10260
rect 83556 10217 83565 10251
rect 83565 10217 83599 10251
rect 83599 10217 83608 10251
rect 83556 10208 83608 10217
rect 84660 10251 84712 10260
rect 84660 10217 84669 10251
rect 84669 10217 84703 10251
rect 84703 10217 84712 10251
rect 84660 10208 84712 10217
rect 27620 10072 27672 10124
rect 29368 10072 29420 10124
rect 41972 10140 42024 10192
rect 44548 10140 44600 10192
rect 37096 10072 37148 10124
rect 37464 10115 37516 10124
rect 37464 10081 37473 10115
rect 37473 10081 37507 10115
rect 37507 10081 37516 10115
rect 37464 10072 37516 10081
rect 37648 10115 37700 10124
rect 37648 10081 37657 10115
rect 37657 10081 37691 10115
rect 37691 10081 37700 10115
rect 37648 10072 37700 10081
rect 37740 10072 37792 10124
rect 38844 10072 38896 10124
rect 27160 10004 27212 10056
rect 27804 10047 27856 10056
rect 27804 10013 27813 10047
rect 27813 10013 27847 10047
rect 27847 10013 27856 10047
rect 27804 10004 27856 10013
rect 27896 10047 27948 10056
rect 27896 10013 27905 10047
rect 27905 10013 27939 10047
rect 27939 10013 27948 10047
rect 27896 10004 27948 10013
rect 32404 10004 32456 10056
rect 32588 10047 32640 10056
rect 32588 10013 32597 10047
rect 32597 10013 32631 10047
rect 32631 10013 32640 10047
rect 32588 10004 32640 10013
rect 32680 10047 32732 10056
rect 32680 10013 32689 10047
rect 32689 10013 32723 10047
rect 32723 10013 32732 10047
rect 32680 10004 32732 10013
rect 33416 10004 33468 10056
rect 35072 10047 35124 10056
rect 35072 10013 35081 10047
rect 35081 10013 35115 10047
rect 35115 10013 35124 10047
rect 35072 10004 35124 10013
rect 24216 9936 24268 9988
rect 27528 9936 27580 9988
rect 27712 9936 27764 9988
rect 30748 9936 30800 9988
rect 7104 9868 7156 9920
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 17316 9868 17368 9920
rect 24032 9868 24084 9920
rect 24124 9868 24176 9920
rect 27988 9868 28040 9920
rect 28080 9868 28132 9920
rect 29000 9868 29052 9920
rect 29644 9868 29696 9920
rect 30288 9911 30340 9920
rect 30288 9877 30297 9911
rect 30297 9877 30331 9911
rect 30331 9877 30340 9911
rect 30288 9868 30340 9877
rect 32220 9868 32272 9920
rect 33416 9911 33468 9920
rect 33416 9877 33425 9911
rect 33425 9877 33459 9911
rect 33459 9877 33468 9911
rect 33416 9868 33468 9877
rect 33876 9936 33928 9988
rect 39120 10004 39172 10056
rect 45100 10072 45152 10124
rect 48964 10140 49016 10192
rect 49700 10183 49752 10192
rect 49700 10149 49709 10183
rect 49709 10149 49743 10183
rect 49743 10149 49752 10183
rect 49700 10140 49752 10149
rect 49884 10183 49936 10192
rect 49884 10149 49893 10183
rect 49893 10149 49927 10183
rect 49927 10149 49936 10183
rect 49884 10140 49936 10149
rect 45284 10072 45336 10124
rect 51264 10140 51316 10192
rect 79416 10183 79468 10192
rect 55496 10072 55548 10124
rect 56140 10115 56192 10124
rect 56140 10081 56149 10115
rect 56149 10081 56183 10115
rect 56183 10081 56192 10115
rect 56140 10072 56192 10081
rect 56508 10072 56560 10124
rect 45836 10047 45888 10056
rect 45836 10013 45845 10047
rect 45845 10013 45879 10047
rect 45879 10013 45888 10047
rect 45836 10004 45888 10013
rect 48228 10004 48280 10056
rect 48412 10047 48464 10056
rect 48412 10013 48421 10047
rect 48421 10013 48455 10047
rect 48455 10013 48464 10047
rect 48412 10004 48464 10013
rect 49976 10047 50028 10056
rect 49976 10013 49985 10047
rect 49985 10013 50019 10047
rect 50019 10013 50028 10047
rect 49976 10004 50028 10013
rect 50896 10004 50948 10056
rect 51632 10047 51684 10056
rect 51632 10013 51641 10047
rect 51641 10013 51675 10047
rect 51675 10013 51684 10047
rect 51632 10004 51684 10013
rect 35348 9868 35400 9920
rect 36084 9868 36136 9920
rect 37004 9868 37056 9920
rect 37096 9868 37148 9920
rect 39212 9868 39264 9920
rect 40040 9868 40092 9920
rect 40408 9868 40460 9920
rect 47124 9936 47176 9988
rect 50252 9936 50304 9988
rect 50344 9936 50396 9988
rect 42616 9911 42668 9920
rect 42616 9877 42625 9911
rect 42625 9877 42659 9911
rect 42659 9877 42668 9911
rect 42616 9868 42668 9877
rect 43168 9911 43220 9920
rect 43168 9877 43177 9911
rect 43177 9877 43211 9911
rect 43211 9877 43220 9911
rect 43168 9868 43220 9877
rect 44088 9868 44140 9920
rect 50620 9868 50672 9920
rect 50712 9868 50764 9920
rect 53380 10004 53432 10056
rect 55864 10004 55916 10056
rect 53472 9936 53524 9988
rect 54484 9936 54536 9988
rect 54576 9936 54628 9988
rect 55128 9868 55180 9920
rect 55864 9868 55916 9920
rect 56784 10004 56836 10056
rect 57704 10115 57756 10124
rect 57704 10081 57713 10115
rect 57713 10081 57747 10115
rect 57747 10081 57756 10115
rect 57704 10072 57756 10081
rect 57888 10072 57940 10124
rect 56600 9936 56652 9988
rect 57060 9936 57112 9988
rect 57428 9936 57480 9988
rect 57796 10004 57848 10056
rect 58624 10004 58676 10056
rect 59452 10072 59504 10124
rect 60740 10072 60792 10124
rect 68928 10115 68980 10124
rect 68928 10081 68937 10115
rect 68937 10081 68971 10115
rect 68971 10081 68980 10115
rect 68928 10072 68980 10081
rect 72056 10115 72108 10124
rect 72056 10081 72065 10115
rect 72065 10081 72099 10115
rect 72099 10081 72108 10115
rect 72056 10072 72108 10081
rect 72240 10072 72292 10124
rect 59820 10047 59872 10056
rect 59820 10013 59829 10047
rect 59829 10013 59863 10047
rect 59863 10013 59872 10047
rect 59820 10004 59872 10013
rect 60464 10047 60516 10056
rect 60464 10013 60473 10047
rect 60473 10013 60507 10047
rect 60507 10013 60516 10047
rect 60464 10004 60516 10013
rect 60556 10004 60608 10056
rect 62028 10047 62080 10056
rect 62028 10013 62037 10047
rect 62037 10013 62071 10047
rect 62071 10013 62080 10047
rect 62028 10004 62080 10013
rect 62764 10004 62816 10056
rect 70860 10047 70912 10056
rect 70860 10013 70869 10047
rect 70869 10013 70903 10047
rect 70903 10013 70912 10047
rect 70860 10004 70912 10013
rect 71412 10047 71464 10056
rect 71412 10013 71421 10047
rect 71421 10013 71455 10047
rect 71455 10013 71464 10047
rect 71412 10004 71464 10013
rect 72424 10047 72476 10056
rect 72424 10013 72433 10047
rect 72433 10013 72467 10047
rect 72467 10013 72476 10047
rect 72424 10004 72476 10013
rect 72608 10047 72660 10056
rect 72608 10013 72617 10047
rect 72617 10013 72651 10047
rect 72651 10013 72660 10047
rect 72608 10004 72660 10013
rect 73896 10004 73948 10056
rect 74080 10047 74132 10056
rect 74080 10013 74089 10047
rect 74089 10013 74123 10047
rect 74123 10013 74132 10047
rect 74080 10004 74132 10013
rect 74356 10047 74408 10056
rect 60280 9936 60332 9988
rect 74356 10013 74365 10047
rect 74365 10013 74399 10047
rect 74399 10013 74408 10047
rect 74356 10004 74408 10013
rect 76564 10004 76616 10056
rect 77300 10047 77352 10056
rect 77300 10013 77309 10047
rect 77309 10013 77343 10047
rect 77343 10013 77352 10047
rect 77300 10004 77352 10013
rect 77392 9979 77444 9988
rect 77392 9945 77401 9979
rect 77401 9945 77435 9979
rect 77435 9945 77444 9979
rect 77392 9936 77444 9945
rect 79416 10149 79425 10183
rect 79425 10149 79459 10183
rect 79459 10149 79468 10183
rect 79416 10140 79468 10149
rect 78036 10004 78088 10056
rect 78404 10004 78456 10056
rect 85212 10140 85264 10192
rect 85120 10072 85172 10124
rect 85948 10072 86000 10124
rect 87236 10072 87288 10124
rect 93492 10208 93544 10260
rect 95884 10251 95936 10260
rect 95884 10217 95893 10251
rect 95893 10217 95927 10251
rect 95927 10217 95936 10251
rect 95884 10208 95936 10217
rect 92388 10140 92440 10192
rect 79508 10004 79560 10056
rect 81072 10004 81124 10056
rect 82912 10047 82964 10056
rect 82912 10013 82921 10047
rect 82921 10013 82955 10047
rect 82955 10013 82964 10047
rect 82912 10004 82964 10013
rect 90364 10072 90416 10124
rect 92756 10072 92808 10124
rect 97540 10183 97592 10192
rect 97540 10149 97549 10183
rect 97549 10149 97583 10183
rect 97583 10149 97592 10183
rect 97540 10140 97592 10149
rect 91928 10047 91980 10056
rect 60924 9868 60976 9920
rect 61292 9868 61344 9920
rect 66260 9911 66312 9920
rect 66260 9877 66269 9911
rect 66269 9877 66303 9911
rect 66303 9877 66312 9911
rect 66260 9868 66312 9877
rect 73620 9911 73672 9920
rect 73620 9877 73629 9911
rect 73629 9877 73663 9911
rect 73663 9877 73672 9911
rect 73620 9868 73672 9877
rect 76288 9868 76340 9920
rect 78496 9868 78548 9920
rect 86960 9911 87012 9920
rect 86960 9877 86969 9911
rect 86969 9877 87003 9911
rect 87003 9877 87012 9911
rect 86960 9868 87012 9877
rect 87236 9911 87288 9920
rect 87236 9877 87245 9911
rect 87245 9877 87279 9911
rect 87279 9877 87288 9911
rect 91928 10013 91937 10047
rect 91937 10013 91971 10047
rect 91971 10013 91980 10047
rect 91928 10004 91980 10013
rect 92664 10004 92716 10056
rect 93308 10004 93360 10056
rect 94228 10047 94280 10056
rect 94228 10013 94237 10047
rect 94237 10013 94271 10047
rect 94271 10013 94280 10047
rect 94228 10004 94280 10013
rect 98276 10208 98328 10260
rect 98368 10251 98420 10260
rect 98368 10217 98377 10251
rect 98377 10217 98411 10251
rect 98411 10217 98420 10251
rect 98368 10208 98420 10217
rect 99564 10251 99616 10260
rect 99564 10217 99573 10251
rect 99573 10217 99607 10251
rect 99607 10217 99616 10251
rect 107660 10251 107712 10260
rect 99564 10208 99616 10217
rect 98920 10115 98972 10124
rect 98920 10081 98929 10115
rect 98929 10081 98963 10115
rect 98963 10081 98972 10115
rect 98920 10072 98972 10081
rect 107660 10217 107669 10251
rect 107669 10217 107703 10251
rect 107703 10217 107712 10251
rect 107660 10208 107712 10217
rect 108948 10251 109000 10260
rect 108948 10217 108957 10251
rect 108957 10217 108991 10251
rect 108991 10217 109000 10251
rect 108948 10208 109000 10217
rect 109684 10208 109736 10260
rect 110972 10208 111024 10260
rect 111340 10208 111392 10260
rect 116952 10208 117004 10260
rect 117136 10251 117188 10260
rect 117136 10217 117145 10251
rect 117145 10217 117179 10251
rect 117179 10217 117188 10251
rect 117136 10208 117188 10217
rect 119528 10251 119580 10260
rect 119528 10217 119537 10251
rect 119537 10217 119571 10251
rect 119571 10217 119580 10251
rect 119528 10208 119580 10217
rect 119620 10208 119672 10260
rect 122104 10208 122156 10260
rect 123116 10251 123168 10260
rect 123116 10217 123125 10251
rect 123125 10217 123159 10251
rect 123159 10217 123168 10251
rect 123116 10208 123168 10217
rect 124956 10251 125008 10260
rect 124956 10217 124965 10251
rect 124965 10217 124999 10251
rect 124999 10217 125008 10251
rect 124956 10208 125008 10217
rect 126612 10208 126664 10260
rect 127348 10251 127400 10260
rect 127348 10217 127357 10251
rect 127357 10217 127391 10251
rect 127391 10217 127400 10251
rect 127348 10208 127400 10217
rect 127440 10208 127492 10260
rect 106740 10140 106792 10192
rect 100852 10115 100904 10124
rect 100852 10081 100861 10115
rect 100861 10081 100895 10115
rect 100895 10081 100904 10115
rect 100852 10072 100904 10081
rect 102232 10115 102284 10124
rect 102232 10081 102241 10115
rect 102241 10081 102275 10115
rect 102275 10081 102284 10115
rect 102232 10072 102284 10081
rect 107660 10072 107712 10124
rect 110052 10072 110104 10124
rect 111248 10072 111300 10124
rect 101588 10047 101640 10056
rect 101588 10013 101597 10047
rect 101597 10013 101631 10047
rect 101631 10013 101640 10047
rect 101588 10004 101640 10013
rect 101772 10004 101824 10056
rect 112536 10072 112588 10124
rect 115572 10115 115624 10124
rect 112260 10004 112312 10056
rect 112904 10047 112956 10056
rect 112904 10013 112913 10047
rect 112913 10013 112947 10047
rect 112947 10013 112956 10047
rect 112904 10004 112956 10013
rect 109040 9936 109092 9988
rect 110052 9936 110104 9988
rect 114652 10004 114704 10056
rect 115572 10081 115581 10115
rect 115581 10081 115615 10115
rect 115615 10081 115624 10115
rect 115572 10072 115624 10081
rect 115940 10004 115992 10056
rect 127532 10140 127584 10192
rect 128360 10208 128412 10260
rect 129556 10208 129608 10260
rect 132960 10208 133012 10260
rect 134064 10208 134116 10260
rect 135076 10208 135128 10260
rect 137468 10251 137520 10260
rect 137468 10217 137477 10251
rect 137477 10217 137511 10251
rect 137511 10217 137520 10251
rect 137468 10208 137520 10217
rect 116584 10115 116636 10124
rect 116584 10081 116593 10115
rect 116593 10081 116627 10115
rect 116627 10081 116636 10115
rect 116584 10072 116636 10081
rect 117964 10072 118016 10124
rect 121184 10047 121236 10056
rect 121184 10013 121193 10047
rect 121193 10013 121227 10047
rect 121227 10013 121236 10047
rect 121184 10004 121236 10013
rect 122104 10004 122156 10056
rect 129004 10115 129056 10124
rect 129004 10081 129013 10115
rect 129013 10081 129047 10115
rect 129047 10081 129056 10115
rect 129004 10072 129056 10081
rect 129740 10072 129792 10124
rect 130660 10072 130712 10124
rect 132408 10115 132460 10124
rect 132408 10081 132417 10115
rect 132417 10081 132451 10115
rect 132451 10081 132460 10115
rect 132408 10072 132460 10081
rect 133420 10115 133472 10124
rect 133420 10081 133429 10115
rect 133429 10081 133463 10115
rect 133463 10081 133472 10115
rect 133420 10072 133472 10081
rect 136272 10115 136324 10124
rect 136272 10081 136281 10115
rect 136281 10081 136315 10115
rect 136315 10081 136324 10115
rect 147220 10140 147272 10192
rect 136272 10072 136324 10081
rect 140780 10072 140832 10124
rect 142160 10072 142212 10124
rect 122748 10047 122800 10056
rect 122748 10013 122757 10047
rect 122757 10013 122791 10047
rect 122791 10013 122800 10047
rect 122748 10004 122800 10013
rect 127348 10004 127400 10056
rect 128084 10004 128136 10056
rect 87236 9868 87288 9877
rect 93124 9868 93176 9920
rect 93400 9868 93452 9920
rect 98368 9868 98420 9920
rect 102140 9868 102192 9920
rect 103336 9868 103388 9920
rect 104256 9868 104308 9920
rect 104624 9911 104676 9920
rect 104624 9877 104633 9911
rect 104633 9877 104667 9911
rect 104667 9877 104676 9911
rect 104624 9868 104676 9877
rect 106188 9868 106240 9920
rect 114560 9868 114612 9920
rect 115848 9868 115900 9920
rect 120908 9936 120960 9988
rect 129924 10004 129976 10056
rect 133512 10047 133564 10056
rect 133512 10013 133521 10047
rect 133521 10013 133555 10047
rect 133555 10013 133564 10047
rect 133512 10004 133564 10013
rect 134800 10047 134852 10056
rect 134800 10013 134809 10047
rect 134809 10013 134843 10047
rect 134843 10013 134852 10047
rect 134800 10004 134852 10013
rect 138020 10047 138072 10056
rect 138020 10013 138029 10047
rect 138029 10013 138063 10047
rect 138063 10013 138072 10047
rect 139124 10047 139176 10056
rect 138020 10004 138072 10013
rect 139124 10013 139133 10047
rect 139133 10013 139167 10047
rect 139167 10013 139176 10047
rect 139124 10004 139176 10013
rect 140412 10047 140464 10056
rect 140412 10013 140421 10047
rect 140421 10013 140455 10047
rect 140455 10013 140464 10047
rect 140412 10004 140464 10013
rect 140872 10004 140924 10056
rect 152096 10251 152148 10260
rect 152096 10217 152105 10251
rect 152105 10217 152139 10251
rect 152139 10217 152148 10251
rect 152096 10208 152148 10217
rect 153200 10208 153252 10260
rect 155316 10251 155368 10260
rect 155316 10217 155325 10251
rect 155325 10217 155359 10251
rect 155359 10217 155368 10251
rect 155316 10208 155368 10217
rect 155960 10208 156012 10260
rect 158720 10208 158772 10260
rect 159548 10208 159600 10260
rect 162676 10251 162728 10260
rect 162676 10217 162685 10251
rect 162685 10217 162719 10251
rect 162719 10217 162728 10251
rect 162676 10208 162728 10217
rect 164332 10208 164384 10260
rect 165620 10251 165672 10260
rect 165620 10217 165629 10251
rect 165629 10217 165663 10251
rect 165663 10217 165672 10251
rect 165620 10208 165672 10217
rect 166724 10208 166776 10260
rect 151268 10140 151320 10192
rect 162308 10140 162360 10192
rect 157984 10115 158036 10124
rect 157984 10081 157993 10115
rect 157993 10081 158027 10115
rect 158027 10081 158036 10115
rect 157984 10072 158036 10081
rect 159364 10115 159416 10124
rect 159364 10081 159373 10115
rect 159373 10081 159407 10115
rect 159407 10081 159416 10115
rect 159364 10072 159416 10081
rect 160468 10115 160520 10124
rect 160468 10081 160477 10115
rect 160477 10081 160511 10115
rect 160511 10081 160520 10115
rect 160468 10072 160520 10081
rect 160560 10072 160612 10124
rect 162860 10115 162912 10124
rect 162860 10081 162869 10115
rect 162869 10081 162903 10115
rect 162903 10081 162912 10115
rect 162860 10072 162912 10081
rect 159548 10047 159600 10056
rect 120724 9868 120776 9920
rect 121092 9868 121144 9920
rect 126244 9911 126296 9920
rect 126244 9877 126253 9911
rect 126253 9877 126287 9911
rect 126287 9877 126296 9911
rect 126244 9868 126296 9877
rect 137836 9936 137888 9988
rect 139032 9936 139084 9988
rect 141056 9936 141108 9988
rect 130200 9868 130252 9920
rect 144184 9911 144236 9920
rect 144184 9877 144193 9911
rect 144193 9877 144227 9911
rect 144227 9877 144236 9911
rect 144184 9868 144236 9877
rect 144552 9911 144604 9920
rect 144552 9877 144561 9911
rect 144561 9877 144595 9911
rect 144595 9877 144604 9911
rect 147864 9936 147916 9988
rect 146668 9911 146720 9920
rect 144552 9868 144604 9877
rect 146668 9877 146677 9911
rect 146677 9877 146711 9911
rect 146711 9877 146720 9911
rect 146668 9868 146720 9877
rect 146944 9911 146996 9920
rect 146944 9877 146953 9911
rect 146953 9877 146987 9911
rect 146987 9877 146996 9911
rect 146944 9868 146996 9877
rect 147128 9911 147180 9920
rect 147128 9877 147137 9911
rect 147137 9877 147171 9911
rect 147171 9877 147180 9911
rect 147128 9868 147180 9877
rect 148140 9911 148192 9920
rect 148140 9877 148149 9911
rect 148149 9877 148183 9911
rect 148183 9877 148192 9911
rect 148140 9868 148192 9877
rect 148784 9936 148836 9988
rect 159548 10013 159557 10047
rect 159557 10013 159591 10047
rect 159591 10013 159600 10047
rect 159548 10004 159600 10013
rect 161572 10047 161624 10056
rect 161572 10013 161581 10047
rect 161581 10013 161615 10047
rect 161615 10013 161624 10047
rect 161572 10004 161624 10013
rect 163964 10047 164016 10056
rect 163964 10013 163973 10047
rect 163973 10013 164007 10047
rect 164007 10013 164016 10047
rect 163964 10004 164016 10013
rect 149980 9868 150032 9920
rect 151084 9911 151136 9920
rect 151084 9877 151093 9911
rect 151093 9877 151127 9911
rect 151127 9877 151136 9911
rect 151084 9868 151136 9877
rect 151636 9868 151688 9920
rect 153200 9868 153252 9920
rect 154856 9911 154908 9920
rect 154856 9877 154865 9911
rect 154865 9877 154899 9911
rect 154899 9877 154908 9911
rect 154856 9868 154908 9877
rect 154948 9868 155000 9920
rect 56667 9766 56719 9818
rect 56731 9766 56783 9818
rect 56795 9766 56847 9818
rect 56859 9766 56911 9818
rect 113088 9766 113140 9818
rect 113152 9766 113204 9818
rect 113216 9766 113268 9818
rect 113280 9766 113332 9818
rect 7104 9707 7156 9716
rect 7104 9673 7113 9707
rect 7113 9673 7147 9707
rect 7147 9673 7156 9707
rect 7104 9664 7156 9673
rect 8024 9664 8076 9716
rect 24216 9664 24268 9716
rect 25136 9664 25188 9716
rect 26792 9664 26844 9716
rect 27620 9707 27672 9716
rect 27620 9673 27629 9707
rect 27629 9673 27663 9707
rect 27663 9673 27672 9707
rect 27620 9664 27672 9673
rect 27804 9664 27856 9716
rect 28816 9664 28868 9716
rect 31392 9664 31444 9716
rect 2964 9596 3016 9648
rect 6092 9639 6144 9648
rect 3332 9528 3384 9580
rect 4528 9528 4580 9580
rect 6092 9605 6101 9639
rect 6101 9605 6135 9639
rect 6135 9605 6144 9639
rect 6092 9596 6144 9605
rect 15292 9639 15344 9648
rect 15292 9605 15301 9639
rect 15301 9605 15335 9639
rect 15335 9605 15344 9639
rect 15292 9596 15344 9605
rect 15568 9596 15620 9648
rect 7012 9528 7064 9580
rect 14372 9528 14424 9580
rect 3884 9460 3936 9512
rect 5908 9460 5960 9512
rect 2596 9392 2648 9444
rect 6920 9392 6972 9444
rect 1124 9324 1176 9376
rect 4068 9324 4120 9376
rect 4712 9324 4764 9376
rect 6368 9324 6420 9376
rect 10324 9460 10376 9512
rect 8852 9392 8904 9444
rect 17500 9460 17552 9512
rect 18604 9460 18656 9512
rect 19892 9528 19944 9580
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 20812 9596 20864 9648
rect 21456 9596 21508 9648
rect 22744 9596 22796 9648
rect 32588 9664 32640 9716
rect 33416 9664 33468 9716
rect 41788 9664 41840 9716
rect 41972 9664 42024 9716
rect 46756 9664 46808 9716
rect 48320 9664 48372 9716
rect 33324 9596 33376 9648
rect 33508 9596 33560 9648
rect 34428 9596 34480 9648
rect 34612 9596 34664 9648
rect 24860 9571 24912 9580
rect 24860 9537 24869 9571
rect 24869 9537 24903 9571
rect 24903 9537 24912 9571
rect 24860 9528 24912 9537
rect 25136 9528 25188 9580
rect 25320 9571 25372 9580
rect 25320 9537 25329 9571
rect 25329 9537 25363 9571
rect 25363 9537 25372 9571
rect 25320 9528 25372 9537
rect 20628 9460 20680 9512
rect 20720 9460 20772 9512
rect 21364 9460 21416 9512
rect 21824 9460 21876 9512
rect 23112 9460 23164 9512
rect 23204 9460 23256 9512
rect 26332 9460 26384 9512
rect 26976 9528 27028 9580
rect 27344 9528 27396 9580
rect 27436 9528 27488 9580
rect 30196 9528 30248 9580
rect 30288 9528 30340 9580
rect 31484 9571 31536 9580
rect 31484 9537 31493 9571
rect 31493 9537 31527 9571
rect 31527 9537 31536 9571
rect 31484 9528 31536 9537
rect 31944 9528 31996 9580
rect 35624 9596 35676 9648
rect 35716 9596 35768 9648
rect 39120 9596 39172 9648
rect 34980 9528 35032 9580
rect 36820 9571 36872 9580
rect 36820 9537 36829 9571
rect 36829 9537 36863 9571
rect 36863 9537 36872 9571
rect 36820 9528 36872 9537
rect 36912 9528 36964 9580
rect 38476 9528 38528 9580
rect 39212 9528 39264 9580
rect 39304 9528 39356 9580
rect 40224 9528 40276 9580
rect 15200 9324 15252 9376
rect 22836 9392 22888 9444
rect 34612 9460 34664 9512
rect 35532 9460 35584 9512
rect 40592 9460 40644 9512
rect 41052 9528 41104 9580
rect 41328 9596 41380 9648
rect 42616 9596 42668 9648
rect 42984 9596 43036 9648
rect 43904 9596 43956 9648
rect 41880 9571 41932 9580
rect 41328 9460 41380 9512
rect 19248 9324 19300 9376
rect 19340 9324 19392 9376
rect 21088 9324 21140 9376
rect 21916 9324 21968 9376
rect 22008 9324 22060 9376
rect 27436 9392 27488 9444
rect 29828 9392 29880 9444
rect 23020 9324 23072 9376
rect 25872 9324 25924 9376
rect 26056 9367 26108 9376
rect 26056 9333 26065 9367
rect 26065 9333 26099 9367
rect 26099 9333 26108 9367
rect 26056 9324 26108 9333
rect 26332 9324 26384 9376
rect 26424 9324 26476 9376
rect 29276 9324 29328 9376
rect 29368 9324 29420 9376
rect 31944 9392 31996 9444
rect 41880 9537 41889 9571
rect 41889 9537 41923 9571
rect 41923 9537 41932 9571
rect 41880 9528 41932 9537
rect 41972 9528 42024 9580
rect 42432 9571 42484 9580
rect 42432 9537 42441 9571
rect 42441 9537 42475 9571
rect 42475 9537 42484 9571
rect 46572 9571 46624 9580
rect 42432 9528 42484 9537
rect 46572 9537 46581 9571
rect 46581 9537 46615 9571
rect 46615 9537 46624 9571
rect 46572 9528 46624 9537
rect 48412 9596 48464 9648
rect 49976 9664 50028 9716
rect 50252 9664 50304 9716
rect 51356 9664 51408 9716
rect 50160 9596 50212 9648
rect 51172 9596 51224 9648
rect 47124 9571 47176 9580
rect 41788 9460 41840 9512
rect 46296 9460 46348 9512
rect 47124 9537 47133 9571
rect 47133 9537 47167 9571
rect 47167 9537 47176 9571
rect 47124 9528 47176 9537
rect 50528 9528 50580 9580
rect 51080 9571 51132 9580
rect 51080 9537 51089 9571
rect 51089 9537 51123 9571
rect 51123 9537 51132 9571
rect 51080 9528 51132 9537
rect 51264 9528 51316 9580
rect 52092 9596 52144 9648
rect 52184 9596 52236 9648
rect 54668 9639 54720 9648
rect 53196 9528 53248 9580
rect 49516 9460 49568 9512
rect 50620 9460 50672 9512
rect 51632 9460 51684 9512
rect 53840 9528 53892 9580
rect 54668 9605 54677 9639
rect 54677 9605 54711 9639
rect 54711 9605 54720 9639
rect 54668 9596 54720 9605
rect 54852 9596 54904 9648
rect 55680 9596 55732 9648
rect 56140 9596 56192 9648
rect 54944 9528 54996 9580
rect 55128 9571 55180 9580
rect 55128 9537 55137 9571
rect 55137 9537 55171 9571
rect 55171 9537 55180 9571
rect 55128 9528 55180 9537
rect 55864 9528 55916 9580
rect 56784 9528 56836 9580
rect 53472 9460 53524 9512
rect 55588 9460 55640 9512
rect 57704 9596 57756 9648
rect 57888 9664 57940 9716
rect 59084 9596 59136 9648
rect 59360 9664 59412 9716
rect 60556 9664 60608 9716
rect 60740 9664 60792 9716
rect 62028 9664 62080 9716
rect 64236 9707 64288 9716
rect 64236 9673 64245 9707
rect 64245 9673 64279 9707
rect 64279 9673 64288 9707
rect 64236 9664 64288 9673
rect 71688 9664 71740 9716
rect 78496 9664 78548 9716
rect 85120 9707 85172 9716
rect 85120 9673 85129 9707
rect 85129 9673 85163 9707
rect 85163 9673 85172 9707
rect 85120 9664 85172 9673
rect 86960 9664 87012 9716
rect 93308 9707 93360 9716
rect 61660 9596 61712 9648
rect 63500 9596 63552 9648
rect 68836 9596 68888 9648
rect 70860 9639 70912 9648
rect 70860 9605 70869 9639
rect 70869 9605 70903 9639
rect 70903 9605 70912 9639
rect 70860 9596 70912 9605
rect 71780 9596 71832 9648
rect 72792 9596 72844 9648
rect 73988 9596 74040 9648
rect 74448 9596 74500 9648
rect 57888 9528 57940 9580
rect 58808 9528 58860 9580
rect 59360 9571 59412 9580
rect 59360 9537 59369 9571
rect 59369 9537 59403 9571
rect 59403 9537 59412 9571
rect 59360 9528 59412 9537
rect 59912 9528 59964 9580
rect 57980 9460 58032 9512
rect 30840 9367 30892 9376
rect 30840 9333 30849 9367
rect 30849 9333 30883 9367
rect 30883 9333 30892 9367
rect 30840 9324 30892 9333
rect 31484 9324 31536 9376
rect 31668 9324 31720 9376
rect 34428 9324 34480 9376
rect 37924 9324 37976 9376
rect 39028 9367 39080 9376
rect 39028 9333 39037 9367
rect 39037 9333 39071 9367
rect 39071 9333 39080 9367
rect 39028 9324 39080 9333
rect 40224 9367 40276 9376
rect 40224 9333 40233 9367
rect 40233 9333 40267 9367
rect 40267 9333 40276 9367
rect 40224 9324 40276 9333
rect 40316 9324 40368 9376
rect 41512 9324 41564 9376
rect 47308 9392 47360 9444
rect 48320 9392 48372 9444
rect 42616 9324 42668 9376
rect 42800 9367 42852 9376
rect 42800 9333 42809 9367
rect 42809 9333 42843 9367
rect 42843 9333 42852 9367
rect 42800 9324 42852 9333
rect 44456 9324 44508 9376
rect 46664 9324 46716 9376
rect 50436 9324 50488 9376
rect 51356 9392 51408 9444
rect 53748 9392 53800 9444
rect 54300 9392 54352 9444
rect 55036 9392 55088 9444
rect 56140 9392 56192 9444
rect 51632 9324 51684 9376
rect 52276 9324 52328 9376
rect 52460 9324 52512 9376
rect 56508 9324 56560 9376
rect 56876 9324 56928 9376
rect 57336 9324 57388 9376
rect 57520 9324 57572 9376
rect 57796 9392 57848 9444
rect 60372 9392 60424 9444
rect 60832 9528 60884 9580
rect 62488 9528 62540 9580
rect 69112 9528 69164 9580
rect 70584 9528 70636 9580
rect 74356 9571 74408 9580
rect 74356 9537 74365 9571
rect 74365 9537 74399 9571
rect 74399 9537 74408 9571
rect 74356 9528 74408 9537
rect 80244 9596 80296 9648
rect 82820 9596 82872 9648
rect 87144 9596 87196 9648
rect 93308 9673 93317 9707
rect 93317 9673 93351 9707
rect 93351 9673 93360 9707
rect 93308 9664 93360 9673
rect 93400 9664 93452 9716
rect 93492 9664 93544 9716
rect 106188 9664 106240 9716
rect 108580 9664 108632 9716
rect 121000 9664 121052 9716
rect 97632 9596 97684 9648
rect 100852 9596 100904 9648
rect 104624 9596 104676 9648
rect 104992 9596 105044 9648
rect 111156 9639 111208 9648
rect 76932 9528 76984 9580
rect 80612 9528 80664 9580
rect 61936 9460 61988 9512
rect 66996 9460 67048 9512
rect 74540 9503 74592 9512
rect 74540 9469 74549 9503
rect 74549 9469 74583 9503
rect 74583 9469 74592 9503
rect 74540 9460 74592 9469
rect 80796 9503 80848 9512
rect 80796 9469 80805 9503
rect 80805 9469 80839 9503
rect 80839 9469 80848 9503
rect 80796 9460 80848 9469
rect 83188 9528 83240 9580
rect 84568 9528 84620 9580
rect 86960 9528 87012 9580
rect 87512 9528 87564 9580
rect 88524 9528 88576 9580
rect 92020 9528 92072 9580
rect 92756 9571 92808 9580
rect 92756 9537 92765 9571
rect 92765 9537 92799 9571
rect 92799 9537 92808 9571
rect 92756 9528 92808 9537
rect 94320 9528 94372 9580
rect 97908 9571 97960 9580
rect 83464 9460 83516 9512
rect 86500 9460 86552 9512
rect 89904 9503 89956 9512
rect 89904 9469 89913 9503
rect 89913 9469 89947 9503
rect 89947 9469 89956 9503
rect 89904 9460 89956 9469
rect 90272 9503 90324 9512
rect 90272 9469 90281 9503
rect 90281 9469 90315 9503
rect 90315 9469 90324 9503
rect 90272 9460 90324 9469
rect 91652 9460 91704 9512
rect 92848 9460 92900 9512
rect 96620 9460 96672 9512
rect 97908 9537 97917 9571
rect 97917 9537 97951 9571
rect 97951 9537 97960 9571
rect 97908 9528 97960 9537
rect 101036 9528 101088 9580
rect 104716 9571 104768 9580
rect 98184 9460 98236 9512
rect 99748 9460 99800 9512
rect 62212 9392 62264 9444
rect 83096 9392 83148 9444
rect 95700 9392 95752 9444
rect 103336 9460 103388 9512
rect 100944 9392 100996 9444
rect 59084 9324 59136 9376
rect 59544 9324 59596 9376
rect 60464 9324 60516 9376
rect 62948 9324 63000 9376
rect 63040 9324 63092 9376
rect 68468 9324 68520 9376
rect 76472 9367 76524 9376
rect 76472 9333 76481 9367
rect 76481 9333 76515 9367
rect 76515 9333 76524 9367
rect 76472 9324 76524 9333
rect 76564 9324 76616 9376
rect 88524 9367 88576 9376
rect 88524 9333 88533 9367
rect 88533 9333 88567 9367
rect 88567 9333 88576 9367
rect 88524 9324 88576 9333
rect 90180 9324 90232 9376
rect 91192 9324 91244 9376
rect 94320 9367 94372 9376
rect 94320 9333 94329 9367
rect 94329 9333 94363 9367
rect 94363 9333 94372 9367
rect 94320 9324 94372 9333
rect 99656 9324 99708 9376
rect 104716 9537 104725 9571
rect 104725 9537 104759 9571
rect 104759 9537 104768 9571
rect 104716 9528 104768 9537
rect 106004 9528 106056 9580
rect 108212 9528 108264 9580
rect 109592 9571 109644 9580
rect 109592 9537 109601 9571
rect 109601 9537 109635 9571
rect 109635 9537 109644 9571
rect 109592 9528 109644 9537
rect 111156 9605 111165 9639
rect 111165 9605 111199 9639
rect 111199 9605 111208 9639
rect 111156 9596 111208 9605
rect 113456 9596 113508 9648
rect 113548 9596 113600 9648
rect 119252 9596 119304 9648
rect 122748 9664 122800 9716
rect 129188 9664 129240 9716
rect 132408 9664 132460 9716
rect 141056 9707 141108 9716
rect 115204 9571 115256 9580
rect 115204 9537 115213 9571
rect 115213 9537 115247 9571
rect 115247 9537 115256 9571
rect 115204 9528 115256 9537
rect 117412 9528 117464 9580
rect 125324 9596 125376 9648
rect 126888 9639 126940 9648
rect 126888 9605 126897 9639
rect 126897 9605 126931 9639
rect 126931 9605 126940 9639
rect 126888 9596 126940 9605
rect 127808 9639 127860 9648
rect 127808 9605 127817 9639
rect 127817 9605 127851 9639
rect 127851 9605 127860 9639
rect 127808 9596 127860 9605
rect 133144 9639 133196 9648
rect 133144 9605 133153 9639
rect 133153 9605 133187 9639
rect 133187 9605 133196 9639
rect 133144 9596 133196 9605
rect 133328 9596 133380 9648
rect 135168 9639 135220 9648
rect 135168 9605 135177 9639
rect 135177 9605 135211 9639
rect 135211 9605 135220 9639
rect 135168 9596 135220 9605
rect 141056 9673 141065 9707
rect 141065 9673 141099 9707
rect 141099 9673 141108 9707
rect 141056 9664 141108 9673
rect 144552 9664 144604 9716
rect 148232 9707 148284 9716
rect 148232 9673 148241 9707
rect 148241 9673 148275 9707
rect 148275 9673 148284 9707
rect 148232 9664 148284 9673
rect 148784 9664 148836 9716
rect 120448 9571 120500 9580
rect 120448 9537 120457 9571
rect 120457 9537 120491 9571
rect 120491 9537 120500 9571
rect 120448 9528 120500 9537
rect 121460 9571 121512 9580
rect 121460 9537 121469 9571
rect 121469 9537 121503 9571
rect 121503 9537 121512 9571
rect 121460 9528 121512 9537
rect 122196 9528 122248 9580
rect 123576 9528 123628 9580
rect 108304 9460 108356 9512
rect 108488 9460 108540 9512
rect 113916 9460 113968 9512
rect 107936 9392 107988 9444
rect 115296 9435 115348 9444
rect 115296 9401 115305 9435
rect 115305 9401 115339 9435
rect 115339 9401 115348 9435
rect 115296 9392 115348 9401
rect 115572 9460 115624 9512
rect 118792 9460 118844 9512
rect 119896 9503 119948 9512
rect 119896 9469 119905 9503
rect 119905 9469 119939 9503
rect 119939 9469 119948 9503
rect 119896 9460 119948 9469
rect 121000 9460 121052 9512
rect 122472 9503 122524 9512
rect 120724 9392 120776 9444
rect 122472 9469 122481 9503
rect 122481 9469 122515 9503
rect 122515 9469 122524 9503
rect 122472 9460 122524 9469
rect 124588 9460 124640 9512
rect 127072 9528 127124 9580
rect 129464 9528 129516 9580
rect 131120 9571 131172 9580
rect 131120 9537 131129 9571
rect 131129 9537 131163 9571
rect 131163 9537 131172 9571
rect 131120 9528 131172 9537
rect 132592 9528 132644 9580
rect 136640 9528 136692 9580
rect 138112 9596 138164 9648
rect 140228 9596 140280 9648
rect 141608 9596 141660 9648
rect 142068 9596 142120 9648
rect 142436 9596 142488 9648
rect 147496 9596 147548 9648
rect 147772 9596 147824 9648
rect 151820 9639 151872 9648
rect 138388 9528 138440 9580
rect 138756 9528 138808 9580
rect 142344 9528 142396 9580
rect 143172 9571 143224 9580
rect 143172 9537 143181 9571
rect 143181 9537 143215 9571
rect 143215 9537 143224 9571
rect 143172 9528 143224 9537
rect 148048 9528 148100 9580
rect 148140 9528 148192 9580
rect 148784 9571 148836 9580
rect 148784 9537 148793 9571
rect 148793 9537 148827 9571
rect 148827 9537 148836 9571
rect 148784 9528 148836 9537
rect 150164 9571 150216 9580
rect 150164 9537 150173 9571
rect 150173 9537 150207 9571
rect 150207 9537 150216 9571
rect 150164 9528 150216 9537
rect 151820 9605 151829 9639
rect 151829 9605 151863 9639
rect 151863 9605 151872 9639
rect 151820 9596 151872 9605
rect 157156 9596 157208 9648
rect 158812 9596 158864 9648
rect 160468 9596 160520 9648
rect 154120 9528 154172 9580
rect 154948 9528 155000 9580
rect 156236 9528 156288 9580
rect 159272 9528 159324 9580
rect 163136 9528 163188 9580
rect 164332 9571 164384 9580
rect 108488 9324 108540 9376
rect 121276 9367 121328 9376
rect 121276 9333 121285 9367
rect 121285 9333 121319 9367
rect 121319 9333 121328 9367
rect 121276 9324 121328 9333
rect 123300 9392 123352 9444
rect 127164 9460 127216 9512
rect 129832 9460 129884 9512
rect 130752 9503 130804 9512
rect 130752 9469 130761 9503
rect 130761 9469 130795 9503
rect 130795 9469 130804 9503
rect 130752 9460 130804 9469
rect 131028 9460 131080 9512
rect 134064 9460 134116 9512
rect 138480 9460 138532 9512
rect 132132 9392 132184 9444
rect 134800 9392 134852 9444
rect 127532 9367 127584 9376
rect 127532 9333 127541 9367
rect 127541 9333 127575 9367
rect 127575 9333 127584 9367
rect 127532 9324 127584 9333
rect 133604 9324 133656 9376
rect 139032 9392 139084 9444
rect 141516 9460 141568 9512
rect 142896 9460 142948 9512
rect 144276 9460 144328 9512
rect 145932 9460 145984 9512
rect 148600 9460 148652 9512
rect 149336 9460 149388 9512
rect 155684 9503 155736 9512
rect 155684 9469 155693 9503
rect 155693 9469 155727 9503
rect 155727 9469 155736 9503
rect 155684 9460 155736 9469
rect 157156 9460 157208 9512
rect 157892 9460 157944 9512
rect 160468 9460 160520 9512
rect 163228 9503 163280 9512
rect 163228 9469 163237 9503
rect 163237 9469 163271 9503
rect 163271 9469 163280 9503
rect 163228 9460 163280 9469
rect 164332 9537 164341 9571
rect 164341 9537 164375 9571
rect 164375 9537 164384 9571
rect 164332 9528 164384 9537
rect 165804 9528 165856 9580
rect 166908 9571 166960 9580
rect 166908 9537 166917 9571
rect 166917 9537 166951 9571
rect 166951 9537 166960 9571
rect 166908 9528 166960 9537
rect 141792 9392 141844 9444
rect 145104 9392 145156 9444
rect 135812 9324 135864 9376
rect 138112 9324 138164 9376
rect 138204 9324 138256 9376
rect 142252 9324 142304 9376
rect 143540 9324 143592 9376
rect 149520 9392 149572 9444
rect 150900 9392 150952 9444
rect 163412 9392 163464 9444
rect 145656 9324 145708 9376
rect 151544 9324 151596 9376
rect 151728 9324 151780 9376
rect 153752 9324 153804 9376
rect 156236 9367 156288 9376
rect 156236 9333 156245 9367
rect 156245 9333 156279 9367
rect 156279 9333 156288 9367
rect 156236 9324 156288 9333
rect 157248 9367 157300 9376
rect 157248 9333 157257 9367
rect 157257 9333 157291 9367
rect 157291 9333 157300 9367
rect 157248 9324 157300 9333
rect 159548 9367 159600 9376
rect 159548 9333 159557 9367
rect 159557 9333 159591 9367
rect 159591 9333 159600 9367
rect 159548 9324 159600 9333
rect 160284 9324 160336 9376
rect 160836 9324 160888 9376
rect 164884 9324 164936 9376
rect 28456 9222 28508 9274
rect 28520 9222 28572 9274
rect 28584 9222 28636 9274
rect 28648 9222 28700 9274
rect 84878 9222 84930 9274
rect 84942 9222 84994 9274
rect 85006 9222 85058 9274
rect 85070 9222 85122 9274
rect 141299 9222 141351 9274
rect 141363 9222 141415 9274
rect 141427 9222 141479 9274
rect 141491 9222 141543 9274
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 4620 9120 4672 9172
rect 8852 9120 8904 9172
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 19892 9163 19944 9172
rect 19892 9129 19901 9163
rect 19901 9129 19935 9163
rect 19935 9129 19944 9163
rect 19892 9120 19944 9129
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 20536 9120 20588 9172
rect 5632 9052 5684 9104
rect 4068 8984 4120 9036
rect 5448 8984 5500 9036
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 5172 8916 5224 8968
rect 7748 8984 7800 9036
rect 15200 8984 15252 9036
rect 15384 8916 15436 8968
rect 16120 8916 16172 8968
rect 21548 9052 21600 9104
rect 17592 8984 17644 9036
rect 22008 9120 22060 9172
rect 24860 9163 24912 9172
rect 24860 9129 24869 9163
rect 24869 9129 24903 9163
rect 24903 9129 24912 9163
rect 24860 9120 24912 9129
rect 25320 9163 25372 9172
rect 25320 9129 25329 9163
rect 25329 9129 25363 9163
rect 25363 9129 25372 9163
rect 25320 9120 25372 9129
rect 25412 9120 25464 9172
rect 25964 9120 26016 9172
rect 28172 9120 28224 9172
rect 28816 9120 28868 9172
rect 30288 9120 30340 9172
rect 22192 9052 22244 9104
rect 31668 9095 31720 9104
rect 31668 9061 31677 9095
rect 31677 9061 31711 9095
rect 31711 9061 31720 9095
rect 31668 9052 31720 9061
rect 22836 9027 22888 9036
rect 8300 8891 8352 8900
rect 8300 8857 8309 8891
rect 8309 8857 8343 8891
rect 8343 8857 8352 8891
rect 8300 8848 8352 8857
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 19524 8916 19576 8968
rect 17960 8848 18012 8900
rect 18144 8848 18196 8900
rect 21456 8848 21508 8900
rect 21916 8916 21968 8968
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 27528 8984 27580 9036
rect 27620 8984 27672 9036
rect 23296 8848 23348 8900
rect 1492 8780 1544 8832
rect 4620 8780 4672 8832
rect 5448 8780 5500 8832
rect 12532 8780 12584 8832
rect 17040 8780 17092 8832
rect 17224 8823 17276 8832
rect 17224 8789 17233 8823
rect 17233 8789 17267 8823
rect 17267 8789 17276 8823
rect 17224 8780 17276 8789
rect 19524 8823 19576 8832
rect 19524 8789 19533 8823
rect 19533 8789 19567 8823
rect 19567 8789 19576 8823
rect 19524 8780 19576 8789
rect 21732 8780 21784 8832
rect 21824 8780 21876 8832
rect 22192 8780 22244 8832
rect 24400 8916 24452 8968
rect 25780 8916 25832 8968
rect 26056 8959 26108 8968
rect 26056 8925 26065 8959
rect 26065 8925 26099 8959
rect 26099 8925 26108 8959
rect 26056 8916 26108 8925
rect 23664 8848 23716 8900
rect 23848 8780 23900 8832
rect 24952 8780 25004 8832
rect 25136 8780 25188 8832
rect 25504 8848 25556 8900
rect 26148 8848 26200 8900
rect 28080 8916 28132 8968
rect 28356 8916 28408 8968
rect 34152 8984 34204 9036
rect 34336 9120 34388 9172
rect 34612 9052 34664 9104
rect 38108 9052 38160 9104
rect 38292 9120 38344 9172
rect 38844 9120 38896 9172
rect 39212 9163 39264 9172
rect 39212 9129 39221 9163
rect 39221 9129 39255 9163
rect 39255 9129 39264 9163
rect 39212 9120 39264 9129
rect 39580 9120 39632 9172
rect 40500 9120 40552 9172
rect 40868 9120 40920 9172
rect 41972 9120 42024 9172
rect 42432 9163 42484 9172
rect 42432 9129 42441 9163
rect 42441 9129 42475 9163
rect 42475 9129 42484 9163
rect 42432 9120 42484 9129
rect 42616 9120 42668 9172
rect 39856 9052 39908 9104
rect 39948 9052 40000 9104
rect 42984 9052 43036 9104
rect 43352 9120 43404 9172
rect 51632 9120 51684 9172
rect 53656 9120 53708 9172
rect 55128 9120 55180 9172
rect 55956 9120 56008 9172
rect 57796 9120 57848 9172
rect 57980 9120 58032 9172
rect 58348 9120 58400 9172
rect 59360 9120 59412 9172
rect 59912 9163 59964 9172
rect 59912 9129 59921 9163
rect 59921 9129 59955 9163
rect 59955 9129 59964 9163
rect 59912 9120 59964 9129
rect 60096 9120 60148 9172
rect 61384 9120 61436 9172
rect 74356 9163 74408 9172
rect 74356 9129 74365 9163
rect 74365 9129 74399 9163
rect 74399 9129 74408 9163
rect 74356 9120 74408 9129
rect 74448 9120 74500 9172
rect 76932 9120 76984 9172
rect 80612 9120 80664 9172
rect 83188 9163 83240 9172
rect 83188 9129 83197 9163
rect 83197 9129 83231 9163
rect 83231 9129 83240 9163
rect 83188 9120 83240 9129
rect 85396 9120 85448 9172
rect 86960 9163 87012 9172
rect 86960 9129 86969 9163
rect 86969 9129 87003 9163
rect 87003 9129 87012 9163
rect 86960 9120 87012 9129
rect 92020 9120 92072 9172
rect 93952 9120 94004 9172
rect 96804 9163 96856 9172
rect 46940 9052 46992 9104
rect 47124 9095 47176 9104
rect 47124 9061 47133 9095
rect 47133 9061 47167 9095
rect 47167 9061 47176 9095
rect 47124 9052 47176 9061
rect 47308 9052 47360 9104
rect 34888 8984 34940 9036
rect 35072 8984 35124 9036
rect 29184 8916 29236 8968
rect 31852 8916 31904 8968
rect 31944 8916 31996 8968
rect 36636 8984 36688 9036
rect 36820 9027 36872 9036
rect 36820 8993 36829 9027
rect 36829 8993 36863 9027
rect 36863 8993 36872 9027
rect 36820 8984 36872 8993
rect 37004 9027 37056 9036
rect 37004 8993 37013 9027
rect 37013 8993 37047 9027
rect 37047 8993 37056 9027
rect 37004 8984 37056 8993
rect 37280 8984 37332 9036
rect 36452 8916 36504 8968
rect 39028 8916 39080 8968
rect 40132 8984 40184 9036
rect 40592 8984 40644 9036
rect 41236 8984 41288 9036
rect 41512 8984 41564 9036
rect 41880 9027 41932 9036
rect 41880 8993 41889 9027
rect 41889 8993 41923 9027
rect 41923 8993 41932 9027
rect 41880 8984 41932 8993
rect 41972 8984 42024 9036
rect 46204 8984 46256 9036
rect 46572 8984 46624 9036
rect 47952 8984 48004 9036
rect 49056 8984 49108 9036
rect 50712 8984 50764 9036
rect 26608 8780 26660 8832
rect 26976 8780 27028 8832
rect 27528 8780 27580 8832
rect 27620 8780 27672 8832
rect 33508 8780 33560 8832
rect 34796 8780 34848 8832
rect 34888 8780 34940 8832
rect 38936 8780 38988 8832
rect 40592 8848 40644 8900
rect 41236 8848 41288 8900
rect 41604 8916 41656 8968
rect 42800 8959 42852 8968
rect 42064 8848 42116 8900
rect 40316 8780 40368 8832
rect 42156 8780 42208 8832
rect 42432 8848 42484 8900
rect 42800 8925 42809 8959
rect 42809 8925 42843 8959
rect 42843 8925 42852 8959
rect 42800 8916 42852 8925
rect 42892 8916 42944 8968
rect 43352 8959 43404 8968
rect 43352 8925 43361 8959
rect 43361 8925 43395 8959
rect 43395 8925 43404 8959
rect 43352 8916 43404 8925
rect 46664 8916 46716 8968
rect 47032 8916 47084 8968
rect 53196 8984 53248 9036
rect 54852 9052 54904 9104
rect 43904 8848 43956 8900
rect 48136 8848 48188 8900
rect 48228 8848 48280 8900
rect 43536 8780 43588 8832
rect 48044 8780 48096 8832
rect 48412 8823 48464 8832
rect 48412 8789 48421 8823
rect 48421 8789 48455 8823
rect 48455 8789 48464 8823
rect 48412 8780 48464 8789
rect 48688 8848 48740 8900
rect 52092 8916 52144 8968
rect 54116 8916 54168 8968
rect 54668 8984 54720 9036
rect 60740 9052 60792 9104
rect 62764 9052 62816 9104
rect 83464 9052 83516 9104
rect 55864 8984 55916 9036
rect 56140 8984 56192 9036
rect 55496 8916 55548 8968
rect 56508 8916 56560 8968
rect 56784 8916 56836 8968
rect 51540 8848 51592 8900
rect 50160 8780 50212 8832
rect 50528 8823 50580 8832
rect 50528 8789 50537 8823
rect 50537 8789 50571 8823
rect 50571 8789 50580 8823
rect 50528 8780 50580 8789
rect 52368 8780 52420 8832
rect 53288 8848 53340 8900
rect 55772 8848 55824 8900
rect 55864 8848 55916 8900
rect 56324 8848 56376 8900
rect 57612 8916 57664 8968
rect 58348 8959 58400 8968
rect 58348 8925 58357 8959
rect 58357 8925 58391 8959
rect 58391 8925 58400 8959
rect 58348 8916 58400 8925
rect 61568 8984 61620 9036
rect 63316 8984 63368 9036
rect 60924 8916 60976 8968
rect 61384 8916 61436 8968
rect 63408 8959 63460 8968
rect 63408 8925 63417 8959
rect 63417 8925 63451 8959
rect 63451 8925 63460 8959
rect 63408 8916 63460 8925
rect 72424 8984 72476 9036
rect 73620 8984 73672 9036
rect 74816 8984 74868 9036
rect 76012 8984 76064 9036
rect 76288 9027 76340 9036
rect 76288 8993 76297 9027
rect 76297 8993 76331 9027
rect 76331 8993 76340 9027
rect 76288 8984 76340 8993
rect 80060 9027 80112 9036
rect 80060 8993 80069 9027
rect 80069 8993 80103 9027
rect 80103 8993 80112 9027
rect 80060 8984 80112 8993
rect 84292 8984 84344 9036
rect 87236 8984 87288 9036
rect 89812 9052 89864 9104
rect 96804 9129 96813 9163
rect 96813 9129 96847 9163
rect 96847 9129 96856 9163
rect 96804 9120 96856 9129
rect 98184 9163 98236 9172
rect 98184 9129 98193 9163
rect 98193 9129 98227 9163
rect 98227 9129 98236 9163
rect 98184 9120 98236 9129
rect 99748 9120 99800 9172
rect 67364 8848 67416 8900
rect 81992 8891 82044 8900
rect 81992 8857 82001 8891
rect 82001 8857 82035 8891
rect 82035 8857 82044 8891
rect 81992 8848 82044 8857
rect 59176 8780 59228 8832
rect 59452 8823 59504 8832
rect 59452 8789 59461 8823
rect 59461 8789 59495 8823
rect 59495 8789 59504 8823
rect 59452 8780 59504 8789
rect 60188 8780 60240 8832
rect 60648 8780 60700 8832
rect 64788 8780 64840 8832
rect 86132 8780 86184 8832
rect 93124 9027 93176 9036
rect 93124 8993 93133 9027
rect 93133 8993 93167 9027
rect 93167 8993 93176 9027
rect 93124 8984 93176 8993
rect 97908 8984 97960 9036
rect 99564 8984 99616 9036
rect 99932 9120 99984 9172
rect 108120 9120 108172 9172
rect 108304 9163 108356 9172
rect 108304 9129 108313 9163
rect 108313 9129 108347 9163
rect 108347 9129 108356 9163
rect 108304 9120 108356 9129
rect 121460 9120 121512 9172
rect 124588 9163 124640 9172
rect 124588 9129 124597 9163
rect 124597 9129 124631 9163
rect 124631 9129 124640 9163
rect 124588 9120 124640 9129
rect 127072 9163 127124 9172
rect 127072 9129 127081 9163
rect 127081 9129 127115 9163
rect 127115 9129 127124 9163
rect 127072 9120 127124 9129
rect 133972 9120 134024 9172
rect 143356 9120 143408 9172
rect 143448 9120 143500 9172
rect 145656 9120 145708 9172
rect 145932 9163 145984 9172
rect 145932 9129 145941 9163
rect 145941 9129 145975 9163
rect 145975 9129 145984 9163
rect 145932 9120 145984 9129
rect 146116 9120 146168 9172
rect 100116 9052 100168 9104
rect 100576 9052 100628 9104
rect 101956 9052 102008 9104
rect 105360 8984 105412 9036
rect 106556 8984 106608 9036
rect 89904 8959 89956 8968
rect 89904 8925 89913 8959
rect 89913 8925 89947 8959
rect 89947 8925 89956 8959
rect 89904 8916 89956 8925
rect 94320 8959 94372 8968
rect 89536 8780 89588 8832
rect 94320 8925 94329 8959
rect 94329 8925 94363 8959
rect 94363 8925 94372 8959
rect 94320 8916 94372 8925
rect 92020 8780 92072 8832
rect 92756 8823 92808 8832
rect 92756 8789 92765 8823
rect 92765 8789 92799 8823
rect 92799 8789 92808 8823
rect 92756 8780 92808 8789
rect 99012 8916 99064 8968
rect 99656 8916 99708 8968
rect 100484 8916 100536 8968
rect 100576 8916 100628 8968
rect 103980 8916 104032 8968
rect 112260 9027 112312 9036
rect 112260 8993 112269 9027
rect 112269 8993 112303 9027
rect 112303 8993 112312 9027
rect 112260 8984 112312 8993
rect 113916 9027 113968 9036
rect 113916 8993 113925 9027
rect 113925 8993 113959 9027
rect 113959 8993 113968 9027
rect 113916 8984 113968 8993
rect 115296 8916 115348 8968
rect 115572 9027 115624 9036
rect 115572 8993 115581 9027
rect 115581 8993 115615 9027
rect 115615 8993 115624 9027
rect 115572 8984 115624 8993
rect 115664 8984 115716 9036
rect 120724 9052 120776 9104
rect 119160 8984 119212 9036
rect 119436 8984 119488 9036
rect 117504 8916 117556 8968
rect 118792 8959 118844 8968
rect 118792 8925 118801 8959
rect 118801 8925 118835 8959
rect 118835 8925 118844 8959
rect 118792 8916 118844 8925
rect 121276 8959 121328 8968
rect 121276 8925 121285 8959
rect 121285 8925 121319 8959
rect 121319 8925 121328 8959
rect 121276 8916 121328 8925
rect 124588 8984 124640 9036
rect 124772 9052 124824 9104
rect 130752 9052 130804 9104
rect 136180 9052 136232 9104
rect 147772 9052 147824 9104
rect 147956 9095 148008 9104
rect 147956 9061 147965 9095
rect 147965 9061 147999 9095
rect 147999 9061 148008 9095
rect 147956 9052 148008 9061
rect 125784 8984 125836 9036
rect 127532 9027 127584 9036
rect 127532 8993 127541 9027
rect 127541 8993 127575 9027
rect 127575 8993 127584 9027
rect 127532 8984 127584 8993
rect 130292 8984 130344 9036
rect 131120 9027 131172 9036
rect 131120 8993 131129 9027
rect 131129 8993 131163 9027
rect 131163 8993 131172 9027
rect 131120 8984 131172 8993
rect 138020 9027 138072 9036
rect 138020 8993 138029 9027
rect 138029 8993 138063 9027
rect 138063 8993 138072 9027
rect 138020 8984 138072 8993
rect 140412 8984 140464 9036
rect 103336 8891 103388 8900
rect 103336 8857 103345 8891
rect 103345 8857 103379 8891
rect 103379 8857 103388 8891
rect 103336 8848 103388 8857
rect 104164 8848 104216 8900
rect 96252 8823 96304 8832
rect 96252 8789 96261 8823
rect 96261 8789 96295 8823
rect 96295 8789 96304 8823
rect 96252 8780 96304 8789
rect 96620 8823 96672 8832
rect 96620 8789 96629 8823
rect 96629 8789 96663 8823
rect 96663 8789 96672 8823
rect 97264 8823 97316 8832
rect 96620 8780 96672 8789
rect 97264 8789 97273 8823
rect 97273 8789 97307 8823
rect 97307 8789 97316 8823
rect 97264 8780 97316 8789
rect 100484 8780 100536 8832
rect 101036 8823 101088 8832
rect 101036 8789 101045 8823
rect 101045 8789 101079 8823
rect 101079 8789 101088 8823
rect 101036 8780 101088 8789
rect 102876 8823 102928 8832
rect 102876 8789 102885 8823
rect 102885 8789 102919 8823
rect 102919 8789 102928 8823
rect 102876 8780 102928 8789
rect 104716 8780 104768 8832
rect 106280 8780 106332 8832
rect 106464 8823 106516 8832
rect 106464 8789 106473 8823
rect 106473 8789 106507 8823
rect 106507 8789 106516 8823
rect 106464 8780 106516 8789
rect 106648 8848 106700 8900
rect 118516 8848 118568 8900
rect 121184 8848 121236 8900
rect 126704 8848 126756 8900
rect 131396 8959 131448 8968
rect 131396 8925 131405 8959
rect 131405 8925 131439 8959
rect 131439 8925 131448 8959
rect 131396 8916 131448 8925
rect 140688 8916 140740 8968
rect 139860 8848 139912 8900
rect 142804 8984 142856 9036
rect 143816 8984 143868 9036
rect 144184 8984 144236 9036
rect 148784 9027 148836 9036
rect 109592 8780 109644 8832
rect 115296 8823 115348 8832
rect 115296 8789 115305 8823
rect 115305 8789 115339 8823
rect 115339 8789 115348 8823
rect 115296 8780 115348 8789
rect 117504 8823 117556 8832
rect 117504 8789 117513 8823
rect 117513 8789 117547 8823
rect 117547 8789 117556 8823
rect 117504 8780 117556 8789
rect 120448 8780 120500 8832
rect 121000 8780 121052 8832
rect 123576 8823 123628 8832
rect 123576 8789 123585 8823
rect 123585 8789 123619 8823
rect 123619 8789 123628 8823
rect 123576 8780 123628 8789
rect 125324 8780 125376 8832
rect 125692 8780 125744 8832
rect 127164 8780 127216 8832
rect 129740 8823 129792 8832
rect 129740 8789 129749 8823
rect 129749 8789 129783 8823
rect 129783 8789 129792 8823
rect 129740 8780 129792 8789
rect 140872 8823 140924 8832
rect 140872 8789 140881 8823
rect 140881 8789 140915 8823
rect 140915 8789 140924 8823
rect 143172 8916 143224 8968
rect 146024 8916 146076 8968
rect 145840 8848 145892 8900
rect 146576 8848 146628 8900
rect 148784 8993 148793 9027
rect 148793 8993 148827 9027
rect 148827 8993 148836 9027
rect 148784 8984 148836 8993
rect 149336 9027 149388 9036
rect 149336 8993 149345 9027
rect 149345 8993 149379 9027
rect 149379 8993 149388 9027
rect 149336 8984 149388 8993
rect 152004 9052 152056 9104
rect 154948 9120 155000 9172
rect 157156 9163 157208 9172
rect 157156 9129 157165 9163
rect 157165 9129 157199 9163
rect 157199 9129 157208 9163
rect 157156 9120 157208 9129
rect 165804 9163 165856 9172
rect 165804 9129 165813 9163
rect 165813 9129 165847 9163
rect 165847 9129 165856 9163
rect 165804 9120 165856 9129
rect 156144 9052 156196 9104
rect 158260 9052 158312 9104
rect 160836 9052 160888 9104
rect 162032 9052 162084 9104
rect 140872 8780 140924 8789
rect 141976 8780 142028 8832
rect 143264 8780 143316 8832
rect 143356 8780 143408 8832
rect 146300 8823 146352 8832
rect 146300 8789 146309 8823
rect 146309 8789 146343 8823
rect 146343 8789 146352 8823
rect 146300 8780 146352 8789
rect 149152 8780 149204 8832
rect 151820 8984 151872 9036
rect 153844 8984 153896 9036
rect 156052 9027 156104 9036
rect 156052 8993 156061 9027
rect 156061 8993 156095 9027
rect 156095 8993 156104 9027
rect 156052 8984 156104 8993
rect 158628 9027 158680 9036
rect 158628 8993 158637 9027
rect 158637 8993 158671 9027
rect 158671 8993 158680 9027
rect 158628 8984 158680 8993
rect 160468 9027 160520 9036
rect 160468 8993 160477 9027
rect 160477 8993 160511 9027
rect 160511 8993 160520 9027
rect 160468 8984 160520 8993
rect 161204 8984 161256 9036
rect 166724 9052 166776 9104
rect 151820 8848 151872 8900
rect 151728 8780 151780 8832
rect 153660 8823 153712 8832
rect 153660 8789 153669 8823
rect 153669 8789 153703 8823
rect 153703 8789 153712 8823
rect 153660 8780 153712 8789
rect 153844 8780 153896 8832
rect 155960 8959 156012 8968
rect 155960 8925 155969 8959
rect 155969 8925 156003 8959
rect 156003 8925 156012 8959
rect 155960 8916 156012 8925
rect 157248 8959 157300 8968
rect 157248 8925 157257 8959
rect 157257 8925 157291 8959
rect 157291 8925 157300 8959
rect 157248 8916 157300 8925
rect 158536 8959 158588 8968
rect 158536 8925 158545 8959
rect 158545 8925 158579 8959
rect 158579 8925 158588 8959
rect 158536 8916 158588 8925
rect 164424 8916 164476 8968
rect 163228 8848 163280 8900
rect 159272 8780 159324 8832
rect 162308 8823 162360 8832
rect 162308 8789 162317 8823
rect 162317 8789 162351 8823
rect 162351 8789 162360 8823
rect 162308 8780 162360 8789
rect 166908 8823 166960 8832
rect 166908 8789 166917 8823
rect 166917 8789 166951 8823
rect 166951 8789 166960 8823
rect 166908 8780 166960 8789
rect 56667 8678 56719 8730
rect 56731 8678 56783 8730
rect 56795 8678 56847 8730
rect 56859 8678 56911 8730
rect 113088 8678 113140 8730
rect 113152 8678 113204 8730
rect 113216 8678 113268 8730
rect 113280 8678 113332 8730
rect 1860 8576 1912 8628
rect 5172 8576 5224 8628
rect 5540 8619 5592 8628
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 4068 8508 4120 8560
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 5264 8508 5316 8560
rect 22284 8576 22336 8628
rect 8852 8508 8904 8560
rect 17592 8508 17644 8560
rect 17684 8508 17736 8560
rect 5540 8440 5592 8492
rect 2228 8304 2280 8356
rect 9956 8440 10008 8492
rect 14832 8483 14884 8492
rect 13360 8372 13412 8424
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 15108 8440 15160 8492
rect 15660 8440 15712 8492
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16672 8440 16724 8492
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 18604 8508 18656 8560
rect 21640 8508 21692 8560
rect 21732 8508 21784 8560
rect 24400 8576 24452 8628
rect 25688 8576 25740 8628
rect 25964 8576 26016 8628
rect 26056 8576 26108 8628
rect 27528 8576 27580 8628
rect 33600 8576 33652 8628
rect 34428 8576 34480 8628
rect 40960 8576 41012 8628
rect 41512 8619 41564 8628
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 17132 8304 17184 8356
rect 9220 8236 9272 8288
rect 15108 8236 15160 8288
rect 18328 8372 18380 8424
rect 17408 8347 17460 8356
rect 17408 8313 17417 8347
rect 17417 8313 17451 8347
rect 17451 8313 17460 8347
rect 17408 8304 17460 8313
rect 17960 8304 18012 8356
rect 19616 8347 19668 8356
rect 19616 8313 19625 8347
rect 19625 8313 19659 8347
rect 19659 8313 19668 8347
rect 19616 8304 19668 8313
rect 21824 8483 21876 8492
rect 20904 8415 20956 8424
rect 20904 8381 20913 8415
rect 20913 8381 20947 8415
rect 20947 8381 20956 8415
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 22928 8440 22980 8492
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 21456 8415 21508 8424
rect 20904 8372 20956 8381
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 33232 8508 33284 8560
rect 34152 8508 34204 8560
rect 36912 8508 36964 8560
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 25596 8483 25648 8492
rect 25596 8449 25605 8483
rect 25605 8449 25639 8483
rect 25639 8449 25648 8483
rect 25596 8440 25648 8449
rect 25780 8440 25832 8492
rect 25136 8372 25188 8424
rect 22100 8347 22152 8356
rect 22100 8313 22109 8347
rect 22109 8313 22143 8347
rect 22143 8313 22152 8347
rect 22100 8304 22152 8313
rect 23020 8347 23072 8356
rect 23020 8313 23029 8347
rect 23029 8313 23063 8347
rect 23063 8313 23072 8347
rect 23020 8304 23072 8313
rect 23940 8347 23992 8356
rect 23940 8313 23949 8347
rect 23949 8313 23983 8347
rect 23983 8313 23992 8347
rect 23940 8304 23992 8313
rect 26608 8440 26660 8492
rect 34428 8440 34480 8492
rect 34796 8483 34848 8492
rect 34796 8449 34805 8483
rect 34805 8449 34839 8483
rect 34839 8449 34848 8483
rect 34796 8440 34848 8449
rect 34888 8440 34940 8492
rect 35532 8483 35584 8492
rect 35532 8449 35541 8483
rect 35541 8449 35575 8483
rect 35575 8449 35584 8483
rect 35532 8440 35584 8449
rect 36728 8483 36780 8492
rect 36728 8449 36737 8483
rect 36737 8449 36771 8483
rect 36771 8449 36780 8483
rect 36728 8440 36780 8449
rect 41512 8585 41521 8619
rect 41521 8585 41555 8619
rect 41555 8585 41564 8619
rect 41512 8576 41564 8585
rect 45928 8576 45980 8628
rect 46112 8576 46164 8628
rect 47492 8576 47544 8628
rect 47584 8576 47636 8628
rect 48228 8576 48280 8628
rect 48504 8576 48556 8628
rect 49332 8576 49384 8628
rect 49792 8576 49844 8628
rect 50252 8576 50304 8628
rect 51540 8576 51592 8628
rect 51724 8576 51776 8628
rect 42432 8508 42484 8560
rect 42616 8508 42668 8560
rect 43076 8508 43128 8560
rect 26700 8372 26752 8424
rect 29184 8372 29236 8424
rect 29276 8372 29328 8424
rect 17592 8236 17644 8288
rect 25780 8236 25832 8288
rect 33784 8304 33836 8356
rect 34336 8372 34388 8424
rect 37188 8372 37240 8424
rect 38292 8440 38344 8492
rect 39396 8440 39448 8492
rect 39856 8440 39908 8492
rect 40960 8440 41012 8492
rect 41604 8440 41656 8492
rect 41696 8440 41748 8492
rect 43536 8440 43588 8492
rect 39212 8372 39264 8424
rect 40684 8372 40736 8424
rect 40776 8372 40828 8424
rect 48320 8508 48372 8560
rect 48412 8508 48464 8560
rect 39764 8304 39816 8356
rect 40040 8304 40092 8356
rect 46480 8440 46532 8492
rect 45560 8372 45612 8424
rect 48780 8440 48832 8492
rect 49976 8508 50028 8560
rect 52644 8576 52696 8628
rect 53196 8576 53248 8628
rect 54024 8576 54076 8628
rect 55772 8576 55824 8628
rect 57796 8576 57848 8628
rect 57888 8576 57940 8628
rect 58532 8576 58584 8628
rect 59268 8576 59320 8628
rect 59452 8619 59504 8628
rect 59452 8585 59461 8619
rect 59461 8585 59495 8619
rect 59495 8585 59504 8619
rect 59452 8576 59504 8585
rect 52368 8508 52420 8560
rect 56784 8508 56836 8560
rect 46756 8372 46808 8424
rect 46848 8372 46900 8424
rect 49884 8372 49936 8424
rect 45744 8279 45796 8288
rect 45744 8245 45753 8279
rect 45753 8245 45787 8279
rect 45787 8245 45796 8279
rect 45744 8236 45796 8245
rect 45928 8304 45980 8356
rect 47860 8304 47912 8356
rect 48412 8304 48464 8356
rect 52000 8440 52052 8492
rect 52736 8483 52788 8492
rect 50160 8372 50212 8424
rect 52368 8372 52420 8424
rect 52736 8449 52745 8483
rect 52745 8449 52779 8483
rect 52779 8449 52788 8483
rect 52736 8440 52788 8449
rect 54760 8440 54812 8492
rect 53012 8372 53064 8424
rect 54852 8372 54904 8424
rect 55680 8440 55732 8492
rect 55956 8440 56008 8492
rect 56048 8440 56100 8492
rect 56232 8440 56284 8492
rect 58256 8508 58308 8560
rect 57428 8440 57480 8492
rect 57612 8440 57664 8492
rect 58992 8483 59044 8492
rect 58992 8449 59001 8483
rect 59001 8449 59035 8483
rect 59035 8449 59044 8483
rect 58992 8440 59044 8449
rect 59084 8440 59136 8492
rect 63040 8576 63092 8628
rect 63408 8576 63460 8628
rect 74080 8576 74132 8628
rect 74356 8576 74408 8628
rect 80152 8619 80204 8628
rect 80152 8585 80161 8619
rect 80161 8585 80195 8619
rect 80195 8585 80204 8619
rect 80152 8576 80204 8585
rect 85856 8576 85908 8628
rect 88340 8576 88392 8628
rect 90272 8576 90324 8628
rect 60004 8508 60056 8560
rect 60188 8483 60240 8492
rect 60188 8449 60197 8483
rect 60197 8449 60231 8483
rect 60231 8449 60240 8483
rect 60188 8440 60240 8449
rect 60372 8440 60424 8492
rect 60556 8440 60608 8492
rect 58348 8372 58400 8424
rect 59176 8372 59228 8424
rect 59820 8372 59872 8424
rect 65064 8508 65116 8560
rect 66260 8508 66312 8560
rect 76564 8508 76616 8560
rect 90456 8508 90508 8560
rect 60832 8440 60884 8492
rect 64420 8483 64472 8492
rect 62856 8415 62908 8424
rect 62856 8381 62865 8415
rect 62865 8381 62899 8415
rect 62899 8381 62908 8415
rect 62856 8372 62908 8381
rect 63868 8415 63920 8424
rect 63868 8381 63877 8415
rect 63877 8381 63911 8415
rect 63911 8381 63920 8415
rect 63868 8372 63920 8381
rect 64420 8449 64429 8483
rect 64429 8449 64463 8483
rect 64463 8449 64472 8483
rect 64420 8440 64472 8449
rect 83464 8483 83516 8492
rect 83464 8449 83473 8483
rect 83473 8449 83507 8483
rect 83507 8449 83516 8483
rect 83464 8440 83516 8449
rect 87604 8440 87656 8492
rect 68100 8372 68152 8424
rect 71780 8415 71832 8424
rect 71780 8381 71789 8415
rect 71789 8381 71823 8415
rect 71823 8381 71832 8415
rect 71780 8372 71832 8381
rect 81992 8415 82044 8424
rect 50712 8304 50764 8356
rect 50528 8236 50580 8288
rect 51080 8236 51132 8288
rect 51632 8304 51684 8356
rect 52184 8304 52236 8356
rect 53288 8304 53340 8356
rect 54944 8347 54996 8356
rect 51816 8236 51868 8288
rect 51908 8236 51960 8288
rect 54392 8279 54444 8288
rect 54392 8245 54401 8279
rect 54401 8245 54435 8279
rect 54435 8245 54444 8279
rect 54392 8236 54444 8245
rect 54944 8313 54953 8347
rect 54953 8313 54987 8347
rect 54987 8313 54996 8347
rect 54944 8304 54996 8313
rect 55312 8304 55364 8356
rect 56784 8304 56836 8356
rect 64328 8304 64380 8356
rect 81992 8381 82001 8415
rect 82001 8381 82035 8415
rect 82035 8381 82044 8415
rect 81992 8372 82044 8381
rect 83004 8415 83056 8424
rect 83004 8381 83013 8415
rect 83013 8381 83047 8415
rect 83047 8381 83056 8415
rect 83004 8372 83056 8381
rect 87236 8372 87288 8424
rect 87972 8372 88024 8424
rect 89260 8483 89312 8492
rect 89260 8449 89269 8483
rect 89269 8449 89303 8483
rect 89303 8449 89312 8483
rect 91652 8483 91704 8492
rect 89260 8440 89312 8449
rect 86868 8304 86920 8356
rect 90456 8372 90508 8424
rect 91652 8449 91661 8483
rect 91661 8449 91695 8483
rect 91695 8449 91704 8483
rect 91652 8440 91704 8449
rect 92848 8483 92900 8492
rect 92848 8449 92857 8483
rect 92857 8449 92891 8483
rect 92891 8449 92900 8483
rect 92848 8440 92900 8449
rect 98276 8576 98328 8628
rect 94964 8508 95016 8560
rect 94596 8440 94648 8492
rect 92112 8372 92164 8424
rect 91100 8304 91152 8356
rect 95608 8347 95660 8356
rect 95608 8313 95617 8347
rect 95617 8313 95651 8347
rect 95651 8313 95660 8347
rect 95608 8304 95660 8313
rect 98000 8440 98052 8492
rect 103336 8576 103388 8628
rect 108396 8576 108448 8628
rect 102692 8508 102744 8560
rect 119896 8576 119948 8628
rect 121276 8576 121328 8628
rect 124680 8619 124732 8628
rect 124680 8585 124689 8619
rect 124689 8585 124723 8619
rect 124723 8585 124732 8619
rect 124680 8576 124732 8585
rect 128084 8619 128136 8628
rect 128084 8585 128093 8619
rect 128093 8585 128127 8619
rect 128127 8585 128136 8619
rect 128084 8576 128136 8585
rect 141608 8576 141660 8628
rect 142252 8576 142304 8628
rect 145104 8576 145156 8628
rect 146300 8576 146352 8628
rect 152740 8576 152792 8628
rect 153936 8576 153988 8628
rect 157156 8576 157208 8628
rect 161664 8576 161716 8628
rect 164792 8576 164844 8628
rect 96620 8372 96672 8424
rect 100300 8440 100352 8492
rect 102876 8440 102928 8492
rect 103980 8440 104032 8492
rect 104624 8483 104676 8492
rect 55864 8236 55916 8288
rect 56140 8236 56192 8288
rect 57244 8236 57296 8288
rect 57428 8236 57480 8288
rect 60832 8236 60884 8288
rect 61016 8279 61068 8288
rect 61016 8245 61025 8279
rect 61025 8245 61059 8279
rect 61059 8245 61068 8279
rect 61016 8236 61068 8245
rect 79416 8236 79468 8288
rect 83832 8279 83884 8288
rect 83832 8245 83841 8279
rect 83841 8245 83875 8279
rect 83875 8245 83884 8279
rect 83832 8236 83884 8245
rect 87512 8279 87564 8288
rect 87512 8245 87521 8279
rect 87521 8245 87555 8279
rect 87555 8245 87564 8279
rect 87512 8236 87564 8245
rect 98000 8279 98052 8288
rect 98000 8245 98009 8279
rect 98009 8245 98043 8279
rect 98043 8245 98052 8279
rect 98000 8236 98052 8245
rect 99380 8236 99432 8288
rect 104624 8449 104633 8483
rect 104633 8449 104667 8483
rect 104667 8449 104676 8483
rect 104624 8440 104676 8449
rect 106464 8440 106516 8492
rect 107108 8483 107160 8492
rect 107108 8449 107117 8483
rect 107117 8449 107151 8483
rect 107151 8449 107160 8483
rect 107108 8440 107160 8449
rect 108488 8483 108540 8492
rect 108488 8449 108497 8483
rect 108497 8449 108531 8483
rect 108531 8449 108540 8483
rect 108488 8440 108540 8449
rect 120908 8508 120960 8560
rect 115848 8440 115900 8492
rect 118516 8440 118568 8492
rect 121184 8440 121236 8492
rect 121368 8483 121420 8492
rect 121368 8449 121377 8483
rect 121377 8449 121411 8483
rect 121411 8449 121420 8483
rect 121368 8440 121420 8449
rect 125692 8483 125744 8492
rect 125692 8449 125701 8483
rect 125701 8449 125735 8483
rect 125735 8449 125744 8483
rect 125692 8440 125744 8449
rect 127072 8508 127124 8560
rect 138112 8508 138164 8560
rect 131028 8483 131080 8492
rect 100300 8347 100352 8356
rect 100300 8313 100309 8347
rect 100309 8313 100343 8347
rect 100343 8313 100352 8347
rect 100300 8304 100352 8313
rect 101220 8304 101272 8356
rect 113456 8372 113508 8424
rect 116584 8372 116636 8424
rect 119896 8415 119948 8424
rect 119896 8381 119905 8415
rect 119905 8381 119939 8415
rect 119939 8381 119948 8415
rect 119896 8372 119948 8381
rect 120908 8415 120960 8424
rect 120908 8381 120917 8415
rect 120917 8381 120951 8415
rect 120951 8381 120960 8415
rect 120908 8372 120960 8381
rect 121000 8372 121052 8424
rect 125968 8372 126020 8424
rect 126704 8415 126756 8424
rect 126704 8381 126713 8415
rect 126713 8381 126747 8415
rect 126747 8381 126756 8415
rect 126704 8372 126756 8381
rect 102324 8236 102376 8288
rect 108580 8236 108632 8288
rect 109776 8236 109828 8288
rect 112260 8279 112312 8288
rect 112260 8245 112269 8279
rect 112269 8245 112303 8279
rect 112303 8245 112312 8279
rect 112260 8236 112312 8245
rect 129556 8415 129608 8424
rect 129556 8381 129565 8415
rect 129565 8381 129599 8415
rect 129599 8381 129608 8415
rect 129556 8372 129608 8381
rect 131028 8449 131037 8483
rect 131037 8449 131071 8483
rect 131071 8449 131080 8483
rect 131028 8440 131080 8449
rect 139216 8440 139268 8492
rect 141792 8415 141844 8424
rect 115848 8236 115900 8288
rect 116492 8236 116544 8288
rect 131212 8236 131264 8288
rect 141792 8381 141801 8415
rect 141801 8381 141835 8415
rect 141835 8381 141844 8415
rect 141792 8372 141844 8381
rect 142436 8440 142488 8492
rect 143356 8440 143408 8492
rect 143908 8483 143960 8492
rect 143908 8449 143917 8483
rect 143917 8449 143951 8483
rect 143951 8449 143960 8483
rect 143908 8440 143960 8449
rect 146852 8508 146904 8560
rect 153016 8508 153068 8560
rect 154212 8508 154264 8560
rect 155316 8508 155368 8560
rect 157524 8508 157576 8560
rect 159364 8508 159416 8560
rect 160100 8508 160152 8560
rect 162400 8508 162452 8560
rect 162768 8508 162820 8560
rect 165160 8508 165212 8560
rect 146208 8440 146260 8492
rect 146392 8483 146444 8492
rect 146392 8449 146396 8483
rect 146396 8449 146430 8483
rect 146430 8449 146444 8483
rect 147772 8483 147824 8492
rect 146392 8440 146444 8449
rect 147772 8449 147781 8483
rect 147781 8449 147815 8483
rect 147815 8449 147824 8483
rect 147772 8440 147824 8449
rect 151176 8440 151228 8492
rect 152464 8440 152516 8492
rect 153200 8440 153252 8492
rect 140596 8304 140648 8356
rect 142804 8304 142856 8356
rect 143264 8304 143316 8356
rect 149244 8415 149296 8424
rect 149244 8381 149253 8415
rect 149253 8381 149287 8415
rect 149287 8381 149296 8415
rect 149244 8372 149296 8381
rect 150532 8415 150584 8424
rect 150532 8381 150541 8415
rect 150541 8381 150575 8415
rect 150575 8381 150584 8415
rect 150532 8372 150584 8381
rect 153108 8372 153160 8424
rect 154856 8440 154908 8492
rect 156052 8483 156104 8492
rect 156052 8449 156061 8483
rect 156061 8449 156095 8483
rect 156095 8449 156104 8483
rect 156052 8440 156104 8449
rect 158996 8440 159048 8492
rect 160744 8483 160796 8492
rect 155408 8372 155460 8424
rect 159456 8415 159508 8424
rect 159456 8381 159465 8415
rect 159465 8381 159499 8415
rect 159499 8381 159508 8415
rect 159456 8372 159508 8381
rect 160744 8449 160753 8483
rect 160753 8449 160787 8483
rect 160787 8449 160796 8483
rect 160744 8440 160796 8449
rect 163780 8440 163832 8492
rect 164700 8440 164752 8492
rect 165620 8483 165672 8492
rect 165620 8449 165629 8483
rect 165629 8449 165663 8483
rect 165663 8449 165672 8483
rect 165620 8440 165672 8449
rect 161112 8372 161164 8424
rect 166172 8372 166224 8424
rect 145196 8304 145248 8356
rect 150900 8304 150952 8356
rect 154304 8347 154356 8356
rect 154304 8313 154313 8347
rect 154313 8313 154347 8347
rect 154347 8313 154356 8347
rect 154304 8304 154356 8313
rect 155040 8304 155092 8356
rect 156512 8304 156564 8356
rect 158536 8347 158588 8356
rect 158536 8313 158545 8347
rect 158545 8313 158579 8347
rect 158579 8313 158588 8347
rect 158536 8304 158588 8313
rect 159732 8304 159784 8356
rect 162124 8304 162176 8356
rect 164608 8304 164660 8356
rect 133052 8236 133104 8288
rect 145012 8279 145064 8288
rect 145012 8245 145021 8279
rect 145021 8245 145055 8279
rect 145055 8245 145064 8279
rect 145012 8236 145064 8245
rect 151176 8279 151228 8288
rect 151176 8245 151185 8279
rect 151185 8245 151219 8279
rect 151219 8245 151228 8279
rect 151176 8236 151228 8245
rect 28456 8134 28508 8186
rect 28520 8134 28572 8186
rect 28584 8134 28636 8186
rect 28648 8134 28700 8186
rect 84878 8134 84930 8186
rect 84942 8134 84994 8186
rect 85006 8134 85058 8186
rect 85070 8134 85122 8186
rect 141299 8134 141351 8186
rect 141363 8134 141415 8186
rect 141427 8134 141479 8186
rect 141491 8134 141543 8186
rect 756 8032 808 8084
rect 8024 8032 8076 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 17684 8032 17736 8084
rect 18144 8032 18196 8084
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 20352 8032 20404 8084
rect 21824 8075 21876 8084
rect 21824 8041 21833 8075
rect 21833 8041 21867 8075
rect 21867 8041 21876 8075
rect 21824 8032 21876 8041
rect 23664 8032 23716 8084
rect 25136 8075 25188 8084
rect 25136 8041 25145 8075
rect 25145 8041 25179 8075
rect 25179 8041 25188 8075
rect 25136 8032 25188 8041
rect 25596 8075 25648 8084
rect 25596 8041 25605 8075
rect 25605 8041 25639 8075
rect 25639 8041 25648 8075
rect 25596 8032 25648 8041
rect 26056 8032 26108 8084
rect 26516 8032 26568 8084
rect 34612 8032 34664 8084
rect 34796 8075 34848 8084
rect 34796 8041 34805 8075
rect 34805 8041 34839 8075
rect 34839 8041 34848 8075
rect 34796 8032 34848 8041
rect 35532 8075 35584 8084
rect 35532 8041 35541 8075
rect 35541 8041 35575 8075
rect 35575 8041 35584 8075
rect 35532 8032 35584 8041
rect 35900 8032 35952 8084
rect 39212 8032 39264 8084
rect 39396 8075 39448 8084
rect 39396 8041 39405 8075
rect 39405 8041 39439 8075
rect 39439 8041 39448 8075
rect 39396 8032 39448 8041
rect 40040 8032 40092 8084
rect 40776 8032 40828 8084
rect 3608 7964 3660 8016
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 6092 7964 6144 8016
rect 12256 7964 12308 8016
rect 14096 7964 14148 8016
rect 25504 7964 25556 8016
rect 25872 8007 25924 8016
rect 25872 7973 25881 8007
rect 25881 7973 25915 8007
rect 25915 7973 25924 8007
rect 25872 7964 25924 7973
rect 26148 7964 26200 8016
rect 41236 8007 41288 8016
rect 41236 7973 41245 8007
rect 41245 7973 41279 8007
rect 41279 7973 41288 8007
rect 41236 7964 41288 7973
rect 41604 8032 41656 8084
rect 44732 8032 44784 8084
rect 44824 8032 44876 8084
rect 49792 8032 49844 8084
rect 49976 8075 50028 8084
rect 49976 8041 49985 8075
rect 49985 8041 50019 8075
rect 50019 8041 50028 8075
rect 49976 8032 50028 8041
rect 50160 8032 50212 8084
rect 51908 8032 51960 8084
rect 52736 8075 52788 8084
rect 52736 8041 52745 8075
rect 52745 8041 52779 8075
rect 52779 8041 52788 8075
rect 53012 8075 53064 8084
rect 52736 8032 52788 8041
rect 53012 8041 53021 8075
rect 53021 8041 53055 8075
rect 53055 8041 53064 8075
rect 53012 8032 53064 8041
rect 55680 8075 55732 8084
rect 55680 8041 55689 8075
rect 55689 8041 55723 8075
rect 55723 8041 55732 8075
rect 55680 8032 55732 8041
rect 15844 7896 15896 7948
rect 16120 7939 16172 7948
rect 16120 7905 16129 7939
rect 16129 7905 16163 7939
rect 16163 7905 16172 7939
rect 16120 7896 16172 7905
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 14832 7871 14884 7880
rect 3608 7692 3660 7744
rect 14832 7837 14841 7871
rect 14841 7837 14875 7871
rect 14875 7837 14884 7871
rect 14832 7828 14884 7837
rect 17592 7828 17644 7880
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 21640 7896 21692 7948
rect 22284 7896 22336 7948
rect 23388 7896 23440 7948
rect 21732 7828 21784 7880
rect 22100 7871 22152 7880
rect 22100 7837 22109 7871
rect 22109 7837 22143 7871
rect 22143 7837 22152 7871
rect 22100 7828 22152 7837
rect 23940 7828 23992 7880
rect 5540 7735 5592 7744
rect 5540 7701 5549 7735
rect 5549 7701 5583 7735
rect 5583 7701 5592 7735
rect 5540 7692 5592 7701
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 14096 7692 14148 7744
rect 14464 7692 14516 7744
rect 19156 7692 19208 7744
rect 19800 7692 19852 7744
rect 20812 7760 20864 7812
rect 20996 7692 21048 7744
rect 25596 7828 25648 7880
rect 25780 7871 25832 7880
rect 25780 7837 25789 7871
rect 25789 7837 25823 7871
rect 25823 7837 25832 7871
rect 25780 7828 25832 7837
rect 24860 7760 24912 7812
rect 27528 7828 27580 7880
rect 35532 7828 35584 7880
rect 36728 7871 36780 7880
rect 36728 7837 36737 7871
rect 36737 7837 36771 7871
rect 36771 7837 36780 7871
rect 36728 7828 36780 7837
rect 24768 7692 24820 7744
rect 33784 7760 33836 7812
rect 33876 7760 33928 7812
rect 34428 7760 34480 7812
rect 37188 7828 37240 7880
rect 38752 7828 38804 7880
rect 38936 7896 38988 7948
rect 39672 7896 39724 7948
rect 39764 7896 39816 7948
rect 27620 7692 27672 7744
rect 35164 7692 35216 7744
rect 36268 7692 36320 7744
rect 37464 7692 37516 7744
rect 39580 7692 39632 7744
rect 41144 7828 41196 7880
rect 41328 7896 41380 7948
rect 42708 7896 42760 7948
rect 44824 7896 44876 7948
rect 45744 7939 45796 7948
rect 45744 7905 45753 7939
rect 45753 7905 45787 7939
rect 45787 7905 45796 7939
rect 45744 7896 45796 7905
rect 45836 7896 45888 7948
rect 47492 7964 47544 8016
rect 48872 7964 48924 8016
rect 41420 7828 41472 7880
rect 42064 7828 42116 7880
rect 46388 7828 46440 7880
rect 46940 7896 46992 7948
rect 49056 7896 49108 7948
rect 50068 7964 50120 8016
rect 50252 7964 50304 8016
rect 56876 8032 56928 8084
rect 57060 8032 57112 8084
rect 58992 8075 59044 8084
rect 40868 7692 40920 7744
rect 40960 7692 41012 7744
rect 41144 7692 41196 7744
rect 41604 7692 41656 7744
rect 46940 7760 46992 7812
rect 47584 7828 47636 7880
rect 48780 7871 48832 7880
rect 47768 7760 47820 7812
rect 48504 7760 48556 7812
rect 48780 7837 48789 7871
rect 48789 7837 48823 7871
rect 48823 7837 48832 7871
rect 48780 7828 48832 7837
rect 49516 7896 49568 7948
rect 56048 7896 56100 7948
rect 49976 7828 50028 7880
rect 50528 7828 50580 7880
rect 49516 7760 49568 7812
rect 49608 7760 49660 7812
rect 51356 7828 51408 7880
rect 51540 7871 51592 7880
rect 51540 7837 51549 7871
rect 51549 7837 51583 7871
rect 51583 7837 51592 7871
rect 51540 7828 51592 7837
rect 51724 7871 51776 7880
rect 51724 7837 51733 7871
rect 51733 7837 51767 7871
rect 51767 7837 51776 7871
rect 51724 7828 51776 7837
rect 52092 7871 52144 7880
rect 52092 7837 52101 7871
rect 52101 7837 52135 7871
rect 52135 7837 52144 7871
rect 52092 7828 52144 7837
rect 52276 7828 52328 7880
rect 54024 7828 54076 7880
rect 54392 7871 54444 7880
rect 54392 7837 54401 7871
rect 54401 7837 54435 7871
rect 54435 7837 54444 7871
rect 54392 7828 54444 7837
rect 54576 7871 54628 7880
rect 54576 7837 54585 7871
rect 54585 7837 54619 7871
rect 54619 7837 54628 7871
rect 54576 7828 54628 7837
rect 42340 7692 42392 7744
rect 47308 7692 47360 7744
rect 47584 7735 47636 7744
rect 47584 7701 47593 7735
rect 47593 7701 47627 7735
rect 47627 7701 47636 7735
rect 47584 7692 47636 7701
rect 47676 7692 47728 7744
rect 50160 7692 50212 7744
rect 50252 7692 50304 7744
rect 55588 7760 55640 7812
rect 55864 7760 55916 7812
rect 57336 7896 57388 7948
rect 57520 7896 57572 7948
rect 57980 7939 58032 7948
rect 57980 7905 57989 7939
rect 57989 7905 58023 7939
rect 58023 7905 58032 7939
rect 57980 7896 58032 7905
rect 58440 7896 58492 7948
rect 58348 7871 58400 7880
rect 58348 7837 58357 7871
rect 58357 7837 58391 7871
rect 58391 7837 58400 7871
rect 58348 7828 58400 7837
rect 58992 8041 59001 8075
rect 59001 8041 59035 8075
rect 59035 8041 59044 8075
rect 58992 8032 59044 8041
rect 60188 8075 60240 8084
rect 60188 8041 60197 8075
rect 60197 8041 60231 8075
rect 60231 8041 60240 8075
rect 60188 8032 60240 8041
rect 60556 8075 60608 8084
rect 60556 8041 60565 8075
rect 60565 8041 60599 8075
rect 60599 8041 60608 8075
rect 60556 8032 60608 8041
rect 62856 8032 62908 8084
rect 71780 8032 71832 8084
rect 87236 8075 87288 8084
rect 87236 8041 87245 8075
rect 87245 8041 87279 8075
rect 87279 8041 87288 8075
rect 87236 8032 87288 8041
rect 92848 8032 92900 8084
rect 102876 8032 102928 8084
rect 107108 8075 107160 8084
rect 107108 8041 107117 8075
rect 107117 8041 107151 8075
rect 107151 8041 107160 8075
rect 107108 8032 107160 8041
rect 108488 8075 108540 8084
rect 108488 8041 108497 8075
rect 108497 8041 108531 8075
rect 108531 8041 108540 8075
rect 108488 8032 108540 8041
rect 124956 8032 125008 8084
rect 125692 8032 125744 8084
rect 129556 8075 129608 8084
rect 61016 7939 61068 7948
rect 59360 7828 59412 7880
rect 60648 7828 60700 7880
rect 57060 7760 57112 7812
rect 61016 7905 61025 7939
rect 61025 7905 61059 7939
rect 61059 7905 61068 7939
rect 61016 7896 61068 7905
rect 62120 7939 62172 7948
rect 62120 7905 62129 7939
rect 62129 7905 62163 7939
rect 62163 7905 62172 7939
rect 62120 7896 62172 7905
rect 68008 7896 68060 7948
rect 71780 7939 71832 7948
rect 71780 7905 71789 7939
rect 71789 7905 71823 7939
rect 71823 7905 71832 7939
rect 71780 7896 71832 7905
rect 72792 7939 72844 7948
rect 72792 7905 72801 7939
rect 72801 7905 72835 7939
rect 72835 7905 72844 7939
rect 72792 7896 72844 7905
rect 79416 7939 79468 7948
rect 79416 7905 79425 7939
rect 79425 7905 79459 7939
rect 79459 7905 79468 7939
rect 79416 7896 79468 7905
rect 80428 7939 80480 7948
rect 80428 7905 80437 7939
rect 80437 7905 80471 7939
rect 80471 7905 80480 7939
rect 80428 7896 80480 7905
rect 81992 7896 82044 7948
rect 83372 7896 83424 7948
rect 83832 7896 83884 7948
rect 89260 7964 89312 8016
rect 87512 7939 87564 7948
rect 87512 7905 87521 7939
rect 87521 7905 87555 7939
rect 87555 7905 87564 7939
rect 87512 7896 87564 7905
rect 88340 7896 88392 7948
rect 90272 7896 90324 7948
rect 91100 7939 91152 7948
rect 91100 7905 91109 7939
rect 91109 7905 91143 7939
rect 91143 7905 91152 7939
rect 91100 7896 91152 7905
rect 98460 7896 98512 7948
rect 72884 7828 72936 7880
rect 80888 7871 80940 7880
rect 50804 7692 50856 7744
rect 52276 7692 52328 7744
rect 52368 7692 52420 7744
rect 55772 7692 55824 7744
rect 56232 7692 56284 7744
rect 56508 7692 56560 7744
rect 57244 7692 57296 7744
rect 59084 7692 59136 7744
rect 64420 7760 64472 7812
rect 71136 7760 71188 7812
rect 67732 7692 67784 7744
rect 68836 7735 68888 7744
rect 68836 7701 68845 7735
rect 68845 7701 68879 7735
rect 68879 7701 68888 7735
rect 68836 7692 68888 7701
rect 80888 7837 80897 7871
rect 80897 7837 80931 7871
rect 80931 7837 80940 7871
rect 80888 7828 80940 7837
rect 84752 7871 84804 7880
rect 84752 7837 84761 7871
rect 84761 7837 84795 7871
rect 84795 7837 84804 7871
rect 84752 7828 84804 7837
rect 80152 7692 80204 7744
rect 83464 7692 83516 7744
rect 91284 7828 91336 7880
rect 100392 7896 100444 7948
rect 103336 7939 103388 7948
rect 103336 7905 103345 7939
rect 103345 7905 103379 7939
rect 103379 7905 103388 7939
rect 103336 7896 103388 7905
rect 103796 7896 103848 7948
rect 112260 7939 112312 7948
rect 112260 7905 112269 7939
rect 112269 7905 112303 7939
rect 112303 7905 112312 7939
rect 112260 7896 112312 7905
rect 91652 7760 91704 7812
rect 106556 7760 106608 7812
rect 114100 7896 114152 7948
rect 116124 7828 116176 7880
rect 119896 7896 119948 7948
rect 126244 7896 126296 7948
rect 127532 7896 127584 7948
rect 129556 8041 129565 8075
rect 129565 8041 129599 8075
rect 129599 8041 129608 8075
rect 129556 8032 129608 8041
rect 146392 8032 146444 8084
rect 147036 8032 147088 8084
rect 152464 8075 152516 8084
rect 152464 8041 152473 8075
rect 152473 8041 152507 8075
rect 152507 8041 152516 8075
rect 152464 8032 152516 8041
rect 154856 8032 154908 8084
rect 166172 8075 166224 8084
rect 166172 8041 166181 8075
rect 166181 8041 166215 8075
rect 166215 8041 166224 8075
rect 166172 8032 166224 8041
rect 131212 7964 131264 8016
rect 129740 7939 129792 7948
rect 129740 7905 129749 7939
rect 129749 7905 129783 7939
rect 129783 7905 129792 7939
rect 129740 7896 129792 7905
rect 129832 7896 129884 7948
rect 133052 7939 133104 7948
rect 133052 7905 133061 7939
rect 133061 7905 133095 7939
rect 133095 7905 133104 7939
rect 133052 7896 133104 7905
rect 149428 7964 149480 8016
rect 156788 8007 156840 8016
rect 156788 7973 156797 8007
rect 156797 7973 156831 8007
rect 156831 7973 156840 8007
rect 156788 7964 156840 7973
rect 164792 8007 164844 8016
rect 164792 7973 164801 8007
rect 164801 7973 164835 8007
rect 164835 7973 164844 8007
rect 164792 7964 164844 7973
rect 140872 7896 140924 7948
rect 141792 7939 141844 7948
rect 141792 7905 141801 7939
rect 141801 7905 141835 7939
rect 141835 7905 141844 7939
rect 141792 7896 141844 7905
rect 142804 7939 142856 7948
rect 142804 7905 142813 7939
rect 142813 7905 142847 7939
rect 142847 7905 142856 7939
rect 142804 7896 142856 7905
rect 145012 7939 145064 7948
rect 145012 7905 145021 7939
rect 145021 7905 145055 7939
rect 145055 7905 145064 7939
rect 145012 7896 145064 7905
rect 145104 7896 145156 7948
rect 147128 7896 147180 7948
rect 150900 7939 150952 7948
rect 150900 7905 150909 7939
rect 150909 7905 150943 7939
rect 150943 7905 150952 7939
rect 150900 7896 150952 7905
rect 153476 7896 153528 7948
rect 159364 7939 159416 7948
rect 56667 7590 56719 7642
rect 56731 7590 56783 7642
rect 56795 7590 56847 7642
rect 56859 7590 56911 7642
rect 5540 7488 5592 7540
rect 14464 7488 14516 7540
rect 19156 7488 19208 7540
rect 27528 7488 27580 7540
rect 27620 7488 27672 7540
rect 33968 7488 34020 7540
rect 34612 7488 34664 7540
rect 40592 7488 40644 7540
rect 40684 7488 40736 7540
rect 42248 7488 42300 7540
rect 4068 7420 4120 7472
rect 18696 7463 18748 7472
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 4528 7284 4580 7336
rect 9588 7352 9640 7404
rect 13912 7352 13964 7404
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8024 7284 8076 7336
rect 14280 7284 14332 7336
rect 15200 7327 15252 7336
rect 15200 7293 15209 7327
rect 15209 7293 15243 7327
rect 15243 7293 15252 7327
rect 15200 7284 15252 7293
rect 16028 7327 16080 7336
rect 16028 7293 16037 7327
rect 16037 7293 16071 7327
rect 16071 7293 16080 7327
rect 16028 7284 16080 7293
rect 18696 7429 18705 7463
rect 18705 7429 18739 7463
rect 18739 7429 18748 7463
rect 18696 7420 18748 7429
rect 19248 7420 19300 7472
rect 19800 7420 19852 7472
rect 19892 7352 19944 7404
rect 19156 7284 19208 7336
rect 19248 7284 19300 7336
rect 20628 7284 20680 7336
rect 20996 7420 21048 7472
rect 21364 7420 21416 7472
rect 34152 7463 34204 7472
rect 21916 7352 21968 7404
rect 25044 7395 25096 7404
rect 23572 7284 23624 7336
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 24676 7327 24728 7336
rect 23664 7284 23716 7293
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 25044 7361 25053 7395
rect 25053 7361 25087 7395
rect 25087 7361 25096 7395
rect 25044 7352 25096 7361
rect 28908 7352 28960 7404
rect 34152 7429 34161 7463
rect 34161 7429 34195 7463
rect 34195 7429 34204 7463
rect 34152 7420 34204 7429
rect 34244 7420 34296 7472
rect 35900 7352 35952 7404
rect 36268 7395 36320 7404
rect 36268 7361 36277 7395
rect 36277 7361 36311 7395
rect 36311 7361 36320 7395
rect 36268 7352 36320 7361
rect 8208 7216 8260 7268
rect 18696 7216 18748 7268
rect 18972 7216 19024 7268
rect 9588 7148 9640 7200
rect 13912 7148 13964 7200
rect 20812 7216 20864 7268
rect 21732 7216 21784 7268
rect 26424 7284 26476 7336
rect 26516 7327 26568 7336
rect 26516 7293 26525 7327
rect 26525 7293 26559 7327
rect 26559 7293 26568 7327
rect 26516 7284 26568 7293
rect 26700 7284 26752 7336
rect 27620 7284 27672 7336
rect 34428 7284 34480 7336
rect 34796 7284 34848 7336
rect 35256 7284 35308 7336
rect 32496 7216 32548 7268
rect 21272 7148 21324 7200
rect 21548 7148 21600 7200
rect 23112 7191 23164 7200
rect 23112 7157 23121 7191
rect 23121 7157 23155 7191
rect 23155 7157 23164 7191
rect 23112 7148 23164 7157
rect 23204 7148 23256 7200
rect 28816 7148 28868 7200
rect 28908 7148 28960 7200
rect 33692 7148 33744 7200
rect 33968 7191 34020 7200
rect 33968 7157 33977 7191
rect 33977 7157 34011 7191
rect 34011 7157 34020 7191
rect 33968 7148 34020 7157
rect 34612 7148 34664 7200
rect 36360 7148 36412 7200
rect 37188 7352 37240 7404
rect 37280 7327 37332 7336
rect 37280 7293 37289 7327
rect 37289 7293 37323 7327
rect 37323 7293 37332 7327
rect 37280 7284 37332 7293
rect 37464 7284 37516 7336
rect 38476 7352 38528 7404
rect 39488 7352 39540 7404
rect 39672 7420 39724 7472
rect 42616 7488 42668 7540
rect 45560 7488 45612 7540
rect 45744 7488 45796 7540
rect 71688 7488 71740 7540
rect 83372 7531 83424 7540
rect 83372 7497 83381 7531
rect 83381 7497 83415 7531
rect 83415 7497 83424 7531
rect 83372 7488 83424 7497
rect 97172 7692 97224 7744
rect 102324 7735 102376 7744
rect 102324 7701 102333 7735
rect 102333 7701 102367 7735
rect 102367 7701 102376 7735
rect 102324 7692 102376 7701
rect 104348 7692 104400 7744
rect 104624 7692 104676 7744
rect 116216 7760 116268 7812
rect 116584 7760 116636 7812
rect 133420 7828 133472 7880
rect 134248 7871 134300 7880
rect 134248 7837 134257 7871
rect 134257 7837 134291 7871
rect 134291 7837 134300 7871
rect 134248 7828 134300 7837
rect 146392 7871 146444 7880
rect 120816 7760 120868 7812
rect 121368 7760 121420 7812
rect 122472 7760 122524 7812
rect 118792 7692 118844 7744
rect 118976 7735 119028 7744
rect 118976 7701 118985 7735
rect 118985 7701 119019 7735
rect 119019 7701 119028 7735
rect 118976 7692 119028 7701
rect 121460 7692 121512 7744
rect 127072 7735 127124 7744
rect 127072 7701 127081 7735
rect 127081 7701 127115 7735
rect 127115 7701 127124 7735
rect 127072 7692 127124 7701
rect 127992 7692 128044 7744
rect 131028 7692 131080 7744
rect 146392 7837 146401 7871
rect 146401 7837 146435 7871
rect 146435 7837 146444 7871
rect 146392 7828 146444 7837
rect 143908 7760 143960 7812
rect 145380 7760 145432 7812
rect 146484 7692 146536 7744
rect 150440 7828 150492 7880
rect 150992 7871 151044 7880
rect 150992 7837 151001 7871
rect 151001 7837 151035 7871
rect 151035 7837 151044 7871
rect 150992 7828 151044 7837
rect 149428 7692 149480 7744
rect 152924 7735 152976 7744
rect 152924 7701 152933 7735
rect 152933 7701 152967 7735
rect 152967 7701 152976 7735
rect 156144 7828 156196 7880
rect 159364 7905 159373 7939
rect 159373 7905 159407 7939
rect 159407 7905 159416 7939
rect 159364 7896 159416 7905
rect 161112 7939 161164 7948
rect 161112 7905 161121 7939
rect 161121 7905 161155 7939
rect 161155 7905 161164 7939
rect 161112 7896 161164 7905
rect 162124 7939 162176 7948
rect 162124 7905 162133 7939
rect 162133 7905 162167 7939
rect 162167 7905 162176 7939
rect 162124 7896 162176 7905
rect 166724 7939 166776 7948
rect 166724 7905 166733 7939
rect 166733 7905 166767 7939
rect 166767 7905 166776 7939
rect 166724 7896 166776 7905
rect 158720 7828 158772 7880
rect 159732 7871 159784 7880
rect 159732 7837 159741 7871
rect 159741 7837 159775 7871
rect 159775 7837 159784 7871
rect 159732 7828 159784 7837
rect 161940 7828 161992 7880
rect 164608 7871 164660 7880
rect 157524 7760 157576 7812
rect 154948 7735 155000 7744
rect 152924 7692 152976 7701
rect 154948 7701 154957 7735
rect 154957 7701 154991 7735
rect 154991 7701 155000 7735
rect 154948 7692 155000 7701
rect 160744 7735 160796 7744
rect 160744 7701 160753 7735
rect 160753 7701 160787 7735
rect 160787 7701 160796 7735
rect 160744 7692 160796 7701
rect 163412 7735 163464 7744
rect 163412 7701 163421 7735
rect 163421 7701 163455 7735
rect 163455 7701 163464 7735
rect 164608 7837 164617 7871
rect 164617 7837 164651 7871
rect 164651 7837 164660 7871
rect 164608 7828 164660 7837
rect 163412 7692 163464 7701
rect 165620 7692 165672 7744
rect 96436 7624 96488 7676
rect 113088 7590 113140 7642
rect 113152 7590 113204 7642
rect 113216 7590 113268 7642
rect 113280 7590 113332 7642
rect 100392 7488 100444 7540
rect 108488 7488 108540 7540
rect 108580 7488 108632 7540
rect 142436 7531 142488 7540
rect 40592 7352 40644 7404
rect 38660 7284 38712 7336
rect 39304 7284 39356 7336
rect 39396 7284 39448 7336
rect 37004 7216 37056 7268
rect 40684 7284 40736 7336
rect 41788 7352 41840 7404
rect 42248 7352 42300 7404
rect 39948 7216 40000 7268
rect 41420 7284 41472 7336
rect 41604 7327 41656 7336
rect 41604 7293 41613 7327
rect 41613 7293 41647 7327
rect 41647 7293 41656 7327
rect 41604 7284 41656 7293
rect 41696 7284 41748 7336
rect 42156 7284 42208 7336
rect 42616 7284 42668 7336
rect 44272 7327 44324 7336
rect 44272 7293 44281 7327
rect 44281 7293 44315 7327
rect 44315 7293 44324 7327
rect 44272 7284 44324 7293
rect 44548 7352 44600 7404
rect 47860 7420 47912 7472
rect 46756 7352 46808 7404
rect 46940 7352 46992 7404
rect 47768 7352 47820 7404
rect 48504 7420 48556 7472
rect 48872 7420 48924 7472
rect 49792 7420 49844 7472
rect 50804 7420 50856 7472
rect 51448 7420 51500 7472
rect 51632 7420 51684 7472
rect 52000 7420 52052 7472
rect 52736 7420 52788 7472
rect 53564 7420 53616 7472
rect 54392 7420 54444 7472
rect 54852 7463 54904 7472
rect 54852 7429 54861 7463
rect 54861 7429 54895 7463
rect 54895 7429 54904 7463
rect 54852 7420 54904 7429
rect 55588 7352 55640 7404
rect 48136 7327 48188 7336
rect 48136 7293 48145 7327
rect 48145 7293 48179 7327
rect 48179 7293 48188 7327
rect 48136 7284 48188 7293
rect 48872 7284 48924 7336
rect 54852 7284 54904 7336
rect 56140 7352 56192 7404
rect 56784 7352 56836 7404
rect 56968 7352 57020 7404
rect 57428 7352 57480 7404
rect 59820 7395 59872 7404
rect 59820 7361 59829 7395
rect 59829 7361 59863 7395
rect 59863 7361 59872 7395
rect 59820 7352 59872 7361
rect 61016 7420 61068 7472
rect 90456 7463 90508 7472
rect 90456 7429 90465 7463
rect 90465 7429 90499 7463
rect 90499 7429 90508 7463
rect 90456 7420 90508 7429
rect 91284 7463 91336 7472
rect 91284 7429 91293 7463
rect 91293 7429 91327 7463
rect 91327 7429 91336 7463
rect 91284 7420 91336 7429
rect 94320 7420 94372 7472
rect 98644 7420 98696 7472
rect 63868 7352 63920 7404
rect 68836 7395 68888 7404
rect 68836 7361 68845 7395
rect 68845 7361 68879 7395
rect 68879 7361 68888 7395
rect 68836 7352 68888 7361
rect 70124 7395 70176 7404
rect 70124 7361 70133 7395
rect 70133 7361 70167 7395
rect 70167 7361 70176 7395
rect 70124 7352 70176 7361
rect 81348 7395 81400 7404
rect 81348 7361 81357 7395
rect 81357 7361 81391 7395
rect 81391 7361 81400 7395
rect 81348 7352 81400 7361
rect 57980 7284 58032 7336
rect 59084 7284 59136 7336
rect 69848 7327 69900 7336
rect 40868 7216 40920 7268
rect 42432 7216 42484 7268
rect 42800 7216 42852 7268
rect 37188 7148 37240 7200
rect 38568 7148 38620 7200
rect 43536 7148 43588 7200
rect 44180 7148 44232 7200
rect 44272 7148 44324 7200
rect 44916 7191 44968 7200
rect 44916 7157 44925 7191
rect 44925 7157 44959 7191
rect 44959 7157 44968 7191
rect 44916 7148 44968 7157
rect 45100 7216 45152 7268
rect 46940 7148 46992 7200
rect 47032 7148 47084 7200
rect 51908 7148 51960 7200
rect 52092 7191 52144 7200
rect 52092 7157 52101 7191
rect 52101 7157 52135 7191
rect 52135 7157 52144 7191
rect 52092 7148 52144 7157
rect 55496 7148 55548 7200
rect 56048 7216 56100 7268
rect 56968 7216 57020 7268
rect 69848 7293 69857 7327
rect 69857 7293 69891 7327
rect 69891 7293 69900 7327
rect 69848 7284 69900 7293
rect 79784 7327 79836 7336
rect 79784 7293 79793 7327
rect 79793 7293 79827 7327
rect 79827 7293 79836 7327
rect 79784 7284 79836 7293
rect 80796 7327 80848 7336
rect 80796 7293 80805 7327
rect 80805 7293 80839 7327
rect 80839 7293 80848 7327
rect 80796 7284 80848 7293
rect 87604 7284 87656 7336
rect 87788 7327 87840 7336
rect 87788 7293 87797 7327
rect 87797 7293 87831 7327
rect 87831 7293 87840 7327
rect 87788 7284 87840 7293
rect 89076 7327 89128 7336
rect 89076 7293 89085 7327
rect 89085 7293 89119 7327
rect 89119 7293 89128 7327
rect 89076 7284 89128 7293
rect 102324 7352 102376 7404
rect 103980 7395 104032 7404
rect 103980 7361 103989 7395
rect 103989 7361 104023 7395
rect 104023 7361 104032 7395
rect 103980 7352 104032 7361
rect 109316 7352 109368 7404
rect 114100 7352 114152 7404
rect 115940 7352 115992 7404
rect 96528 7284 96580 7336
rect 96896 7284 96948 7336
rect 104532 7284 104584 7336
rect 113272 7284 113324 7336
rect 113456 7284 113508 7336
rect 115756 7327 115808 7336
rect 115756 7293 115765 7327
rect 115765 7293 115799 7327
rect 115799 7293 115808 7327
rect 115756 7284 115808 7293
rect 142436 7497 142445 7531
rect 142445 7497 142479 7531
rect 142479 7497 142488 7531
rect 142436 7488 142488 7497
rect 145012 7488 145064 7540
rect 147036 7531 147088 7540
rect 147036 7497 147045 7531
rect 147045 7497 147079 7531
rect 147079 7497 147088 7531
rect 147036 7488 147088 7497
rect 147128 7488 147180 7540
rect 149244 7488 149296 7540
rect 150440 7531 150492 7540
rect 116952 7420 117004 7472
rect 150440 7497 150449 7531
rect 150449 7497 150483 7531
rect 150483 7497 150492 7531
rect 150440 7488 150492 7497
rect 156144 7531 156196 7540
rect 156144 7497 156153 7531
rect 156153 7497 156187 7531
rect 156187 7497 156196 7531
rect 156144 7488 156196 7497
rect 158720 7531 158772 7540
rect 158720 7497 158729 7531
rect 158729 7497 158763 7531
rect 158763 7497 158772 7531
rect 158720 7488 158772 7497
rect 159456 7531 159508 7540
rect 159456 7497 159465 7531
rect 159465 7497 159499 7531
rect 159499 7497 159508 7531
rect 159456 7488 159508 7497
rect 163412 7488 163464 7540
rect 117136 7395 117188 7404
rect 117136 7361 117145 7395
rect 117145 7361 117179 7395
rect 117179 7361 117188 7395
rect 117136 7352 117188 7361
rect 118976 7395 119028 7404
rect 118976 7361 118985 7395
rect 118985 7361 119019 7395
rect 119019 7361 119028 7395
rect 118976 7352 119028 7361
rect 120632 7352 120684 7404
rect 122932 7395 122984 7404
rect 122932 7361 122941 7395
rect 122941 7361 122975 7395
rect 122975 7361 122984 7395
rect 122932 7352 122984 7361
rect 121368 7327 121420 7336
rect 121368 7293 121377 7327
rect 121377 7293 121411 7327
rect 121411 7293 121420 7327
rect 121368 7284 121420 7293
rect 125416 7327 125468 7336
rect 56600 7148 56652 7200
rect 57612 7191 57664 7200
rect 57612 7157 57621 7191
rect 57621 7157 57655 7191
rect 57655 7157 57664 7191
rect 57612 7148 57664 7157
rect 58348 7191 58400 7200
rect 58348 7157 58357 7191
rect 58357 7157 58391 7191
rect 58391 7157 58400 7191
rect 58348 7148 58400 7157
rect 60280 7191 60332 7200
rect 60280 7157 60289 7191
rect 60289 7157 60323 7191
rect 60323 7157 60332 7191
rect 60280 7148 60332 7157
rect 81900 7191 81952 7200
rect 81900 7157 81909 7191
rect 81909 7157 81943 7191
rect 81943 7157 81952 7191
rect 81900 7148 81952 7157
rect 104348 7148 104400 7200
rect 125416 7293 125425 7327
rect 125425 7293 125459 7327
rect 125459 7293 125468 7327
rect 125416 7284 125468 7293
rect 152924 7420 152976 7472
rect 126888 7395 126940 7404
rect 126888 7361 126897 7395
rect 126897 7361 126931 7395
rect 126931 7361 126940 7395
rect 126888 7352 126940 7361
rect 133236 7352 133288 7404
rect 144368 7395 144420 7404
rect 144368 7361 144377 7395
rect 144377 7361 144411 7395
rect 144411 7361 144420 7395
rect 144368 7352 144420 7361
rect 149336 7395 149388 7404
rect 149336 7361 149345 7395
rect 149345 7361 149379 7395
rect 149379 7361 149388 7395
rect 149336 7352 149388 7361
rect 155868 7395 155920 7404
rect 155868 7361 155877 7395
rect 155877 7361 155911 7395
rect 155911 7361 155920 7395
rect 155868 7352 155920 7361
rect 160928 7352 160980 7404
rect 164976 7395 165028 7404
rect 164976 7361 164985 7395
rect 164985 7361 165019 7395
rect 165019 7361 165028 7395
rect 164976 7352 165028 7361
rect 127440 7284 127492 7336
rect 129832 7284 129884 7336
rect 132224 7327 132276 7336
rect 132224 7293 132233 7327
rect 132233 7293 132267 7327
rect 132267 7293 132276 7327
rect 132224 7284 132276 7293
rect 133420 7327 133472 7336
rect 133420 7293 133429 7327
rect 133429 7293 133463 7327
rect 133463 7293 133472 7327
rect 133420 7284 133472 7293
rect 142804 7327 142856 7336
rect 142804 7293 142813 7327
rect 142813 7293 142847 7327
rect 142847 7293 142856 7327
rect 142804 7284 142856 7293
rect 143816 7327 143868 7336
rect 143816 7293 143825 7327
rect 143825 7293 143859 7327
rect 143859 7293 143868 7327
rect 143816 7284 143868 7293
rect 148048 7327 148100 7336
rect 148048 7293 148057 7327
rect 148057 7293 148091 7327
rect 148091 7293 148100 7327
rect 148048 7284 148100 7293
rect 149520 7327 149572 7336
rect 149520 7293 149529 7327
rect 149529 7293 149563 7327
rect 149563 7293 149572 7327
rect 149520 7284 149572 7293
rect 155224 7284 155276 7336
rect 155316 7327 155368 7336
rect 155316 7293 155325 7327
rect 155325 7293 155359 7327
rect 155359 7293 155368 7327
rect 159916 7327 159968 7336
rect 155316 7284 155368 7293
rect 159916 7293 159925 7327
rect 159925 7293 159959 7327
rect 159959 7293 159968 7327
rect 159916 7284 159968 7293
rect 160836 7284 160888 7336
rect 163320 7284 163372 7336
rect 164240 7284 164292 7336
rect 134892 7191 134944 7200
rect 134892 7157 134901 7191
rect 134901 7157 134935 7191
rect 134935 7157 134944 7191
rect 134892 7148 134944 7157
rect 141792 7191 141844 7200
rect 141792 7157 141801 7191
rect 141801 7157 141835 7191
rect 141835 7157 141844 7191
rect 141792 7148 141844 7157
rect 153016 7191 153068 7200
rect 153016 7157 153025 7191
rect 153025 7157 153059 7191
rect 153059 7157 153068 7191
rect 153016 7148 153068 7157
rect 163504 7191 163556 7200
rect 163504 7157 163513 7191
rect 163513 7157 163547 7191
rect 163547 7157 163556 7191
rect 163504 7148 163556 7157
rect 28456 7046 28508 7098
rect 28520 7046 28572 7098
rect 28584 7046 28636 7098
rect 28648 7046 28700 7098
rect 84878 7046 84930 7098
rect 84942 7046 84994 7098
rect 85006 7046 85058 7098
rect 85070 7046 85122 7098
rect 141299 7046 141351 7098
rect 141363 7046 141415 7098
rect 141427 7046 141479 7098
rect 141491 7046 141543 7098
rect 4804 6944 4856 6996
rect 5724 6919 5776 6928
rect 5724 6885 5733 6919
rect 5733 6885 5767 6919
rect 5767 6885 5776 6919
rect 5724 6876 5776 6885
rect 9772 6876 9824 6928
rect 14096 6944 14148 6996
rect 15476 6944 15528 6996
rect 23664 6987 23716 6996
rect 23664 6953 23673 6987
rect 23673 6953 23707 6987
rect 23707 6953 23716 6987
rect 23664 6944 23716 6953
rect 23848 6944 23900 6996
rect 26240 6944 26292 6996
rect 26516 6944 26568 6996
rect 26608 6944 26660 6996
rect 28816 6944 28868 6996
rect 33784 6944 33836 6996
rect 36452 6944 36504 6996
rect 36912 6944 36964 6996
rect 38292 6944 38344 6996
rect 38476 6987 38528 6996
rect 38476 6953 38485 6987
rect 38485 6953 38519 6987
rect 38519 6953 38528 6987
rect 38476 6944 38528 6953
rect 38844 6944 38896 6996
rect 39396 6987 39448 6996
rect 39396 6953 39405 6987
rect 39405 6953 39439 6987
rect 39439 6953 39448 6987
rect 39396 6944 39448 6953
rect 39488 6944 39540 6996
rect 41420 6944 41472 6996
rect 3608 6808 3660 6860
rect 6368 6851 6420 6860
rect 4252 6740 4304 6792
rect 6368 6817 6377 6851
rect 6377 6817 6411 6851
rect 6411 6817 6420 6851
rect 6368 6808 6420 6817
rect 7932 6808 7984 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 13360 6808 13412 6860
rect 14280 6851 14332 6860
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 14280 6808 14332 6817
rect 15292 6808 15344 6860
rect 19524 6808 19576 6860
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 20904 6808 20956 6860
rect 21364 6808 21416 6860
rect 23664 6808 23716 6860
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 26792 6808 26844 6860
rect 21088 6740 21140 6792
rect 16488 6715 16540 6724
rect 16488 6681 16497 6715
rect 16497 6681 16531 6715
rect 16531 6681 16540 6715
rect 16488 6672 16540 6681
rect 10876 6647 10928 6656
rect 10876 6613 10885 6647
rect 10885 6613 10919 6647
rect 10919 6613 10928 6647
rect 10876 6604 10928 6613
rect 21272 6647 21324 6656
rect 21272 6613 21281 6647
rect 21281 6613 21315 6647
rect 21315 6613 21324 6647
rect 22468 6740 22520 6792
rect 26240 6740 26292 6792
rect 29276 6808 29328 6860
rect 27988 6783 28040 6792
rect 27988 6749 27997 6783
rect 27997 6749 28031 6783
rect 28031 6749 28040 6783
rect 27988 6740 28040 6749
rect 28172 6740 28224 6792
rect 33784 6740 33836 6792
rect 33968 6783 34020 6792
rect 33968 6749 33977 6783
rect 33977 6749 34011 6783
rect 34011 6749 34020 6783
rect 33968 6740 34020 6749
rect 35440 6808 35492 6860
rect 35532 6808 35584 6860
rect 36360 6808 36412 6860
rect 34704 6740 34756 6792
rect 36084 6740 36136 6792
rect 36268 6783 36320 6792
rect 36268 6749 36277 6783
rect 36277 6749 36311 6783
rect 36311 6749 36320 6783
rect 36268 6740 36320 6749
rect 36728 6808 36780 6860
rect 41788 6944 41840 6996
rect 40316 6808 40368 6860
rect 40592 6808 40644 6860
rect 41696 6876 41748 6928
rect 45100 6944 45152 6996
rect 45468 6944 45520 6996
rect 46664 6944 46716 6996
rect 46756 6944 46808 6996
rect 47124 6944 47176 6996
rect 48872 6944 48924 6996
rect 48964 6944 49016 6996
rect 50252 6944 50304 6996
rect 50344 6944 50396 6996
rect 51448 6944 51500 6996
rect 52460 6944 52512 6996
rect 52736 6944 52788 6996
rect 54116 6944 54168 6996
rect 55128 6944 55180 6996
rect 57336 6987 57388 6996
rect 57336 6953 57345 6987
rect 57345 6953 57379 6987
rect 57379 6953 57388 6987
rect 57336 6944 57388 6953
rect 57520 6944 57572 6996
rect 57704 6944 57756 6996
rect 59084 6944 59136 6996
rect 68836 6987 68888 6996
rect 68836 6953 68845 6987
rect 68845 6953 68879 6987
rect 68879 6953 68888 6987
rect 68836 6944 68888 6953
rect 70124 6987 70176 6996
rect 70124 6953 70133 6987
rect 70133 6953 70167 6987
rect 70167 6953 70176 6987
rect 70124 6944 70176 6953
rect 88156 6944 88208 6996
rect 95332 6944 95384 6996
rect 42156 6876 42208 6928
rect 41420 6808 41472 6860
rect 42524 6808 42576 6860
rect 42616 6808 42668 6860
rect 37280 6783 37332 6792
rect 37280 6749 37289 6783
rect 37289 6749 37323 6783
rect 37323 6749 37332 6783
rect 37280 6740 37332 6749
rect 38016 6740 38068 6792
rect 39764 6783 39816 6792
rect 39764 6749 39773 6783
rect 39773 6749 39807 6783
rect 39807 6749 39816 6783
rect 39764 6740 39816 6749
rect 39948 6740 40000 6792
rect 41236 6740 41288 6792
rect 41604 6740 41656 6792
rect 41972 6740 42024 6792
rect 42248 6740 42300 6792
rect 21640 6672 21692 6724
rect 24768 6672 24820 6724
rect 25136 6672 25188 6724
rect 25044 6647 25096 6656
rect 21272 6604 21324 6613
rect 25044 6613 25053 6647
rect 25053 6613 25087 6647
rect 25087 6613 25096 6647
rect 25044 6604 25096 6613
rect 27804 6604 27856 6656
rect 27988 6604 28040 6656
rect 28264 6604 28316 6656
rect 28356 6604 28408 6656
rect 36636 6672 36688 6724
rect 36912 6672 36964 6724
rect 37004 6672 37056 6724
rect 42524 6672 42576 6724
rect 50712 6876 50764 6928
rect 50896 6876 50948 6928
rect 55680 6876 55732 6928
rect 56508 6876 56560 6928
rect 57428 6876 57480 6928
rect 57980 6876 58032 6928
rect 83188 6919 83240 6928
rect 83188 6885 83197 6919
rect 83197 6885 83231 6919
rect 83231 6885 83240 6919
rect 83188 6876 83240 6885
rect 87788 6919 87840 6928
rect 87788 6885 87797 6919
rect 87797 6885 87831 6919
rect 87831 6885 87840 6919
rect 87788 6876 87840 6885
rect 43628 6808 43680 6860
rect 45560 6808 45612 6860
rect 43720 6783 43772 6792
rect 43720 6749 43729 6783
rect 43729 6749 43763 6783
rect 43763 6749 43772 6783
rect 43720 6740 43772 6749
rect 44916 6783 44968 6792
rect 44916 6749 44925 6783
rect 44925 6749 44959 6783
rect 44959 6749 44968 6783
rect 44916 6740 44968 6749
rect 45376 6740 45428 6792
rect 46940 6740 46992 6792
rect 47400 6740 47452 6792
rect 48136 6740 48188 6792
rect 49792 6740 49844 6792
rect 51264 6783 51316 6792
rect 51264 6749 51273 6783
rect 51273 6749 51307 6783
rect 51307 6749 51316 6783
rect 51264 6740 51316 6749
rect 52184 6808 52236 6860
rect 52276 6808 52328 6860
rect 53196 6808 53248 6860
rect 56140 6808 56192 6860
rect 57336 6808 57388 6860
rect 42892 6672 42944 6724
rect 35440 6604 35492 6656
rect 38016 6647 38068 6656
rect 38016 6613 38025 6647
rect 38025 6613 38059 6647
rect 38059 6613 38068 6647
rect 38016 6604 38068 6613
rect 38844 6647 38896 6656
rect 38844 6613 38853 6647
rect 38853 6613 38887 6647
rect 38887 6613 38896 6647
rect 38844 6604 38896 6613
rect 38936 6604 38988 6656
rect 41420 6604 41472 6656
rect 41512 6604 41564 6656
rect 50528 6672 50580 6724
rect 50620 6672 50672 6724
rect 51448 6672 51500 6724
rect 54760 6740 54812 6792
rect 56232 6740 56284 6792
rect 56324 6740 56376 6792
rect 58256 6808 58308 6860
rect 60280 6808 60332 6860
rect 60464 6808 60516 6860
rect 57612 6783 57664 6792
rect 57612 6749 57621 6783
rect 57621 6749 57655 6783
rect 57655 6749 57664 6783
rect 57612 6740 57664 6749
rect 57888 6740 57940 6792
rect 58164 6783 58216 6792
rect 58164 6749 58173 6783
rect 58173 6749 58207 6783
rect 58207 6749 58216 6783
rect 58164 6740 58216 6749
rect 58532 6740 58584 6792
rect 63408 6808 63460 6860
rect 65432 6808 65484 6860
rect 73252 6808 73304 6860
rect 79784 6808 79836 6860
rect 81900 6851 81952 6860
rect 81900 6817 81909 6851
rect 81909 6817 81943 6851
rect 81943 6817 81952 6851
rect 81900 6808 81952 6817
rect 87604 6808 87656 6860
rect 88432 6808 88484 6860
rect 95608 6808 95660 6860
rect 74724 6740 74776 6792
rect 82820 6740 82872 6792
rect 45836 6604 45888 6656
rect 46480 6604 46532 6656
rect 48504 6647 48556 6656
rect 48504 6613 48513 6647
rect 48513 6613 48547 6647
rect 48547 6613 48556 6647
rect 72056 6672 72108 6724
rect 91376 6740 91428 6792
rect 102324 6876 102376 6928
rect 103980 6919 104032 6928
rect 103980 6885 103989 6919
rect 103989 6885 104023 6919
rect 104023 6885 104032 6919
rect 103980 6876 104032 6885
rect 104072 6876 104124 6928
rect 110880 6876 110932 6928
rect 113456 6944 113508 6996
rect 113548 6944 113600 6996
rect 118976 6987 119028 6996
rect 118976 6953 118985 6987
rect 118985 6953 119019 6987
rect 119019 6953 119028 6987
rect 118976 6944 119028 6953
rect 121368 6987 121420 6996
rect 121368 6953 121377 6987
rect 121377 6953 121411 6987
rect 121411 6953 121420 6987
rect 121368 6944 121420 6953
rect 132224 6987 132276 6996
rect 132224 6953 132233 6987
rect 132233 6953 132267 6987
rect 132267 6953 132276 6987
rect 132224 6944 132276 6953
rect 155224 6987 155276 6996
rect 155224 6953 155233 6987
rect 155233 6953 155267 6987
rect 155267 6953 155276 6987
rect 155224 6944 155276 6953
rect 163320 6987 163372 6996
rect 163320 6953 163329 6987
rect 163329 6953 163363 6987
rect 163363 6953 163372 6987
rect 163320 6944 163372 6953
rect 109500 6808 109552 6860
rect 112260 6808 112312 6860
rect 102140 6740 102192 6792
rect 96252 6672 96304 6724
rect 108672 6740 108724 6792
rect 106372 6672 106424 6724
rect 114652 6783 114704 6792
rect 114652 6749 114661 6783
rect 114661 6749 114695 6783
rect 114695 6749 114704 6783
rect 114652 6740 114704 6749
rect 114836 6808 114888 6860
rect 117780 6808 117832 6860
rect 125416 6851 125468 6860
rect 118608 6740 118660 6792
rect 121828 6783 121880 6792
rect 121828 6749 121837 6783
rect 121837 6749 121871 6783
rect 121871 6749 121880 6783
rect 121828 6740 121880 6749
rect 113640 6672 113692 6724
rect 125416 6817 125425 6851
rect 125425 6817 125459 6851
rect 125459 6817 125468 6851
rect 125416 6808 125468 6817
rect 127440 6851 127492 6860
rect 127440 6817 127449 6851
rect 127449 6817 127483 6851
rect 127483 6817 127492 6851
rect 127440 6808 127492 6817
rect 129832 6851 129884 6860
rect 129832 6817 129841 6851
rect 129841 6817 129875 6851
rect 129875 6817 129884 6851
rect 129832 6808 129884 6817
rect 136180 6919 136232 6928
rect 136180 6885 136189 6919
rect 136189 6885 136223 6919
rect 136223 6885 136232 6919
rect 136180 6876 136232 6885
rect 142896 6876 142948 6928
rect 153752 6876 153804 6928
rect 162400 6919 162452 6928
rect 162400 6885 162409 6919
rect 162409 6885 162443 6919
rect 162443 6885 162452 6919
rect 162400 6876 162452 6885
rect 164884 6876 164936 6928
rect 141792 6851 141844 6860
rect 128544 6783 128596 6792
rect 128544 6749 128553 6783
rect 128553 6749 128587 6783
rect 128587 6749 128596 6783
rect 128544 6740 128596 6749
rect 123024 6672 123076 6724
rect 141792 6817 141801 6851
rect 141801 6817 141835 6851
rect 141835 6817 141844 6851
rect 141792 6808 141844 6817
rect 146944 6808 146996 6860
rect 148048 6808 148100 6860
rect 151820 6851 151872 6860
rect 151820 6817 151829 6851
rect 151829 6817 151863 6851
rect 151863 6817 151872 6851
rect 151820 6808 151872 6817
rect 156144 6808 156196 6860
rect 159916 6808 159968 6860
rect 163504 6851 163556 6860
rect 163504 6817 163513 6851
rect 163513 6817 163547 6851
rect 163547 6817 163556 6851
rect 163504 6808 163556 6817
rect 131120 6783 131172 6792
rect 131120 6749 131129 6783
rect 131129 6749 131163 6783
rect 131163 6749 131172 6783
rect 131120 6740 131172 6749
rect 134892 6783 134944 6792
rect 134892 6749 134901 6783
rect 134901 6749 134935 6783
rect 134935 6749 134944 6783
rect 134892 6740 134944 6749
rect 135996 6783 136048 6792
rect 135996 6749 136005 6783
rect 136005 6749 136039 6783
rect 136039 6749 136048 6783
rect 135996 6740 136048 6749
rect 142896 6783 142948 6792
rect 142896 6749 142905 6783
rect 142905 6749 142939 6783
rect 142939 6749 142948 6783
rect 142896 6740 142948 6749
rect 150808 6740 150860 6792
rect 152096 6783 152148 6792
rect 152096 6749 152105 6783
rect 152105 6749 152139 6783
rect 152139 6749 152148 6783
rect 152096 6740 152148 6749
rect 153016 6783 153068 6792
rect 153016 6749 153025 6783
rect 153025 6749 153059 6783
rect 153059 6749 153068 6783
rect 153016 6740 153068 6749
rect 153752 6740 153804 6792
rect 161480 6740 161532 6792
rect 162400 6672 162452 6724
rect 164240 6740 164292 6792
rect 48504 6604 48556 6613
rect 52368 6604 52420 6656
rect 56324 6604 56376 6656
rect 56416 6647 56468 6656
rect 56416 6613 56425 6647
rect 56425 6613 56459 6647
rect 56459 6613 56468 6647
rect 56416 6604 56468 6613
rect 56968 6604 57020 6656
rect 59452 6604 59504 6656
rect 59820 6647 59872 6656
rect 59820 6613 59829 6647
rect 59829 6613 59863 6647
rect 59863 6613 59872 6647
rect 59820 6604 59872 6613
rect 64512 6604 64564 6656
rect 69940 6604 69992 6656
rect 70124 6604 70176 6656
rect 79140 6604 79192 6656
rect 81348 6604 81400 6656
rect 81992 6604 82044 6656
rect 88524 6604 88576 6656
rect 100576 6604 100628 6656
rect 103060 6604 103112 6656
rect 108948 6604 109000 6656
rect 113456 6604 113508 6656
rect 115756 6647 115808 6656
rect 115756 6613 115765 6647
rect 115765 6613 115799 6647
rect 115799 6613 115808 6647
rect 115756 6604 115808 6613
rect 117136 6647 117188 6656
rect 117136 6613 117145 6647
rect 117145 6613 117179 6647
rect 117179 6613 117188 6647
rect 117136 6604 117188 6613
rect 120632 6647 120684 6656
rect 120632 6613 120641 6647
rect 120641 6613 120675 6647
rect 120675 6613 120684 6647
rect 120632 6604 120684 6613
rect 124220 6604 124272 6656
rect 126980 6604 127032 6656
rect 133236 6604 133288 6656
rect 144368 6604 144420 6656
rect 145196 6604 145248 6656
rect 149336 6647 149388 6656
rect 149336 6613 149345 6647
rect 149345 6613 149379 6647
rect 149379 6613 149388 6647
rect 149336 6604 149388 6613
rect 155500 6647 155552 6656
rect 155500 6613 155509 6647
rect 155509 6613 155543 6647
rect 155543 6613 155552 6647
rect 155500 6604 155552 6613
rect 155868 6604 155920 6656
rect 164516 6604 164568 6656
rect 164976 6604 165028 6656
rect 56667 6502 56719 6554
rect 56731 6502 56783 6554
rect 56795 6502 56847 6554
rect 56859 6502 56911 6554
rect 113088 6502 113140 6554
rect 113152 6502 113204 6554
rect 113216 6502 113268 6554
rect 113280 6502 113332 6554
rect 4252 6443 4304 6452
rect 4252 6409 4261 6443
rect 4261 6409 4295 6443
rect 4295 6409 4304 6443
rect 4252 6400 4304 6409
rect 21916 6400 21968 6452
rect 3700 6332 3752 6384
rect 8208 6332 8260 6384
rect 10692 6332 10744 6384
rect 9220 6264 9272 6316
rect 15108 6264 15160 6316
rect 21088 6307 21140 6316
rect 3240 6239 3292 6248
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 5816 6196 5868 6248
rect 8024 6196 8076 6248
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 15936 6196 15988 6248
rect 19524 6239 19576 6248
rect 19524 6205 19533 6239
rect 19533 6205 19567 6239
rect 19567 6205 19576 6239
rect 19524 6196 19576 6205
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 22008 6264 22060 6316
rect 24952 6264 25004 6316
rect 22652 6196 22704 6248
rect 25596 6196 25648 6248
rect 26240 6264 26292 6316
rect 26516 6307 26568 6316
rect 26516 6273 26525 6307
rect 26525 6273 26559 6307
rect 26559 6273 26568 6307
rect 26516 6264 26568 6273
rect 27804 6332 27856 6384
rect 31116 6400 31168 6452
rect 36176 6400 36228 6452
rect 36268 6400 36320 6452
rect 36636 6400 36688 6452
rect 39580 6400 39632 6452
rect 39764 6443 39816 6452
rect 39764 6409 39773 6443
rect 39773 6409 39807 6443
rect 39807 6409 39816 6443
rect 39764 6400 39816 6409
rect 39856 6400 39908 6452
rect 40868 6400 40920 6452
rect 41144 6400 41196 6452
rect 43536 6400 43588 6452
rect 43720 6400 43772 6452
rect 47676 6400 47728 6452
rect 47768 6400 47820 6452
rect 50712 6400 50764 6452
rect 50804 6400 50856 6452
rect 51264 6400 51316 6452
rect 51448 6400 51500 6452
rect 52368 6400 52420 6452
rect 52736 6400 52788 6452
rect 54024 6400 54076 6452
rect 57612 6400 57664 6452
rect 60280 6400 60332 6452
rect 81900 6400 81952 6452
rect 87788 6400 87840 6452
rect 89536 6400 89588 6452
rect 98000 6400 98052 6452
rect 104440 6400 104492 6452
rect 104716 6400 104768 6452
rect 29828 6307 29880 6316
rect 29828 6273 29837 6307
rect 29837 6273 29871 6307
rect 29871 6273 29880 6307
rect 29828 6264 29880 6273
rect 30380 6264 30432 6316
rect 30840 6264 30892 6316
rect 34704 6264 34756 6316
rect 35072 6264 35124 6316
rect 31116 6196 31168 6248
rect 33692 6196 33744 6248
rect 35992 6264 36044 6316
rect 36084 6264 36136 6316
rect 37280 6264 37332 6316
rect 37464 6332 37516 6384
rect 41328 6332 41380 6384
rect 41420 6332 41472 6384
rect 42984 6332 43036 6384
rect 43168 6332 43220 6384
rect 37832 6264 37884 6316
rect 38936 6264 38988 6316
rect 41144 6264 41196 6316
rect 4896 6128 4948 6180
rect 3424 6060 3476 6112
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 24308 6060 24360 6112
rect 29092 6060 29144 6112
rect 29276 6128 29328 6180
rect 39488 6196 39540 6248
rect 41604 6264 41656 6316
rect 41696 6307 41748 6316
rect 41696 6273 41705 6307
rect 41705 6273 41739 6307
rect 41739 6273 41748 6307
rect 41696 6264 41748 6273
rect 41880 6264 41932 6316
rect 42156 6264 42208 6316
rect 42800 6264 42852 6316
rect 43444 6332 43496 6384
rect 52276 6332 52328 6384
rect 54668 6332 54720 6384
rect 55496 6375 55548 6384
rect 55496 6341 55505 6375
rect 55505 6341 55539 6375
rect 55539 6341 55548 6375
rect 55496 6332 55548 6341
rect 47216 6307 47268 6316
rect 41328 6196 41380 6248
rect 43536 6196 43588 6248
rect 45468 6196 45520 6248
rect 45652 6239 45704 6248
rect 45652 6205 45661 6239
rect 45661 6205 45695 6239
rect 45695 6205 45704 6239
rect 45652 6196 45704 6205
rect 45836 6196 45888 6248
rect 45928 6196 45980 6248
rect 46480 6196 46532 6248
rect 47216 6273 47225 6307
rect 47225 6273 47259 6307
rect 47259 6273 47268 6307
rect 47216 6264 47268 6273
rect 47308 6264 47360 6316
rect 50160 6264 50212 6316
rect 50712 6264 50764 6316
rect 46848 6196 46900 6248
rect 51172 6264 51224 6316
rect 51632 6264 51684 6316
rect 52460 6264 52512 6316
rect 52644 6307 52696 6316
rect 52644 6273 52653 6307
rect 52653 6273 52687 6307
rect 52687 6273 52696 6307
rect 52644 6264 52696 6273
rect 58532 6332 58584 6384
rect 43352 6128 43404 6180
rect 48044 6128 48096 6180
rect 48136 6128 48188 6180
rect 50712 6128 50764 6180
rect 51448 6128 51500 6180
rect 51908 6196 51960 6248
rect 52368 6196 52420 6248
rect 56416 6264 56468 6316
rect 57428 6264 57480 6316
rect 55036 6196 55088 6248
rect 59268 6307 59320 6316
rect 59268 6273 59277 6307
rect 59277 6273 59311 6307
rect 59311 6273 59320 6307
rect 59268 6264 59320 6273
rect 59452 6332 59504 6384
rect 89996 6332 90048 6384
rect 92020 6332 92072 6384
rect 104348 6332 104400 6384
rect 104624 6332 104676 6384
rect 106280 6332 106332 6384
rect 63868 6264 63920 6316
rect 64512 6307 64564 6316
rect 64512 6273 64521 6307
rect 64521 6273 64555 6307
rect 64555 6273 64564 6307
rect 64512 6264 64564 6273
rect 66076 6307 66128 6316
rect 66076 6273 66085 6307
rect 66085 6273 66119 6307
rect 66119 6273 66128 6307
rect 66076 6264 66128 6273
rect 69940 6307 69992 6316
rect 69940 6273 69949 6307
rect 69949 6273 69983 6307
rect 69983 6273 69992 6307
rect 69940 6264 69992 6273
rect 71780 6264 71832 6316
rect 91836 6307 91888 6316
rect 65524 6239 65576 6248
rect 55864 6128 55916 6180
rect 57612 6128 57664 6180
rect 57796 6128 57848 6180
rect 65524 6205 65533 6239
rect 65533 6205 65567 6239
rect 65567 6205 65576 6239
rect 65524 6196 65576 6205
rect 70952 6239 71004 6248
rect 70952 6205 70961 6239
rect 70961 6205 70995 6239
rect 70995 6205 71004 6239
rect 70952 6196 71004 6205
rect 87512 6239 87564 6248
rect 87512 6205 87521 6239
rect 87521 6205 87555 6239
rect 87555 6205 87564 6239
rect 87512 6196 87564 6205
rect 90272 6239 90324 6248
rect 90272 6205 90281 6239
rect 90281 6205 90315 6239
rect 90315 6205 90324 6239
rect 90272 6196 90324 6205
rect 91192 6196 91244 6248
rect 91836 6273 91845 6307
rect 91845 6273 91879 6307
rect 91879 6273 91888 6307
rect 91836 6264 91888 6273
rect 97264 6264 97316 6316
rect 36084 6103 36136 6112
rect 36084 6069 36093 6103
rect 36093 6069 36127 6103
rect 36127 6069 36136 6103
rect 36084 6060 36136 6069
rect 36176 6060 36228 6112
rect 51264 6060 51316 6112
rect 51356 6060 51408 6112
rect 75736 6128 75788 6180
rect 101680 6196 101732 6248
rect 103336 6196 103388 6248
rect 104808 6196 104860 6248
rect 106280 6196 106332 6248
rect 103520 6128 103572 6180
rect 107476 6196 107528 6248
rect 130016 6332 130068 6384
rect 134892 6332 134944 6384
rect 141792 6332 141844 6384
rect 142804 6375 142856 6384
rect 142804 6341 142813 6375
rect 142813 6341 142847 6375
rect 142847 6341 142856 6375
rect 142804 6332 142856 6341
rect 150808 6375 150860 6384
rect 150808 6341 150817 6375
rect 150817 6341 150851 6375
rect 150851 6341 150860 6375
rect 150808 6332 150860 6341
rect 153016 6332 153068 6384
rect 157248 6332 157300 6384
rect 159456 6400 159508 6452
rect 161480 6443 161532 6452
rect 161480 6409 161489 6443
rect 161489 6409 161523 6443
rect 161523 6409 161532 6443
rect 161480 6400 161532 6409
rect 163504 6400 163556 6452
rect 164792 6332 164844 6384
rect 108304 6196 108356 6248
rect 113456 6196 113508 6248
rect 115756 6196 115808 6248
rect 121460 6196 121512 6248
rect 123024 6264 123076 6316
rect 145748 6264 145800 6316
rect 122840 6196 122892 6248
rect 128912 6196 128964 6248
rect 148416 6239 148468 6248
rect 148416 6205 148425 6239
rect 148425 6205 148459 6239
rect 148459 6205 148468 6239
rect 148416 6196 148468 6205
rect 150072 6264 150124 6316
rect 153476 6264 153528 6316
rect 154856 6307 154908 6316
rect 154856 6273 154865 6307
rect 154865 6273 154899 6307
rect 154899 6273 154908 6307
rect 154856 6264 154908 6273
rect 164976 6307 165028 6316
rect 164976 6273 164985 6307
rect 164985 6273 165019 6307
rect 165019 6273 165028 6307
rect 164976 6264 165028 6273
rect 153384 6239 153436 6248
rect 153384 6205 153393 6239
rect 153393 6205 153427 6239
rect 153427 6205 153436 6239
rect 153384 6196 153436 6205
rect 154580 6196 154632 6248
rect 158260 6239 158312 6248
rect 158260 6205 158269 6239
rect 158269 6205 158303 6239
rect 158303 6205 158312 6239
rect 158260 6196 158312 6205
rect 163504 6196 163556 6248
rect 114836 6128 114888 6180
rect 75828 6060 75880 6112
rect 28456 5958 28508 6010
rect 28520 5958 28572 6010
rect 28584 5958 28636 6010
rect 28648 5958 28700 6010
rect 84878 5958 84930 6010
rect 84942 5958 84994 6010
rect 85006 5958 85058 6010
rect 85070 5958 85122 6010
rect 9220 5899 9272 5908
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 12348 5899 12400 5908
rect 12348 5865 12357 5899
rect 12357 5865 12391 5899
rect 12391 5865 12400 5899
rect 12348 5856 12400 5865
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 19524 5899 19576 5908
rect 3792 5788 3844 5840
rect 3424 5763 3476 5772
rect 3424 5729 3433 5763
rect 3433 5729 3467 5763
rect 3467 5729 3476 5763
rect 3424 5720 3476 5729
rect 4160 5720 4212 5772
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 5356 5627 5408 5636
rect 5356 5593 5365 5627
rect 5365 5593 5399 5627
rect 5399 5593 5408 5627
rect 5356 5584 5408 5593
rect 14740 5788 14792 5840
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 19524 5865 19533 5899
rect 19533 5865 19567 5899
rect 19567 5865 19576 5899
rect 19524 5856 19576 5865
rect 21088 5856 21140 5908
rect 24952 5856 25004 5908
rect 25596 5899 25648 5908
rect 25596 5865 25605 5899
rect 25605 5865 25639 5899
rect 25639 5865 25648 5899
rect 25596 5856 25648 5865
rect 26792 5856 26844 5908
rect 28816 5856 28868 5908
rect 30380 5856 30432 5908
rect 21180 5788 21232 5840
rect 12348 5652 12400 5704
rect 21364 5720 21416 5772
rect 22008 5652 22060 5704
rect 17132 5584 17184 5636
rect 24032 5695 24084 5704
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 3700 5516 3752 5568
rect 5724 5516 5776 5568
rect 8024 5559 8076 5568
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 21180 5516 21232 5568
rect 24860 5584 24912 5636
rect 26516 5788 26568 5840
rect 33692 5899 33744 5908
rect 33692 5865 33701 5899
rect 33701 5865 33735 5899
rect 33735 5865 33744 5899
rect 33692 5856 33744 5865
rect 35348 5856 35400 5908
rect 36084 5856 36136 5908
rect 37924 5856 37976 5908
rect 38016 5856 38068 5908
rect 42708 5856 42760 5908
rect 28080 5720 28132 5772
rect 26424 5695 26476 5704
rect 26424 5661 26433 5695
rect 26433 5661 26467 5695
rect 26467 5661 26476 5695
rect 26424 5652 26476 5661
rect 27988 5652 28040 5704
rect 35072 5788 35124 5840
rect 35256 5788 35308 5840
rect 42984 5831 43036 5840
rect 42984 5797 42993 5831
rect 42993 5797 43027 5831
rect 43027 5797 43036 5831
rect 42984 5788 43036 5797
rect 44364 5856 44416 5908
rect 45928 5856 45980 5908
rect 48596 5856 48648 5908
rect 49792 5856 49844 5908
rect 51080 5856 51132 5908
rect 51264 5856 51316 5908
rect 56968 5856 57020 5908
rect 57244 5856 57296 5908
rect 57428 5899 57480 5908
rect 57428 5865 57437 5899
rect 57437 5865 57471 5899
rect 57471 5865 57480 5899
rect 57428 5856 57480 5865
rect 59728 5856 59780 5908
rect 64512 5899 64564 5908
rect 64512 5865 64521 5899
rect 64521 5865 64555 5899
rect 64555 5865 64564 5899
rect 64512 5856 64564 5865
rect 69940 5899 69992 5908
rect 69940 5865 69949 5899
rect 69949 5865 69983 5899
rect 69983 5865 69992 5899
rect 69940 5856 69992 5865
rect 90272 5899 90324 5908
rect 90272 5865 90281 5899
rect 90281 5865 90315 5899
rect 90315 5865 90324 5899
rect 90272 5856 90324 5865
rect 34980 5720 35032 5772
rect 35348 5720 35400 5772
rect 36636 5720 36688 5772
rect 37096 5720 37148 5772
rect 37280 5720 37332 5772
rect 37832 5720 37884 5772
rect 37924 5720 37976 5772
rect 40500 5720 40552 5772
rect 41696 5720 41748 5772
rect 34152 5695 34204 5704
rect 34152 5661 34161 5695
rect 34161 5661 34195 5695
rect 34195 5661 34204 5695
rect 34152 5652 34204 5661
rect 34244 5584 34296 5636
rect 34796 5584 34848 5636
rect 35900 5584 35952 5636
rect 36268 5652 36320 5704
rect 39856 5652 39908 5704
rect 40316 5652 40368 5704
rect 47492 5720 47544 5772
rect 47860 5720 47912 5772
rect 51172 5763 51224 5772
rect 42156 5652 42208 5704
rect 44548 5652 44600 5704
rect 45284 5627 45336 5636
rect 45284 5593 45293 5627
rect 45293 5593 45327 5627
rect 45327 5593 45336 5627
rect 45284 5584 45336 5593
rect 46296 5652 46348 5704
rect 50068 5652 50120 5704
rect 51172 5729 51181 5763
rect 51181 5729 51215 5763
rect 51215 5729 51224 5763
rect 51172 5720 51224 5729
rect 52644 5763 52696 5772
rect 52644 5729 52653 5763
rect 52653 5729 52687 5763
rect 52687 5729 52696 5763
rect 52644 5720 52696 5729
rect 52736 5720 52788 5772
rect 54668 5720 54720 5772
rect 55128 5695 55180 5704
rect 47400 5584 47452 5636
rect 47492 5584 47544 5636
rect 54852 5584 54904 5636
rect 55128 5661 55137 5695
rect 55137 5661 55171 5695
rect 55171 5661 55180 5695
rect 55128 5652 55180 5661
rect 65432 5788 65484 5840
rect 100944 6060 100996 6112
rect 107752 6060 107804 6112
rect 117688 6060 117740 6112
rect 124128 6060 124180 6112
rect 148876 6128 148928 6180
rect 150256 6128 150308 6180
rect 157432 6128 157484 6180
rect 164884 6128 164936 6180
rect 165160 6171 165212 6180
rect 165160 6137 165169 6171
rect 165169 6137 165203 6171
rect 165203 6137 165212 6171
rect 165160 6128 165212 6137
rect 156328 6103 156380 6112
rect 156328 6069 156337 6103
rect 156337 6069 156371 6103
rect 156371 6069 156380 6103
rect 156328 6060 156380 6069
rect 163596 6103 163648 6112
rect 163596 6069 163605 6103
rect 163605 6069 163639 6103
rect 163639 6069 163648 6103
rect 163596 6060 163648 6069
rect 93216 5924 93268 5976
rect 141299 5958 141351 6010
rect 141363 5958 141415 6010
rect 141427 5958 141479 6010
rect 141491 5958 141543 6010
rect 116124 5856 116176 5908
rect 116216 5856 116268 5908
rect 128912 5899 128964 5908
rect 55496 5584 55548 5636
rect 56600 5652 56652 5704
rect 57520 5652 57572 5704
rect 59820 5720 59872 5772
rect 66812 5720 66864 5772
rect 87512 5763 87564 5772
rect 87512 5729 87521 5763
rect 87521 5729 87555 5763
rect 87555 5729 87564 5763
rect 87512 5720 87564 5729
rect 88708 5763 88760 5772
rect 88708 5729 88717 5763
rect 88717 5729 88751 5763
rect 88751 5729 88760 5763
rect 88708 5720 88760 5729
rect 63316 5652 63368 5704
rect 106648 5788 106700 5840
rect 106740 5788 106792 5840
rect 107660 5720 107712 5772
rect 104440 5652 104492 5704
rect 112720 5720 112772 5772
rect 118332 5720 118384 5772
rect 128912 5865 128921 5899
rect 128921 5865 128955 5899
rect 128955 5865 128964 5899
rect 128912 5856 128964 5865
rect 148416 5899 148468 5908
rect 148416 5865 148425 5899
rect 148425 5865 148459 5899
rect 148459 5865 148468 5899
rect 148416 5856 148468 5865
rect 153384 5856 153436 5908
rect 130016 5763 130068 5772
rect 130016 5729 130025 5763
rect 130025 5729 130059 5763
rect 130059 5729 130068 5763
rect 130016 5720 130068 5729
rect 148876 5788 148928 5840
rect 157432 5856 157484 5908
rect 157524 5856 157576 5908
rect 159272 5899 159324 5908
rect 159272 5865 159281 5899
rect 159281 5865 159315 5899
rect 159315 5865 159324 5899
rect 159272 5856 159324 5865
rect 163504 5899 163556 5908
rect 163504 5865 163513 5899
rect 163513 5865 163547 5899
rect 163547 5865 163556 5899
rect 163504 5856 163556 5865
rect 154672 5788 154724 5840
rect 153844 5720 153896 5772
rect 156420 5720 156472 5772
rect 163596 5763 163648 5772
rect 163596 5729 163605 5763
rect 163605 5729 163639 5763
rect 163639 5729 163648 5763
rect 163596 5720 163648 5729
rect 164700 5763 164752 5772
rect 164700 5729 164709 5763
rect 164709 5729 164743 5763
rect 164743 5729 164752 5763
rect 164700 5720 164752 5729
rect 26516 5516 26568 5568
rect 30380 5516 30432 5568
rect 36452 5516 36504 5568
rect 38200 5516 38252 5568
rect 41880 5516 41932 5568
rect 41972 5516 42024 5568
rect 42340 5516 42392 5568
rect 42432 5516 42484 5568
rect 46848 5516 46900 5568
rect 47216 5516 47268 5568
rect 55036 5516 55088 5568
rect 55128 5516 55180 5568
rect 55956 5516 56008 5568
rect 56140 5516 56192 5568
rect 58348 5584 58400 5636
rect 69112 5584 69164 5636
rect 91284 5584 91336 5636
rect 58992 5516 59044 5568
rect 59268 5516 59320 5568
rect 64420 5516 64472 5568
rect 66076 5516 66128 5568
rect 71044 5516 71096 5568
rect 71780 5516 71832 5568
rect 90732 5559 90784 5568
rect 90732 5525 90741 5559
rect 90741 5525 90775 5559
rect 90775 5525 90784 5559
rect 90732 5516 90784 5525
rect 91836 5516 91888 5568
rect 101404 5584 101456 5636
rect 104072 5584 104124 5636
rect 99104 5516 99156 5568
rect 56667 5414 56719 5466
rect 56731 5414 56783 5466
rect 56795 5414 56847 5466
rect 56859 5414 56911 5466
rect 8024 5312 8076 5364
rect 6460 5244 6512 5296
rect 43536 5312 43588 5364
rect 43628 5312 43680 5364
rect 45652 5312 45704 5364
rect 45836 5312 45888 5364
rect 46112 5312 46164 5364
rect 51080 5312 51132 5364
rect 51356 5312 51408 5364
rect 57244 5312 57296 5364
rect 63868 5312 63920 5364
rect 67088 5312 67140 5364
rect 92940 5312 92992 5364
rect 99104 5380 99156 5432
rect 102232 5516 102284 5568
rect 108764 5584 108816 5636
rect 104532 5516 104584 5568
rect 121460 5652 121512 5704
rect 121828 5695 121880 5704
rect 121828 5661 121837 5695
rect 121837 5661 121871 5695
rect 121871 5661 121880 5695
rect 121828 5652 121880 5661
rect 122840 5695 122892 5704
rect 122840 5661 122849 5695
rect 122849 5661 122883 5695
rect 122883 5661 122892 5695
rect 122840 5652 122892 5661
rect 123116 5584 123168 5636
rect 110972 5559 111024 5568
rect 110972 5525 110981 5559
rect 110981 5525 111015 5559
rect 111015 5525 111024 5559
rect 110972 5516 111024 5525
rect 114652 5516 114704 5568
rect 114836 5516 114888 5568
rect 116860 5516 116912 5568
rect 123024 5516 123076 5568
rect 123760 5516 123812 5568
rect 153476 5652 153528 5704
rect 126060 5516 126112 5568
rect 130936 5559 130988 5568
rect 130936 5525 130945 5559
rect 130945 5525 130979 5559
rect 130979 5525 130988 5559
rect 130936 5516 130988 5525
rect 150072 5559 150124 5568
rect 150072 5525 150081 5559
rect 150081 5525 150115 5559
rect 150115 5525 150124 5559
rect 150072 5516 150124 5525
rect 152004 5559 152056 5568
rect 152004 5525 152013 5559
rect 152013 5525 152047 5559
rect 152047 5525 152056 5559
rect 152004 5516 152056 5525
rect 154580 5516 154632 5568
rect 154856 5559 154908 5568
rect 154856 5525 154865 5559
rect 154865 5525 154899 5559
rect 154899 5525 154908 5559
rect 154856 5516 154908 5525
rect 156328 5652 156380 5704
rect 157340 5695 157392 5704
rect 157340 5661 157349 5695
rect 157349 5661 157383 5695
rect 157383 5661 157392 5695
rect 157340 5652 157392 5661
rect 158076 5652 158128 5704
rect 159180 5695 159232 5704
rect 159180 5661 159189 5695
rect 159189 5661 159223 5695
rect 159223 5661 159232 5695
rect 159180 5652 159232 5661
rect 165068 5695 165120 5704
rect 165068 5661 165077 5695
rect 165077 5661 165111 5695
rect 165111 5661 165120 5695
rect 165068 5652 165120 5661
rect 155776 5516 155828 5568
rect 164976 5516 165028 5568
rect 18880 5287 18932 5296
rect 3240 5176 3292 5228
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 16028 5176 16080 5228
rect 18052 5176 18104 5228
rect 18880 5253 18889 5287
rect 18889 5253 18923 5287
rect 18923 5253 18932 5287
rect 18880 5244 18932 5253
rect 21272 5244 21324 5296
rect 23296 5244 23348 5296
rect 21456 5219 21508 5228
rect 21456 5185 21465 5219
rect 21465 5185 21499 5219
rect 21499 5185 21508 5219
rect 21456 5176 21508 5185
rect 26424 5244 26476 5296
rect 34428 5244 34480 5296
rect 46020 5244 46072 5296
rect 4436 5151 4488 5160
rect 4436 5117 4445 5151
rect 4445 5117 4479 5151
rect 4479 5117 4488 5151
rect 4436 5108 4488 5117
rect 15016 5108 15068 5160
rect 20720 5108 20772 5160
rect 22560 5108 22612 5160
rect 8208 5040 8260 5092
rect 29184 5176 29236 5228
rect 29276 5176 29328 5228
rect 25320 5151 25372 5160
rect 25320 5117 25329 5151
rect 25329 5117 25363 5151
rect 25363 5117 25372 5151
rect 25320 5108 25372 5117
rect 29644 5108 29696 5160
rect 34060 5108 34112 5160
rect 34888 5176 34940 5228
rect 34980 5176 35032 5228
rect 40776 5176 40828 5228
rect 40868 5176 40920 5228
rect 41328 5176 41380 5228
rect 41420 5176 41472 5228
rect 43076 5176 43128 5228
rect 46388 5219 46440 5228
rect 46388 5185 46397 5219
rect 46397 5185 46431 5219
rect 46431 5185 46440 5219
rect 46388 5176 46440 5185
rect 46664 5244 46716 5296
rect 67640 5244 67692 5296
rect 48044 5176 48096 5228
rect 48504 5176 48556 5228
rect 49700 5176 49752 5228
rect 52828 5176 52880 5228
rect 53656 5176 53708 5228
rect 55404 5176 55456 5228
rect 55772 5176 55824 5228
rect 57060 5176 57112 5228
rect 57336 5176 57388 5228
rect 59544 5176 59596 5228
rect 63316 5176 63368 5228
rect 66536 5176 66588 5228
rect 91100 5176 91152 5228
rect 92296 5176 92348 5228
rect 43352 5108 43404 5160
rect 46204 5108 46256 5160
rect 49332 5108 49384 5160
rect 62672 5108 62724 5160
rect 63408 5108 63460 5160
rect 70492 5108 70544 5160
rect 86776 5151 86828 5160
rect 86776 5117 86785 5151
rect 86785 5117 86819 5151
rect 86819 5117 86828 5151
rect 86776 5108 86828 5117
rect 87788 5151 87840 5160
rect 87788 5117 87797 5151
rect 87797 5117 87831 5151
rect 87831 5117 87840 5151
rect 87788 5108 87840 5117
rect 89444 5108 89496 5160
rect 90824 5151 90876 5160
rect 90824 5117 90833 5151
rect 90833 5117 90867 5151
rect 90867 5117 90876 5151
rect 90824 5108 90876 5117
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 23388 4972 23440 5024
rect 31576 4972 31628 5024
rect 31668 4972 31720 5024
rect 35072 4972 35124 5024
rect 36452 4972 36504 5024
rect 36544 4972 36596 5024
rect 43352 4972 43404 5024
rect 43536 4972 43588 5024
rect 50988 4972 51040 5024
rect 51264 4972 51316 5024
rect 53748 4972 53800 5024
rect 56048 4972 56100 5024
rect 56324 4972 56376 5024
rect 57060 5040 57112 5092
rect 57980 5040 58032 5092
rect 58992 5040 59044 5092
rect 65064 5040 65116 5092
rect 90364 5040 90416 5092
rect 113088 5414 113140 5466
rect 113152 5414 113204 5466
rect 113216 5414 113268 5466
rect 113280 5414 113332 5466
rect 102140 5312 102192 5364
rect 100760 5176 100812 5228
rect 106464 5312 106516 5364
rect 121920 5312 121972 5364
rect 127624 5312 127676 5364
rect 145840 5355 145892 5364
rect 145840 5321 145849 5355
rect 145849 5321 145883 5355
rect 145883 5321 145892 5355
rect 145840 5312 145892 5321
rect 166908 5312 166960 5364
rect 109776 5244 109828 5296
rect 104440 5176 104492 5228
rect 105636 5176 105688 5228
rect 105820 5219 105872 5228
rect 105820 5185 105829 5219
rect 105829 5185 105863 5219
rect 105863 5185 105872 5219
rect 105820 5176 105872 5185
rect 106188 5176 106240 5228
rect 107936 5176 107988 5228
rect 103060 5151 103112 5160
rect 103060 5117 103069 5151
rect 103069 5117 103103 5151
rect 103103 5117 103112 5151
rect 103060 5108 103112 5117
rect 104072 5151 104124 5160
rect 104072 5117 104081 5151
rect 104081 5117 104115 5151
rect 104115 5117 104124 5151
rect 104072 5108 104124 5117
rect 106004 5108 106056 5160
rect 112904 5244 112956 5296
rect 110236 5219 110288 5228
rect 110236 5185 110245 5219
rect 110245 5185 110279 5219
rect 110279 5185 110288 5219
rect 110236 5176 110288 5185
rect 115388 5176 115440 5228
rect 117136 5176 117188 5228
rect 124680 5176 124732 5228
rect 128360 5176 128412 5228
rect 146300 5176 146352 5228
rect 152004 5176 152056 5228
rect 152924 5219 152976 5228
rect 152924 5185 152933 5219
rect 152933 5185 152967 5219
rect 152967 5185 152976 5219
rect 152924 5176 152976 5185
rect 154856 5176 154908 5228
rect 156604 5219 156656 5228
rect 156604 5185 156613 5219
rect 156613 5185 156647 5219
rect 156647 5185 156656 5219
rect 156604 5176 156656 5185
rect 158260 5219 158312 5228
rect 158260 5185 158269 5219
rect 158269 5185 158303 5219
rect 158303 5185 158312 5219
rect 158260 5176 158312 5185
rect 159548 5219 159600 5228
rect 159548 5185 159557 5219
rect 159557 5185 159591 5219
rect 159591 5185 159600 5219
rect 159548 5176 159600 5185
rect 164700 5176 164752 5228
rect 110328 5151 110380 5160
rect 110328 5117 110337 5151
rect 110337 5117 110371 5151
rect 110371 5117 110380 5151
rect 110328 5108 110380 5117
rect 153936 5151 153988 5160
rect 153936 5117 153945 5151
rect 153945 5117 153979 5151
rect 153979 5117 153988 5151
rect 153936 5108 153988 5117
rect 155316 5151 155368 5160
rect 155316 5117 155325 5151
rect 155325 5117 155359 5151
rect 155359 5117 155368 5151
rect 155316 5108 155368 5117
rect 156512 5151 156564 5160
rect 156512 5117 156521 5151
rect 156521 5117 156555 5151
rect 156555 5117 156564 5151
rect 156512 5108 156564 5117
rect 158812 5108 158864 5160
rect 103796 5040 103848 5092
rect 106096 5040 106148 5092
rect 110420 5040 110472 5092
rect 115296 5040 115348 5092
rect 62488 4972 62540 5024
rect 64420 4972 64472 5024
rect 70676 4972 70728 5024
rect 91836 5015 91888 5024
rect 91836 4981 91845 5015
rect 91845 4981 91879 5015
rect 91879 4981 91888 5015
rect 91836 4972 91888 4981
rect 106188 4972 106240 5024
rect 116216 4972 116268 5024
rect 28456 4870 28508 4922
rect 28520 4870 28572 4922
rect 28584 4870 28636 4922
rect 28648 4870 28700 4922
rect 84878 4870 84930 4922
rect 84942 4870 84994 4922
rect 85006 4870 85058 4922
rect 85070 4870 85122 4922
rect 141299 4870 141351 4922
rect 141363 4870 141415 4922
rect 141427 4870 141479 4922
rect 141491 4870 141543 4922
rect 3240 4768 3292 4820
rect 3700 4768 3752 4820
rect 7380 4768 7432 4820
rect 16028 4811 16080 4820
rect 16028 4777 16037 4811
rect 16037 4777 16071 4811
rect 16071 4777 16080 4811
rect 16028 4768 16080 4777
rect 4160 4632 4212 4684
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 17408 4768 17460 4820
rect 21456 4768 21508 4820
rect 22560 4811 22612 4820
rect 21364 4632 21416 4684
rect 22560 4777 22569 4811
rect 22569 4777 22603 4811
rect 22603 4777 22612 4811
rect 22560 4768 22612 4777
rect 25320 4768 25372 4820
rect 27896 4768 27948 4820
rect 29736 4768 29788 4820
rect 36544 4768 36596 4820
rect 26148 4700 26200 4752
rect 30380 4700 30432 4752
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 5908 4539 5960 4548
rect 5908 4505 5917 4539
rect 5917 4505 5951 4539
rect 5951 4505 5960 4539
rect 5908 4496 5960 4505
rect 12256 4496 12308 4548
rect 3884 4428 3936 4480
rect 5816 4428 5868 4480
rect 8484 4428 8536 4480
rect 16672 4471 16724 4480
rect 16672 4437 16681 4471
rect 16681 4437 16715 4471
rect 16715 4437 16724 4471
rect 16672 4428 16724 4437
rect 17960 4428 18012 4480
rect 22284 4428 22336 4480
rect 26976 4632 27028 4684
rect 30472 4632 30524 4684
rect 28172 4564 28224 4616
rect 26424 4496 26476 4548
rect 34520 4700 34572 4752
rect 34888 4700 34940 4752
rect 35164 4700 35216 4752
rect 36452 4700 36504 4752
rect 36820 4700 36872 4752
rect 37004 4700 37056 4752
rect 38936 4700 38988 4752
rect 39212 4700 39264 4752
rect 46204 4700 46256 4752
rect 46388 4768 46440 4820
rect 49700 4811 49752 4820
rect 49700 4777 49709 4811
rect 49709 4777 49743 4811
rect 49743 4777 49752 4811
rect 49700 4768 49752 4777
rect 50068 4768 50120 4820
rect 49332 4700 49384 4752
rect 50528 4768 50580 4820
rect 52828 4768 52880 4820
rect 53656 4811 53708 4820
rect 53656 4777 53665 4811
rect 53665 4777 53699 4811
rect 53699 4777 53708 4811
rect 53656 4768 53708 4777
rect 55220 4768 55272 4820
rect 55496 4768 55548 4820
rect 57428 4768 57480 4820
rect 57612 4768 57664 4820
rect 81624 4768 81676 4820
rect 86776 4768 86828 4820
rect 56968 4700 57020 4752
rect 57336 4700 57388 4752
rect 60464 4700 60516 4752
rect 60740 4700 60792 4752
rect 39856 4632 39908 4684
rect 41512 4632 41564 4684
rect 41604 4632 41656 4684
rect 45652 4632 45704 4684
rect 30748 4564 30800 4616
rect 31484 4564 31536 4616
rect 30840 4496 30892 4548
rect 31852 4496 31904 4548
rect 24952 4471 25004 4480
rect 24952 4437 24961 4471
rect 24961 4437 24995 4471
rect 24995 4437 25004 4471
rect 24952 4428 25004 4437
rect 25044 4428 25096 4480
rect 32496 4428 32548 4480
rect 34428 4564 34480 4616
rect 36820 4564 36872 4616
rect 36912 4564 36964 4616
rect 40040 4564 40092 4616
rect 40224 4607 40276 4616
rect 40224 4573 40233 4607
rect 40233 4573 40267 4607
rect 40267 4573 40276 4607
rect 40224 4564 40276 4573
rect 40868 4564 40920 4616
rect 45560 4564 45612 4616
rect 36636 4496 36688 4548
rect 36728 4496 36780 4548
rect 41420 4496 41472 4548
rect 41512 4496 41564 4548
rect 44916 4496 44968 4548
rect 45192 4496 45244 4548
rect 33968 4428 34020 4480
rect 34060 4428 34112 4480
rect 45744 4428 45796 4480
rect 46112 4632 46164 4684
rect 46388 4632 46440 4684
rect 46572 4675 46624 4684
rect 46572 4641 46581 4675
rect 46581 4641 46615 4675
rect 46615 4641 46624 4675
rect 46572 4632 46624 4641
rect 46848 4632 46900 4684
rect 47676 4632 47728 4684
rect 56324 4632 56376 4684
rect 57612 4632 57664 4684
rect 63684 4632 63736 4684
rect 87788 4675 87840 4684
rect 87788 4641 87797 4675
rect 87797 4641 87831 4675
rect 87831 4641 87840 4675
rect 92756 4768 92808 4820
rect 104440 4811 104492 4820
rect 104440 4777 104449 4811
rect 104449 4777 104483 4811
rect 104483 4777 104492 4811
rect 104440 4768 104492 4777
rect 118884 4768 118936 4820
rect 121920 4811 121972 4820
rect 121920 4777 121929 4811
rect 121929 4777 121963 4811
rect 121963 4777 121972 4811
rect 121920 4768 121972 4777
rect 129188 4811 129240 4820
rect 129188 4777 129197 4811
rect 129197 4777 129231 4811
rect 129231 4777 129240 4811
rect 129188 4768 129240 4777
rect 130200 4811 130252 4820
rect 130200 4777 130209 4811
rect 130209 4777 130243 4811
rect 130243 4777 130252 4811
rect 130200 4768 130252 4777
rect 131304 4768 131356 4820
rect 146668 4768 146720 4820
rect 150164 4811 150216 4820
rect 150164 4777 150173 4811
rect 150173 4777 150207 4811
rect 150207 4777 150216 4811
rect 150164 4768 150216 4777
rect 151728 4811 151780 4820
rect 151728 4777 151737 4811
rect 151737 4777 151771 4811
rect 151771 4777 151780 4811
rect 151728 4768 151780 4777
rect 152924 4768 152976 4820
rect 153660 4768 153712 4820
rect 156052 4768 156104 4820
rect 156604 4811 156656 4820
rect 156604 4777 156613 4811
rect 156613 4777 156647 4811
rect 156647 4777 156656 4811
rect 156604 4768 156656 4777
rect 158260 4811 158312 4820
rect 158260 4777 158269 4811
rect 158269 4777 158303 4811
rect 158303 4777 158312 4811
rect 158260 4768 158312 4777
rect 163964 4768 164016 4820
rect 90548 4700 90600 4752
rect 87788 4632 87840 4641
rect 46480 4564 46532 4616
rect 46204 4496 46256 4548
rect 46480 4428 46532 4480
rect 46664 4496 46716 4548
rect 48044 4539 48096 4548
rect 48044 4505 48053 4539
rect 48053 4505 48087 4539
rect 48087 4505 48096 4539
rect 48044 4496 48096 4505
rect 48228 4539 48280 4548
rect 48228 4505 48237 4539
rect 48237 4505 48271 4539
rect 48271 4505 48280 4539
rect 48228 4496 48280 4505
rect 48964 4564 49016 4616
rect 54760 4564 54812 4616
rect 55588 4564 55640 4616
rect 55772 4607 55824 4616
rect 55772 4573 55781 4607
rect 55781 4573 55815 4607
rect 55815 4573 55824 4607
rect 55772 4564 55824 4573
rect 49240 4471 49292 4480
rect 49240 4437 49249 4471
rect 49249 4437 49283 4471
rect 49283 4437 49292 4471
rect 49240 4428 49292 4437
rect 61292 4564 61344 4616
rect 90364 4607 90416 4616
rect 90364 4573 90373 4607
rect 90373 4573 90407 4607
rect 90407 4573 90416 4607
rect 90364 4564 90416 4573
rect 100392 4700 100444 4752
rect 103060 4632 103112 4684
rect 103796 4700 103848 4752
rect 110788 4700 110840 4752
rect 107016 4632 107068 4684
rect 109592 4632 109644 4684
rect 117044 4632 117096 4684
rect 100576 4564 100628 4616
rect 110328 4564 110380 4616
rect 49976 4428 50028 4480
rect 50620 4428 50672 4480
rect 51632 4428 51684 4480
rect 52092 4428 52144 4480
rect 55128 4428 55180 4480
rect 55496 4428 55548 4480
rect 57520 4496 57572 4548
rect 60648 4496 60700 4548
rect 61384 4496 61436 4548
rect 91100 4496 91152 4548
rect 92204 4496 92256 4548
rect 113456 4496 113508 4548
rect 113548 4496 113600 4548
rect 117136 4496 117188 4548
rect 56048 4428 56100 4480
rect 57612 4428 57664 4480
rect 57704 4428 57756 4480
rect 66444 4428 66496 4480
rect 92296 4471 92348 4480
rect 92296 4437 92305 4471
rect 92305 4437 92339 4471
rect 92339 4437 92348 4471
rect 92296 4428 92348 4437
rect 94964 4428 95016 4480
rect 100392 4428 100444 4480
rect 105912 4471 105964 4480
rect 105912 4437 105921 4471
rect 105921 4437 105955 4471
rect 105955 4437 105964 4471
rect 105912 4428 105964 4437
rect 110236 4471 110288 4480
rect 110236 4437 110245 4471
rect 110245 4437 110279 4471
rect 110279 4437 110288 4471
rect 110236 4428 110288 4437
rect 115388 4471 115440 4480
rect 115388 4437 115397 4471
rect 115397 4437 115431 4471
rect 115431 4437 115440 4471
rect 115388 4428 115440 4437
rect 130476 4496 130528 4548
rect 122748 4428 122800 4480
rect 128360 4428 128412 4480
rect 129372 4428 129424 4480
rect 130844 4428 130896 4480
rect 146300 4496 146352 4548
rect 147404 4496 147456 4548
rect 152188 4632 152240 4684
rect 155316 4632 155368 4684
rect 156328 4632 156380 4684
rect 149612 4496 149664 4548
rect 132684 4428 132736 4480
rect 155132 4496 155184 4548
rect 153292 4428 153344 4480
rect 154856 4471 154908 4480
rect 154856 4437 154865 4471
rect 154865 4437 154899 4471
rect 154899 4437 154908 4471
rect 154856 4428 154908 4437
rect 156420 4428 156472 4480
rect 159548 4471 159600 4480
rect 159548 4437 159557 4471
rect 159557 4437 159591 4471
rect 159591 4437 159600 4471
rect 159548 4428 159600 4437
rect 163596 4471 163648 4480
rect 163596 4437 163605 4471
rect 163605 4437 163639 4471
rect 163639 4437 163648 4471
rect 163596 4428 163648 4437
rect 164700 4471 164752 4480
rect 164700 4437 164709 4471
rect 164709 4437 164743 4471
rect 164743 4437 164752 4471
rect 164700 4428 164752 4437
rect 56667 4326 56719 4378
rect 56731 4326 56783 4378
rect 56795 4326 56847 4378
rect 56859 4326 56911 4378
rect 113088 4326 113140 4378
rect 113152 4326 113204 4378
rect 113216 4326 113268 4378
rect 113280 4326 113332 4378
rect 3976 4267 4028 4276
rect 3976 4233 3985 4267
rect 3985 4233 4019 4267
rect 4019 4233 4028 4267
rect 3976 4224 4028 4233
rect 4068 4224 4120 4276
rect 9864 4224 9916 4276
rect 12072 4224 12124 4276
rect 31576 4224 31628 4276
rect 31668 4224 31720 4276
rect 31852 4224 31904 4276
rect 32220 4224 32272 4276
rect 34980 4224 35032 4276
rect 35164 4224 35216 4276
rect 9220 4156 9272 4208
rect 1308 4088 1360 4140
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 7012 4020 7064 4072
rect 8024 4088 8076 4140
rect 10140 4088 10192 4140
rect 14372 4088 14424 4140
rect 5356 3952 5408 4004
rect 8392 4020 8444 4072
rect 16304 4020 16356 4072
rect 16396 4020 16448 4072
rect 19616 4088 19668 4140
rect 21088 4063 21140 4072
rect 21088 4029 21097 4063
rect 21097 4029 21131 4063
rect 21131 4029 21140 4063
rect 21088 4020 21140 4029
rect 21364 4088 21416 4140
rect 24124 4088 24176 4140
rect 25412 4088 25464 4140
rect 29828 4156 29880 4208
rect 31116 4156 31168 4208
rect 36360 4156 36412 4208
rect 36636 4224 36688 4276
rect 48228 4224 48280 4276
rect 36728 4156 36780 4208
rect 36820 4156 36872 4208
rect 39672 4156 39724 4208
rect 40040 4156 40092 4208
rect 41512 4156 41564 4208
rect 26332 4088 26384 4140
rect 27804 4088 27856 4140
rect 32680 4131 32732 4140
rect 25504 4020 25556 4072
rect 3148 3884 3200 3936
rect 9312 3952 9364 4004
rect 9404 3952 9456 4004
rect 7932 3884 7984 3936
rect 16580 3884 16632 3936
rect 16764 3884 16816 3936
rect 18052 3884 18104 3936
rect 18420 3884 18472 3936
rect 20260 3884 20312 3936
rect 20444 3884 20496 3936
rect 21364 3884 21416 3936
rect 22008 3884 22060 3936
rect 23940 3884 23992 3936
rect 24216 3952 24268 4004
rect 25688 4020 25740 4072
rect 32680 4097 32689 4131
rect 32689 4097 32723 4131
rect 32723 4097 32732 4131
rect 32680 4088 32732 4097
rect 33232 4088 33284 4140
rect 42800 4156 42852 4208
rect 41972 4088 42024 4140
rect 42524 4088 42576 4140
rect 42616 4088 42668 4140
rect 45928 4156 45980 4208
rect 46020 4156 46072 4208
rect 48596 4156 48648 4208
rect 49792 4156 49844 4208
rect 49976 4224 50028 4276
rect 53196 4224 53248 4276
rect 51264 4156 51316 4208
rect 51540 4156 51592 4208
rect 55036 4224 55088 4276
rect 55128 4224 55180 4276
rect 55588 4156 55640 4208
rect 55772 4224 55824 4276
rect 56968 4224 57020 4276
rect 57060 4224 57112 4276
rect 61476 4224 61528 4276
rect 64604 4224 64656 4276
rect 57704 4156 57756 4208
rect 43352 4088 43404 4140
rect 44548 4088 44600 4140
rect 44824 4088 44876 4140
rect 47492 4088 47544 4140
rect 47952 4131 48004 4140
rect 47952 4097 47961 4131
rect 47961 4097 47995 4131
rect 47995 4097 48004 4131
rect 47952 4088 48004 4097
rect 48228 4088 48280 4140
rect 49608 4131 49660 4140
rect 40776 4020 40828 4072
rect 41052 4063 41104 4072
rect 41052 4029 41061 4063
rect 41061 4029 41095 4063
rect 41095 4029 41104 4063
rect 41052 4020 41104 4029
rect 26700 3952 26752 4004
rect 30748 3884 30800 3936
rect 31300 3952 31352 4004
rect 49608 4097 49617 4131
rect 49617 4097 49651 4131
rect 49651 4097 49660 4131
rect 49608 4088 49660 4097
rect 49700 4088 49752 4140
rect 51448 4020 51500 4072
rect 51632 4088 51684 4140
rect 51816 4020 51868 4072
rect 52000 4063 52052 4072
rect 52000 4029 52009 4063
rect 52009 4029 52043 4063
rect 52043 4029 52052 4063
rect 52000 4020 52052 4029
rect 52368 4088 52420 4140
rect 54300 4088 54352 4140
rect 55312 4131 55364 4140
rect 55312 4097 55321 4131
rect 55321 4097 55355 4131
rect 55355 4097 55364 4131
rect 55312 4088 55364 4097
rect 55496 4088 55548 4140
rect 56232 4088 56284 4140
rect 56324 4088 56376 4140
rect 60556 4088 60608 4140
rect 54760 4020 54812 4072
rect 55772 4020 55824 4072
rect 68284 4156 68336 4208
rect 61108 4131 61160 4140
rect 61108 4097 61117 4131
rect 61117 4097 61151 4131
rect 61151 4097 61160 4131
rect 61108 4088 61160 4097
rect 62212 4131 62264 4140
rect 62212 4097 62221 4131
rect 62221 4097 62255 4131
rect 62255 4097 62264 4131
rect 62212 4088 62264 4097
rect 62764 4131 62816 4140
rect 62764 4097 62773 4131
rect 62773 4097 62807 4131
rect 62807 4097 62816 4131
rect 62764 4088 62816 4097
rect 62948 4088 63000 4140
rect 63224 4131 63276 4140
rect 63224 4097 63233 4131
rect 63233 4097 63267 4131
rect 63267 4097 63276 4131
rect 63224 4088 63276 4097
rect 63316 4131 63368 4140
rect 63316 4097 63325 4131
rect 63325 4097 63359 4131
rect 63359 4097 63368 4131
rect 63316 4088 63368 4097
rect 68744 4088 68796 4140
rect 41512 3952 41564 4004
rect 45284 3952 45336 4004
rect 39948 3884 40000 3936
rect 40040 3884 40092 3936
rect 49424 3952 49476 4004
rect 50068 3952 50120 4004
rect 56048 3952 56100 4004
rect 64420 4020 64472 4072
rect 70032 4131 70084 4140
rect 70032 4097 70041 4131
rect 70041 4097 70075 4131
rect 70075 4097 70084 4131
rect 70032 4088 70084 4097
rect 70216 4088 70268 4140
rect 70584 4088 70636 4140
rect 70952 4131 71004 4140
rect 70952 4097 70961 4131
rect 70961 4097 70995 4131
rect 70995 4097 71004 4131
rect 70952 4088 71004 4097
rect 71044 4131 71096 4140
rect 71044 4097 71053 4131
rect 71053 4097 71087 4131
rect 71087 4097 71096 4131
rect 71964 4131 72016 4140
rect 71044 4088 71096 4097
rect 71964 4097 71973 4131
rect 71973 4097 72007 4131
rect 72007 4097 72016 4131
rect 71964 4088 72016 4097
rect 72056 4131 72108 4140
rect 72056 4097 72065 4131
rect 72065 4097 72099 4131
rect 72099 4097 72108 4131
rect 72056 4088 72108 4097
rect 76012 4088 76064 4140
rect 105912 4224 105964 4276
rect 113548 4224 113600 4276
rect 114008 4224 114060 4276
rect 115388 4224 115440 4276
rect 125876 4224 125928 4276
rect 153476 4267 153528 4276
rect 153476 4233 153485 4267
rect 153485 4233 153519 4267
rect 153519 4233 153528 4267
rect 153476 4224 153528 4233
rect 88892 4156 88944 4208
rect 76380 4088 76432 4140
rect 89168 4131 89220 4140
rect 89168 4097 89177 4131
rect 89177 4097 89211 4131
rect 89211 4097 89220 4131
rect 89168 4088 89220 4097
rect 91100 4088 91152 4140
rect 92296 4088 92348 4140
rect 100484 4088 100536 4140
rect 102232 4088 102284 4140
rect 106464 4088 106516 4140
rect 106648 4131 106700 4140
rect 106648 4097 106657 4131
rect 106657 4097 106691 4131
rect 106691 4097 106700 4131
rect 107752 4131 107804 4140
rect 106648 4088 106700 4097
rect 107752 4097 107761 4131
rect 107761 4097 107795 4131
rect 107795 4097 107804 4131
rect 107752 4088 107804 4097
rect 107844 4131 107896 4140
rect 107844 4097 107853 4131
rect 107853 4097 107887 4131
rect 107887 4097 107896 4131
rect 107844 4088 107896 4097
rect 109040 4088 109092 4140
rect 70400 4020 70452 4072
rect 71228 4020 71280 4072
rect 71320 4020 71372 4072
rect 77852 4020 77904 4072
rect 89996 4020 90048 4072
rect 91928 4020 91980 4072
rect 100300 4020 100352 4072
rect 108212 4020 108264 4072
rect 108396 4020 108448 4072
rect 113640 4088 113692 4140
rect 114836 4088 114888 4140
rect 117044 4156 117096 4208
rect 138664 4156 138716 4208
rect 115848 4131 115900 4140
rect 115848 4097 115857 4131
rect 115857 4097 115891 4131
rect 115891 4097 115900 4131
rect 115848 4088 115900 4097
rect 120080 4088 120132 4140
rect 121644 4088 121696 4140
rect 124588 4131 124640 4140
rect 124588 4097 124597 4131
rect 124597 4097 124631 4131
rect 124631 4097 124640 4131
rect 124588 4088 124640 4097
rect 125600 4131 125652 4140
rect 125600 4097 125609 4131
rect 125609 4097 125643 4131
rect 125643 4097 125652 4131
rect 125600 4088 125652 4097
rect 125968 4088 126020 4140
rect 126888 4131 126940 4140
rect 126888 4097 126897 4131
rect 126897 4097 126931 4131
rect 126931 4097 126940 4131
rect 126888 4088 126940 4097
rect 127164 4088 127216 4140
rect 130200 4131 130252 4140
rect 130200 4097 130209 4131
rect 130209 4097 130243 4131
rect 130243 4097 130252 4131
rect 130200 4088 130252 4097
rect 130292 4131 130344 4140
rect 130292 4097 130301 4131
rect 130301 4097 130335 4131
rect 130335 4097 130344 4131
rect 131304 4131 131356 4140
rect 130292 4088 130344 4097
rect 131304 4097 131313 4131
rect 131313 4097 131347 4131
rect 131347 4097 131356 4131
rect 131304 4088 131356 4097
rect 131396 4131 131448 4140
rect 131396 4097 131405 4131
rect 131405 4097 131439 4131
rect 131439 4097 131448 4131
rect 131396 4088 131448 4097
rect 109316 4020 109368 4072
rect 61384 3952 61436 4004
rect 45652 3884 45704 3936
rect 47768 3884 47820 3936
rect 47952 3927 48004 3936
rect 47952 3893 47961 3927
rect 47961 3893 47995 3927
rect 47995 3893 48004 3927
rect 47952 3884 48004 3893
rect 48504 3884 48556 3936
rect 55496 3884 55548 3936
rect 55772 3884 55824 3936
rect 58532 3884 58584 3936
rect 58716 3884 58768 3936
rect 64052 3884 64104 3936
rect 64604 3884 64656 3936
rect 70124 3884 70176 3936
rect 70308 3884 70360 3936
rect 70584 3884 70636 3936
rect 74540 3952 74592 4004
rect 84660 3952 84712 4004
rect 100484 3952 100536 4004
rect 83004 3884 83056 3936
rect 89260 3927 89312 3936
rect 89260 3893 89269 3927
rect 89269 3893 89303 3927
rect 89303 3893 89312 3927
rect 89260 3884 89312 3893
rect 100208 3884 100260 3936
rect 104256 3952 104308 4004
rect 107568 3952 107620 4004
rect 109224 3952 109276 4004
rect 111616 3952 111668 4004
rect 108856 3884 108908 3936
rect 108948 3884 109000 3936
rect 114744 3952 114796 4004
rect 114928 3952 114980 4004
rect 121736 4020 121788 4072
rect 129832 4020 129884 4072
rect 148232 4131 148284 4140
rect 148232 4097 148241 4131
rect 148241 4097 148275 4131
rect 148275 4097 148284 4131
rect 148232 4088 148284 4097
rect 150164 4088 150216 4140
rect 155040 4131 155092 4140
rect 155040 4097 155049 4131
rect 155049 4097 155083 4131
rect 155083 4097 155092 4131
rect 155040 4088 155092 4097
rect 156052 4131 156104 4140
rect 156052 4097 156061 4131
rect 156061 4097 156095 4131
rect 156095 4097 156104 4131
rect 156052 4088 156104 4097
rect 156236 4088 156288 4140
rect 149060 4020 149112 4072
rect 155960 4020 156012 4072
rect 158536 4131 158588 4140
rect 158536 4097 158545 4131
rect 158545 4097 158579 4131
rect 158579 4097 158588 4131
rect 158536 4088 158588 4097
rect 160560 4088 160612 4140
rect 161756 4088 161808 4140
rect 162492 4088 162544 4140
rect 164884 4088 164936 4140
rect 165528 4131 165580 4140
rect 165528 4097 165537 4131
rect 165537 4097 165571 4131
rect 165571 4097 165580 4131
rect 165528 4088 165580 4097
rect 165620 4131 165672 4140
rect 165620 4097 165629 4131
rect 165629 4097 165663 4131
rect 165663 4097 165672 4131
rect 165620 4088 165672 4097
rect 158720 4020 158772 4072
rect 160284 4063 160336 4072
rect 160284 4029 160293 4063
rect 160293 4029 160327 4063
rect 160327 4029 160336 4063
rect 160284 4020 160336 4029
rect 161572 4020 161624 4072
rect 162308 4063 162360 4072
rect 162308 4029 162317 4063
rect 162317 4029 162351 4063
rect 162351 4029 162360 4063
rect 162308 4020 162360 4029
rect 113548 3884 113600 3936
rect 114836 3884 114888 3936
rect 115020 3884 115072 3936
rect 117596 3884 117648 3936
rect 122288 3884 122340 3936
rect 134892 3952 134944 4004
rect 144092 3952 144144 4004
rect 158168 3952 158220 4004
rect 126428 3927 126480 3936
rect 126428 3893 126437 3927
rect 126437 3893 126471 3927
rect 126471 3893 126480 3927
rect 126428 3884 126480 3893
rect 151084 3884 151136 3936
rect 28456 3782 28508 3834
rect 28520 3782 28572 3834
rect 28584 3782 28636 3834
rect 28648 3782 28700 3834
rect 84878 3782 84930 3834
rect 84942 3782 84994 3834
rect 85006 3782 85058 3834
rect 85070 3782 85122 3834
rect 141299 3782 141351 3834
rect 141363 3782 141415 3834
rect 141427 3782 141479 3834
rect 141491 3782 141543 3834
rect 3608 3680 3660 3732
rect 6368 3680 6420 3732
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 7196 3723 7248 3732
rect 7196 3689 7205 3723
rect 7205 3689 7239 3723
rect 7239 3689 7248 3723
rect 7196 3680 7248 3689
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 9220 3680 9272 3732
rect 9680 3680 9732 3732
rect 11704 3680 11756 3732
rect 16304 3680 16356 3732
rect 4068 3612 4120 3664
rect 8668 3612 8720 3664
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 6644 3476 6696 3528
rect 9220 3544 9272 3596
rect 4896 3408 4948 3460
rect 7012 3451 7064 3460
rect 7012 3417 7021 3451
rect 7021 3417 7055 3451
rect 7055 3417 7064 3451
rect 7012 3408 7064 3417
rect 7748 3408 7800 3460
rect 10048 3408 10100 3460
rect 14372 3544 14424 3596
rect 11520 3451 11572 3460
rect 11520 3417 11529 3451
rect 11529 3417 11563 3451
rect 11563 3417 11572 3451
rect 11520 3408 11572 3417
rect 3976 3340 4028 3392
rect 10692 3340 10744 3392
rect 11980 3383 12032 3392
rect 11980 3349 11989 3383
rect 11989 3349 12023 3383
rect 12023 3349 12032 3383
rect 11980 3340 12032 3349
rect 15292 3612 15344 3664
rect 16672 3612 16724 3664
rect 19616 3680 19668 3732
rect 19892 3680 19944 3732
rect 25044 3723 25096 3732
rect 25044 3689 25053 3723
rect 25053 3689 25087 3723
rect 25087 3689 25096 3723
rect 25044 3680 25096 3689
rect 24032 3612 24084 3664
rect 24124 3612 24176 3664
rect 24860 3612 24912 3664
rect 15660 3544 15712 3596
rect 17960 3544 18012 3596
rect 19340 3544 19392 3596
rect 21916 3587 21968 3596
rect 18328 3476 18380 3528
rect 20720 3476 20772 3528
rect 21088 3519 21140 3528
rect 21088 3485 21097 3519
rect 21097 3485 21131 3519
rect 21131 3485 21140 3519
rect 21088 3476 21140 3485
rect 21916 3553 21925 3587
rect 21925 3553 21959 3587
rect 21959 3553 21968 3587
rect 21916 3544 21968 3553
rect 24492 3544 24544 3596
rect 26332 3723 26384 3732
rect 26332 3689 26341 3723
rect 26341 3689 26375 3723
rect 26375 3689 26384 3723
rect 26332 3680 26384 3689
rect 27988 3723 28040 3732
rect 27988 3689 27997 3723
rect 27997 3689 28031 3723
rect 28031 3689 28040 3723
rect 27988 3680 28040 3689
rect 28080 3680 28132 3732
rect 28908 3680 28960 3732
rect 29644 3723 29696 3732
rect 29644 3689 29653 3723
rect 29653 3689 29687 3723
rect 29687 3689 29696 3723
rect 29644 3680 29696 3689
rect 30012 3680 30064 3732
rect 47676 3680 47728 3732
rect 48044 3723 48096 3732
rect 48044 3689 48053 3723
rect 48053 3689 48087 3723
rect 48087 3689 48096 3723
rect 48044 3680 48096 3689
rect 48136 3680 48188 3732
rect 49608 3723 49660 3732
rect 49608 3689 49617 3723
rect 49617 3689 49651 3723
rect 49651 3689 49660 3723
rect 49608 3680 49660 3689
rect 50160 3680 50212 3732
rect 51724 3723 51776 3732
rect 51724 3689 51733 3723
rect 51733 3689 51767 3723
rect 51767 3689 51776 3723
rect 51724 3680 51776 3689
rect 51908 3680 51960 3732
rect 25412 3612 25464 3664
rect 26976 3612 27028 3664
rect 27252 3612 27304 3664
rect 32496 3612 32548 3664
rect 32680 3655 32732 3664
rect 32680 3621 32689 3655
rect 32689 3621 32723 3655
rect 32723 3621 32732 3655
rect 32680 3612 32732 3621
rect 32956 3612 33008 3664
rect 41236 3612 41288 3664
rect 25504 3544 25556 3596
rect 35808 3544 35860 3596
rect 35900 3544 35952 3596
rect 36360 3544 36412 3596
rect 37372 3544 37424 3596
rect 41972 3544 42024 3596
rect 42064 3544 42116 3596
rect 42984 3544 43036 3596
rect 43076 3544 43128 3596
rect 44456 3587 44508 3596
rect 14556 3408 14608 3460
rect 17316 3408 17368 3460
rect 20904 3408 20956 3460
rect 21088 3340 21140 3392
rect 21824 3408 21876 3460
rect 22008 3340 22060 3392
rect 25044 3476 25096 3528
rect 27988 3476 28040 3528
rect 25504 3408 25556 3460
rect 27068 3408 27120 3460
rect 25688 3340 25740 3392
rect 25872 3383 25924 3392
rect 25872 3349 25881 3383
rect 25881 3349 25915 3383
rect 25915 3349 25924 3383
rect 25872 3340 25924 3349
rect 37464 3519 37516 3528
rect 37464 3485 37473 3519
rect 37473 3485 37507 3519
rect 37507 3485 37516 3519
rect 37464 3476 37516 3485
rect 38108 3476 38160 3528
rect 39856 3476 39908 3528
rect 39948 3476 40000 3528
rect 29552 3408 29604 3460
rect 41052 3408 41104 3460
rect 29644 3340 29696 3392
rect 34612 3340 34664 3392
rect 34704 3340 34756 3392
rect 41420 3408 41472 3460
rect 41604 3476 41656 3528
rect 43536 3476 43588 3528
rect 44456 3553 44465 3587
rect 44465 3553 44499 3587
rect 44499 3553 44508 3587
rect 44456 3544 44508 3553
rect 44548 3544 44600 3596
rect 45468 3544 45520 3596
rect 45652 3612 45704 3664
rect 46296 3612 46348 3664
rect 49424 3612 49476 3664
rect 52000 3612 52052 3664
rect 41880 3408 41932 3460
rect 42340 3408 42392 3460
rect 45836 3519 45888 3528
rect 45836 3485 45845 3519
rect 45845 3485 45879 3519
rect 45879 3485 45888 3519
rect 45836 3476 45888 3485
rect 46112 3519 46164 3528
rect 46112 3485 46121 3519
rect 46121 3485 46155 3519
rect 46155 3485 46164 3519
rect 46112 3476 46164 3485
rect 51080 3544 51132 3596
rect 54760 3612 54812 3664
rect 55312 3680 55364 3732
rect 57244 3680 57296 3732
rect 58256 3723 58308 3732
rect 58256 3689 58265 3723
rect 58265 3689 58299 3723
rect 58299 3689 58308 3723
rect 58256 3680 58308 3689
rect 58716 3723 58768 3732
rect 58716 3689 58725 3723
rect 58725 3689 58759 3723
rect 58759 3689 58768 3723
rect 58716 3680 58768 3689
rect 55680 3612 55732 3664
rect 56416 3612 56468 3664
rect 60648 3680 60700 3732
rect 60740 3680 60792 3732
rect 83740 3680 83792 3732
rect 89168 3723 89220 3732
rect 89168 3689 89177 3723
rect 89177 3689 89211 3723
rect 89211 3689 89220 3723
rect 89168 3680 89220 3689
rect 92572 3680 92624 3732
rect 61108 3612 61160 3664
rect 63592 3612 63644 3664
rect 63868 3655 63920 3664
rect 63868 3621 63877 3655
rect 63877 3621 63911 3655
rect 63911 3621 63920 3655
rect 63868 3612 63920 3621
rect 68836 3612 68888 3664
rect 52368 3587 52420 3596
rect 46756 3476 46808 3528
rect 48872 3519 48924 3528
rect 44088 3408 44140 3460
rect 45468 3408 45520 3460
rect 41236 3340 41288 3392
rect 43444 3340 43496 3392
rect 43536 3340 43588 3392
rect 46204 3408 46256 3460
rect 46296 3408 46348 3460
rect 48596 3408 48648 3460
rect 48872 3485 48881 3519
rect 48881 3485 48915 3519
rect 48915 3485 48924 3519
rect 48872 3476 48924 3485
rect 52368 3553 52377 3587
rect 52377 3553 52411 3587
rect 52411 3553 52420 3587
rect 52368 3544 52420 3553
rect 51816 3476 51868 3528
rect 54024 3476 54076 3528
rect 57152 3544 57204 3596
rect 60556 3544 60608 3596
rect 63040 3544 63092 3596
rect 63224 3544 63276 3596
rect 65248 3544 65300 3596
rect 56324 3476 56376 3528
rect 48964 3408 49016 3460
rect 54484 3408 54536 3460
rect 55864 3408 55916 3460
rect 56692 3408 56744 3460
rect 60096 3476 60148 3528
rect 62764 3476 62816 3528
rect 62948 3476 63000 3528
rect 69020 3544 69072 3596
rect 48412 3340 48464 3392
rect 52184 3340 52236 3392
rect 53288 3340 53340 3392
rect 55956 3340 56008 3392
rect 56968 3383 57020 3392
rect 56968 3349 56977 3383
rect 56977 3349 57011 3383
rect 57011 3349 57020 3383
rect 56968 3340 57020 3349
rect 57060 3340 57112 3392
rect 62028 3408 62080 3460
rect 62212 3408 62264 3460
rect 64236 3408 64288 3460
rect 60372 3340 60424 3392
rect 60464 3340 60516 3392
rect 62488 3383 62540 3392
rect 62488 3349 62497 3383
rect 62497 3349 62531 3383
rect 62531 3349 62540 3383
rect 62488 3340 62540 3349
rect 62764 3340 62816 3392
rect 67640 3519 67692 3528
rect 67640 3485 67649 3519
rect 67649 3485 67683 3519
rect 67683 3485 67692 3519
rect 67640 3476 67692 3485
rect 70584 3612 70636 3664
rect 71780 3655 71832 3664
rect 71780 3621 71789 3655
rect 71789 3621 71823 3655
rect 71823 3621 71832 3655
rect 71780 3612 71832 3621
rect 71964 3612 72016 3664
rect 72700 3612 72752 3664
rect 67456 3408 67508 3460
rect 72148 3544 72200 3596
rect 72884 3612 72936 3664
rect 72976 3612 73028 3664
rect 78220 3612 78272 3664
rect 89444 3655 89496 3664
rect 89444 3621 89453 3655
rect 89453 3621 89487 3655
rect 89487 3621 89496 3655
rect 89444 3612 89496 3621
rect 91100 3612 91152 3664
rect 91744 3612 91796 3664
rect 73068 3544 73120 3596
rect 88432 3544 88484 3596
rect 66076 3340 66128 3392
rect 66352 3340 66404 3392
rect 68744 3340 68796 3392
rect 69112 3340 69164 3392
rect 70400 3340 70452 3392
rect 71136 3476 71188 3528
rect 72332 3476 72384 3528
rect 73344 3476 73396 3528
rect 78956 3476 79008 3528
rect 70952 3408 71004 3460
rect 71596 3408 71648 3460
rect 72056 3408 72108 3460
rect 72424 3408 72476 3460
rect 81900 3408 81952 3460
rect 73344 3340 73396 3392
rect 73712 3383 73764 3392
rect 73712 3349 73721 3383
rect 73721 3349 73755 3383
rect 73755 3349 73764 3383
rect 73712 3340 73764 3349
rect 73804 3340 73856 3392
rect 85948 3340 86000 3392
rect 88340 3383 88392 3392
rect 88340 3349 88349 3383
rect 88349 3349 88383 3383
rect 88383 3349 88392 3383
rect 88340 3340 88392 3349
rect 88800 3383 88852 3392
rect 88800 3349 88809 3383
rect 88809 3349 88843 3383
rect 88843 3349 88852 3383
rect 88800 3340 88852 3349
rect 89996 3340 90048 3392
rect 90456 3383 90508 3392
rect 90456 3349 90465 3383
rect 90465 3349 90499 3383
rect 90499 3349 90508 3383
rect 90456 3340 90508 3349
rect 93216 3680 93268 3732
rect 100576 3680 100628 3732
rect 100024 3612 100076 3664
rect 107936 3612 107988 3664
rect 100300 3544 100352 3596
rect 108120 3544 108172 3596
rect 108396 3680 108448 3732
rect 113548 3680 113600 3732
rect 113640 3680 113692 3732
rect 115756 3680 115808 3732
rect 117504 3680 117556 3732
rect 124956 3723 125008 3732
rect 124956 3689 124965 3723
rect 124965 3689 124999 3723
rect 124999 3689 125008 3723
rect 124956 3680 125008 3689
rect 125692 3680 125744 3732
rect 131028 3680 131080 3732
rect 133512 3723 133564 3732
rect 133512 3689 133521 3723
rect 133521 3689 133555 3723
rect 133555 3689 133564 3723
rect 133512 3680 133564 3689
rect 143356 3680 143408 3732
rect 108948 3612 109000 3664
rect 139952 3612 140004 3664
rect 146024 3655 146076 3664
rect 146024 3621 146033 3655
rect 146033 3621 146067 3655
rect 146067 3621 146076 3655
rect 146024 3612 146076 3621
rect 149980 3655 150032 3664
rect 149980 3621 149989 3655
rect 149989 3621 150023 3655
rect 150023 3621 150032 3655
rect 149980 3612 150032 3621
rect 150164 3612 150216 3664
rect 152556 3612 152608 3664
rect 164424 3680 164476 3732
rect 165528 3723 165580 3732
rect 165528 3689 165537 3723
rect 165537 3689 165571 3723
rect 165571 3689 165580 3723
rect 165528 3680 165580 3689
rect 166724 3612 166776 3664
rect 126612 3544 126664 3596
rect 130200 3544 130252 3596
rect 131580 3544 131632 3596
rect 144736 3544 144788 3596
rect 162308 3544 162360 3596
rect 102324 3519 102376 3528
rect 102324 3485 102333 3519
rect 102333 3485 102367 3519
rect 102367 3485 102376 3519
rect 102324 3476 102376 3485
rect 102968 3476 103020 3528
rect 108028 3476 108080 3528
rect 108212 3476 108264 3528
rect 109224 3476 109276 3528
rect 109408 3476 109460 3528
rect 114008 3476 114060 3528
rect 94228 3408 94280 3460
rect 102232 3408 102284 3460
rect 106464 3408 106516 3460
rect 106740 3408 106792 3460
rect 107936 3408 107988 3460
rect 108856 3408 108908 3460
rect 108948 3408 109000 3460
rect 121736 3476 121788 3528
rect 124956 3476 125008 3528
rect 126428 3476 126480 3528
rect 129740 3476 129792 3528
rect 131948 3476 132000 3528
rect 133788 3476 133840 3528
rect 137100 3476 137152 3528
rect 148140 3476 148192 3528
rect 115020 3408 115072 3460
rect 91468 3340 91520 3392
rect 92296 3383 92348 3392
rect 92296 3349 92305 3383
rect 92305 3349 92339 3383
rect 92339 3349 92348 3383
rect 92296 3340 92348 3349
rect 100024 3340 100076 3392
rect 103336 3383 103388 3392
rect 103336 3349 103345 3383
rect 103345 3349 103379 3383
rect 103379 3349 103388 3383
rect 103336 3340 103388 3349
rect 103428 3340 103480 3392
rect 107568 3340 107620 3392
rect 107752 3340 107804 3392
rect 109868 3340 109920 3392
rect 114836 3383 114888 3392
rect 114836 3349 114845 3383
rect 114845 3349 114879 3383
rect 114879 3349 114888 3383
rect 114836 3340 114888 3349
rect 115848 3340 115900 3392
rect 117964 3340 118016 3392
rect 120080 3340 120132 3392
rect 121276 3340 121328 3392
rect 121644 3383 121696 3392
rect 121644 3349 121653 3383
rect 121653 3349 121687 3383
rect 121687 3349 121696 3383
rect 121644 3340 121696 3349
rect 123484 3340 123536 3392
rect 124588 3383 124640 3392
rect 124588 3349 124597 3383
rect 124597 3349 124631 3383
rect 124631 3349 124640 3383
rect 124588 3340 124640 3349
rect 125600 3340 125652 3392
rect 126336 3340 126388 3392
rect 126888 3340 126940 3392
rect 128636 3340 128688 3392
rect 131304 3340 131356 3392
rect 132316 3340 132368 3392
rect 137284 3383 137336 3392
rect 137284 3349 137293 3383
rect 137293 3349 137327 3383
rect 137327 3349 137336 3383
rect 137284 3340 137336 3349
rect 138756 3383 138808 3392
rect 138756 3349 138765 3383
rect 138765 3349 138799 3383
rect 138799 3349 138808 3383
rect 138756 3340 138808 3349
rect 142988 3408 143040 3460
rect 144828 3340 144880 3392
rect 149060 3340 149112 3392
rect 151084 3408 151136 3460
rect 151636 3451 151688 3460
rect 151636 3417 151645 3451
rect 151645 3417 151679 3451
rect 151679 3417 151688 3451
rect 151636 3408 151688 3417
rect 152004 3340 152056 3392
rect 163228 3476 163280 3528
rect 155040 3408 155092 3460
rect 157248 3408 157300 3460
rect 158720 3408 158772 3460
rect 159916 3408 159968 3460
rect 153568 3340 153620 3392
rect 156052 3340 156104 3392
rect 156972 3340 157024 3392
rect 159456 3340 159508 3392
rect 160560 3340 160612 3392
rect 161756 3340 161808 3392
rect 162492 3340 162544 3392
rect 164424 3340 164476 3392
rect 164608 3340 164660 3392
rect 56667 3238 56719 3290
rect 56731 3238 56783 3290
rect 56795 3238 56847 3290
rect 56859 3238 56911 3290
rect 113088 3238 113140 3290
rect 113152 3238 113204 3290
rect 113216 3238 113268 3290
rect 113280 3238 113332 3290
rect 3884 3136 3936 3188
rect 11612 3136 11664 3188
rect 11704 3136 11756 3188
rect 21640 3136 21692 3188
rect 22468 3136 22520 3188
rect 6368 3068 6420 3120
rect 3700 3000 3752 3052
rect 4528 3000 4580 3052
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 7840 3000 7892 3052
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10140 3068 10192 3120
rect 17316 3068 17368 3120
rect 17868 3068 17920 3120
rect 10232 3000 10284 3052
rect 11980 3000 12032 3052
rect 13268 3043 13320 3052
rect 13268 3009 13277 3043
rect 13277 3009 13311 3043
rect 13311 3009 13320 3043
rect 13268 3000 13320 3009
rect 16028 3000 16080 3052
rect 17960 3000 18012 3052
rect 18420 3043 18472 3052
rect 756 2864 808 2916
rect 4896 2907 4948 2916
rect 4896 2873 4905 2907
rect 4905 2873 4939 2907
rect 4939 2873 4948 2907
rect 4896 2864 4948 2873
rect 4988 2864 5040 2916
rect 6184 2932 6236 2984
rect 17132 2932 17184 2984
rect 5540 2839 5592 2848
rect 5540 2805 5549 2839
rect 5549 2805 5583 2839
rect 5583 2805 5592 2839
rect 5540 2796 5592 2805
rect 6276 2864 6328 2916
rect 7380 2907 7432 2916
rect 7380 2873 7389 2907
rect 7389 2873 7423 2907
rect 7423 2873 7432 2907
rect 7380 2864 7432 2873
rect 7472 2864 7524 2916
rect 9680 2796 9732 2848
rect 9864 2864 9916 2916
rect 15384 2864 15436 2916
rect 18420 3009 18429 3043
rect 18429 3009 18463 3043
rect 18463 3009 18472 3043
rect 18420 3000 18472 3009
rect 18604 3000 18656 3052
rect 25320 3136 25372 3188
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 21548 3000 21600 3052
rect 21732 3000 21784 3052
rect 23112 3000 23164 3052
rect 18972 2932 19024 2984
rect 18696 2864 18748 2916
rect 19708 2864 19760 2916
rect 20352 2932 20404 2984
rect 10232 2796 10284 2848
rect 12440 2796 12492 2848
rect 14188 2796 14240 2848
rect 17960 2796 18012 2848
rect 18328 2796 18380 2848
rect 18512 2796 18564 2848
rect 19340 2796 19392 2848
rect 23480 2796 23532 2848
rect 23756 2932 23808 2984
rect 25412 3000 25464 3052
rect 25228 2932 25280 2984
rect 25964 3068 26016 3120
rect 28908 3136 28960 3188
rect 29552 3136 29604 3188
rect 30380 3136 30432 3188
rect 33232 3136 33284 3188
rect 33324 3136 33376 3188
rect 39488 3136 39540 3188
rect 39580 3136 39632 3188
rect 41512 3136 41564 3188
rect 41604 3136 41656 3188
rect 44088 3136 44140 3188
rect 44824 3179 44876 3188
rect 44824 3145 44833 3179
rect 44833 3145 44867 3179
rect 44867 3145 44876 3179
rect 44824 3136 44876 3145
rect 44916 3136 44968 3188
rect 46296 3136 46348 3188
rect 46480 3179 46532 3188
rect 46480 3145 46489 3179
rect 46489 3145 46523 3179
rect 46523 3145 46532 3179
rect 46480 3136 46532 3145
rect 46664 3136 46716 3188
rect 47124 3136 47176 3188
rect 47584 3179 47636 3188
rect 47584 3145 47593 3179
rect 47593 3145 47627 3179
rect 47627 3145 47636 3179
rect 47584 3136 47636 3145
rect 27436 3043 27488 3052
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 29644 3000 29696 3052
rect 26148 2864 26200 2916
rect 27344 2864 27396 2916
rect 28172 2932 28224 2984
rect 30288 2864 30340 2916
rect 30748 3068 30800 3120
rect 36544 3068 36596 3120
rect 30932 3043 30984 3052
rect 30932 3009 30941 3043
rect 30941 3009 30975 3043
rect 30975 3009 30984 3043
rect 30932 3000 30984 3009
rect 31208 3000 31260 3052
rect 31944 3000 31996 3052
rect 33692 3000 33744 3052
rect 36728 3043 36780 3052
rect 36728 3009 36737 3043
rect 36737 3009 36771 3043
rect 36771 3009 36780 3043
rect 37004 3068 37056 3120
rect 39028 3068 39080 3120
rect 36728 3000 36780 3009
rect 37832 3000 37884 3052
rect 39948 3068 40000 3120
rect 40040 3068 40092 3120
rect 41052 3068 41104 3120
rect 31668 2932 31720 2984
rect 31852 2932 31904 2984
rect 32588 2932 32640 2984
rect 36360 2932 36412 2984
rect 39672 3000 39724 3052
rect 38016 2932 38068 2984
rect 38752 2932 38804 2984
rect 38936 2975 38988 2984
rect 38936 2941 38945 2975
rect 38945 2941 38979 2975
rect 38979 2941 38988 2975
rect 38936 2932 38988 2941
rect 39028 2932 39080 2984
rect 39580 2932 39632 2984
rect 40132 3000 40184 3052
rect 40316 3043 40368 3052
rect 40316 3009 40325 3043
rect 40325 3009 40359 3043
rect 40359 3009 40368 3043
rect 40316 3000 40368 3009
rect 40776 3000 40828 3052
rect 43076 3068 43128 3120
rect 43444 3068 43496 3120
rect 49332 3136 49384 3188
rect 49516 3136 49568 3188
rect 41696 3000 41748 3052
rect 42340 3000 42392 3052
rect 39948 2932 40000 2984
rect 43352 3000 43404 3052
rect 43536 3000 43588 3052
rect 43812 3000 43864 3052
rect 44824 3000 44876 3052
rect 44916 3000 44968 3052
rect 48044 3068 48096 3120
rect 53104 3068 53156 3120
rect 53196 3068 53248 3120
rect 55220 3136 55272 3188
rect 55680 3068 55732 3120
rect 56140 3136 56192 3188
rect 56968 3136 57020 3188
rect 60464 3136 60516 3188
rect 60556 3136 60608 3188
rect 61108 3136 61160 3188
rect 62304 3179 62356 3188
rect 62304 3145 62313 3179
rect 62313 3145 62347 3179
rect 62347 3145 62356 3179
rect 62304 3136 62356 3145
rect 62672 3136 62724 3188
rect 64420 3179 64472 3188
rect 64420 3145 64429 3179
rect 64429 3145 64463 3179
rect 64463 3145 64472 3179
rect 64420 3136 64472 3145
rect 64512 3136 64564 3188
rect 70124 3136 70176 3188
rect 70400 3136 70452 3188
rect 71780 3136 71832 3188
rect 73528 3179 73580 3188
rect 73528 3145 73537 3179
rect 73537 3145 73571 3179
rect 73571 3145 73580 3179
rect 73528 3136 73580 3145
rect 88432 3179 88484 3188
rect 88432 3145 88441 3179
rect 88441 3145 88475 3179
rect 88475 3145 88484 3179
rect 88432 3136 88484 3145
rect 88800 3136 88852 3188
rect 93308 3136 93360 3188
rect 104440 3136 104492 3188
rect 108948 3136 109000 3188
rect 109040 3136 109092 3188
rect 133236 3179 133288 3188
rect 57980 3068 58032 3120
rect 58992 3068 59044 3120
rect 65708 3068 65760 3120
rect 65984 3068 66036 3120
rect 45560 3043 45612 3052
rect 45560 3009 45569 3043
rect 45569 3009 45603 3043
rect 45603 3009 45612 3043
rect 45560 3000 45612 3009
rect 45744 3000 45796 3052
rect 42708 2975 42760 2984
rect 42708 2941 42717 2975
rect 42717 2941 42751 2975
rect 42751 2941 42760 2975
rect 42708 2932 42760 2941
rect 25688 2796 25740 2848
rect 25780 2796 25832 2848
rect 26516 2796 26568 2848
rect 27620 2796 27672 2848
rect 34704 2796 34756 2848
rect 34796 2796 34848 2848
rect 35624 2796 35676 2848
rect 36360 2796 36412 2848
rect 36728 2796 36780 2848
rect 38200 2796 38252 2848
rect 38292 2796 38344 2848
rect 39856 2796 39908 2848
rect 40500 2796 40552 2848
rect 41696 2864 41748 2916
rect 41880 2864 41932 2916
rect 41972 2864 42024 2916
rect 46572 2932 46624 2984
rect 47216 3000 47268 3052
rect 47584 3000 47636 3052
rect 48228 3000 48280 3052
rect 48780 3043 48832 3052
rect 48780 3009 48789 3043
rect 48789 3009 48823 3043
rect 48823 3009 48832 3043
rect 48780 3000 48832 3009
rect 49056 3000 49108 3052
rect 49148 3000 49200 3052
rect 50712 3000 50764 3052
rect 50804 3000 50856 3052
rect 53472 3000 53524 3052
rect 53656 3000 53708 3052
rect 54944 3000 54996 3052
rect 55128 3043 55180 3052
rect 55128 3009 55137 3043
rect 55137 3009 55171 3043
rect 55171 3009 55180 3043
rect 55128 3000 55180 3009
rect 55864 3000 55916 3052
rect 56324 3000 56376 3052
rect 57060 3000 57112 3052
rect 57244 3000 57296 3052
rect 45652 2864 45704 2916
rect 45836 2864 45888 2916
rect 49148 2864 49200 2916
rect 49332 2932 49384 2984
rect 51080 2864 51132 2916
rect 51264 2932 51316 2984
rect 51724 2864 51776 2916
rect 52184 2864 52236 2916
rect 55312 2864 55364 2916
rect 55496 2932 55548 2984
rect 57428 2932 57480 2984
rect 58440 2932 58492 2984
rect 58808 3000 58860 3052
rect 58900 3000 58952 3052
rect 59636 2932 59688 2984
rect 60464 3000 60516 3052
rect 60556 3000 60608 3052
rect 60648 2932 60700 2984
rect 60924 2932 60976 2984
rect 62396 3000 62448 3052
rect 63500 3000 63552 3052
rect 63776 3000 63828 3052
rect 63960 2932 64012 2984
rect 64512 3000 64564 3052
rect 68376 3000 68428 3052
rect 65340 2975 65392 2984
rect 65340 2941 65349 2975
rect 65349 2941 65383 2975
rect 65383 2941 65392 2975
rect 65340 2932 65392 2941
rect 66720 2975 66772 2984
rect 66720 2941 66729 2975
rect 66729 2941 66763 2975
rect 66763 2941 66772 2975
rect 66720 2932 66772 2941
rect 70216 3000 70268 3052
rect 70584 3000 70636 3052
rect 71136 3000 71188 3052
rect 71688 3000 71740 3052
rect 72056 3068 72108 3120
rect 86684 3068 86736 3120
rect 101588 3068 101640 3120
rect 74264 3000 74316 3052
rect 87328 3043 87380 3052
rect 87328 3009 87337 3043
rect 87337 3009 87371 3043
rect 87371 3009 87380 3043
rect 87328 3000 87380 3009
rect 88432 3000 88484 3052
rect 90272 3000 90324 3052
rect 90732 3000 90784 3052
rect 91836 3043 91888 3052
rect 91836 3009 91845 3043
rect 91845 3009 91879 3043
rect 91879 3009 91888 3043
rect 91836 3000 91888 3009
rect 102140 3000 102192 3052
rect 68560 2932 68612 2984
rect 71320 2932 71372 2984
rect 73620 2932 73672 2984
rect 76104 2932 76156 2984
rect 76564 2932 76616 2984
rect 80980 2932 81032 2984
rect 83096 2975 83148 2984
rect 83096 2941 83105 2975
rect 83105 2941 83139 2975
rect 83139 2941 83148 2975
rect 83096 2932 83148 2941
rect 86316 2975 86368 2984
rect 86316 2941 86325 2975
rect 86325 2941 86359 2975
rect 86359 2941 86368 2975
rect 86316 2932 86368 2941
rect 88156 2932 88208 2984
rect 103060 2932 103112 2984
rect 103520 3068 103572 3120
rect 107844 3111 107896 3120
rect 107844 3077 107853 3111
rect 107853 3077 107887 3111
rect 107887 3077 107896 3111
rect 107844 3068 107896 3077
rect 108120 3068 108172 3120
rect 107476 3000 107528 3052
rect 107752 3043 107804 3052
rect 107752 3009 107761 3043
rect 107761 3009 107795 3043
rect 107795 3009 107804 3043
rect 107752 3000 107804 3009
rect 108856 3068 108908 3120
rect 109408 3000 109460 3052
rect 109592 3043 109644 3052
rect 109592 3009 109601 3043
rect 109601 3009 109635 3043
rect 109635 3009 109644 3043
rect 109592 3000 109644 3009
rect 109776 3000 109828 3052
rect 111524 3000 111576 3052
rect 112812 3000 112864 3052
rect 114560 3000 114612 3052
rect 117228 3000 117280 3052
rect 119436 3000 119488 3052
rect 104164 2932 104216 2984
rect 104348 2975 104400 2984
rect 104348 2941 104357 2975
rect 104357 2941 104391 2975
rect 104391 2941 104400 2975
rect 104348 2932 104400 2941
rect 105452 2932 105504 2984
rect 108580 2932 108632 2984
rect 109132 2932 109184 2984
rect 120080 2932 120132 2984
rect 122472 3043 122524 3052
rect 122472 3009 122481 3043
rect 122481 3009 122515 3043
rect 122515 3009 122524 3043
rect 122472 3000 122524 3009
rect 126888 3000 126940 3052
rect 128176 3000 128228 3052
rect 125784 2932 125836 2984
rect 127992 2975 128044 2984
rect 127992 2941 128001 2975
rect 128001 2941 128035 2975
rect 128035 2941 128044 2975
rect 127992 2932 128044 2941
rect 133236 3145 133245 3179
rect 133245 3145 133279 3179
rect 133279 3145 133288 3179
rect 133236 3136 133288 3145
rect 134248 3179 134300 3188
rect 134248 3145 134257 3179
rect 134257 3145 134291 3179
rect 134291 3145 134300 3179
rect 134248 3136 134300 3145
rect 138572 3136 138624 3188
rect 144920 3136 144972 3188
rect 145380 3179 145432 3188
rect 145380 3145 145389 3179
rect 145389 3145 145423 3179
rect 145423 3145 145432 3179
rect 145380 3136 145432 3145
rect 149060 3136 149112 3188
rect 150348 3136 150400 3188
rect 154304 3179 154356 3188
rect 154304 3145 154313 3179
rect 154313 3145 154347 3179
rect 154347 3145 154356 3179
rect 154304 3136 154356 3145
rect 154948 3136 155000 3188
rect 156604 3136 156656 3188
rect 159732 3136 159784 3188
rect 160744 3179 160796 3188
rect 160744 3145 160753 3179
rect 160753 3145 160787 3179
rect 160787 3145 160796 3179
rect 160744 3136 160796 3145
rect 164332 3136 164384 3188
rect 165068 3179 165120 3188
rect 165068 3145 165077 3179
rect 165077 3145 165111 3179
rect 165111 3145 165120 3179
rect 165068 3136 165120 3145
rect 144460 3068 144512 3120
rect 161112 3068 161164 3120
rect 133052 3000 133104 3052
rect 134156 3043 134208 3052
rect 134156 3009 134165 3043
rect 134165 3009 134199 3043
rect 134199 3009 134208 3043
rect 134156 3000 134208 3009
rect 136640 3043 136692 3052
rect 136640 3009 136649 3043
rect 136649 3009 136683 3043
rect 136683 3009 136692 3043
rect 136640 3000 136692 3009
rect 136824 3000 136876 3052
rect 138020 3000 138072 3052
rect 139860 3000 139912 3052
rect 145564 3000 145616 3052
rect 149060 3043 149112 3052
rect 149060 3009 149069 3043
rect 149069 3009 149103 3043
rect 149103 3009 149112 3043
rect 149060 3000 149112 3009
rect 139400 2932 139452 2984
rect 141148 2932 141200 2984
rect 143172 2975 143224 2984
rect 143172 2941 143181 2975
rect 143181 2941 143215 2975
rect 143215 2941 143224 2975
rect 143172 2932 143224 2941
rect 143724 2932 143776 2984
rect 154396 3000 154448 3052
rect 155224 3043 155276 3052
rect 155224 3009 155233 3043
rect 155233 3009 155267 3043
rect 155267 3009 155276 3043
rect 155224 3000 155276 3009
rect 156236 3043 156288 3052
rect 156236 3009 156245 3043
rect 156245 3009 156279 3043
rect 156279 3009 156288 3043
rect 156236 3000 156288 3009
rect 160652 3043 160704 3052
rect 156696 2932 156748 2984
rect 158260 2975 158312 2984
rect 158260 2941 158269 2975
rect 158269 2941 158303 2975
rect 158303 2941 158312 2975
rect 158260 2932 158312 2941
rect 55772 2864 55824 2916
rect 56140 2864 56192 2916
rect 58072 2864 58124 2916
rect 42984 2796 43036 2848
rect 48964 2796 49016 2848
rect 54208 2796 54260 2848
rect 54576 2839 54628 2848
rect 54576 2805 54585 2839
rect 54585 2805 54619 2839
rect 54619 2805 54628 2839
rect 54576 2796 54628 2805
rect 55404 2796 55456 2848
rect 55496 2796 55548 2848
rect 57336 2796 57388 2848
rect 57704 2796 57756 2848
rect 58992 2864 59044 2916
rect 59452 2864 59504 2916
rect 58808 2796 58860 2848
rect 62764 2864 62816 2916
rect 63500 2864 63552 2916
rect 67180 2864 67232 2916
rect 67364 2864 67416 2916
rect 63224 2796 63276 2848
rect 64604 2796 64656 2848
rect 67732 2796 67784 2848
rect 69572 2839 69624 2848
rect 69572 2805 69581 2839
rect 69581 2805 69615 2839
rect 69615 2805 69624 2839
rect 69572 2796 69624 2805
rect 70492 2864 70544 2916
rect 70952 2864 71004 2916
rect 74908 2864 74960 2916
rect 105268 2864 105320 2916
rect 72424 2796 72476 2848
rect 73804 2796 73856 2848
rect 74264 2796 74316 2848
rect 77300 2796 77352 2848
rect 87420 2839 87472 2848
rect 87420 2805 87429 2839
rect 87429 2805 87463 2839
rect 87463 2805 87472 2839
rect 87420 2796 87472 2805
rect 88524 2796 88576 2848
rect 90364 2796 90416 2848
rect 100116 2796 100168 2848
rect 103244 2839 103296 2848
rect 103244 2805 103253 2839
rect 103253 2805 103287 2839
rect 103287 2805 103296 2839
rect 103244 2796 103296 2805
rect 103888 2839 103940 2848
rect 103888 2805 103897 2839
rect 103897 2805 103931 2839
rect 103931 2805 103940 2839
rect 103888 2796 103940 2805
rect 104256 2796 104308 2848
rect 108856 2864 108908 2916
rect 110328 2864 110380 2916
rect 111432 2864 111484 2916
rect 111616 2864 111668 2916
rect 114560 2864 114612 2916
rect 118700 2864 118752 2916
rect 122380 2864 122432 2916
rect 123852 2864 123904 2916
rect 110696 2796 110748 2848
rect 110880 2796 110932 2848
rect 111064 2796 111116 2848
rect 116124 2796 116176 2848
rect 116216 2796 116268 2848
rect 122656 2796 122708 2848
rect 134524 2864 134576 2916
rect 139676 2864 139728 2916
rect 142620 2864 142672 2916
rect 151360 2864 151412 2916
rect 152004 2864 152056 2916
rect 126888 2796 126940 2848
rect 127900 2796 127952 2848
rect 135444 2796 135496 2848
rect 136732 2839 136784 2848
rect 136732 2805 136741 2839
rect 136741 2805 136775 2839
rect 136775 2805 136784 2839
rect 136732 2796 136784 2805
rect 136916 2796 136968 2848
rect 140964 2796 141016 2848
rect 142252 2796 142304 2848
rect 145748 2796 145800 2848
rect 149152 2839 149204 2848
rect 149152 2805 149161 2839
rect 149161 2805 149195 2839
rect 149195 2805 149204 2839
rect 149152 2796 149204 2805
rect 149244 2796 149296 2848
rect 150900 2796 150952 2848
rect 158812 2864 158864 2916
rect 160652 3009 160661 3043
rect 160661 3009 160695 3043
rect 160695 3009 160704 3043
rect 160652 3000 160704 3009
rect 164148 3000 164200 3052
rect 165068 3000 165120 3052
rect 162032 2975 162084 2984
rect 162032 2941 162041 2975
rect 162041 2941 162075 2975
rect 162075 2941 162084 2975
rect 162032 2932 162084 2941
rect 160192 2864 160244 2916
rect 159824 2796 159876 2848
rect 164608 2796 164660 2848
rect 28456 2694 28508 2746
rect 28520 2694 28572 2746
rect 28584 2694 28636 2746
rect 28648 2694 28700 2746
rect 84878 2694 84930 2746
rect 84942 2694 84994 2746
rect 85006 2694 85058 2746
rect 85070 2694 85122 2746
rect 141299 2694 141351 2746
rect 141363 2694 141415 2746
rect 141427 2694 141479 2746
rect 141491 2694 141543 2746
rect 3700 2635 3752 2644
rect 3700 2601 3709 2635
rect 3709 2601 3743 2635
rect 3743 2601 3752 2635
rect 3700 2592 3752 2601
rect 4712 2635 4764 2644
rect 4712 2601 4721 2635
rect 4721 2601 4755 2635
rect 4755 2601 4764 2635
rect 4712 2592 4764 2601
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 12164 2592 12216 2644
rect 572 2524 624 2576
rect 9496 2524 9548 2576
rect 18328 2567 18380 2576
rect 18328 2533 18337 2567
rect 18337 2533 18371 2567
rect 18371 2533 18380 2567
rect 18328 2524 18380 2533
rect 20536 2524 20588 2576
rect 21732 2524 21784 2576
rect 23020 2592 23072 2644
rect 23756 2635 23808 2644
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 25136 2592 25188 2644
rect 25412 2635 25464 2644
rect 25412 2601 25421 2635
rect 25421 2601 25455 2635
rect 25455 2601 25464 2635
rect 25412 2592 25464 2601
rect 27436 2592 27488 2644
rect 28264 2592 28316 2644
rect 28816 2592 28868 2644
rect 29644 2635 29696 2644
rect 29644 2601 29653 2635
rect 29653 2601 29687 2635
rect 29687 2601 29696 2635
rect 29644 2592 29696 2601
rect 30932 2635 30984 2644
rect 30932 2601 30941 2635
rect 30941 2601 30975 2635
rect 30975 2601 30984 2635
rect 30932 2592 30984 2601
rect 35072 2592 35124 2644
rect 35348 2592 35400 2644
rect 38016 2592 38068 2644
rect 38384 2592 38436 2644
rect 39672 2592 39724 2644
rect 26056 2524 26108 2576
rect 26516 2524 26568 2576
rect 5540 2456 5592 2508
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 9772 2456 9824 2508
rect 10692 2499 10744 2508
rect 10692 2465 10701 2499
rect 10701 2465 10735 2499
rect 10735 2465 10744 2499
rect 10692 2456 10744 2465
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 18512 2431 18564 2440
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 7840 2252 7892 2304
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 19616 2388 19668 2440
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 21088 2388 21140 2440
rect 13268 2320 13320 2372
rect 10324 2252 10376 2304
rect 19616 2295 19668 2304
rect 19616 2261 19625 2295
rect 19625 2261 19659 2295
rect 19659 2261 19668 2295
rect 19616 2252 19668 2261
rect 19708 2252 19760 2304
rect 22192 2295 22244 2304
rect 22192 2261 22201 2295
rect 22201 2261 22235 2295
rect 22235 2261 22244 2295
rect 22192 2252 22244 2261
rect 23480 2456 23532 2508
rect 23940 2456 23992 2508
rect 25780 2431 25832 2440
rect 25780 2397 25789 2431
rect 25789 2397 25823 2431
rect 25823 2397 25832 2431
rect 25780 2388 25832 2397
rect 26148 2431 26200 2440
rect 26148 2397 26157 2431
rect 26157 2397 26191 2431
rect 26191 2397 26200 2431
rect 26148 2388 26200 2397
rect 27344 2431 27396 2440
rect 27344 2397 27353 2431
rect 27353 2397 27387 2431
rect 27387 2397 27396 2431
rect 27344 2388 27396 2397
rect 35716 2456 35768 2508
rect 35808 2456 35860 2508
rect 37004 2456 37056 2508
rect 39948 2524 40000 2576
rect 40224 2635 40276 2644
rect 40224 2601 40233 2635
rect 40233 2601 40267 2635
rect 40267 2601 40276 2635
rect 40224 2592 40276 2601
rect 41328 2592 41380 2644
rect 41880 2592 41932 2644
rect 42432 2592 42484 2644
rect 44088 2592 44140 2644
rect 44180 2592 44232 2644
rect 45560 2635 45612 2644
rect 45560 2601 45569 2635
rect 45569 2601 45603 2635
rect 45603 2601 45612 2635
rect 45560 2592 45612 2601
rect 40500 2524 40552 2576
rect 38752 2456 38804 2508
rect 32680 2388 32732 2440
rect 32772 2388 32824 2440
rect 35256 2388 35308 2440
rect 35532 2388 35584 2440
rect 36268 2388 36320 2440
rect 36360 2388 36412 2440
rect 36636 2388 36688 2440
rect 38660 2388 38712 2440
rect 38936 2431 38988 2440
rect 38936 2397 38945 2431
rect 38945 2397 38979 2431
rect 38979 2397 38988 2431
rect 39120 2431 39172 2440
rect 38936 2388 38988 2397
rect 39120 2397 39129 2431
rect 39129 2397 39163 2431
rect 39163 2397 39172 2431
rect 39120 2388 39172 2397
rect 39396 2388 39448 2440
rect 40500 2388 40552 2440
rect 40868 2456 40920 2508
rect 41972 2456 42024 2508
rect 41144 2388 41196 2440
rect 43904 2456 43956 2508
rect 44272 2456 44324 2508
rect 26516 2252 26568 2304
rect 30840 2252 30892 2304
rect 31852 2252 31904 2304
rect 35348 2252 35400 2304
rect 35624 2252 35676 2304
rect 44180 2388 44232 2440
rect 45836 2524 45888 2576
rect 46204 2592 46256 2644
rect 46480 2592 46532 2644
rect 46572 2592 46624 2644
rect 47032 2592 47084 2644
rect 47216 2592 47268 2644
rect 47768 2592 47820 2644
rect 48872 2592 48924 2644
rect 49056 2635 49108 2644
rect 49056 2601 49065 2635
rect 49065 2601 49099 2635
rect 49099 2601 49108 2635
rect 49056 2592 49108 2601
rect 49148 2592 49200 2644
rect 50804 2592 50856 2644
rect 50896 2592 50948 2644
rect 51724 2592 51776 2644
rect 52828 2635 52880 2644
rect 52828 2601 52837 2635
rect 52837 2601 52871 2635
rect 52871 2601 52880 2635
rect 52828 2592 52880 2601
rect 53288 2635 53340 2644
rect 53288 2601 53297 2635
rect 53297 2601 53331 2635
rect 53331 2601 53340 2635
rect 53288 2592 53340 2601
rect 53656 2635 53708 2644
rect 53656 2601 53665 2635
rect 53665 2601 53699 2635
rect 53699 2601 53708 2635
rect 53656 2592 53708 2601
rect 55220 2635 55272 2644
rect 55220 2601 55229 2635
rect 55229 2601 55263 2635
rect 55263 2601 55272 2635
rect 55220 2592 55272 2601
rect 55680 2592 55732 2644
rect 56232 2592 56284 2644
rect 57060 2592 57112 2644
rect 57152 2592 57204 2644
rect 58808 2592 58860 2644
rect 60740 2592 60792 2644
rect 60924 2635 60976 2644
rect 60924 2601 60933 2635
rect 60933 2601 60967 2635
rect 60967 2601 60976 2635
rect 60924 2592 60976 2601
rect 61292 2635 61344 2644
rect 61292 2601 61301 2635
rect 61301 2601 61335 2635
rect 61335 2601 61344 2635
rect 61292 2592 61344 2601
rect 62580 2592 62632 2644
rect 62856 2592 62908 2644
rect 63500 2635 63552 2644
rect 63500 2601 63509 2635
rect 63509 2601 63543 2635
rect 63543 2601 63552 2635
rect 63500 2592 63552 2601
rect 63684 2635 63736 2644
rect 63684 2601 63693 2635
rect 63693 2601 63727 2635
rect 63727 2601 63736 2635
rect 63684 2592 63736 2601
rect 64512 2635 64564 2644
rect 64512 2601 64521 2635
rect 64521 2601 64555 2635
rect 64555 2601 64564 2635
rect 64512 2592 64564 2601
rect 66536 2635 66588 2644
rect 66536 2601 66545 2635
rect 66545 2601 66579 2635
rect 66579 2601 66588 2635
rect 66536 2592 66588 2601
rect 67548 2635 67600 2644
rect 67548 2601 67557 2635
rect 67557 2601 67591 2635
rect 67591 2601 67600 2635
rect 67548 2592 67600 2601
rect 68560 2635 68612 2644
rect 68560 2601 68569 2635
rect 68569 2601 68603 2635
rect 68603 2601 68612 2635
rect 68560 2592 68612 2601
rect 70216 2592 70268 2644
rect 70584 2592 70636 2644
rect 71136 2592 71188 2644
rect 71688 2592 71740 2644
rect 71872 2635 71924 2644
rect 71872 2601 71881 2635
rect 71881 2601 71915 2635
rect 71915 2601 71924 2635
rect 71872 2592 71924 2601
rect 72148 2592 72200 2644
rect 74264 2635 74316 2644
rect 74264 2601 74273 2635
rect 74273 2601 74307 2635
rect 74307 2601 74316 2635
rect 74264 2592 74316 2601
rect 74724 2592 74776 2644
rect 79692 2592 79744 2644
rect 80888 2592 80940 2644
rect 81992 2635 82044 2644
rect 81992 2601 82001 2635
rect 82001 2601 82035 2635
rect 82035 2601 82044 2635
rect 81992 2592 82044 2601
rect 83464 2635 83516 2644
rect 83464 2601 83473 2635
rect 83473 2601 83507 2635
rect 83507 2601 83516 2635
rect 83464 2592 83516 2601
rect 83556 2592 83608 2644
rect 86960 2635 87012 2644
rect 61476 2524 61528 2576
rect 85764 2524 85816 2576
rect 86960 2601 86969 2635
rect 86969 2601 87003 2635
rect 87003 2601 87012 2635
rect 86960 2592 87012 2601
rect 87328 2635 87380 2644
rect 87328 2601 87337 2635
rect 87337 2601 87371 2635
rect 87371 2601 87380 2635
rect 87328 2592 87380 2601
rect 87604 2635 87656 2644
rect 87604 2601 87613 2635
rect 87613 2601 87647 2635
rect 87647 2601 87656 2635
rect 87604 2592 87656 2601
rect 88432 2635 88484 2644
rect 88432 2601 88441 2635
rect 88441 2601 88475 2635
rect 88475 2601 88484 2635
rect 88432 2592 88484 2601
rect 90272 2635 90324 2644
rect 90272 2601 90281 2635
rect 90281 2601 90315 2635
rect 90315 2601 90324 2635
rect 90272 2592 90324 2601
rect 102140 2592 102192 2644
rect 102968 2592 103020 2644
rect 103244 2592 103296 2644
rect 104164 2635 104216 2644
rect 104164 2601 104173 2635
rect 104173 2601 104207 2635
rect 104207 2601 104216 2635
rect 104164 2592 104216 2601
rect 108488 2635 108540 2644
rect 108488 2601 108497 2635
rect 108497 2601 108531 2635
rect 108531 2601 108540 2635
rect 108488 2592 108540 2601
rect 109500 2635 109552 2644
rect 109500 2601 109509 2635
rect 109509 2601 109543 2635
rect 109543 2601 109552 2635
rect 109500 2592 109552 2601
rect 109592 2592 109644 2644
rect 110328 2592 110380 2644
rect 110420 2592 110472 2644
rect 110788 2592 110840 2644
rect 111524 2635 111576 2644
rect 111524 2601 111533 2635
rect 111533 2601 111567 2635
rect 111567 2601 111576 2635
rect 111524 2592 111576 2601
rect 112720 2635 112772 2644
rect 112720 2601 112729 2635
rect 112729 2601 112763 2635
rect 112763 2601 112772 2635
rect 112720 2592 112772 2601
rect 113456 2592 113508 2644
rect 114560 2635 114612 2644
rect 114560 2601 114569 2635
rect 114569 2601 114603 2635
rect 114603 2601 114612 2635
rect 114560 2592 114612 2601
rect 117228 2635 117280 2644
rect 117228 2601 117237 2635
rect 117237 2601 117271 2635
rect 117271 2601 117280 2635
rect 117228 2592 117280 2601
rect 117688 2592 117740 2644
rect 118516 2592 118568 2644
rect 119804 2592 119856 2644
rect 120816 2635 120868 2644
rect 120816 2601 120825 2635
rect 120825 2601 120859 2635
rect 120859 2601 120868 2635
rect 120816 2592 120868 2601
rect 122380 2635 122432 2644
rect 122380 2601 122389 2635
rect 122389 2601 122423 2635
rect 122423 2601 122432 2635
rect 122380 2592 122432 2601
rect 123760 2635 123812 2644
rect 123760 2601 123769 2635
rect 123769 2601 123803 2635
rect 123803 2601 123812 2635
rect 123760 2592 123812 2601
rect 124220 2592 124272 2644
rect 126060 2635 126112 2644
rect 126060 2601 126069 2635
rect 126069 2601 126103 2635
rect 126103 2601 126112 2635
rect 126060 2592 126112 2601
rect 126888 2635 126940 2644
rect 126888 2601 126897 2635
rect 126897 2601 126931 2635
rect 126931 2601 126940 2635
rect 126888 2592 126940 2601
rect 126980 2592 127032 2644
rect 88340 2524 88392 2576
rect 118056 2524 118108 2576
rect 46296 2456 46348 2508
rect 45744 2388 45796 2440
rect 46204 2388 46256 2440
rect 48412 2456 48464 2508
rect 46480 2388 46532 2440
rect 50620 2456 50672 2508
rect 50712 2456 50764 2508
rect 48596 2388 48648 2440
rect 50252 2431 50304 2440
rect 50252 2397 50261 2431
rect 50261 2397 50295 2431
rect 50295 2397 50304 2431
rect 50252 2388 50304 2397
rect 44824 2320 44876 2372
rect 45376 2320 45428 2372
rect 46848 2320 46900 2372
rect 47124 2320 47176 2372
rect 47584 2320 47636 2372
rect 52644 2456 52696 2508
rect 54024 2499 54076 2508
rect 54024 2465 54033 2499
rect 54033 2465 54067 2499
rect 54067 2465 54076 2499
rect 54024 2456 54076 2465
rect 54208 2456 54260 2508
rect 51172 2388 51224 2440
rect 51356 2388 51408 2440
rect 51540 2388 51592 2440
rect 52092 2388 52144 2440
rect 53288 2388 53340 2440
rect 54576 2431 54628 2440
rect 54576 2397 54585 2431
rect 54585 2397 54619 2431
rect 54619 2397 54628 2431
rect 54576 2388 54628 2397
rect 55680 2456 55732 2508
rect 57244 2456 57296 2508
rect 57336 2456 57388 2508
rect 59728 2456 59780 2508
rect 59820 2456 59872 2508
rect 60556 2456 60608 2508
rect 61016 2456 61068 2508
rect 61384 2456 61436 2508
rect 61752 2456 61804 2508
rect 63224 2456 63276 2508
rect 63316 2456 63368 2508
rect 56048 2388 56100 2440
rect 56508 2388 56560 2440
rect 56968 2388 57020 2440
rect 57612 2388 57664 2440
rect 59360 2388 59412 2440
rect 61108 2431 61160 2440
rect 61108 2397 61117 2431
rect 61117 2397 61151 2431
rect 61151 2397 61160 2431
rect 61108 2388 61160 2397
rect 61660 2388 61712 2440
rect 63500 2388 63552 2440
rect 69756 2456 69808 2508
rect 72884 2456 72936 2508
rect 42616 2252 42668 2304
rect 51264 2320 51316 2372
rect 60004 2320 60056 2372
rect 51356 2252 51408 2304
rect 51448 2252 51500 2304
rect 51816 2252 51868 2304
rect 51908 2252 51960 2304
rect 56048 2252 56100 2304
rect 60556 2252 60608 2304
rect 62212 2252 62264 2304
rect 62396 2252 62448 2304
rect 63500 2252 63552 2304
rect 64972 2252 65024 2304
rect 67548 2252 67600 2304
rect 68008 2252 68060 2304
rect 70400 2252 70452 2304
rect 71320 2320 71372 2372
rect 73436 2252 73488 2304
rect 76564 2431 76616 2440
rect 76564 2397 76573 2431
rect 76573 2397 76607 2431
rect 76607 2397 76616 2431
rect 76564 2388 76616 2397
rect 76656 2431 76708 2440
rect 76656 2397 76665 2431
rect 76665 2397 76699 2431
rect 76699 2397 76708 2431
rect 80796 2456 80848 2508
rect 76656 2388 76708 2397
rect 79324 2431 79376 2440
rect 79324 2397 79333 2431
rect 79333 2397 79367 2431
rect 79367 2397 79376 2431
rect 79324 2388 79376 2397
rect 80428 2388 80480 2440
rect 91376 2499 91428 2508
rect 91376 2465 91385 2499
rect 91385 2465 91419 2499
rect 91419 2465 91428 2499
rect 91376 2456 91428 2465
rect 102876 2456 102928 2508
rect 86960 2388 87012 2440
rect 75736 2320 75788 2372
rect 80888 2320 80940 2372
rect 74632 2252 74684 2304
rect 75000 2252 75052 2304
rect 88800 2320 88852 2372
rect 84476 2252 84528 2304
rect 88616 2295 88668 2304
rect 88616 2261 88625 2295
rect 88625 2261 88659 2295
rect 88659 2261 88668 2295
rect 88616 2252 88668 2261
rect 92020 2388 92072 2440
rect 103888 2456 103940 2508
rect 103244 2320 103296 2372
rect 108120 2388 108172 2440
rect 89904 2252 89956 2304
rect 100760 2252 100812 2304
rect 107844 2320 107896 2372
rect 104992 2295 105044 2304
rect 104992 2261 105001 2295
rect 105001 2261 105035 2295
rect 105035 2261 105044 2295
rect 104992 2252 105044 2261
rect 107752 2295 107804 2304
rect 107752 2261 107761 2295
rect 107761 2261 107795 2295
rect 107795 2261 107804 2295
rect 107752 2252 107804 2261
rect 107936 2252 107988 2304
rect 108580 2456 108632 2508
rect 118240 2456 118292 2508
rect 120724 2524 120776 2576
rect 161572 2592 161624 2644
rect 161940 2592 161992 2644
rect 164332 2592 164384 2644
rect 151820 2524 151872 2576
rect 155868 2567 155920 2576
rect 155868 2533 155877 2567
rect 155877 2533 155911 2567
rect 155911 2533 155920 2567
rect 155868 2524 155920 2533
rect 157340 2567 157392 2576
rect 157340 2533 157349 2567
rect 157349 2533 157383 2567
rect 157383 2533 157392 2567
rect 157340 2524 157392 2533
rect 159548 2524 159600 2576
rect 160192 2567 160244 2576
rect 160192 2533 160201 2567
rect 160201 2533 160235 2567
rect 160235 2533 160244 2567
rect 160192 2524 160244 2533
rect 111524 2388 111576 2440
rect 114284 2388 114336 2440
rect 116768 2388 116820 2440
rect 118976 2320 119028 2372
rect 120264 2320 120316 2372
rect 120908 2388 120960 2440
rect 124220 2388 124272 2440
rect 125600 2388 125652 2440
rect 127532 2388 127584 2440
rect 109592 2252 109644 2304
rect 111248 2252 111300 2304
rect 112260 2252 112312 2304
rect 113916 2252 113968 2304
rect 114284 2252 114336 2304
rect 114468 2252 114520 2304
rect 115112 2252 115164 2304
rect 115940 2252 115992 2304
rect 116768 2295 116820 2304
rect 116768 2261 116777 2295
rect 116777 2261 116811 2295
rect 116811 2261 116820 2295
rect 116768 2252 116820 2261
rect 117412 2295 117464 2304
rect 117412 2261 117421 2295
rect 117421 2261 117455 2295
rect 117455 2261 117464 2295
rect 117412 2252 117464 2261
rect 118516 2252 118568 2304
rect 118608 2252 118660 2304
rect 119160 2252 119212 2304
rect 119344 2295 119396 2304
rect 119344 2261 119353 2295
rect 119353 2261 119387 2295
rect 119387 2261 119396 2295
rect 119344 2252 119396 2261
rect 120908 2252 120960 2304
rect 124220 2295 124272 2304
rect 124220 2261 124229 2295
rect 124229 2261 124263 2295
rect 124263 2261 124272 2295
rect 124220 2252 124272 2261
rect 125324 2252 125376 2304
rect 125600 2252 125652 2304
rect 127164 2252 127216 2304
rect 142896 2499 142948 2508
rect 142896 2465 142905 2499
rect 142905 2465 142939 2499
rect 142939 2465 142948 2499
rect 142896 2456 142948 2465
rect 145196 2456 145248 2508
rect 146484 2456 146536 2508
rect 147772 2499 147824 2508
rect 147772 2465 147781 2499
rect 147781 2465 147815 2499
rect 147815 2465 147824 2499
rect 147772 2456 147824 2465
rect 149336 2456 149388 2508
rect 149428 2456 149480 2508
rect 152096 2456 152148 2508
rect 164516 2456 164568 2508
rect 130108 2388 130160 2440
rect 131120 2388 131172 2440
rect 134248 2388 134300 2440
rect 131028 2320 131080 2372
rect 135996 2388 136048 2440
rect 128176 2252 128228 2304
rect 129004 2252 129056 2304
rect 133052 2252 133104 2304
rect 134156 2295 134208 2304
rect 134156 2261 134165 2295
rect 134165 2261 134199 2295
rect 134199 2261 134208 2295
rect 134156 2252 134208 2261
rect 137468 2388 137520 2440
rect 138664 2431 138716 2440
rect 138664 2397 138673 2431
rect 138673 2397 138707 2431
rect 138707 2397 138716 2431
rect 138664 2388 138716 2397
rect 139308 2388 139360 2440
rect 139584 2388 139636 2440
rect 138020 2363 138072 2372
rect 136640 2252 136692 2304
rect 137652 2295 137704 2304
rect 137652 2261 137661 2295
rect 137661 2261 137695 2295
rect 137695 2261 137704 2295
rect 137652 2252 137704 2261
rect 138020 2329 138029 2363
rect 138029 2329 138063 2363
rect 138063 2329 138072 2363
rect 138020 2320 138072 2329
rect 140872 2320 140924 2372
rect 140780 2252 140832 2304
rect 146300 2431 146352 2440
rect 146300 2397 146309 2431
rect 146309 2397 146343 2431
rect 146343 2397 146352 2431
rect 146300 2388 146352 2397
rect 147036 2388 147088 2440
rect 150900 2431 150952 2440
rect 147772 2320 147824 2372
rect 145196 2252 145248 2304
rect 145564 2252 145616 2304
rect 145932 2252 145984 2304
rect 149060 2252 149112 2304
rect 149888 2252 149940 2304
rect 150900 2397 150909 2431
rect 150909 2397 150943 2431
rect 150943 2397 150952 2431
rect 150900 2388 150952 2397
rect 151820 2388 151872 2440
rect 155500 2388 155552 2440
rect 151176 2320 151228 2372
rect 156236 2388 156288 2440
rect 158444 2388 158496 2440
rect 159364 2431 159416 2440
rect 159364 2397 159373 2431
rect 159373 2397 159407 2431
rect 159407 2397 159416 2431
rect 159364 2388 159416 2397
rect 161020 2388 161072 2440
rect 162216 2388 162268 2440
rect 164608 2431 164660 2440
rect 164608 2397 164617 2431
rect 164617 2397 164651 2431
rect 164651 2397 164660 2431
rect 164608 2388 164660 2397
rect 161572 2320 161624 2372
rect 165804 2320 165856 2372
rect 150716 2252 150768 2304
rect 154396 2252 154448 2304
rect 154764 2252 154816 2304
rect 155224 2295 155276 2304
rect 155224 2261 155233 2295
rect 155233 2261 155267 2295
rect 155267 2261 155276 2295
rect 155224 2252 155276 2261
rect 157708 2295 157760 2304
rect 157708 2261 157717 2295
rect 157717 2261 157751 2295
rect 157751 2261 157760 2295
rect 157708 2252 157760 2261
rect 160284 2252 160336 2304
rect 160652 2295 160704 2304
rect 160652 2261 160661 2295
rect 160661 2261 160695 2295
rect 160695 2261 160704 2295
rect 160652 2252 160704 2261
rect 164148 2252 164200 2304
rect 56667 2150 56719 2202
rect 56731 2150 56783 2202
rect 56795 2150 56847 2202
rect 56859 2150 56911 2202
rect 113088 2150 113140 2202
rect 113152 2150 113204 2202
rect 113216 2150 113268 2202
rect 113280 2150 113332 2202
rect 6276 2091 6328 2100
rect 6276 2057 6285 2091
rect 6285 2057 6319 2091
rect 6319 2057 6328 2091
rect 6276 2048 6328 2057
rect 7288 2048 7340 2100
rect 12164 2048 12216 2100
rect 18512 2048 18564 2100
rect 19616 2048 19668 2100
rect 42616 2048 42668 2100
rect 42800 2091 42852 2100
rect 42800 2057 42809 2091
rect 42809 2057 42843 2091
rect 42843 2057 42852 2091
rect 42800 2048 42852 2057
rect 2964 1980 3016 2032
rect 3056 1912 3108 1964
rect 3240 1887 3292 1896
rect 3240 1853 3249 1887
rect 3249 1853 3283 1887
rect 3283 1853 3292 1887
rect 3240 1844 3292 1853
rect 5172 1912 5224 1964
rect 2780 1776 2832 1828
rect 7196 1844 7248 1896
rect 8392 1912 8444 1964
rect 9220 1887 9272 1896
rect 9220 1853 9229 1887
rect 9229 1853 9263 1887
rect 9263 1853 9272 1887
rect 9220 1844 9272 1853
rect 10324 1980 10376 2032
rect 32496 1980 32548 2032
rect 32680 1980 32732 2032
rect 38476 1980 38528 2032
rect 38568 1980 38620 2032
rect 41328 1980 41380 2032
rect 41420 1980 41472 2032
rect 10784 1955 10836 1964
rect 10784 1921 10793 1955
rect 10793 1921 10827 1955
rect 10827 1921 10836 1955
rect 10784 1912 10836 1921
rect 15384 1912 15436 1964
rect 11152 1887 11204 1896
rect 11152 1853 11161 1887
rect 11161 1853 11195 1887
rect 11195 1853 11204 1887
rect 11152 1844 11204 1853
rect 15108 1887 15160 1896
rect 15108 1853 15117 1887
rect 15117 1853 15151 1887
rect 15151 1853 15160 1887
rect 15108 1844 15160 1853
rect 19800 1844 19852 1896
rect 21272 1912 21324 1964
rect 22560 1844 22612 1896
rect 23664 1887 23716 1896
rect 23664 1853 23673 1887
rect 23673 1853 23707 1887
rect 23707 1853 23716 1887
rect 23664 1844 23716 1853
rect 25044 1912 25096 1964
rect 26240 1912 26292 1964
rect 26792 1912 26844 1964
rect 4068 1708 4120 1760
rect 11796 1776 11848 1828
rect 13820 1776 13872 1828
rect 5172 1751 5224 1760
rect 5172 1717 5181 1751
rect 5181 1717 5215 1751
rect 5215 1717 5224 1751
rect 5172 1708 5224 1717
rect 7564 1708 7616 1760
rect 8668 1708 8720 1760
rect 21272 1751 21324 1760
rect 21272 1717 21281 1751
rect 21281 1717 21315 1751
rect 21315 1717 21324 1751
rect 21272 1708 21324 1717
rect 22560 1751 22612 1760
rect 22560 1717 22569 1751
rect 22569 1717 22603 1751
rect 22603 1717 22612 1751
rect 22560 1708 22612 1717
rect 22744 1776 22796 1828
rect 26332 1844 26384 1896
rect 26608 1844 26660 1896
rect 28816 1912 28868 1964
rect 28264 1844 28316 1896
rect 30104 1955 30156 1964
rect 30104 1921 30113 1955
rect 30113 1921 30147 1955
rect 30147 1921 30156 1955
rect 30472 1955 30524 1964
rect 30104 1912 30156 1921
rect 30472 1921 30481 1955
rect 30481 1921 30515 1955
rect 30515 1921 30524 1955
rect 30472 1912 30524 1921
rect 36636 1912 36688 1964
rect 36728 1912 36780 1964
rect 41604 1912 41656 1964
rect 43536 2048 43588 2100
rect 44180 2091 44232 2100
rect 44180 2057 44189 2091
rect 44189 2057 44223 2091
rect 44223 2057 44232 2091
rect 44180 2048 44232 2057
rect 44272 2048 44324 2100
rect 47308 2048 47360 2100
rect 47584 2048 47636 2100
rect 49056 2048 49108 2100
rect 51080 2048 51132 2100
rect 51264 2048 51316 2100
rect 52460 2048 52512 2100
rect 53104 2048 53156 2100
rect 55496 2048 55548 2100
rect 47216 1980 47268 2032
rect 47676 1980 47728 2032
rect 43628 1912 43680 1964
rect 44180 1912 44232 1964
rect 45100 1912 45152 1964
rect 46112 1955 46164 1964
rect 46112 1921 46121 1955
rect 46121 1921 46155 1955
rect 46155 1921 46164 1955
rect 46112 1912 46164 1921
rect 46480 1912 46532 1964
rect 46848 1912 46900 1964
rect 47584 1912 47636 1964
rect 48136 1912 48188 1964
rect 48688 1912 48740 1964
rect 49424 1980 49476 2032
rect 50252 1980 50304 2032
rect 53840 1980 53892 2032
rect 54116 1980 54168 2032
rect 60004 2048 60056 2100
rect 60372 2091 60424 2100
rect 60372 2057 60381 2091
rect 60381 2057 60415 2091
rect 60415 2057 60424 2091
rect 60372 2048 60424 2057
rect 55864 1980 55916 2032
rect 51908 1912 51960 1964
rect 53656 1955 53708 1964
rect 33600 1844 33652 1896
rect 35348 1844 35400 1896
rect 37004 1844 37056 1896
rect 37280 1844 37332 1896
rect 41052 1844 41104 1896
rect 41144 1844 41196 1896
rect 50712 1844 50764 1896
rect 26240 1708 26292 1760
rect 29000 1708 29052 1760
rect 33508 1776 33560 1828
rect 36452 1776 36504 1828
rect 51448 1844 51500 1896
rect 52184 1887 52236 1896
rect 52184 1853 52193 1887
rect 52193 1853 52227 1887
rect 52227 1853 52236 1887
rect 52184 1844 52236 1853
rect 53656 1921 53665 1955
rect 53665 1921 53699 1955
rect 53699 1921 53708 1955
rect 53656 1912 53708 1921
rect 55220 1955 55272 1964
rect 55220 1921 55229 1955
rect 55229 1921 55263 1955
rect 55263 1921 55272 1955
rect 55220 1912 55272 1921
rect 55956 1912 56008 1964
rect 56324 1980 56376 2032
rect 60832 2048 60884 2100
rect 63776 2048 63828 2100
rect 64696 2048 64748 2100
rect 65064 2048 65116 2100
rect 66812 2091 66864 2100
rect 66812 2057 66821 2091
rect 66821 2057 66855 2091
rect 66855 2057 66864 2091
rect 66812 2048 66864 2057
rect 66904 2048 66956 2100
rect 67732 2048 67784 2100
rect 57704 1912 57756 1964
rect 57888 1955 57940 1964
rect 57888 1921 57897 1955
rect 57897 1921 57931 1955
rect 57931 1921 57940 1955
rect 57888 1912 57940 1921
rect 58440 1912 58492 1964
rect 58808 1912 58860 1964
rect 36820 1708 36872 1760
rect 37096 1708 37148 1760
rect 38108 1708 38160 1760
rect 38568 1708 38620 1760
rect 38660 1708 38712 1760
rect 39028 1708 39080 1760
rect 41328 1708 41380 1760
rect 43628 1708 43680 1760
rect 43720 1708 43772 1760
rect 45468 1708 45520 1760
rect 47492 1708 47544 1760
rect 49056 1708 49108 1760
rect 49148 1708 49200 1760
rect 50620 1708 50672 1760
rect 50712 1708 50764 1760
rect 51816 1776 51868 1828
rect 54944 1844 54996 1896
rect 57336 1844 57388 1896
rect 57980 1844 58032 1896
rect 60372 1912 60424 1964
rect 59912 1844 59964 1896
rect 60740 1912 60792 1964
rect 61016 1844 61068 1896
rect 61568 1912 61620 1964
rect 61752 1980 61804 2032
rect 63684 2023 63736 2032
rect 63684 1989 63693 2023
rect 63693 1989 63727 2023
rect 63727 1989 63736 2023
rect 63684 1980 63736 1989
rect 65340 1980 65392 2032
rect 65432 1980 65484 2032
rect 69296 2048 69348 2100
rect 71044 2091 71096 2100
rect 71044 2057 71053 2091
rect 71053 2057 71087 2091
rect 71087 2057 71096 2091
rect 71044 2048 71096 2057
rect 73252 2048 73304 2100
rect 73712 2048 73764 2100
rect 77576 2091 77628 2100
rect 77576 2057 77585 2091
rect 77585 2057 77619 2091
rect 77619 2057 77628 2091
rect 77576 2048 77628 2057
rect 78036 2091 78088 2100
rect 78036 2057 78045 2091
rect 78045 2057 78079 2091
rect 78079 2057 78088 2091
rect 78036 2048 78088 2057
rect 79140 2091 79192 2100
rect 79140 2057 79149 2091
rect 79149 2057 79183 2091
rect 79183 2057 79192 2091
rect 79140 2048 79192 2057
rect 79324 2048 79376 2100
rect 80888 2048 80940 2100
rect 81348 2048 81400 2100
rect 82820 2048 82872 2100
rect 83096 2091 83148 2100
rect 83096 2057 83105 2091
rect 83105 2057 83139 2091
rect 83139 2057 83148 2091
rect 83096 2048 83148 2057
rect 84752 2091 84804 2100
rect 84752 2057 84761 2091
rect 84761 2057 84795 2091
rect 84795 2057 84804 2091
rect 84752 2048 84804 2057
rect 85764 2091 85816 2100
rect 85764 2057 85773 2091
rect 85773 2057 85807 2091
rect 85807 2057 85816 2091
rect 85764 2048 85816 2057
rect 88892 2091 88944 2100
rect 88892 2057 88901 2091
rect 88901 2057 88935 2091
rect 88935 2057 88944 2091
rect 88892 2048 88944 2057
rect 102324 2048 102376 2100
rect 103336 2048 103388 2100
rect 106556 2091 106608 2100
rect 106556 2057 106565 2091
rect 106565 2057 106599 2091
rect 106599 2057 106608 2091
rect 106556 2048 106608 2057
rect 107016 2048 107068 2100
rect 108120 2048 108172 2100
rect 62488 1955 62540 1964
rect 62488 1921 62497 1955
rect 62497 1921 62531 1955
rect 62531 1921 62540 1955
rect 62856 1955 62908 1964
rect 62488 1912 62540 1921
rect 62856 1921 62865 1955
rect 62865 1921 62899 1955
rect 62899 1921 62908 1955
rect 62856 1912 62908 1921
rect 63500 1912 63552 1964
rect 65616 1912 65668 1964
rect 67364 1912 67416 1964
rect 51264 1708 51316 1760
rect 57704 1776 57756 1828
rect 62212 1776 62264 1828
rect 62672 1844 62724 1896
rect 63040 1844 63092 1896
rect 64604 1844 64656 1896
rect 66812 1844 66864 1896
rect 68100 1955 68152 1964
rect 68100 1921 68109 1955
rect 68109 1921 68143 1955
rect 68143 1921 68152 1955
rect 68100 1912 68152 1921
rect 72884 1980 72936 2032
rect 72976 1980 73028 2032
rect 73896 1980 73948 2032
rect 88616 1980 88668 2032
rect 100668 1980 100720 2032
rect 70308 1912 70360 1964
rect 70952 1955 71004 1964
rect 70952 1921 70961 1955
rect 70961 1921 70995 1955
rect 70995 1921 71004 1955
rect 70952 1912 71004 1921
rect 72516 1912 72568 1964
rect 69204 1844 69256 1896
rect 72424 1887 72476 1896
rect 72424 1853 72433 1887
rect 72433 1853 72467 1887
rect 72467 1853 72476 1887
rect 72424 1844 72476 1853
rect 53656 1708 53708 1760
rect 55404 1708 55456 1760
rect 55588 1751 55640 1760
rect 55588 1717 55597 1751
rect 55597 1717 55631 1751
rect 55631 1717 55640 1751
rect 55588 1708 55640 1717
rect 56140 1708 56192 1760
rect 56508 1708 56560 1760
rect 56968 1708 57020 1760
rect 57796 1708 57848 1760
rect 60096 1708 60148 1760
rect 62120 1708 62172 1760
rect 74632 1912 74684 1964
rect 75644 1912 75696 1964
rect 75092 1887 75144 1896
rect 75092 1853 75101 1887
rect 75101 1853 75135 1887
rect 75135 1853 75144 1887
rect 75092 1844 75144 1853
rect 75920 1844 75972 1896
rect 78588 1912 78640 1964
rect 79048 1955 79100 1964
rect 79048 1921 79057 1955
rect 79057 1921 79091 1955
rect 79091 1921 79100 1955
rect 79048 1912 79100 1921
rect 81348 1955 81400 1964
rect 81072 1844 81124 1896
rect 81348 1921 81357 1955
rect 81357 1921 81391 1955
rect 81391 1921 81400 1955
rect 81348 1912 81400 1921
rect 82176 1955 82228 1964
rect 82176 1921 82185 1955
rect 82185 1921 82219 1955
rect 82219 1921 82228 1955
rect 82176 1912 82228 1921
rect 84660 1955 84712 1964
rect 84660 1921 84669 1955
rect 84669 1921 84703 1955
rect 84703 1921 84712 1955
rect 84660 1912 84712 1921
rect 85672 1955 85724 1964
rect 85672 1921 85681 1955
rect 85681 1921 85715 1955
rect 85715 1921 85724 1955
rect 85672 1912 85724 1921
rect 86316 1912 86368 1964
rect 87236 1912 87288 1964
rect 88432 1912 88484 1964
rect 89260 1912 89312 1964
rect 91928 1955 91980 1964
rect 91928 1921 91937 1955
rect 91937 1921 91971 1955
rect 91971 1921 91980 1955
rect 91928 1912 91980 1921
rect 81256 1844 81308 1896
rect 83464 1887 83516 1896
rect 83464 1853 83473 1887
rect 83473 1853 83507 1887
rect 83507 1853 83516 1887
rect 83464 1844 83516 1853
rect 84568 1844 84620 1896
rect 88156 1819 88208 1828
rect 66628 1708 66680 1760
rect 66720 1708 66772 1760
rect 67272 1708 67324 1760
rect 67732 1708 67784 1760
rect 70032 1708 70084 1760
rect 71504 1708 71556 1760
rect 73620 1708 73672 1760
rect 74172 1708 74224 1760
rect 74264 1708 74316 1760
rect 80520 1708 80572 1760
rect 88156 1785 88165 1819
rect 88165 1785 88199 1819
rect 88199 1785 88208 1819
rect 88156 1776 88208 1785
rect 91284 1844 91336 1896
rect 95148 1776 95200 1828
rect 96620 1776 96672 1828
rect 97724 1776 97776 1828
rect 104348 1912 104400 1964
rect 104900 1980 104952 2032
rect 117780 2023 117832 2032
rect 105268 1955 105320 1964
rect 105268 1921 105277 1955
rect 105277 1921 105311 1955
rect 105311 1921 105320 1955
rect 105268 1912 105320 1921
rect 106924 1912 106976 1964
rect 107752 1955 107804 1964
rect 107752 1921 107761 1955
rect 107761 1921 107795 1955
rect 107795 1921 107804 1955
rect 107752 1912 107804 1921
rect 109040 1912 109092 1964
rect 109592 1912 109644 1964
rect 111064 1912 111116 1964
rect 111340 1955 111392 1964
rect 111340 1921 111349 1955
rect 111349 1921 111383 1955
rect 111383 1921 111392 1955
rect 111340 1912 111392 1921
rect 112168 1955 112220 1964
rect 112168 1921 112177 1955
rect 112177 1921 112211 1955
rect 112211 1921 112220 1955
rect 112168 1912 112220 1921
rect 112904 1912 112956 1964
rect 104808 1844 104860 1896
rect 108580 1844 108632 1896
rect 108672 1844 108724 1896
rect 109776 1887 109828 1896
rect 109776 1853 109785 1887
rect 109785 1853 109819 1887
rect 109819 1853 109828 1887
rect 109776 1844 109828 1853
rect 110696 1844 110748 1896
rect 111248 1844 111300 1896
rect 112076 1844 112128 1896
rect 112260 1844 112312 1896
rect 113456 1844 113508 1896
rect 113824 1887 113876 1896
rect 113824 1853 113833 1887
rect 113833 1853 113867 1887
rect 113867 1853 113876 1887
rect 113824 1844 113876 1853
rect 117780 1989 117789 2023
rect 117789 1989 117823 2023
rect 117823 1989 117832 2023
rect 117780 1980 117832 1989
rect 117872 1980 117924 2032
rect 118792 1980 118844 2032
rect 119160 1980 119212 2032
rect 120540 1980 120592 2032
rect 120632 1980 120684 2032
rect 121184 1980 121236 2032
rect 122932 2023 122984 2032
rect 115572 1912 115624 1964
rect 116216 1955 116268 1964
rect 116216 1921 116225 1955
rect 116225 1921 116259 1955
rect 116259 1921 116268 1955
rect 116216 1912 116268 1921
rect 117688 1955 117740 1964
rect 117688 1921 117697 1955
rect 117697 1921 117731 1955
rect 117731 1921 117740 1955
rect 117688 1912 117740 1921
rect 116768 1844 116820 1896
rect 118608 1912 118660 1964
rect 120172 1912 120224 1964
rect 121000 1955 121052 1964
rect 121000 1921 121009 1955
rect 121009 1921 121043 1955
rect 121043 1921 121052 1955
rect 121000 1912 121052 1921
rect 122380 1912 122432 1964
rect 122012 1844 122064 1896
rect 122932 1989 122941 2023
rect 122941 1989 122975 2023
rect 122975 1989 122984 2023
rect 122932 1980 122984 1989
rect 124680 2023 124732 2032
rect 124680 1989 124689 2023
rect 124689 1989 124723 2023
rect 124723 1989 124732 2023
rect 124680 1980 124732 1989
rect 125600 1980 125652 2032
rect 126796 1980 126848 2032
rect 122840 1955 122892 1964
rect 122840 1921 122849 1955
rect 122849 1921 122883 1955
rect 122883 1921 122892 1955
rect 122840 1912 122892 1921
rect 130660 1980 130712 2032
rect 130936 2048 130988 2100
rect 138664 2048 138716 2100
rect 139400 2048 139452 2100
rect 139584 2091 139636 2100
rect 139584 2057 139593 2091
rect 139593 2057 139627 2091
rect 139627 2057 139636 2091
rect 139584 2048 139636 2057
rect 141148 2091 141200 2100
rect 141148 2057 141157 2091
rect 141157 2057 141191 2091
rect 141191 2057 141200 2091
rect 141148 2048 141200 2057
rect 146392 2048 146444 2100
rect 150992 2048 151044 2100
rect 153752 2091 153804 2100
rect 153752 2057 153761 2091
rect 153761 2057 153795 2091
rect 153795 2057 153804 2091
rect 153752 2048 153804 2057
rect 154856 2048 154908 2100
rect 155776 2091 155828 2100
rect 155776 2057 155785 2091
rect 155785 2057 155819 2091
rect 155819 2057 155828 2091
rect 155776 2048 155828 2057
rect 160928 2091 160980 2100
rect 160928 2057 160937 2091
rect 160937 2057 160971 2091
rect 160971 2057 160980 2091
rect 160928 2048 160980 2057
rect 162400 2048 162452 2100
rect 164976 2048 165028 2100
rect 127072 1955 127124 1964
rect 127072 1921 127081 1955
rect 127081 1921 127115 1955
rect 127115 1921 127124 1955
rect 127072 1912 127124 1921
rect 128268 1912 128320 1964
rect 131212 1912 131264 1964
rect 126152 1844 126204 1896
rect 126612 1887 126664 1896
rect 126612 1853 126621 1887
rect 126621 1853 126655 1887
rect 126655 1853 126664 1887
rect 126612 1844 126664 1853
rect 83556 1708 83608 1760
rect 85580 1708 85632 1760
rect 100024 1708 100076 1760
rect 102416 1751 102468 1760
rect 102416 1717 102425 1751
rect 102425 1717 102459 1751
rect 102459 1717 102468 1751
rect 102416 1708 102468 1717
rect 102508 1708 102560 1760
rect 106924 1708 106976 1760
rect 110604 1708 110656 1760
rect 111616 1751 111668 1760
rect 111616 1717 111625 1751
rect 111625 1717 111659 1751
rect 111659 1717 111668 1751
rect 111616 1708 111668 1717
rect 112260 1751 112312 1760
rect 112260 1717 112269 1751
rect 112269 1717 112303 1751
rect 112303 1717 112312 1751
rect 112260 1708 112312 1717
rect 117780 1776 117832 1828
rect 128544 1776 128596 1828
rect 131028 1844 131080 1896
rect 133696 1887 133748 1896
rect 133696 1853 133705 1887
rect 133705 1853 133739 1887
rect 133739 1853 133748 1887
rect 133696 1844 133748 1853
rect 135352 1887 135404 1896
rect 135352 1853 135361 1887
rect 135361 1853 135395 1887
rect 135395 1853 135404 1887
rect 135352 1844 135404 1853
rect 138940 1980 138992 2032
rect 139308 2023 139360 2032
rect 139308 1989 139317 2023
rect 139317 1989 139351 2023
rect 139351 1989 139360 2023
rect 139308 1980 139360 1989
rect 144828 1980 144880 2032
rect 137284 1844 137336 1896
rect 137560 1844 137612 1896
rect 138756 1912 138808 1964
rect 139492 1955 139544 1964
rect 139492 1921 139501 1955
rect 139501 1921 139535 1955
rect 139535 1921 139544 1955
rect 139492 1912 139544 1921
rect 141608 1912 141660 1964
rect 144276 1955 144328 1964
rect 143172 1887 143224 1896
rect 143172 1853 143181 1887
rect 143181 1853 143215 1887
rect 143215 1853 143224 1887
rect 143172 1844 143224 1853
rect 144276 1921 144285 1955
rect 144285 1921 144319 1955
rect 144319 1921 144328 1955
rect 144276 1912 144328 1921
rect 146668 1912 146720 1964
rect 147864 1887 147916 1896
rect 147864 1853 147873 1887
rect 147873 1853 147907 1887
rect 147907 1853 147916 1887
rect 147864 1844 147916 1853
rect 154580 1980 154632 2032
rect 149152 1955 149204 1964
rect 149152 1921 149161 1955
rect 149161 1921 149195 1955
rect 149195 1921 149204 1955
rect 149152 1912 149204 1921
rect 150256 1955 150308 1964
rect 150256 1921 150265 1955
rect 150265 1921 150299 1955
rect 150299 1921 150308 1955
rect 150256 1912 150308 1921
rect 152648 1955 152700 1964
rect 152648 1921 152657 1955
rect 152657 1921 152691 1955
rect 152691 1921 152700 1955
rect 152648 1912 152700 1921
rect 153660 1955 153712 1964
rect 153660 1921 153669 1955
rect 153669 1921 153703 1955
rect 153703 1921 153712 1955
rect 153660 1912 153712 1921
rect 154672 1955 154724 1964
rect 154672 1921 154681 1955
rect 154681 1921 154715 1955
rect 154715 1921 154724 1955
rect 154672 1912 154724 1921
rect 155868 1912 155920 1964
rect 156696 1955 156748 1964
rect 156696 1921 156705 1955
rect 156705 1921 156739 1955
rect 156739 1921 156748 1955
rect 156696 1912 156748 1921
rect 158168 1912 158220 1964
rect 159824 1955 159876 1964
rect 159824 1921 159833 1955
rect 159833 1921 159867 1955
rect 159867 1921 159876 1955
rect 159824 1912 159876 1921
rect 160836 1955 160888 1964
rect 160836 1921 160845 1955
rect 160845 1921 160879 1955
rect 160879 1921 160888 1955
rect 160836 1912 160888 1921
rect 161940 1955 161992 1964
rect 161940 1921 161949 1955
rect 161949 1921 161983 1955
rect 161983 1921 161992 1955
rect 161940 1912 161992 1921
rect 163964 1912 164016 1964
rect 164884 1955 164936 1964
rect 164884 1921 164893 1955
rect 164893 1921 164927 1955
rect 164927 1921 164936 1955
rect 164884 1912 164936 1921
rect 166080 1912 166132 1964
rect 166908 1912 166960 1964
rect 166172 1844 166224 1896
rect 166540 1844 166592 1896
rect 115112 1708 115164 1760
rect 118240 1708 118292 1760
rect 118424 1751 118476 1760
rect 118424 1717 118433 1751
rect 118433 1717 118467 1751
rect 118467 1717 118476 1751
rect 118424 1708 118476 1717
rect 118976 1708 119028 1760
rect 119712 1708 119764 1760
rect 119896 1751 119948 1760
rect 119896 1717 119905 1751
rect 119905 1717 119939 1751
rect 119939 1717 119948 1751
rect 119896 1708 119948 1717
rect 120172 1708 120224 1760
rect 120356 1708 120408 1760
rect 121184 1708 121236 1760
rect 123944 1751 123996 1760
rect 123944 1717 123953 1751
rect 123953 1717 123987 1751
rect 123987 1717 123996 1751
rect 123944 1708 123996 1717
rect 126060 1708 126112 1760
rect 126244 1708 126296 1760
rect 129188 1751 129240 1760
rect 129188 1717 129197 1751
rect 129197 1717 129231 1751
rect 129231 1717 129240 1751
rect 129188 1708 129240 1717
rect 132500 1708 132552 1760
rect 133420 1708 133472 1760
rect 134156 1708 134208 1760
rect 135904 1751 135956 1760
rect 135904 1717 135913 1751
rect 135913 1717 135947 1751
rect 135947 1717 135956 1751
rect 135904 1708 135956 1717
rect 137836 1708 137888 1760
rect 139492 1708 139544 1760
rect 141056 1708 141108 1760
rect 155868 1708 155920 1760
rect 156880 1708 156932 1760
rect 158352 1751 158404 1760
rect 158352 1717 158361 1751
rect 158361 1717 158395 1751
rect 158395 1717 158404 1751
rect 158352 1708 158404 1717
rect 158720 1751 158772 1760
rect 158720 1717 158729 1751
rect 158729 1717 158763 1751
rect 158763 1717 158772 1751
rect 158720 1708 158772 1717
rect 159640 1751 159692 1760
rect 159640 1717 159649 1751
rect 159649 1717 159683 1751
rect 159683 1717 159692 1751
rect 159640 1708 159692 1717
rect 28456 1606 28508 1658
rect 28520 1606 28572 1658
rect 28584 1606 28636 1658
rect 28648 1606 28700 1658
rect 84878 1606 84930 1658
rect 84942 1606 84994 1658
rect 85006 1606 85058 1658
rect 85070 1606 85122 1658
rect 95056 1640 95108 1692
rect 96988 1640 97040 1692
rect 100300 1640 100352 1692
rect 95976 1572 96028 1624
rect 99472 1572 99524 1624
rect 100116 1572 100168 1624
rect 141299 1606 141351 1658
rect 141363 1606 141415 1658
rect 141427 1606 141479 1658
rect 141491 1606 141543 1658
rect 2044 1504 2096 1556
rect 3056 1504 3108 1556
rect 3240 1504 3292 1556
rect 7196 1547 7248 1556
rect 7196 1513 7205 1547
rect 7205 1513 7239 1547
rect 7239 1513 7248 1547
rect 7196 1504 7248 1513
rect 9220 1547 9272 1556
rect 9220 1513 9229 1547
rect 9229 1513 9263 1547
rect 9263 1513 9272 1547
rect 9220 1504 9272 1513
rect 1676 1436 1728 1488
rect 7472 1436 7524 1488
rect 2412 1368 2464 1420
rect 10784 1504 10836 1556
rect 15108 1547 15160 1556
rect 15108 1513 15117 1547
rect 15117 1513 15151 1547
rect 15151 1513 15160 1547
rect 15108 1504 15160 1513
rect 18604 1436 18656 1488
rect 22192 1504 22244 1556
rect 25044 1547 25096 1556
rect 25044 1513 25053 1547
rect 25053 1513 25087 1547
rect 25087 1513 25096 1547
rect 25044 1504 25096 1513
rect 26792 1547 26844 1556
rect 26792 1513 26801 1547
rect 26801 1513 26835 1547
rect 26835 1513 26844 1547
rect 26792 1504 26844 1513
rect 28264 1547 28316 1556
rect 28264 1513 28273 1547
rect 28273 1513 28307 1547
rect 28307 1513 28316 1547
rect 28264 1504 28316 1513
rect 30472 1547 30524 1556
rect 22100 1436 22152 1488
rect 24032 1436 24084 1488
rect 11612 1411 11664 1420
rect 11612 1377 11621 1411
rect 11621 1377 11655 1411
rect 11655 1377 11664 1411
rect 11612 1368 11664 1377
rect 11796 1368 11848 1420
rect 20720 1368 20772 1420
rect 22560 1411 22612 1420
rect 22560 1377 22569 1411
rect 22569 1377 22603 1411
rect 22603 1377 22612 1411
rect 22560 1368 22612 1377
rect 7748 1343 7800 1352
rect 7748 1309 7757 1343
rect 7757 1309 7791 1343
rect 7791 1309 7800 1343
rect 7748 1300 7800 1309
rect 11152 1300 11204 1352
rect 6000 1164 6052 1216
rect 6276 1207 6328 1216
rect 6276 1173 6285 1207
rect 6285 1173 6319 1207
rect 6319 1173 6328 1207
rect 6276 1164 6328 1173
rect 6736 1207 6788 1216
rect 6736 1173 6745 1207
rect 6745 1173 6779 1207
rect 6779 1173 6788 1207
rect 6736 1164 6788 1173
rect 8392 1164 8444 1216
rect 15108 1300 15160 1352
rect 18880 1343 18932 1352
rect 12808 1164 12860 1216
rect 12992 1207 13044 1216
rect 12992 1173 13001 1207
rect 13001 1173 13035 1207
rect 13035 1173 13044 1207
rect 12992 1164 13044 1173
rect 18880 1309 18889 1343
rect 18889 1309 18923 1343
rect 18923 1309 18932 1343
rect 18880 1300 18932 1309
rect 23480 1300 23532 1352
rect 23572 1300 23624 1352
rect 17500 1232 17552 1284
rect 18696 1232 18748 1284
rect 28080 1368 28132 1420
rect 26148 1343 26200 1352
rect 26148 1309 26157 1343
rect 26157 1309 26191 1343
rect 26191 1309 26200 1343
rect 26148 1300 26200 1309
rect 26516 1343 26568 1352
rect 26516 1309 26525 1343
rect 26525 1309 26559 1343
rect 26559 1309 26568 1343
rect 26516 1300 26568 1309
rect 27344 1343 27396 1352
rect 27344 1309 27353 1343
rect 27353 1309 27387 1343
rect 27387 1309 27396 1343
rect 27344 1300 27396 1309
rect 27712 1300 27764 1352
rect 28356 1343 28408 1352
rect 28356 1309 28365 1343
rect 28365 1309 28399 1343
rect 28399 1309 28408 1343
rect 28632 1368 28684 1420
rect 30472 1513 30481 1547
rect 30481 1513 30515 1547
rect 30515 1513 30524 1547
rect 30472 1504 30524 1513
rect 30748 1504 30800 1556
rect 32772 1504 32824 1556
rect 33416 1504 33468 1556
rect 40500 1504 40552 1556
rect 40684 1504 40736 1556
rect 41972 1504 42024 1556
rect 42248 1504 42300 1556
rect 46480 1547 46532 1556
rect 46480 1513 46489 1547
rect 46489 1513 46523 1547
rect 46523 1513 46532 1547
rect 46480 1504 46532 1513
rect 30288 1436 30340 1488
rect 33508 1436 33560 1488
rect 33876 1479 33928 1488
rect 33876 1445 33885 1479
rect 33885 1445 33919 1479
rect 33919 1445 33928 1479
rect 33876 1436 33928 1445
rect 34336 1436 34388 1488
rect 40132 1436 40184 1488
rect 32496 1368 32548 1420
rect 28356 1300 28408 1309
rect 24676 1232 24728 1284
rect 26056 1232 26108 1284
rect 28632 1232 28684 1284
rect 30840 1300 30892 1352
rect 33600 1343 33652 1352
rect 33600 1309 33609 1343
rect 33609 1309 33643 1343
rect 33643 1309 33652 1343
rect 33600 1300 33652 1309
rect 35348 1343 35400 1352
rect 33140 1232 33192 1284
rect 35348 1309 35357 1343
rect 35357 1309 35391 1343
rect 35391 1309 35400 1343
rect 35348 1300 35400 1309
rect 35440 1300 35492 1352
rect 35900 1300 35952 1352
rect 36452 1368 36504 1420
rect 39580 1368 39632 1420
rect 39672 1368 39724 1420
rect 43996 1436 44048 1488
rect 34888 1275 34940 1284
rect 34888 1241 34897 1275
rect 34897 1241 34931 1275
rect 34931 1241 34940 1275
rect 34888 1232 34940 1241
rect 35072 1232 35124 1284
rect 35992 1232 36044 1284
rect 36820 1300 36872 1352
rect 37004 1343 37056 1352
rect 37004 1309 37013 1343
rect 37013 1309 37047 1343
rect 37047 1309 37056 1343
rect 37004 1300 37056 1309
rect 37556 1300 37608 1352
rect 39028 1300 39080 1352
rect 39120 1300 39172 1352
rect 40224 1300 40276 1352
rect 40868 1368 40920 1420
rect 40960 1368 41012 1420
rect 41328 1368 41380 1420
rect 41512 1411 41564 1420
rect 41512 1377 41521 1411
rect 41521 1377 41555 1411
rect 41555 1377 41564 1411
rect 41512 1368 41564 1377
rect 40408 1300 40460 1352
rect 43812 1368 43864 1420
rect 41696 1300 41748 1352
rect 42524 1300 42576 1352
rect 42616 1300 42668 1352
rect 39488 1232 39540 1284
rect 17224 1164 17276 1216
rect 19616 1164 19668 1216
rect 20812 1164 20864 1216
rect 22744 1164 22796 1216
rect 23572 1164 23624 1216
rect 24584 1164 24636 1216
rect 25780 1164 25832 1216
rect 30288 1164 30340 1216
rect 30840 1207 30892 1216
rect 30840 1173 30849 1207
rect 30849 1173 30883 1207
rect 30883 1173 30892 1207
rect 30840 1164 30892 1173
rect 40408 1164 40460 1216
rect 40592 1232 40644 1284
rect 44916 1368 44968 1420
rect 43260 1164 43312 1216
rect 44364 1300 44416 1352
rect 45652 1436 45704 1488
rect 48596 1504 48648 1556
rect 48688 1504 48740 1556
rect 50988 1504 51040 1556
rect 51080 1504 51132 1556
rect 58808 1547 58860 1556
rect 58808 1513 58817 1547
rect 58817 1513 58851 1547
rect 58851 1513 58860 1547
rect 58808 1504 58860 1513
rect 59084 1504 59136 1556
rect 61568 1504 61620 1556
rect 62120 1547 62172 1556
rect 62120 1513 62129 1547
rect 62129 1513 62163 1547
rect 62163 1513 62172 1547
rect 62120 1504 62172 1513
rect 62488 1504 62540 1556
rect 63316 1547 63368 1556
rect 63316 1513 63325 1547
rect 63325 1513 63359 1547
rect 63359 1513 63368 1547
rect 63316 1504 63368 1513
rect 63776 1504 63828 1556
rect 69848 1504 69900 1556
rect 70308 1504 70360 1556
rect 70400 1504 70452 1556
rect 72608 1504 72660 1556
rect 75000 1504 75052 1556
rect 75092 1504 75144 1556
rect 80980 1504 81032 1556
rect 81256 1504 81308 1556
rect 84660 1504 84712 1556
rect 46756 1436 46808 1488
rect 50344 1436 50396 1488
rect 55220 1479 55272 1488
rect 45376 1368 45428 1420
rect 46480 1368 46532 1420
rect 46572 1368 46624 1420
rect 50528 1368 50580 1420
rect 53196 1368 53248 1420
rect 53472 1368 53524 1420
rect 54300 1368 54352 1420
rect 55220 1445 55229 1479
rect 55229 1445 55263 1479
rect 55263 1445 55272 1479
rect 55220 1436 55272 1445
rect 55496 1436 55548 1488
rect 57704 1368 57756 1420
rect 59912 1368 59964 1420
rect 46940 1300 46992 1352
rect 48780 1300 48832 1352
rect 44732 1232 44784 1284
rect 45652 1232 45704 1284
rect 45836 1232 45888 1284
rect 47308 1232 47360 1284
rect 44640 1207 44692 1216
rect 44640 1173 44649 1207
rect 44649 1173 44683 1207
rect 44683 1173 44692 1207
rect 44640 1164 44692 1173
rect 44916 1164 44968 1216
rect 47584 1207 47636 1216
rect 47584 1173 47593 1207
rect 47593 1173 47627 1207
rect 47627 1173 47636 1207
rect 47584 1164 47636 1173
rect 47768 1232 47820 1284
rect 49056 1300 49108 1352
rect 50068 1300 50120 1352
rect 50344 1300 50396 1352
rect 51908 1300 51960 1352
rect 52184 1300 52236 1352
rect 53656 1300 53708 1352
rect 53840 1343 53892 1352
rect 53840 1309 53849 1343
rect 53849 1309 53883 1343
rect 53883 1309 53892 1343
rect 53840 1300 53892 1309
rect 55220 1300 55272 1352
rect 55588 1343 55640 1352
rect 55588 1309 55597 1343
rect 55597 1309 55631 1343
rect 55631 1309 55640 1343
rect 55588 1300 55640 1309
rect 50068 1164 50120 1216
rect 50160 1164 50212 1216
rect 55312 1164 55364 1216
rect 56048 1164 56100 1216
rect 56232 1300 56284 1352
rect 56968 1343 57020 1352
rect 56508 1207 56560 1216
rect 56508 1173 56517 1207
rect 56517 1173 56551 1207
rect 56551 1173 56560 1207
rect 56508 1164 56560 1173
rect 56968 1309 56977 1343
rect 56977 1309 57011 1343
rect 57011 1309 57020 1343
rect 56968 1300 57020 1309
rect 57244 1232 57296 1284
rect 57888 1300 57940 1352
rect 60832 1411 60884 1420
rect 60832 1377 60841 1411
rect 60841 1377 60875 1411
rect 60875 1377 60884 1411
rect 60832 1368 60884 1377
rect 62856 1411 62908 1420
rect 62856 1377 62865 1411
rect 62865 1377 62899 1411
rect 62899 1377 62908 1411
rect 62856 1368 62908 1377
rect 60280 1232 60332 1284
rect 58992 1164 59044 1216
rect 61016 1300 61068 1352
rect 62304 1343 62356 1352
rect 62304 1309 62313 1343
rect 62313 1309 62347 1343
rect 62347 1309 62356 1343
rect 62304 1300 62356 1309
rect 63684 1368 63736 1420
rect 65616 1411 65668 1420
rect 65616 1377 65625 1411
rect 65625 1377 65659 1411
rect 65659 1377 65668 1411
rect 65616 1368 65668 1377
rect 66812 1368 66864 1420
rect 67364 1411 67416 1420
rect 67364 1377 67373 1411
rect 67373 1377 67407 1411
rect 67407 1377 67416 1411
rect 67364 1368 67416 1377
rect 68560 1411 68612 1420
rect 68560 1377 68569 1411
rect 68569 1377 68603 1411
rect 68603 1377 68612 1411
rect 68560 1368 68612 1377
rect 68744 1368 68796 1420
rect 72976 1411 73028 1420
rect 72976 1377 72985 1411
rect 72985 1377 73019 1411
rect 73019 1377 73028 1411
rect 72976 1368 73028 1377
rect 74356 1411 74408 1420
rect 74356 1377 74365 1411
rect 74365 1377 74399 1411
rect 74399 1377 74408 1411
rect 74356 1368 74408 1377
rect 63776 1343 63828 1352
rect 63776 1309 63785 1343
rect 63785 1309 63819 1343
rect 63819 1309 63828 1343
rect 63776 1300 63828 1309
rect 63960 1343 64012 1352
rect 63960 1309 63969 1343
rect 63969 1309 64003 1343
rect 64003 1309 64012 1343
rect 63960 1300 64012 1309
rect 65984 1343 66036 1352
rect 65984 1309 65993 1343
rect 65993 1309 66027 1343
rect 66027 1309 66036 1343
rect 65984 1300 66036 1309
rect 60648 1232 60700 1284
rect 60740 1164 60792 1216
rect 61200 1232 61252 1284
rect 67088 1300 67140 1352
rect 67272 1300 67324 1352
rect 70952 1343 71004 1352
rect 61476 1164 61528 1216
rect 62304 1164 62356 1216
rect 62672 1164 62724 1216
rect 65156 1207 65208 1216
rect 65156 1173 65165 1207
rect 65165 1173 65199 1207
rect 65199 1173 65208 1207
rect 65156 1164 65208 1173
rect 66904 1232 66956 1284
rect 70952 1309 70961 1343
rect 70961 1309 70995 1343
rect 70995 1309 71004 1343
rect 70952 1300 71004 1309
rect 71504 1343 71556 1352
rect 71504 1309 71513 1343
rect 71513 1309 71547 1343
rect 71547 1309 71556 1343
rect 71504 1300 71556 1309
rect 71780 1343 71832 1352
rect 71780 1309 71789 1343
rect 71789 1309 71823 1343
rect 71823 1309 71832 1343
rect 71780 1300 71832 1309
rect 72056 1343 72108 1352
rect 72056 1309 72065 1343
rect 72065 1309 72099 1343
rect 72099 1309 72108 1343
rect 72056 1300 72108 1309
rect 72516 1300 72568 1352
rect 76748 1368 76800 1420
rect 77300 1411 77352 1420
rect 77300 1377 77309 1411
rect 77309 1377 77343 1411
rect 77343 1377 77352 1411
rect 77300 1368 77352 1377
rect 76104 1343 76156 1352
rect 67088 1207 67140 1216
rect 67088 1173 67097 1207
rect 67097 1173 67131 1207
rect 67131 1173 67140 1207
rect 67088 1164 67140 1173
rect 68652 1164 68704 1216
rect 73896 1232 73948 1284
rect 71872 1164 71924 1216
rect 72608 1164 72660 1216
rect 73068 1164 73120 1216
rect 76104 1309 76113 1343
rect 76113 1309 76147 1343
rect 76147 1309 76156 1343
rect 78036 1368 78088 1420
rect 76104 1300 76156 1309
rect 79324 1343 79376 1352
rect 79324 1309 79333 1343
rect 79333 1309 79367 1343
rect 79367 1309 79376 1343
rect 79324 1300 79376 1309
rect 79416 1343 79468 1352
rect 79416 1309 79425 1343
rect 79425 1309 79459 1343
rect 79459 1309 79468 1343
rect 79600 1343 79652 1352
rect 79416 1300 79468 1309
rect 79600 1309 79609 1343
rect 79609 1309 79643 1343
rect 79643 1309 79652 1343
rect 79600 1300 79652 1309
rect 80152 1232 80204 1284
rect 75184 1164 75236 1216
rect 78588 1164 78640 1216
rect 79048 1164 79100 1216
rect 79968 1164 80020 1216
rect 83096 1368 83148 1420
rect 84200 1411 84252 1420
rect 84200 1377 84209 1411
rect 84209 1377 84243 1411
rect 84243 1377 84252 1411
rect 84200 1368 84252 1377
rect 87420 1504 87472 1556
rect 91284 1504 91336 1556
rect 92296 1504 92348 1556
rect 99196 1504 99248 1556
rect 84568 1343 84620 1352
rect 81348 1275 81400 1284
rect 81348 1241 81357 1275
rect 81357 1241 81391 1275
rect 81391 1241 81400 1275
rect 81348 1232 81400 1241
rect 81532 1232 81584 1284
rect 82176 1232 82228 1284
rect 84568 1309 84577 1343
rect 84577 1309 84611 1343
rect 84611 1309 84620 1343
rect 84568 1300 84620 1309
rect 100208 1436 100260 1488
rect 101772 1504 101824 1556
rect 102508 1504 102560 1556
rect 104348 1504 104400 1556
rect 105268 1504 105320 1556
rect 107936 1504 107988 1556
rect 110972 1504 111024 1556
rect 112536 1504 112588 1556
rect 117412 1504 117464 1556
rect 117688 1504 117740 1556
rect 118056 1504 118108 1556
rect 118792 1504 118844 1556
rect 135904 1504 135956 1556
rect 137560 1547 137612 1556
rect 137560 1513 137569 1547
rect 137569 1513 137603 1547
rect 137603 1513 137612 1547
rect 137560 1504 137612 1513
rect 138756 1504 138808 1556
rect 143172 1504 143224 1556
rect 158168 1547 158220 1556
rect 158168 1513 158177 1547
rect 158177 1513 158211 1547
rect 158211 1513 158220 1547
rect 158168 1504 158220 1513
rect 159824 1504 159876 1556
rect 164884 1504 164936 1556
rect 166080 1547 166132 1556
rect 166080 1513 166089 1547
rect 166089 1513 166123 1547
rect 166123 1513 166132 1547
rect 166080 1504 166132 1513
rect 126152 1479 126204 1488
rect 85672 1368 85724 1420
rect 87420 1368 87472 1420
rect 88892 1411 88944 1420
rect 88892 1377 88901 1411
rect 88901 1377 88935 1411
rect 88935 1377 88944 1411
rect 88892 1368 88944 1377
rect 89720 1368 89772 1420
rect 91928 1368 91980 1420
rect 99472 1368 99524 1420
rect 99564 1368 99616 1420
rect 100576 1368 100628 1420
rect 102324 1411 102376 1420
rect 87236 1343 87288 1352
rect 87236 1309 87245 1343
rect 87245 1309 87279 1343
rect 87279 1309 87288 1343
rect 87236 1300 87288 1309
rect 88432 1343 88484 1352
rect 81164 1164 81216 1216
rect 81992 1207 82044 1216
rect 81992 1173 82001 1207
rect 82001 1173 82035 1207
rect 82035 1173 82044 1207
rect 81992 1164 82044 1173
rect 82636 1164 82688 1216
rect 85488 1207 85540 1216
rect 85488 1173 85497 1207
rect 85497 1173 85531 1207
rect 85531 1173 85540 1207
rect 85488 1164 85540 1173
rect 86500 1207 86552 1216
rect 86500 1173 86509 1207
rect 86509 1173 86543 1207
rect 86543 1173 86552 1207
rect 86500 1164 86552 1173
rect 87788 1232 87840 1284
rect 87052 1164 87104 1216
rect 87604 1207 87656 1216
rect 87604 1173 87613 1207
rect 87613 1173 87647 1207
rect 87647 1173 87656 1207
rect 87604 1164 87656 1173
rect 88432 1309 88441 1343
rect 88441 1309 88475 1343
rect 88475 1309 88484 1343
rect 88432 1300 88484 1309
rect 90180 1300 90232 1352
rect 91100 1300 91152 1352
rect 94780 1300 94832 1352
rect 102324 1377 102333 1411
rect 102333 1377 102367 1411
rect 102367 1377 102376 1411
rect 102324 1368 102376 1377
rect 103520 1411 103572 1420
rect 103520 1377 103529 1411
rect 103529 1377 103563 1411
rect 103563 1377 103572 1411
rect 103520 1368 103572 1377
rect 106372 1368 106424 1420
rect 106924 1411 106976 1420
rect 106924 1377 106933 1411
rect 106933 1377 106967 1411
rect 106967 1377 106976 1411
rect 106924 1368 106976 1377
rect 107752 1368 107804 1420
rect 109224 1368 109276 1420
rect 110788 1368 110840 1420
rect 111800 1368 111852 1420
rect 112444 1368 112496 1420
rect 112628 1411 112680 1420
rect 112628 1377 112637 1411
rect 112637 1377 112671 1411
rect 112671 1377 112680 1411
rect 112628 1368 112680 1377
rect 113824 1411 113876 1420
rect 113824 1377 113833 1411
rect 113833 1377 113867 1411
rect 113867 1377 113876 1411
rect 113824 1368 113876 1377
rect 115020 1368 115072 1420
rect 116216 1368 116268 1420
rect 118424 1411 118476 1420
rect 118424 1377 118433 1411
rect 118433 1377 118467 1411
rect 118467 1377 118476 1411
rect 118424 1368 118476 1377
rect 96252 1232 96304 1284
rect 102232 1232 102284 1284
rect 105268 1300 105320 1352
rect 109040 1343 109092 1352
rect 109040 1309 109049 1343
rect 109049 1309 109083 1343
rect 109083 1309 109092 1343
rect 109040 1300 109092 1309
rect 88156 1164 88208 1216
rect 89996 1164 90048 1216
rect 91100 1164 91152 1216
rect 91376 1207 91428 1216
rect 91376 1173 91385 1207
rect 91385 1173 91419 1207
rect 91419 1173 91428 1207
rect 91376 1164 91428 1173
rect 94044 1164 94096 1216
rect 105820 1232 105872 1284
rect 106096 1207 106148 1216
rect 106096 1173 106105 1207
rect 106105 1173 106139 1207
rect 106139 1173 106148 1207
rect 106096 1164 106148 1173
rect 107016 1207 107068 1216
rect 107016 1173 107025 1207
rect 107025 1173 107059 1207
rect 107059 1173 107068 1207
rect 107016 1164 107068 1173
rect 109776 1300 109828 1352
rect 109224 1232 109276 1284
rect 109040 1164 109092 1216
rect 109408 1232 109460 1284
rect 111248 1300 111300 1352
rect 111616 1343 111668 1352
rect 111616 1309 111625 1343
rect 111625 1309 111659 1343
rect 111659 1309 111668 1343
rect 111616 1300 111668 1309
rect 112260 1300 112312 1352
rect 118884 1368 118936 1420
rect 119712 1368 119764 1420
rect 121000 1411 121052 1420
rect 119896 1343 119948 1352
rect 111340 1232 111392 1284
rect 114100 1232 114152 1284
rect 118148 1232 118200 1284
rect 119896 1309 119905 1343
rect 119905 1309 119939 1343
rect 119939 1309 119948 1343
rect 119896 1300 119948 1309
rect 120356 1343 120408 1352
rect 120356 1309 120365 1343
rect 120365 1309 120399 1343
rect 120399 1309 120408 1343
rect 120356 1300 120408 1309
rect 121000 1377 121009 1411
rect 121009 1377 121043 1411
rect 121043 1377 121052 1411
rect 121000 1368 121052 1377
rect 123944 1411 123996 1420
rect 122288 1343 122340 1352
rect 122288 1309 122297 1343
rect 122297 1309 122331 1343
rect 122331 1309 122340 1343
rect 122288 1300 122340 1309
rect 123944 1377 123953 1411
rect 123953 1377 123987 1411
rect 123987 1377 123996 1411
rect 123944 1368 123996 1377
rect 126152 1445 126161 1479
rect 126161 1445 126195 1479
rect 126195 1445 126204 1479
rect 126152 1436 126204 1445
rect 126244 1368 126296 1420
rect 130660 1436 130712 1488
rect 135260 1436 135312 1488
rect 139860 1436 139912 1488
rect 129188 1411 129240 1420
rect 129188 1377 129197 1411
rect 129197 1377 129231 1411
rect 129231 1377 129240 1411
rect 129188 1368 129240 1377
rect 129832 1368 129884 1420
rect 125784 1343 125836 1352
rect 125784 1309 125793 1343
rect 125793 1309 125827 1343
rect 125827 1309 125836 1343
rect 125784 1300 125836 1309
rect 131028 1300 131080 1352
rect 134616 1368 134668 1420
rect 135352 1411 135404 1420
rect 135352 1377 135361 1411
rect 135361 1377 135395 1411
rect 135395 1377 135404 1411
rect 135352 1368 135404 1377
rect 135444 1368 135496 1420
rect 138664 1411 138716 1420
rect 136640 1343 136692 1352
rect 109684 1164 109736 1216
rect 111156 1164 111208 1216
rect 114008 1164 114060 1216
rect 115572 1207 115624 1216
rect 115572 1173 115581 1207
rect 115581 1173 115615 1207
rect 115615 1173 115624 1207
rect 115572 1164 115624 1173
rect 116216 1207 116268 1216
rect 116216 1173 116225 1207
rect 116225 1173 116259 1207
rect 116259 1173 116268 1207
rect 116216 1164 116268 1173
rect 116308 1164 116360 1216
rect 122840 1164 122892 1216
rect 124128 1164 124180 1216
rect 126980 1207 127032 1216
rect 126980 1173 126989 1207
rect 126989 1173 127023 1207
rect 127023 1173 127032 1207
rect 126980 1164 127032 1173
rect 128268 1207 128320 1216
rect 128268 1173 128277 1207
rect 128277 1173 128311 1207
rect 128311 1173 128320 1207
rect 128268 1164 128320 1173
rect 131212 1164 131264 1216
rect 132040 1207 132092 1216
rect 132040 1173 132049 1207
rect 132049 1173 132083 1207
rect 132083 1173 132092 1207
rect 132040 1164 132092 1173
rect 136640 1309 136649 1343
rect 136649 1309 136683 1343
rect 136683 1309 136692 1343
rect 136640 1300 136692 1309
rect 138664 1377 138673 1411
rect 138673 1377 138707 1411
rect 138707 1377 138716 1411
rect 138664 1368 138716 1377
rect 139952 1411 140004 1420
rect 139952 1377 139961 1411
rect 139961 1377 139995 1411
rect 139995 1377 140004 1411
rect 139952 1368 140004 1377
rect 141148 1411 141200 1420
rect 141148 1377 141157 1411
rect 141157 1377 141191 1411
rect 141191 1377 141200 1411
rect 141148 1368 141200 1377
rect 151912 1436 151964 1488
rect 147864 1411 147916 1420
rect 147864 1377 147873 1411
rect 147873 1377 147907 1411
rect 147907 1377 147916 1411
rect 147864 1368 147916 1377
rect 148508 1368 148560 1420
rect 150256 1368 150308 1420
rect 156788 1411 156840 1420
rect 156788 1377 156797 1411
rect 156797 1377 156831 1411
rect 156831 1377 156840 1411
rect 156788 1368 156840 1377
rect 163964 1368 164016 1420
rect 165436 1411 165488 1420
rect 134616 1232 134668 1284
rect 139676 1300 139728 1352
rect 143172 1300 143224 1352
rect 144920 1343 144972 1352
rect 144920 1309 144929 1343
rect 144929 1309 144963 1343
rect 144963 1309 144972 1343
rect 144920 1300 144972 1309
rect 145748 1300 145800 1352
rect 149060 1300 149112 1352
rect 134340 1207 134392 1216
rect 134340 1173 134349 1207
rect 134349 1173 134383 1207
rect 134383 1173 134392 1207
rect 134340 1164 134392 1173
rect 134432 1164 134484 1216
rect 136088 1164 136140 1216
rect 140044 1232 140096 1284
rect 140964 1232 141016 1284
rect 141148 1232 141200 1284
rect 149152 1275 149204 1284
rect 149152 1241 149161 1275
rect 149161 1241 149195 1275
rect 149195 1241 149204 1275
rect 149152 1232 149204 1241
rect 150072 1300 150124 1352
rect 151360 1343 151412 1352
rect 151360 1309 151369 1343
rect 151369 1309 151403 1343
rect 151403 1309 151412 1343
rect 151360 1300 151412 1309
rect 151452 1300 151504 1352
rect 152648 1343 152700 1352
rect 152648 1309 152657 1343
rect 152657 1309 152691 1343
rect 152691 1309 152700 1343
rect 152648 1300 152700 1309
rect 155776 1343 155828 1352
rect 155776 1309 155785 1343
rect 155785 1309 155819 1343
rect 155819 1309 155828 1343
rect 155776 1300 155828 1309
rect 156880 1343 156932 1352
rect 156880 1309 156889 1343
rect 156889 1309 156923 1343
rect 156923 1309 156932 1343
rect 156880 1300 156932 1309
rect 155224 1232 155276 1284
rect 158720 1300 158772 1352
rect 159640 1343 159692 1352
rect 159640 1309 159649 1343
rect 159649 1309 159683 1343
rect 159683 1309 159692 1343
rect 159640 1300 159692 1309
rect 161112 1343 161164 1352
rect 161112 1309 161121 1343
rect 161121 1309 161155 1343
rect 161155 1309 161164 1343
rect 161112 1300 161164 1309
rect 162308 1300 162360 1352
rect 159548 1232 159600 1284
rect 160836 1275 160888 1284
rect 160836 1241 160845 1275
rect 160845 1241 160879 1275
rect 160879 1241 160888 1275
rect 160836 1232 160888 1241
rect 162860 1300 162912 1352
rect 165436 1377 165445 1411
rect 165445 1377 165479 1411
rect 165479 1377 165488 1411
rect 165436 1368 165488 1377
rect 166724 1343 166776 1352
rect 166724 1309 166733 1343
rect 166733 1309 166767 1343
rect 166767 1309 166776 1343
rect 166724 1300 166776 1309
rect 139676 1164 139728 1216
rect 144000 1164 144052 1216
rect 144276 1164 144328 1216
rect 146024 1207 146076 1216
rect 146024 1173 146033 1207
rect 146033 1173 146067 1207
rect 146067 1173 146076 1207
rect 146024 1164 146076 1173
rect 146668 1164 146720 1216
rect 151728 1164 151780 1216
rect 152924 1164 152976 1216
rect 153660 1207 153712 1216
rect 153660 1173 153669 1207
rect 153669 1173 153703 1207
rect 153703 1173 153712 1207
rect 153660 1164 153712 1173
rect 154028 1164 154080 1216
rect 154672 1164 154724 1216
rect 161296 1164 161348 1216
rect 161480 1164 161532 1216
rect 161940 1207 161992 1216
rect 161940 1173 161949 1207
rect 161949 1173 161983 1207
rect 161983 1173 161992 1207
rect 161940 1164 161992 1173
rect 162768 1164 162820 1216
rect 164424 1164 164476 1216
rect 166816 1207 166868 1216
rect 166816 1173 166825 1207
rect 166825 1173 166859 1207
rect 166859 1173 166868 1207
rect 166816 1164 166868 1173
rect 166908 1164 166960 1216
rect 56667 1062 56719 1114
rect 56731 1062 56783 1114
rect 56795 1062 56847 1114
rect 56859 1062 56911 1114
rect 97356 1028 97408 1080
rect 113088 1062 113140 1114
rect 113152 1062 113204 1114
rect 113216 1062 113268 1114
rect 113280 1062 113332 1114
rect 6736 960 6788 1012
rect 5632 824 5684 876
rect 6000 892 6052 944
rect 8116 867 8168 876
rect 8116 833 8125 867
rect 8125 833 8159 867
rect 8159 833 8168 867
rect 8116 824 8168 833
rect 10968 824 11020 876
rect 12992 960 13044 1012
rect 19616 960 19668 1012
rect 19800 1003 19852 1012
rect 19800 969 19809 1003
rect 19809 969 19843 1003
rect 19843 969 19852 1003
rect 19800 960 19852 969
rect 23664 960 23716 1012
rect 24676 960 24728 1012
rect 24952 1003 25004 1012
rect 24952 969 24961 1003
rect 24961 969 24995 1003
rect 24995 969 25004 1003
rect 24952 960 25004 969
rect 25872 1003 25924 1012
rect 25872 969 25881 1003
rect 25881 969 25915 1003
rect 25915 969 25924 1003
rect 25872 960 25924 969
rect 26148 960 26200 1012
rect 27988 960 28040 1012
rect 30196 960 30248 1012
rect 30288 960 30340 1012
rect 31944 960 31996 1012
rect 35716 960 35768 1012
rect 36360 1003 36412 1012
rect 36360 969 36369 1003
rect 36369 969 36403 1003
rect 36403 969 36412 1003
rect 36360 960 36412 969
rect 36452 960 36504 1012
rect 4344 756 4396 808
rect 4896 756 4948 808
rect 9680 756 9732 808
rect 5632 731 5684 740
rect 5632 697 5641 731
rect 5641 697 5675 731
rect 5675 697 5684 731
rect 5632 688 5684 697
rect 7840 688 7892 740
rect 35072 892 35124 944
rect 12440 756 12492 808
rect 10968 663 11020 672
rect 10968 629 10977 663
rect 10977 629 11011 663
rect 11011 629 11020 663
rect 10968 620 11020 629
rect 20628 824 20680 876
rect 22008 824 22060 876
rect 18328 756 18380 808
rect 24032 799 24084 808
rect 24032 765 24041 799
rect 24041 765 24075 799
rect 24075 765 24084 799
rect 24032 756 24084 765
rect 25872 824 25924 876
rect 27896 867 27948 876
rect 27528 799 27580 808
rect 27528 765 27537 799
rect 27537 765 27571 799
rect 27571 765 27580 799
rect 27528 756 27580 765
rect 27896 833 27905 867
rect 27905 833 27939 867
rect 27939 833 27948 867
rect 27896 824 27948 833
rect 30104 824 30156 876
rect 29000 756 29052 808
rect 33416 824 33468 876
rect 33876 867 33928 876
rect 33876 833 33885 867
rect 33885 833 33919 867
rect 33919 833 33928 867
rect 33876 824 33928 833
rect 34704 824 34756 876
rect 37464 892 37516 944
rect 35440 867 35492 876
rect 35440 833 35449 867
rect 35449 833 35483 867
rect 35483 833 35492 867
rect 35440 824 35492 833
rect 37556 824 37608 876
rect 37832 824 37884 876
rect 40776 960 40828 1012
rect 40960 960 41012 1012
rect 42248 960 42300 1012
rect 42340 960 42392 1012
rect 44548 960 44600 1012
rect 44824 1003 44876 1012
rect 44824 969 44833 1003
rect 44833 969 44867 1003
rect 44867 969 44876 1003
rect 44824 960 44876 969
rect 44916 960 44968 1012
rect 47216 960 47268 1012
rect 47860 960 47912 1012
rect 49608 960 49660 1012
rect 50160 960 50212 1012
rect 50436 960 50488 1012
rect 102416 960 102468 1012
rect 27988 688 28040 740
rect 28080 688 28132 740
rect 14280 620 14332 672
rect 18052 663 18104 672
rect 18052 629 18061 663
rect 18061 629 18095 663
rect 18095 629 18104 663
rect 18052 620 18104 629
rect 26516 620 26568 672
rect 28816 620 28868 672
rect 30196 620 30248 672
rect 34704 688 34756 740
rect 34888 688 34940 740
rect 36544 688 36596 740
rect 38292 756 38344 808
rect 40684 892 40736 944
rect 40868 892 40920 944
rect 38936 824 38988 876
rect 41512 867 41564 876
rect 39028 756 39080 808
rect 39304 756 39356 808
rect 40500 756 40552 808
rect 40592 756 40644 808
rect 41512 833 41521 867
rect 41521 833 41555 867
rect 41555 833 41564 867
rect 41512 824 41564 833
rect 36452 620 36504 672
rect 39304 620 39356 672
rect 40408 688 40460 740
rect 40868 688 40920 740
rect 41696 688 41748 740
rect 41604 620 41656 672
rect 41972 892 42024 944
rect 42524 892 42576 944
rect 43076 892 43128 944
rect 65156 892 65208 944
rect 66352 935 66404 944
rect 66352 901 66361 935
rect 66361 901 66395 935
rect 66395 901 66404 935
rect 66352 892 66404 901
rect 42984 824 43036 876
rect 43904 824 43956 876
rect 44088 824 44140 876
rect 44916 824 44968 876
rect 45652 824 45704 876
rect 46296 867 46348 876
rect 46296 833 46305 867
rect 46305 833 46339 867
rect 46339 833 46348 867
rect 46296 824 46348 833
rect 44640 756 44692 808
rect 49424 824 49476 876
rect 50160 824 50212 876
rect 52552 867 52604 876
rect 52552 833 52561 867
rect 52561 833 52595 867
rect 52595 833 52604 867
rect 52552 824 52604 833
rect 53012 824 53064 876
rect 55312 824 55364 876
rect 55496 824 55548 876
rect 57796 824 57848 876
rect 58532 867 58584 876
rect 58532 833 58541 867
rect 58541 833 58575 867
rect 58575 833 58584 867
rect 58532 824 58584 833
rect 47400 756 47452 808
rect 45376 688 45428 740
rect 46112 688 46164 740
rect 49056 688 49108 740
rect 49700 688 49752 740
rect 49792 688 49844 740
rect 50804 756 50856 808
rect 50896 756 50948 808
rect 54484 756 54536 808
rect 56968 756 57020 808
rect 58992 756 59044 808
rect 59728 824 59780 876
rect 60464 867 60516 876
rect 60464 833 60473 867
rect 60473 833 60507 867
rect 60507 833 60516 867
rect 60464 824 60516 833
rect 61476 824 61528 876
rect 63776 867 63828 876
rect 59912 756 59964 808
rect 50160 688 50212 740
rect 52000 688 52052 740
rect 52920 731 52972 740
rect 52920 697 52929 731
rect 52929 697 52963 731
rect 52963 697 52972 731
rect 52920 688 52972 697
rect 53472 620 53524 672
rect 53656 620 53708 672
rect 55220 688 55272 740
rect 56416 688 56468 740
rect 60372 688 60424 740
rect 63776 833 63785 867
rect 63785 833 63819 867
rect 63819 833 63828 867
rect 68744 892 68796 944
rect 68836 892 68888 944
rect 70124 892 70176 944
rect 70676 892 70728 944
rect 70860 892 70912 944
rect 71872 935 71924 944
rect 71872 901 71881 935
rect 71881 901 71915 935
rect 71915 901 71924 935
rect 71872 892 71924 901
rect 75092 892 75144 944
rect 75184 892 75236 944
rect 80520 935 80572 944
rect 63776 824 63828 833
rect 69204 867 69256 876
rect 69204 833 69213 867
rect 69213 833 69247 867
rect 69247 833 69256 867
rect 69204 824 69256 833
rect 71780 824 71832 876
rect 72976 824 73028 876
rect 76656 824 76708 876
rect 79232 824 79284 876
rect 79416 824 79468 876
rect 68928 799 68980 808
rect 61200 688 61252 740
rect 68928 765 68937 799
rect 68937 765 68971 799
rect 68971 765 68980 799
rect 68928 756 68980 765
rect 69848 756 69900 808
rect 74264 756 74316 808
rect 75828 799 75880 808
rect 75828 765 75837 799
rect 75837 765 75871 799
rect 75871 765 75880 799
rect 75828 756 75880 765
rect 77576 799 77628 808
rect 77576 765 77585 799
rect 77585 765 77619 799
rect 77619 765 77628 799
rect 77576 756 77628 765
rect 78680 799 78732 808
rect 78680 765 78689 799
rect 78689 765 78723 799
rect 78723 765 78732 799
rect 78680 756 78732 765
rect 65064 688 65116 740
rect 65616 688 65668 740
rect 68100 688 68152 740
rect 69112 688 69164 740
rect 70216 688 70268 740
rect 75736 688 75788 740
rect 56048 620 56100 672
rect 56232 620 56284 672
rect 57428 620 57480 672
rect 59636 620 59688 672
rect 60464 620 60516 672
rect 60648 620 60700 672
rect 65432 620 65484 672
rect 65524 620 65576 672
rect 79600 688 79652 740
rect 80520 901 80529 935
rect 80529 901 80563 935
rect 80563 901 80572 935
rect 80520 892 80572 901
rect 81072 824 81124 876
rect 83464 824 83516 876
rect 84844 892 84896 944
rect 86316 892 86368 944
rect 89628 892 89680 944
rect 90180 892 90232 944
rect 92020 892 92072 944
rect 88616 824 88668 876
rect 84016 756 84068 808
rect 89352 824 89404 876
rect 93676 892 93728 944
rect 94412 892 94464 944
rect 104992 960 105044 1012
rect 105176 892 105228 944
rect 102600 756 102652 808
rect 104256 824 104308 876
rect 107016 960 107068 1012
rect 107844 1003 107896 1012
rect 107844 969 107853 1003
rect 107853 969 107887 1003
rect 107887 969 107896 1003
rect 107844 960 107896 969
rect 133696 1003 133748 1012
rect 133696 969 133705 1003
rect 133705 969 133739 1003
rect 133739 969 133748 1003
rect 133696 960 133748 969
rect 133880 960 133932 1012
rect 135628 960 135680 1012
rect 136088 1003 136140 1012
rect 136088 969 136097 1003
rect 136097 969 136131 1003
rect 136131 969 136140 1003
rect 136088 960 136140 969
rect 139216 960 139268 1012
rect 140780 960 140832 1012
rect 141056 1003 141108 1012
rect 141056 969 141065 1003
rect 141065 969 141099 1003
rect 141099 969 141108 1003
rect 141056 960 141108 969
rect 143172 1003 143224 1012
rect 143172 969 143181 1003
rect 143181 969 143215 1003
rect 143215 969 143224 1003
rect 143172 960 143224 969
rect 155224 1003 155276 1012
rect 155224 969 155233 1003
rect 155233 969 155267 1003
rect 155267 969 155276 1003
rect 155224 960 155276 969
rect 155776 1003 155828 1012
rect 155776 969 155785 1003
rect 155785 969 155819 1003
rect 155819 969 155828 1003
rect 155776 960 155828 969
rect 104992 756 105044 808
rect 109224 892 109276 944
rect 106096 824 106148 876
rect 110788 892 110840 944
rect 106372 799 106424 808
rect 106372 765 106381 799
rect 106381 765 106415 799
rect 106415 765 106424 799
rect 106372 756 106424 765
rect 82176 731 82228 740
rect 82176 697 82185 731
rect 82185 697 82219 731
rect 82219 697 82228 731
rect 82176 688 82228 697
rect 88984 731 89036 740
rect 88984 697 88993 731
rect 88993 697 89027 731
rect 89027 697 89036 731
rect 88984 688 89036 697
rect 89076 688 89128 740
rect 107936 756 107988 808
rect 109408 756 109460 808
rect 111156 824 111208 876
rect 114008 892 114060 944
rect 116216 935 116268 944
rect 116216 901 116225 935
rect 116225 901 116259 935
rect 116259 901 116268 935
rect 116216 892 116268 901
rect 114928 799 114980 808
rect 111248 688 111300 740
rect 114928 765 114937 799
rect 114937 765 114971 799
rect 114971 765 114980 799
rect 114928 756 114980 765
rect 116308 824 116360 876
rect 118148 824 118200 876
rect 118424 756 118476 808
rect 119344 824 119396 876
rect 122656 867 122708 876
rect 122656 833 122665 867
rect 122665 833 122699 867
rect 122699 833 122708 867
rect 122656 824 122708 833
rect 123944 824 123996 876
rect 125600 867 125652 876
rect 125600 833 125617 867
rect 125617 833 125651 867
rect 125651 833 125652 867
rect 126152 867 126204 876
rect 125600 824 125652 833
rect 126152 833 126161 867
rect 126161 833 126195 867
rect 126195 833 126204 867
rect 126152 824 126204 833
rect 129188 824 129240 876
rect 132960 824 133012 876
rect 133696 824 133748 876
rect 136916 824 136968 876
rect 137652 867 137704 876
rect 137652 833 137661 867
rect 137661 833 137695 867
rect 137695 833 137704 867
rect 137652 824 137704 833
rect 133972 756 134024 808
rect 134064 756 134116 808
rect 139216 799 139268 808
rect 139216 765 139225 799
rect 139225 765 139259 799
rect 139259 765 139268 799
rect 139216 756 139268 765
rect 141056 824 141108 876
rect 140872 756 140924 808
rect 142160 824 142212 876
rect 83280 663 83332 672
rect 83280 629 83289 663
rect 83289 629 83323 663
rect 83323 629 83332 663
rect 83280 620 83332 629
rect 84292 663 84344 672
rect 84292 629 84301 663
rect 84301 629 84335 663
rect 84335 629 84344 663
rect 84292 620 84344 629
rect 86132 663 86184 672
rect 86132 629 86141 663
rect 86141 629 86175 663
rect 86175 629 86184 663
rect 86132 620 86184 629
rect 95608 620 95660 672
rect 103060 620 103112 672
rect 104256 663 104308 672
rect 104256 629 104265 663
rect 104265 629 104299 663
rect 104299 629 104308 663
rect 104256 620 104308 629
rect 106372 620 106424 672
rect 120080 688 120132 740
rect 115572 620 115624 672
rect 125784 688 125836 740
rect 126980 620 127032 672
rect 131764 688 131816 740
rect 137744 731 137796 740
rect 137744 697 137753 731
rect 137753 697 137787 731
rect 137787 697 137796 731
rect 137744 688 137796 697
rect 137928 688 137980 740
rect 146024 824 146076 876
rect 151728 867 151780 876
rect 151728 833 151737 867
rect 151737 833 151771 867
rect 151771 833 151780 867
rect 151728 824 151780 833
rect 158260 960 158312 1012
rect 158352 960 158404 1012
rect 161296 1003 161348 1012
rect 159456 867 159508 876
rect 159456 833 159465 867
rect 159465 833 159499 867
rect 159499 833 159508 867
rect 159456 824 159508 833
rect 161296 969 161305 1003
rect 161305 969 161339 1003
rect 161339 969 161348 1003
rect 161296 960 161348 969
rect 166816 1003 166868 1012
rect 166816 969 166825 1003
rect 166825 969 166859 1003
rect 166859 969 166868 1003
rect 166816 960 166868 969
rect 162032 867 162084 876
rect 162032 833 162041 867
rect 162041 833 162075 867
rect 162075 833 162084 867
rect 162032 824 162084 833
rect 162768 824 162820 876
rect 132132 620 132184 672
rect 132500 663 132552 672
rect 132500 629 132509 663
rect 132509 629 132543 663
rect 132543 629 132552 663
rect 132500 620 132552 629
rect 132960 663 133012 672
rect 132960 629 132969 663
rect 132969 629 133003 663
rect 133003 629 133012 663
rect 132960 620 133012 629
rect 144000 620 144052 672
rect 151912 731 151964 740
rect 151912 697 151921 731
rect 151921 697 151955 731
rect 151955 697 151964 731
rect 151912 688 151964 697
rect 156788 756 156840 808
rect 160468 799 160520 808
rect 160468 765 160477 799
rect 160477 765 160511 799
rect 160511 765 160520 799
rect 160468 756 160520 765
rect 165988 799 166040 808
rect 165988 765 165997 799
rect 165997 765 166031 799
rect 166031 765 166040 799
rect 165988 756 166040 765
rect 28456 518 28508 570
rect 28520 518 28572 570
rect 28584 518 28636 570
rect 28648 518 28700 570
rect 84878 518 84930 570
rect 84942 518 84994 570
rect 85006 518 85058 570
rect 85070 518 85122 570
rect 141299 518 141351 570
rect 141363 518 141415 570
rect 141427 518 141479 570
rect 141491 518 141543 570
rect 8760 416 8812 468
rect 27528 416 27580 468
rect 28816 416 28868 468
rect 32772 416 32824 468
rect 32864 416 32916 468
rect 42340 416 42392 468
rect 42800 416 42852 468
rect 42984 416 43036 468
rect 50896 416 50948 468
rect 52736 416 52788 468
rect 53012 416 53064 468
rect 57152 416 57204 468
rect 57428 416 57480 468
rect 68928 416 68980 468
rect 69112 416 69164 468
rect 72976 416 73028 468
rect 81624 416 81676 468
rect 89076 416 89128 468
rect 101128 416 101180 468
rect 137744 416 137796 468
rect 138296 416 138348 468
rect 140872 416 140924 468
rect 10968 348 11020 400
rect 19248 348 19300 400
rect 23480 348 23532 400
rect 81992 348 82044 400
rect 98552 348 98604 400
rect 114928 348 114980 400
rect 132132 348 132184 400
rect 140320 348 140372 400
rect 17224 280 17276 332
rect 82176 280 82228 332
rect 95056 280 95108 332
rect 21272 212 21324 264
rect 83280 212 83332 264
rect 104808 280 104860 332
rect 114468 280 114520 332
rect 118424 280 118476 332
rect 132040 280 132092 332
rect 132960 280 133012 332
rect 107936 212 107988 264
rect 108120 212 108172 264
rect 160468 212 160520 264
rect 30840 144 30892 196
rect 91376 144 91428 196
rect 106280 144 106332 196
rect 151912 144 151964 196
rect 24032 76 24084 128
rect 36452 119 36504 128
rect 18052 8 18104 60
rect 34336 8 34388 60
rect 34520 8 34572 60
rect 35808 8 35860 60
rect 36452 85 36461 119
rect 36461 85 36495 119
rect 36495 85 36504 119
rect 36452 76 36504 85
rect 36544 76 36596 128
rect 36728 76 36780 128
rect 40960 76 41012 128
rect 41144 8 41196 60
rect 41328 76 41380 128
rect 47400 76 47452 128
rect 47584 76 47636 128
rect 48136 76 48188 128
rect 50160 76 50212 128
rect 50344 76 50396 128
rect 78680 76 78732 128
rect 104256 76 104308 128
rect 134064 76 134116 128
rect 139124 76 139176 128
rect 49976 8 50028 60
rect 75828 8 75880 60
rect 107752 8 107804 60
rect 156788 8 156840 60
<< metal2 >>
rect 33690 13016 33746 13025
rect 754 12200 810 13000
rect 1122 12200 1178 13000
rect 1490 12200 1546 13000
rect 1858 12200 1914 13000
rect 2226 12200 2282 13000
rect 2594 12200 2650 13000
rect 2962 12200 3018 13000
rect 3330 12200 3386 13000
rect 3698 12200 3754 13000
rect 4066 12200 4122 13000
rect 4434 12200 4490 13000
rect 4802 12200 4858 13000
rect 5170 12200 5226 13000
rect 5538 12200 5594 13000
rect 5906 12200 5962 13000
rect 6274 12200 6330 13000
rect 6642 12200 6698 13000
rect 7010 12200 7066 13000
rect 7378 12200 7434 13000
rect 7746 12200 7802 13000
rect 8114 12200 8170 13000
rect 8482 12200 8538 13000
rect 8850 12200 8906 13000
rect 9218 12200 9274 13000
rect 9586 12200 9642 13000
rect 9954 12200 10010 13000
rect 10322 12200 10378 13000
rect 10690 12200 10746 13000
rect 11058 12200 11114 13000
rect 11426 12200 11482 13000
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 768 8090 796 12200
rect 1136 9382 1164 12200
rect 1124 9376 1176 9382
rect 1124 9318 1176 9324
rect 1504 8838 1532 12200
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1872 8634 1900 12200
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 2240 8362 2268 12200
rect 2608 9450 2636 12200
rect 2870 10432 2926 10441
rect 2870 10367 2926 10376
rect 2884 10198 2912 10367
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2976 9654 3004 12200
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 3344 9586 3372 12200
rect 3712 12152 3740 12200
rect 3712 12124 3832 12152
rect 3698 12064 3754 12073
rect 3698 11999 3754 12008
rect 3712 11286 3740 11999
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 3606 10976 3662 10985
rect 3606 10911 3662 10920
rect 3620 9926 3648 10911
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 756 8084 808 8090
rect 756 8026 808 8032
rect 3620 8022 3648 8366
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3620 7750 3648 7822
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 6866 3648 7278
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3712 6390 3740 10610
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3252 5234 3280 6190
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3698 6080 3754 6089
rect 3436 5778 3464 6054
rect 3698 6015 3754 6024
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3712 5574 3740 6015
rect 3804 5846 3832 12124
rect 4080 11642 4108 12200
rect 3988 11614 4108 11642
rect 3988 10674 4016 11614
rect 4160 11552 4212 11558
rect 4066 11520 4122 11529
rect 4160 11494 4212 11500
rect 4066 11455 4122 11464
rect 4080 11082 4108 11455
rect 4172 11150 4200 11494
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10062 4016 10406
rect 4172 10130 4200 11086
rect 4356 10674 4384 11154
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4356 10266 4384 10610
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4448 10010 4476 12200
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4540 11218 4568 12106
rect 4816 11914 4844 12200
rect 4816 11886 4936 11914
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4816 11354 4844 11698
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4816 10674 4844 11290
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4712 10056 4764 10062
rect 4080 9897 4108 9998
rect 4448 9982 4660 10010
rect 4712 9998 4764 10004
rect 4436 9920 4488 9926
rect 4066 9888 4122 9897
rect 4436 9862 4488 9868
rect 4066 9823 4122 9832
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3896 9178 3924 9454
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 4080 9042 4108 9318
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4066 8800 4122 8809
rect 4066 8735 4122 8744
rect 4080 8566 4108 8735
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 4080 7478 4108 8191
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4066 7168 4122 7177
rect 4122 7126 4200 7154
rect 4066 7103 4122 7112
rect 4066 6624 4122 6633
rect 4066 6559 4122 6568
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 4080 5658 4108 6559
rect 4172 5778 4200 7126
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4264 6458 4292 6734
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4080 5630 4200 5658
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3882 5536 3938 5545
rect 3882 5471 3938 5480
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3252 4826 3280 5170
rect 3698 4992 3754 5001
rect 3698 4927 3754 4936
rect 3712 4826 3740 4927
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3896 4486 3924 5471
rect 4172 4690 4200 5630
rect 4448 5166 4476 9862
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4540 7342 4568 9522
rect 4632 9178 4660 9982
rect 4724 9382 4752 9998
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4632 7954 4660 8774
rect 4724 8673 4752 9318
rect 4710 8664 4766 8673
rect 4710 8599 4766 8608
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4802 7712 4858 7721
rect 4802 7647 4858 7656
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4816 7002 4844 7647
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4908 6186 4936 11886
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 9926 5120 10610
rect 5184 10010 5212 12200
rect 5184 9982 5304 10010
rect 5080 9920 5132 9926
rect 5078 9888 5080 9897
rect 5132 9888 5134 9897
rect 5078 9823 5134 9832
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5184 8634 5212 8910
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5276 8566 5304 9982
rect 5552 9330 5580 12200
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5552 9302 5672 9330
rect 5538 9208 5594 9217
rect 5538 9143 5594 9152
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5460 8838 5488 8978
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 5354 5672 5410 5681
rect 5354 5607 5356 5616
rect 5408 5607 5410 5616
rect 5356 5578 5408 5584
rect 5354 5264 5410 5273
rect 5354 5199 5356 5208
rect 5408 5199 5410 5208
rect 5356 5170 5408 5176
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 5460 4729 5488 8774
rect 5552 8634 5580 9143
rect 5644 9110 5672 9302
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5552 8498 5580 8570
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5552 7546 5580 7686
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5552 7177 5580 7278
rect 5538 7168 5594 7177
rect 5538 7103 5594 7112
rect 5736 6934 5764 11222
rect 5920 9518 5948 12200
rect 6288 11778 6316 12200
rect 6288 11750 6500 11778
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6104 11150 6132 11494
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6104 9654 6132 11086
rect 6288 10810 6316 11630
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 6368 9376 6420 9382
rect 6090 9344 6146 9353
rect 6368 9318 6420 9324
rect 6090 9279 6146 9288
rect 6104 8022 6132 9279
rect 6380 9042 6408 9318
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6380 8634 6408 8978
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 6366 6896 6422 6905
rect 6366 6831 6368 6840
rect 6420 6831 6422 6840
rect 6368 6802 6420 6808
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5828 5778 5856 6190
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5446 4720 5502 4729
rect 4160 4684 4212 4690
rect 5446 4655 5502 4664
rect 4160 4626 4212 4632
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3988 4282 4016 4558
rect 4066 4448 4122 4457
rect 4066 4383 4122 4392
rect 4080 4282 4108 4383
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 938 3088 994 3097
rect 938 3023 994 3032
rect 756 2916 808 2922
rect 756 2858 808 2864
rect 572 2576 624 2582
rect 572 2518 624 2524
rect 584 800 612 2518
rect 768 800 796 2858
rect 952 800 980 3023
rect 1320 800 1348 4082
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 4066 3904 4122 3913
rect 2962 2272 3018 2281
rect 2962 2207 3018 2216
rect 2976 2038 3004 2207
rect 2964 2032 3016 2038
rect 2964 1974 3016 1980
rect 3056 1964 3108 1970
rect 3056 1906 3108 1912
rect 2780 1828 2832 1834
rect 2780 1770 2832 1776
rect 2044 1556 2096 1562
rect 2044 1498 2096 1504
rect 1676 1488 1728 1494
rect 1676 1430 1728 1436
rect 1688 800 1716 1430
rect 2056 800 2084 1498
rect 2412 1420 2464 1426
rect 2412 1362 2464 1368
rect 2424 800 2452 1362
rect 2792 800 2820 1770
rect 3068 1562 3096 1906
rect 3056 1556 3108 1562
rect 3056 1498 3108 1504
rect 3160 800 3188 3878
rect 4066 3839 4122 3848
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3240 1896 3292 1902
rect 3240 1838 3292 1844
rect 3252 1562 3280 1838
rect 3240 1556 3292 1562
rect 3240 1498 3292 1504
rect 3620 898 3648 3674
rect 4080 3670 4108 3839
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3712 2650 3740 2994
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3804 1193 3832 2382
rect 3790 1184 3846 1193
rect 3790 1119 3846 1128
rect 3528 870 3648 898
rect 3528 800 3556 870
rect 3896 800 3924 3130
rect 3988 2825 4016 3334
rect 4540 3058 4568 4014
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 3974 2816 4030 2825
rect 3974 2751 4030 2760
rect 4724 2650 4752 2994
rect 4908 2922 4936 3402
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4068 1760 4120 1766
rect 4066 1728 4068 1737
rect 4120 1728 4122 1737
rect 4066 1663 4122 1672
rect 4264 870 4384 898
rect 4264 800 4292 870
rect 4356 814 4384 870
rect 4632 870 4752 898
rect 4344 808 4396 814
rect 570 0 626 800
rect 754 0 810 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4632 800 4660 870
rect 4344 750 4396 756
rect 4618 0 4674 800
rect 4724 796 4752 870
rect 4896 808 4948 814
rect 4724 768 4896 796
rect 5000 800 5028 2858
rect 5172 1964 5224 1970
rect 5172 1906 5224 1912
rect 5184 1766 5212 1906
rect 5172 1760 5224 1766
rect 5170 1728 5172 1737
rect 5224 1728 5226 1737
rect 5170 1663 5226 1672
rect 5368 800 5396 3946
rect 5736 3602 5764 5510
rect 6472 5302 6500 11750
rect 6656 6225 6684 12200
rect 7024 10248 7052 12200
rect 7024 10220 7236 10248
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7024 9586 7052 10066
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7116 9722 7144 9862
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6826 7440 6882 7449
rect 6826 7375 6882 7384
rect 6642 6216 6698 6225
rect 6642 6151 6698 6160
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 5906 4584 5962 4593
rect 5906 4519 5908 4528
rect 5960 4519 5962 4528
rect 5908 4490 5960 4496
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 2514 5580 2790
rect 5828 2514 5856 4422
rect 5906 4176 5962 4185
rect 5906 4111 5962 4120
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5920 1850 5948 4111
rect 6090 4040 6146 4049
rect 6090 3975 6146 3984
rect 5736 1822 5948 1850
rect 5632 876 5684 882
rect 5632 818 5684 824
rect 4896 750 4948 756
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5644 785 5672 818
rect 5736 800 5764 1822
rect 6000 1216 6052 1222
rect 6000 1158 6052 1164
rect 6012 950 6040 1158
rect 6000 944 6052 950
rect 6000 886 6052 892
rect 6104 800 6132 3975
rect 6458 3904 6514 3913
rect 6458 3839 6514 3848
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6182 3360 6238 3369
rect 6182 3295 6238 3304
rect 6196 2990 6224 3295
rect 6380 3126 6408 3674
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6288 2106 6316 2858
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 6276 1216 6328 1222
rect 6276 1158 6328 1164
rect 5630 776 5686 785
rect 5630 711 5632 720
rect 5684 711 5686 720
rect 5632 682 5684 688
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6288 377 6316 1158
rect 6472 800 6500 3839
rect 6642 3768 6698 3777
rect 6642 3703 6644 3712
rect 6696 3703 6698 3712
rect 6644 3674 6696 3680
rect 6656 3534 6684 3674
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6736 1216 6788 1222
rect 6736 1158 6788 1164
rect 6748 1018 6776 1158
rect 6736 1012 6788 1018
rect 6736 954 6788 960
rect 6840 800 6868 7375
rect 6932 5778 6960 9386
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 7208 5545 7236 10220
rect 7392 9489 7420 12200
rect 7654 11248 7710 11257
rect 7654 11183 7656 11192
rect 7708 11183 7710 11192
rect 7656 11154 7708 11160
rect 7378 9480 7434 9489
rect 7378 9415 7434 9424
rect 7760 9042 7788 12200
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8036 11150 8064 11698
rect 8024 11144 8076 11150
rect 8022 11112 8024 11121
rect 8076 11112 8078 11121
rect 8022 11047 8078 11056
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9722 8064 9862
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8036 7342 8064 8026
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7944 6866 7972 7278
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 8128 6497 8156 12200
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8312 10266 8340 10542
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8496 9081 8524 12200
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8482 9072 8538 9081
rect 8482 9007 8538 9016
rect 8298 8936 8354 8945
rect 8298 8871 8300 8880
rect 8352 8871 8354 8880
rect 8300 8842 8352 8848
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8220 7177 8248 7210
rect 8206 7168 8262 7177
rect 8206 7103 8262 7112
rect 8114 6488 8170 6497
rect 8114 6423 8170 6432
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 7746 5808 7802 5817
rect 7746 5743 7748 5752
rect 7800 5743 7802 5752
rect 7748 5714 7800 5720
rect 8036 5574 8064 6190
rect 8024 5568 8076 5574
rect 7194 5536 7250 5545
rect 8024 5510 8076 5516
rect 7194 5471 7250 5480
rect 8036 5370 8064 5510
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8220 5098 8248 6326
rect 8588 6254 8616 11018
rect 8864 9450 8892 12200
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8864 8566 8892 9114
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 9232 8294 9260 12200
rect 9310 10976 9366 10985
rect 9310 10911 9366 10920
rect 9324 10674 9352 10911
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 10266 9352 10610
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9600 8378 9628 12200
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9692 11694 9720 11766
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9692 11218 9720 11494
rect 9784 11286 9812 11494
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 10810 9720 11154
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9680 10192 9732 10198
rect 9678 10160 9680 10169
rect 9732 10160 9734 10169
rect 9678 10095 9734 10104
rect 9968 8498 9996 12200
rect 10336 9518 10364 12200
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9600 8350 9812 8378
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 6866 8984 7686
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9600 7206 9628 7346
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 9232 6089 9260 6258
rect 9218 6080 9274 6089
rect 9218 6015 9274 6024
rect 9232 5914 9260 6015
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7194 4312 7250 4321
rect 7194 4247 7250 4256
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7024 3466 7052 4014
rect 7208 3738 7236 4247
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 7392 2922 7420 4762
rect 8484 4480 8536 4486
rect 9600 4457 9628 7142
rect 9784 6934 9812 8350
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 10704 6390 10732 12200
rect 10876 6656 10928 6662
rect 10874 6624 10876 6633
rect 10928 6624 10930 6633
rect 10874 6559 10930 6568
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5778 10456 6190
rect 11072 5953 11100 12200
rect 11440 11014 11468 12200
rect 11532 11354 11560 12310
rect 11794 12200 11850 13000
rect 12162 12200 12218 13000
rect 12530 12200 12586 13000
rect 12898 12200 12954 13000
rect 13266 12200 13322 13000
rect 13634 12200 13690 13000
rect 14002 12200 14058 13000
rect 14370 12200 14426 13000
rect 14738 12200 14794 13000
rect 15106 12200 15162 13000
rect 15474 12200 15530 13000
rect 15842 12200 15898 13000
rect 16210 12200 16266 13000
rect 16578 12200 16634 13000
rect 16946 12200 17002 13000
rect 17314 12200 17370 13000
rect 17682 12200 17738 13000
rect 18050 12200 18106 13000
rect 18418 12200 18474 13000
rect 18786 12200 18842 13000
rect 19154 12200 19210 13000
rect 19522 12200 19578 13000
rect 19890 12200 19946 13000
rect 20258 12200 20314 13000
rect 20626 12200 20682 13000
rect 20994 12200 21050 13000
rect 21362 12200 21418 13000
rect 21730 12200 21786 13000
rect 22098 12200 22154 13000
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11808 9625 11836 12200
rect 11794 9616 11850 9625
rect 11794 9551 11850 9560
rect 12176 8401 12204 12200
rect 12544 8838 12572 12200
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12636 10674 12664 11018
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 10266 12664 10610
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12162 8392 12218 8401
rect 12162 8327 12218 8336
rect 12256 8016 12308 8022
rect 12912 7993 12940 12200
rect 12256 7958 12308 7964
rect 12898 7984 12954 7993
rect 11058 5944 11114 5953
rect 11058 5879 11114 5888
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10874 5128 10930 5137
rect 10874 5063 10930 5072
rect 8484 4422 8536 4428
rect 9586 4448 9642 4457
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7208 1902 7236 2246
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7196 1896 7248 1902
rect 7196 1838 7248 1844
rect 7208 1562 7236 1838
rect 7196 1556 7248 1562
rect 7196 1498 7248 1504
rect 7300 1306 7328 2042
rect 7484 1494 7512 2858
rect 7564 1760 7616 1766
rect 7564 1702 7616 1708
rect 7472 1488 7524 1494
rect 7472 1430 7524 1436
rect 7208 1278 7328 1306
rect 7208 800 7236 1278
rect 7576 800 7604 1702
rect 7760 1358 7788 3402
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7852 2310 7880 2994
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 6274 368 6330 377
rect 6274 303 6330 312
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7852 746 7880 2246
rect 7944 800 7972 3878
rect 8036 3777 8064 4082
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8022 3768 8078 3777
rect 8022 3703 8024 3712
rect 8076 3703 8078 3712
rect 8024 3674 8076 3680
rect 8404 2122 8432 4014
rect 8496 3058 8524 4422
rect 9586 4383 9642 4392
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 9232 3738 9260 4150
rect 9324 4134 9720 4162
rect 9324 4010 9352 4134
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8496 2650 8524 2994
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8312 2094 8432 2122
rect 8114 912 8170 921
rect 8114 847 8116 856
rect 8168 847 8170 856
rect 8116 818 8168 824
rect 8312 800 8340 2094
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 8404 1222 8432 1906
rect 8680 1766 8708 3606
rect 9232 3602 9260 3674
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9034 2272 9090 2281
rect 9034 2207 9090 2216
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 8392 1216 8444 1222
rect 8392 1158 8444 1164
rect 8404 1057 8432 1158
rect 8390 1048 8446 1057
rect 8390 983 8446 992
rect 8680 870 8800 898
rect 8680 800 8708 870
rect 7840 740 7892 746
rect 7840 682 7892 688
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 8772 474 8800 870
rect 9048 800 9076 2207
rect 9220 1896 9272 1902
rect 9220 1838 9272 1844
rect 9232 1562 9260 1838
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 9416 800 9444 3946
rect 9692 3738 9720 4134
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9678 3360 9734 3369
rect 9678 3295 9734 3304
rect 9692 3210 9720 3295
rect 9508 3182 9720 3210
rect 9508 2582 9536 3182
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9692 814 9720 2790
rect 9784 2514 9812 2994
rect 9876 2922 9904 4218
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9784 2417 9812 2450
rect 9770 2408 9826 2417
rect 9770 2343 9826 2352
rect 10060 1408 10088 3402
rect 10152 3126 10180 4082
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10244 2854 10272 2994
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10138 2544 10194 2553
rect 10704 2514 10732 3334
rect 10138 2479 10194 2488
rect 10692 2508 10744 2514
rect 9784 1380 10088 1408
rect 9680 808 9732 814
rect 8760 468 8812 474
rect 8760 410 8812 416
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9784 800 9812 1380
rect 10152 800 10180 2479
rect 10692 2450 10744 2456
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 2038 10364 2246
rect 10782 2136 10838 2145
rect 10782 2071 10838 2080
rect 10324 2032 10376 2038
rect 10324 1974 10376 1980
rect 10796 1970 10824 2071
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 10796 1562 10824 1906
rect 10784 1556 10836 1562
rect 10784 1498 10836 1504
rect 10506 1320 10562 1329
rect 10506 1255 10562 1264
rect 10520 800 10548 1255
rect 10888 800 10916 5063
rect 12268 4554 12296 7958
rect 12898 7919 12954 7928
rect 13280 7177 13308 12200
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13372 7750 13400 8366
rect 13648 7857 13676 12200
rect 14016 10826 14044 12200
rect 14016 10798 14136 10826
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10266 14044 10610
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14108 8022 14136 10798
rect 14384 9586 14412 12200
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14476 11694 14504 11766
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 13634 7848 13690 7857
rect 13634 7783 13690 7792
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 13266 7168 13322 7177
rect 13266 7103 13322 7112
rect 12438 7032 12494 7041
rect 12438 6967 12494 6976
rect 12452 6633 12480 6967
rect 13372 6866 13400 7686
rect 14108 7410 14136 7686
rect 14476 7546 14504 7686
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 13924 7206 13952 7346
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 14108 7002 14136 7346
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14292 6866 14320 7278
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 12438 6624 12494 6633
rect 12438 6559 12494 6568
rect 12346 6352 12402 6361
rect 12346 6287 12402 6296
rect 12360 5914 12388 6287
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12360 5710 12388 5850
rect 14752 5846 14780 12200
rect 15120 8498 15148 12200
rect 15292 9648 15344 9654
rect 15344 9608 15424 9636
rect 15292 9590 15344 9596
rect 15200 9376 15252 9382
rect 15252 9324 15332 9330
rect 15200 9318 15332 9324
rect 15212 9302 15332 9318
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14844 7886 14872 8434
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 15120 6322 15148 8230
rect 15212 7342 15240 8978
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15304 6866 15332 9302
rect 15396 8974 15424 9608
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15488 7002 15516 12200
rect 15568 9648 15620 9654
rect 15566 9616 15568 9625
rect 15620 9616 15622 9625
rect 15566 9551 15622 9560
rect 15856 8616 15884 12200
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 15856 8588 15976 8616
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15672 7585 15700 8434
rect 15856 8090 15884 8434
rect 15948 8129 15976 8588
rect 15934 8120 15990 8129
rect 15844 8084 15896 8090
rect 15934 8055 15990 8064
rect 15844 8026 15896 8032
rect 15856 7954 15884 8026
rect 16132 7954 16160 8910
rect 16224 8537 16252 12200
rect 16486 11792 16542 11801
rect 16486 11727 16542 11736
rect 16500 11354 16528 11727
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16500 11150 16528 11290
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16592 10470 16620 12200
rect 16960 11218 16988 12200
rect 17328 11558 17356 12200
rect 17696 11626 17724 12200
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 17328 10266 17356 10542
rect 18064 10538 18092 12200
rect 18432 10538 18460 12200
rect 18800 10606 18828 12200
rect 19168 11218 19196 12200
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18708 10266 18736 10406
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 19536 10198 19564 12200
rect 19904 11286 19932 12200
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 20088 11150 20116 11494
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19720 10674 19748 11018
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19720 10266 19748 10610
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19524 10192 19576 10198
rect 17314 10160 17370 10169
rect 19524 10134 19576 10140
rect 20088 10130 20116 11086
rect 20180 10130 20208 11630
rect 17314 10095 17370 10104
rect 20076 10124 20128 10130
rect 17328 10062 17356 10095
rect 20076 10066 20128 10072
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17038 9752 17094 9761
rect 17038 9687 17094 9696
rect 17052 8838 17080 9687
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 16210 8528 16266 8537
rect 16210 8463 16266 8472
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16684 8090 16712 8434
rect 17236 8401 17264 8774
rect 17328 8498 17356 9862
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 17512 9178 17540 9454
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17604 8566 17632 8978
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17684 8560 17736 8566
rect 17972 8514 18000 8842
rect 17684 8502 17736 8508
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17222 8392 17278 8401
rect 17132 8356 17184 8362
rect 17222 8327 17278 8336
rect 17408 8356 17460 8362
rect 17132 8298 17184 8304
rect 17408 8298 17460 8304
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 15658 7576 15714 7585
rect 15658 7511 15714 7520
rect 16028 7336 16080 7342
rect 16026 7304 16028 7313
rect 16080 7304 16082 7313
rect 16026 7239 16082 7248
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 16486 6760 16542 6769
rect 16486 6695 16488 6704
rect 16540 6695 16542 6704
rect 16488 6666 16540 6672
rect 16854 6624 16910 6633
rect 16854 6559 16910 6568
rect 16868 6361 16896 6559
rect 16854 6352 16910 6361
rect 15108 6316 15160 6322
rect 16854 6287 16910 6296
rect 17038 6352 17094 6361
rect 17038 6287 17094 6296
rect 15108 6258 15160 6264
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15948 5914 15976 6190
rect 17052 5953 17080 6287
rect 17038 5944 17094 5953
rect 15936 5908 15988 5914
rect 17038 5879 17094 5888
rect 15936 5850 15988 5856
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 17144 5642 17172 8298
rect 17314 6080 17370 6089
rect 17314 6015 17370 6024
rect 17328 5817 17356 6015
rect 17314 5808 17370 5817
rect 17314 5743 17370 5752
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12530 4448 12586 4457
rect 12530 4383 12586 4392
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11518 3496 11574 3505
rect 11518 3431 11520 3440
rect 11572 3431 11574 3440
rect 11520 3402 11572 3408
rect 11716 3194 11744 3674
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 11164 1358 11192 1838
rect 11242 1456 11298 1465
rect 11624 1426 11652 3130
rect 11992 3058 12020 3334
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11702 2816 11758 2825
rect 11702 2751 11758 2760
rect 11242 1391 11298 1400
rect 11612 1420 11664 1426
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 10968 876 11020 882
rect 10968 818 11020 824
rect 9680 750 9732 756
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 10980 678 11008 818
rect 11256 800 11284 1391
rect 11612 1362 11664 1368
rect 11716 1034 11744 2751
rect 11992 2650 12020 2994
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11796 1828 11848 1834
rect 11796 1770 11848 1776
rect 11808 1426 11836 1770
rect 11796 1420 11848 1426
rect 11796 1362 11848 1368
rect 12084 1034 12112 4218
rect 12544 4185 12572 4383
rect 12530 4176 12586 4185
rect 12530 4111 12586 4120
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14384 3602 14412 4082
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12346 2952 12402 2961
rect 12346 2887 12402 2896
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12176 2106 12204 2586
rect 12164 2100 12216 2106
rect 12164 2042 12216 2048
rect 11624 1006 11744 1034
rect 11992 1006 12112 1034
rect 11624 800 11652 1006
rect 11992 800 12020 1006
rect 12360 800 12388 2887
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 814 12480 2790
rect 13280 2378 13308 2994
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12714 2000 12770 2009
rect 12714 1935 12770 1944
rect 12440 808 12492 814
rect 10968 672 11020 678
rect 10968 614 11020 620
rect 10980 406 11008 614
rect 10968 400 11020 406
rect 10968 342 11020 348
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12728 800 12756 1935
rect 13082 1864 13138 1873
rect 13082 1799 13138 1808
rect 13820 1828 13872 1834
rect 12808 1216 12860 1222
rect 12806 1184 12808 1193
rect 12992 1216 13044 1222
rect 12860 1184 12862 1193
rect 12992 1158 13044 1164
rect 12806 1119 12862 1128
rect 13004 1018 13032 1158
rect 12992 1012 13044 1018
rect 12992 954 13044 960
rect 13096 800 13124 1799
rect 13820 1770 13872 1776
rect 13450 1592 13506 1601
rect 13450 1527 13506 1536
rect 13464 800 13492 1527
rect 13832 800 13860 1770
rect 14200 800 14228 2790
rect 14568 800 14596 3402
rect 15028 2530 15056 5102
rect 16040 4826 16068 5170
rect 17420 4826 17448 8298
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17604 7886 17632 8230
rect 17696 8090 17724 8502
rect 17880 8498 18000 8514
rect 17868 8492 18000 8498
rect 17920 8486 18000 8492
rect 17868 8434 17920 8440
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17972 4622 18000 8298
rect 18064 5234 18092 8910
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18156 8090 18184 8842
rect 18616 8566 18644 9454
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18340 8090 18368 8366
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18616 7886 18644 8502
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18708 7274 18736 7414
rect 18696 7268 18748 7274
rect 18696 7210 18748 7216
rect 18892 5302 18920 7822
rect 19156 7744 19208 7750
rect 19260 7721 19288 9318
rect 19156 7686 19208 7692
rect 19246 7712 19302 7721
rect 19168 7546 19196 7686
rect 19246 7647 19302 7656
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19248 7472 19300 7478
rect 18984 7420 19248 7426
rect 18984 7414 19300 7420
rect 18984 7398 19288 7414
rect 18984 7274 19012 7398
rect 19156 7336 19208 7342
rect 19248 7336 19300 7342
rect 19208 7296 19248 7324
rect 19156 7278 19208 7284
rect 19248 7278 19300 7284
rect 18972 7268 19024 7274
rect 18972 7210 19024 7216
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16316 3738 16344 4014
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 14936 2502 15056 2530
rect 14936 800 14964 2502
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15120 1562 15148 1838
rect 15108 1556 15160 1562
rect 15108 1498 15160 1504
rect 15120 1358 15148 1498
rect 15108 1352 15160 1358
rect 15108 1294 15160 1300
rect 15304 800 15332 3606
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15396 1970 15424 2858
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 15672 800 15700 3538
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15842 2680 15898 2689
rect 15842 2615 15898 2624
rect 15856 2417 15884 2615
rect 15842 2408 15898 2417
rect 15842 2343 15898 2352
rect 16040 800 16068 2994
rect 16408 800 16436 4014
rect 16580 3936 16632 3942
rect 16578 3904 16580 3913
rect 16632 3904 16634 3913
rect 16578 3839 16634 3848
rect 16684 3670 16712 4422
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16776 800 16804 3878
rect 17972 3602 18000 4422
rect 18064 3942 18092 4966
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 17316 3460 17368 3466
rect 17316 3402 17368 3408
rect 17328 3126 17356 3402
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17868 3120 17920 3126
rect 18340 3074 18368 3470
rect 17868 3062 17920 3068
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 17144 800 17172 2926
rect 17500 1284 17552 1290
rect 17500 1226 17552 1232
rect 17224 1216 17276 1222
rect 17224 1158 17276 1164
rect 12440 750 12492 756
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14280 672 14332 678
rect 14280 614 14332 620
rect 14292 105 14320 614
rect 14278 96 14334 105
rect 14278 31 14334 40
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17236 338 17264 1158
rect 17512 800 17540 1226
rect 17880 800 17908 3062
rect 17972 3058 18368 3074
rect 18432 3058 18460 3878
rect 19352 3602 19380 9318
rect 19904 9178 19932 9522
rect 20272 9353 20300 12200
rect 20640 11744 20668 12200
rect 20720 11756 20772 11762
rect 20640 11716 20720 11744
rect 20720 11698 20772 11704
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20824 11082 20852 11630
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20626 9616 20682 9625
rect 20536 9580 20588 9586
rect 20626 9551 20682 9560
rect 20536 9522 20588 9528
rect 20258 9344 20314 9353
rect 20258 9279 20314 9288
rect 20548 9178 20576 9522
rect 20640 9518 20668 9551
rect 20732 9518 20760 10066
rect 20824 9654 20852 11018
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 21008 9466 21036 12200
rect 21376 9518 21404 12200
rect 21638 10704 21694 10713
rect 21638 10639 21640 10648
rect 21692 10639 21694 10648
rect 21640 10610 21692 10616
rect 21744 10441 21772 12200
rect 22112 11286 22140 12200
rect 22388 11762 22416 12718
rect 22466 12200 22522 13000
rect 22834 12200 22890 13000
rect 23202 12200 23258 13000
rect 23296 12572 23348 12578
rect 23296 12514 23348 12520
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22388 11354 22416 11698
rect 22480 11529 22508 12200
rect 22466 11520 22522 11529
rect 22466 11455 22522 11464
rect 22848 11393 22876 12200
rect 23216 12152 23244 12200
rect 23308 12152 23336 12514
rect 23570 12200 23626 13000
rect 23938 12200 23994 13000
rect 24306 12200 24362 13000
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24492 12232 24544 12238
rect 23216 12124 23336 12152
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 22834 11384 22890 11393
rect 22376 11348 22428 11354
rect 22834 11319 22890 11328
rect 22376 11290 22428 11296
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 23400 11150 23428 12038
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23584 10962 23612 12200
rect 23584 10934 23704 10962
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 21730 10432 21786 10441
rect 21730 10367 21786 10376
rect 23584 10062 23612 10746
rect 23388 10056 23440 10062
rect 23386 10024 23388 10033
rect 23572 10056 23624 10062
rect 23440 10024 23442 10033
rect 23572 9998 23624 10004
rect 23386 9959 23442 9968
rect 23676 9897 23704 10934
rect 23952 10305 23980 12200
rect 24216 12096 24268 12102
rect 24320 12084 24348 12200
rect 24492 12174 24544 12180
rect 24504 12084 24532 12174
rect 24320 12056 24532 12084
rect 24216 12038 24268 12044
rect 24228 11286 24256 12038
rect 24596 11762 24624 12242
rect 24674 12200 24730 13000
rect 25042 12200 25098 13000
rect 25410 12200 25466 13000
rect 25778 12200 25834 13000
rect 26146 12200 26202 13000
rect 26240 12640 26292 12646
rect 26240 12582 26292 12588
rect 24688 11937 24716 12200
rect 25056 12073 25084 12200
rect 25042 12064 25098 12073
rect 25042 11999 25098 12008
rect 24674 11928 24730 11937
rect 24674 11863 24730 11872
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24596 11286 24624 11698
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24584 11280 24636 11286
rect 24584 11222 24636 11228
rect 24228 11150 24256 11222
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24320 10538 24348 10950
rect 24688 10810 24716 10950
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24780 10674 24808 10950
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 23938 10296 23994 10305
rect 23938 10231 23994 10240
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 23662 9888 23718 9897
rect 23662 9823 23718 9832
rect 21456 9648 21508 9654
rect 22744 9648 22796 9654
rect 21456 9590 21508 9596
rect 21364 9512 21416 9518
rect 21008 9438 21312 9466
rect 21364 9454 21416 9460
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19536 8838 19564 8910
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19536 6866 19564 8774
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 19536 5914 19564 6190
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19628 4146 19656 8298
rect 19812 7750 19840 8434
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19812 7478 19840 7686
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19904 6866 19932 7346
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19628 3738 19656 4082
rect 20272 3942 20300 9114
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20364 3754 20392 8026
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 20272 3726 20392 3754
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 17960 3052 18368 3058
rect 18012 3046 18368 3052
rect 18420 3052 18472 3058
rect 17960 2994 18012 3000
rect 18604 3052 18656 3058
rect 18420 2994 18472 3000
rect 18524 3012 18604 3040
rect 18524 2938 18552 3012
rect 18604 2994 18656 3000
rect 17972 2910 18552 2938
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18696 2916 18748 2922
rect 17972 2854 18000 2910
rect 18696 2858 18748 2864
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 18340 2582 18368 2790
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18524 2446 18552 2790
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18524 2106 18552 2382
rect 18512 2100 18564 2106
rect 18512 2042 18564 2048
rect 18604 1488 18656 1494
rect 18604 1430 18656 1436
rect 18248 870 18368 898
rect 18248 800 18276 870
rect 18340 814 18368 870
rect 18328 808 18380 814
rect 17224 332 17276 338
rect 17224 274 17276 280
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18052 672 18104 678
rect 18052 614 18104 620
rect 18064 66 18092 614
rect 18052 60 18104 66
rect 18052 2 18104 8
rect 18234 0 18290 800
rect 18616 800 18644 1430
rect 18708 1290 18736 2858
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18892 1358 18920 2382
rect 18880 1352 18932 1358
rect 18880 1294 18932 1300
rect 18696 1284 18748 1290
rect 18696 1226 18748 1232
rect 18984 800 19012 2926
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19352 800 19380 2790
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19628 2310 19656 2382
rect 19720 2310 19748 2858
rect 19616 2304 19668 2310
rect 19616 2246 19668 2252
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 19628 2106 19656 2246
rect 19616 2100 19668 2106
rect 19616 2042 19668 2048
rect 19800 1896 19852 1902
rect 19800 1838 19852 1844
rect 19616 1216 19668 1222
rect 19616 1158 19668 1164
rect 19628 1018 19656 1158
rect 19812 1018 19840 1838
rect 19616 1012 19668 1018
rect 19616 954 19668 960
rect 19800 1012 19852 1018
rect 19800 954 19852 960
rect 19904 898 19932 3674
rect 20272 2446 20300 3726
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20260 2440 20312 2446
rect 20258 2408 20260 2417
rect 20312 2408 20314 2417
rect 20258 2343 20314 2352
rect 20364 1442 20392 2926
rect 19720 870 19932 898
rect 20088 1414 20392 1442
rect 19720 800 19748 870
rect 20088 800 20116 1414
rect 20456 800 20484 3878
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20548 2582 20576 2994
rect 20536 2576 20588 2582
rect 20536 2518 20588 2524
rect 20640 882 20668 7278
rect 20824 7274 20852 7754
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 20916 6866 20944 8366
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 21008 7478 21036 7686
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21100 6798 21128 9318
rect 21284 7290 21312 9438
rect 21468 8906 21496 9590
rect 21560 9574 22048 9602
rect 22796 9596 23244 9602
rect 22744 9590 23244 9596
rect 22756 9574 23244 9590
rect 21560 9110 21588 9574
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21638 9208 21694 9217
rect 21638 9143 21694 9152
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 21652 8566 21680 9143
rect 21836 8838 21864 9454
rect 22020 9382 22048 9574
rect 23216 9518 23244 9574
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22558 9344 22614 9353
rect 21928 8974 21956 9318
rect 22558 9279 22614 9288
rect 22190 9208 22246 9217
rect 22008 9172 22060 9178
rect 22190 9143 22246 9152
rect 22008 9114 22060 9120
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21744 8566 21772 8774
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 21192 7262 21312 7290
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21100 6089 21128 6258
rect 21086 6080 21142 6089
rect 21086 6015 21142 6024
rect 21100 5914 21128 6015
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21192 5846 21220 7262
rect 21272 7200 21324 7206
rect 21376 7188 21404 7414
rect 21324 7160 21404 7188
rect 21272 7142 21324 7148
rect 21376 6866 21404 7160
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20732 3534 20760 5102
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 21100 3534 21128 4014
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20916 2122 20944 3402
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 21100 3233 21128 3334
rect 21086 3224 21142 3233
rect 21086 3159 21142 3168
rect 21088 2440 21140 2446
rect 21086 2408 21088 2417
rect 21140 2408 21142 2417
rect 21086 2343 21142 2352
rect 20732 2094 20944 2122
rect 20732 1426 20760 2094
rect 20720 1420 20772 1426
rect 20720 1362 20772 1368
rect 20812 1216 20864 1222
rect 20812 1158 20864 1164
rect 20628 876 20680 882
rect 20628 818 20680 824
rect 20824 800 20852 1158
rect 21192 800 21220 5510
rect 21284 5302 21312 6598
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21376 5778 21404 6054
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 21272 5296 21324 5302
rect 21272 5238 21324 5244
rect 21376 4690 21404 5714
rect 21468 5234 21496 8366
rect 21836 8090 21864 8434
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21468 4826 21496 5170
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21376 3942 21404 4082
rect 21364 3936 21416 3942
rect 21270 3904 21326 3913
rect 21364 3878 21416 3884
rect 21270 3839 21326 3848
rect 21284 1970 21312 3839
rect 21560 3058 21588 7142
rect 21652 6730 21680 7890
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21744 7274 21772 7822
rect 22020 7426 22048 9114
rect 22204 9110 22232 9143
rect 22192 9104 22244 9110
rect 22192 9046 22244 9052
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22112 7886 22140 8298
rect 22204 8265 22232 8774
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 22190 8256 22246 8265
rect 22190 8191 22246 8200
rect 22296 7954 22324 8570
rect 22572 8537 22600 9279
rect 22848 9042 22876 9386
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22558 8528 22614 8537
rect 22558 8463 22614 8472
rect 22928 8492 22980 8498
rect 23032 8480 23060 9318
rect 23124 8498 23152 9454
rect 23296 8900 23348 8906
rect 23296 8842 23348 8848
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 22980 8452 23060 8480
rect 23112 8492 23164 8498
rect 22928 8434 22980 8440
rect 23112 8434 23164 8440
rect 23020 8356 23072 8362
rect 23020 8298 23072 8304
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 21928 7410 22048 7426
rect 21916 7404 22048 7410
rect 21968 7398 22048 7404
rect 21916 7346 21968 7352
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21928 6458 21956 7346
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22020 5710 22048 6258
rect 22008 5704 22060 5710
rect 22008 5646 22060 5652
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 21652 3998 22140 4026
rect 21652 3194 21680 3998
rect 22008 3936 22060 3942
rect 21730 3904 21786 3913
rect 22008 3878 22060 3884
rect 21730 3839 21786 3848
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21744 3058 21772 3839
rect 21914 3632 21970 3641
rect 21914 3567 21916 3576
rect 21968 3567 21970 3576
rect 21916 3538 21968 3544
rect 22020 3482 22048 3878
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21928 3454 22048 3482
rect 21548 3052 21600 3058
rect 21548 2994 21600 3000
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21546 2816 21602 2825
rect 21546 2751 21602 2760
rect 21560 2417 21588 2751
rect 21744 2582 21772 2994
rect 21732 2576 21784 2582
rect 21732 2518 21784 2524
rect 21546 2408 21602 2417
rect 21546 2343 21602 2352
rect 21272 1964 21324 1970
rect 21272 1906 21324 1912
rect 21272 1760 21324 1766
rect 21272 1702 21324 1708
rect 18328 750 18380 756
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19246 504 19302 513
rect 19246 439 19302 448
rect 19260 406 19288 439
rect 19248 400 19300 406
rect 19248 342 19300 348
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21284 270 21312 1702
rect 21836 1442 21864 3402
rect 21560 1414 21864 1442
rect 21560 800 21588 1414
rect 21928 800 21956 3454
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22020 882 22048 3334
rect 22112 1494 22140 3998
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22204 1562 22232 2246
rect 22192 1556 22244 1562
rect 22192 1498 22244 1504
rect 22100 1488 22152 1494
rect 22100 1430 22152 1436
rect 22008 876 22060 882
rect 22008 818 22060 824
rect 22296 800 22324 4422
rect 22480 3194 22508 6734
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22560 5160 22612 5166
rect 22560 5102 22612 5108
rect 22572 4826 22600 5102
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22560 1896 22612 1902
rect 22560 1838 22612 1844
rect 22572 1766 22600 1838
rect 22560 1760 22612 1766
rect 22560 1702 22612 1708
rect 22572 1426 22600 1702
rect 22560 1420 22612 1426
rect 22560 1362 22612 1368
rect 22664 800 22692 6190
rect 23032 2650 23060 8298
rect 23124 7206 23152 8434
rect 23308 8401 23336 8842
rect 23676 8498 23704 8842
rect 23848 8832 23900 8838
rect 23846 8800 23848 8809
rect 23900 8800 23902 8809
rect 23846 8735 23902 8744
rect 23952 8514 23980 9998
rect 24044 9926 24072 10134
rect 24136 9926 24164 10406
rect 24780 10130 24808 10610
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 24216 9988 24268 9994
rect 24216 9930 24268 9936
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 24228 9722 24256 9930
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 24674 9616 24730 9625
rect 24872 9586 24900 11018
rect 25424 10849 25452 12200
rect 25410 10840 25466 10849
rect 25410 10775 25466 10784
rect 25792 10577 25820 12200
rect 26160 12152 26188 12200
rect 26252 12152 26280 12582
rect 26514 12200 26570 13000
rect 26606 12200 26662 12209
rect 26882 12200 26938 13000
rect 27250 12200 27306 13000
rect 27618 12200 27674 13000
rect 27986 12200 28042 13000
rect 28354 12200 28410 13000
rect 28448 12232 28500 12238
rect 26160 12124 26280 12152
rect 26528 12152 26556 12200
rect 26528 12144 26606 12152
rect 26528 12135 26662 12144
rect 26528 12124 26648 12135
rect 26896 12102 26924 12200
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26608 11756 26660 11762
rect 26608 11698 26660 11704
rect 26146 11656 26202 11665
rect 26146 11591 26202 11600
rect 26056 10804 26108 10810
rect 26056 10746 26108 10752
rect 25872 10668 25924 10674
rect 26068 10656 26096 10746
rect 25924 10628 26096 10656
rect 25872 10610 25924 10616
rect 25778 10568 25834 10577
rect 25778 10503 25834 10512
rect 25884 10198 25912 10610
rect 26160 10470 26188 11591
rect 26620 11286 26648 11698
rect 27264 11694 27292 12200
rect 27632 12170 27660 12200
rect 27620 12164 27672 12170
rect 27620 12106 27672 12112
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27896 12096 27948 12102
rect 27896 12038 27948 12044
rect 27252 11688 27304 11694
rect 27252 11630 27304 11636
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27068 11552 27120 11558
rect 27068 11494 27120 11500
rect 26608 11280 26660 11286
rect 26608 11222 26660 11228
rect 27080 11218 27108 11494
rect 27068 11212 27120 11218
rect 27068 11154 27120 11160
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27264 10674 27292 10950
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 26882 10432 26938 10441
rect 27066 10432 27122 10441
rect 26882 10367 26938 10376
rect 26988 10390 27066 10418
rect 25136 10192 25188 10198
rect 25136 10134 25188 10140
rect 25872 10192 25924 10198
rect 25872 10134 25924 10140
rect 25148 9722 25176 10134
rect 26896 9761 26924 10367
rect 26988 10198 27016 10390
rect 27066 10367 27122 10376
rect 26976 10192 27028 10198
rect 26976 10134 27028 10140
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 26882 9752 26938 9761
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 26792 9716 26844 9722
rect 26882 9687 26938 9696
rect 26792 9658 26844 9664
rect 25318 9616 25374 9625
rect 24674 9551 24730 9560
rect 24860 9580 24912 9586
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24412 8634 24440 8910
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 23664 8492 23716 8498
rect 23952 8486 24072 8514
rect 23664 8434 23716 8440
rect 23294 8392 23350 8401
rect 23294 8327 23350 8336
rect 23676 8090 23704 8434
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23388 7948 23440 7954
rect 23308 7908 23388 7936
rect 23202 7440 23258 7449
rect 23202 7375 23258 7384
rect 23216 7206 23244 7375
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23204 7200 23256 7206
rect 23204 7142 23256 7148
rect 23308 5302 23336 7908
rect 23388 7890 23440 7896
rect 23952 7886 23980 8298
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23584 7398 23888 7426
rect 23584 7342 23612 7398
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 23676 7002 23704 7278
rect 23860 7002 23888 7398
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 23676 6866 23704 6938
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 24044 5710 24072 8486
rect 24688 7342 24716 9551
rect 24860 9522 24912 9528
rect 25136 9580 25188 9586
rect 25318 9551 25320 9560
rect 25136 9522 25188 9528
rect 25372 9551 25374 9560
rect 25320 9522 25372 9528
rect 24872 9178 24900 9522
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 25148 8838 25176 9522
rect 25332 9178 25360 9522
rect 26332 9512 26384 9518
rect 26384 9472 26464 9500
rect 26332 9454 26384 9460
rect 26436 9382 26464 9472
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25412 9172 25464 9178
rect 25884 9160 25912 9318
rect 25964 9172 26016 9178
rect 25884 9132 25964 9160
rect 25412 9114 25464 9120
rect 25964 9114 26016 9120
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24768 7744 24820 7750
rect 24872 7721 24900 7754
rect 24768 7686 24820 7692
rect 24858 7712 24914 7721
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24306 7032 24362 7041
rect 24306 6967 24362 6976
rect 24320 6118 24348 6967
rect 24780 6730 24808 7686
rect 24858 7647 24914 7656
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24964 6322 24992 8774
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25148 8090 25176 8366
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 25056 6662 25084 7346
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24952 6316 25004 6322
rect 24952 6258 25004 6264
rect 24308 6112 24360 6118
rect 24308 6054 24360 6060
rect 24964 5914 24992 6258
rect 24952 5908 25004 5914
rect 24952 5850 25004 5856
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 23296 5296 23348 5302
rect 23296 5238 23348 5244
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 22744 1828 22796 1834
rect 22744 1770 22796 1776
rect 22756 1222 22784 1770
rect 23124 1442 23152 2994
rect 23032 1414 23152 1442
rect 22744 1216 22796 1222
rect 22744 1158 22796 1164
rect 23032 800 23060 1414
rect 23400 800 23428 4966
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 24136 4026 24164 4082
rect 23860 3998 24164 4026
rect 24216 4004 24268 4010
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23492 2514 23520 2790
rect 23768 2650 23796 2926
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23480 2508 23532 2514
rect 23480 2450 23532 2456
rect 23664 1896 23716 1902
rect 23664 1838 23716 1844
rect 23480 1352 23532 1358
rect 23480 1294 23532 1300
rect 23572 1352 23624 1358
rect 23572 1294 23624 1300
rect 21272 264 21324 270
rect 21272 206 21324 212
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23492 406 23520 1294
rect 23584 1222 23612 1294
rect 23572 1216 23624 1222
rect 23572 1158 23624 1164
rect 23676 1018 23704 1838
rect 23860 1442 23888 3998
rect 24216 3946 24268 3952
rect 23940 3936 23992 3942
rect 24228 3890 24256 3946
rect 23992 3884 24256 3890
rect 23940 3878 24256 3884
rect 23952 3862 24256 3878
rect 24872 3670 24900 5578
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 24032 3664 24084 3670
rect 24032 3606 24084 3612
rect 24124 3664 24176 3670
rect 24124 3606 24176 3612
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 23938 3224 23994 3233
rect 23938 3159 23994 3168
rect 23952 2514 23980 3159
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 24044 1494 24072 3606
rect 23768 1414 23888 1442
rect 24032 1488 24084 1494
rect 24032 1430 24084 1436
rect 23664 1012 23716 1018
rect 23664 954 23716 960
rect 23768 800 23796 1414
rect 24032 808 24084 814
rect 23480 400 23532 406
rect 23480 342 23532 348
rect 23754 0 23810 800
rect 24136 800 24164 3606
rect 24492 3596 24544 3602
rect 24492 3538 24544 3544
rect 24504 800 24532 3538
rect 24858 3224 24914 3233
rect 24858 3159 24914 3168
rect 24676 1284 24728 1290
rect 24676 1226 24728 1232
rect 24584 1216 24636 1222
rect 24584 1158 24636 1164
rect 24032 750 24084 756
rect 24044 134 24072 750
rect 24032 128 24084 134
rect 24032 70 24084 76
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24596 241 24624 1158
rect 24688 1018 24716 1226
rect 24676 1012 24728 1018
rect 24676 954 24728 960
rect 24872 800 24900 3159
rect 24964 1018 24992 4422
rect 25056 3738 25084 4422
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 25056 3534 25084 3674
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 25148 2650 25176 6666
rect 25240 2990 25268 8434
rect 25320 5160 25372 5166
rect 25320 5102 25372 5108
rect 25332 4826 25360 5102
rect 25320 4820 25372 4826
rect 25320 4762 25372 4768
rect 25424 4146 25452 9114
rect 26068 8974 26096 9318
rect 25780 8968 25832 8974
rect 25780 8910 25832 8916
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 25504 8900 25556 8906
rect 25504 8842 25556 8848
rect 25516 8022 25544 8842
rect 25688 8628 25740 8634
rect 25608 8588 25688 8616
rect 25608 8498 25636 8588
rect 25688 8570 25740 8576
rect 25792 8498 25820 8910
rect 26068 8634 26096 8910
rect 26148 8900 26200 8906
rect 26148 8842 26200 8848
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25608 8090 25636 8434
rect 25780 8288 25832 8294
rect 25700 8236 25780 8242
rect 25700 8230 25832 8236
rect 25976 8242 26004 8570
rect 25700 8214 25820 8230
rect 25976 8214 26096 8242
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25504 8016 25556 8022
rect 25504 7958 25556 7964
rect 25700 7970 25728 8214
rect 26068 8090 26096 8214
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26160 8022 26188 8842
rect 25872 8016 25924 8022
rect 25700 7942 25820 7970
rect 25872 7958 25924 7964
rect 26148 8016 26200 8022
rect 26148 7958 26200 7964
rect 25792 7886 25820 7942
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 25608 7041 25636 7822
rect 25884 7392 25912 7958
rect 25884 7364 26004 7392
rect 25976 7324 26004 7364
rect 25976 7296 26096 7324
rect 25594 7032 25650 7041
rect 25594 6967 25650 6976
rect 25596 6248 25648 6254
rect 25596 6190 25648 6196
rect 25608 5914 25636 6190
rect 25596 5908 25648 5914
rect 25596 5850 25648 5856
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25688 4072 25740 4078
rect 25688 4014 25740 4020
rect 25412 3664 25464 3670
rect 25412 3606 25464 3612
rect 25424 3233 25452 3606
rect 25516 3602 25544 4014
rect 25700 3618 25728 4014
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25608 3590 25728 3618
rect 25504 3460 25556 3466
rect 25504 3402 25556 3408
rect 25410 3224 25466 3233
rect 25320 3188 25372 3194
rect 25410 3159 25466 3168
rect 25320 3130 25372 3136
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25136 2644 25188 2650
rect 25136 2586 25188 2592
rect 25044 1964 25096 1970
rect 25044 1906 25096 1912
rect 25056 1562 25084 1906
rect 25332 1578 25360 3130
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25424 2650 25452 2994
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 25516 1714 25544 3402
rect 25608 2938 25636 3590
rect 26068 3482 26096 7296
rect 26240 6996 26292 7002
rect 26240 6938 26292 6944
rect 26252 6798 26280 6938
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 26148 4752 26200 4758
rect 26148 4694 26200 4700
rect 25700 3454 26096 3482
rect 25700 3398 25728 3454
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 25872 3392 25924 3398
rect 25872 3334 25924 3340
rect 25608 2910 25728 2938
rect 25700 2854 25728 2910
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25792 2446 25820 2790
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 25516 1686 25636 1714
rect 25044 1556 25096 1562
rect 25044 1498 25096 1504
rect 25240 1550 25360 1578
rect 24952 1012 25004 1018
rect 24952 954 25004 960
rect 25240 800 25268 1550
rect 25608 800 25636 1686
rect 25792 1222 25820 2382
rect 25780 1216 25832 1222
rect 25780 1158 25832 1164
rect 25884 1018 25912 3334
rect 25964 3120 26016 3126
rect 25964 3062 26016 3068
rect 25872 1012 25924 1018
rect 25872 954 25924 960
rect 25884 882 25912 954
rect 25872 876 25924 882
rect 25872 818 25924 824
rect 25976 800 26004 3062
rect 26160 2922 26188 4694
rect 26148 2916 26200 2922
rect 26148 2858 26200 2864
rect 26056 2576 26108 2582
rect 26056 2518 26108 2524
rect 26068 1290 26096 2518
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26160 1358 26188 2382
rect 26252 1970 26280 6258
rect 26344 4146 26372 9318
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26620 8498 26648 8774
rect 26608 8492 26660 8498
rect 26608 8434 26660 8440
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 26422 8256 26478 8265
rect 26422 8191 26478 8200
rect 26436 7721 26464 8191
rect 26516 8084 26568 8090
rect 26712 8072 26740 8366
rect 26568 8044 26740 8072
rect 26516 8026 26568 8032
rect 26422 7712 26478 7721
rect 26422 7647 26478 7656
rect 26436 7398 26740 7426
rect 26436 7342 26464 7398
rect 26712 7342 26740 7398
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 26516 7336 26568 7342
rect 26516 7278 26568 7284
rect 26700 7336 26752 7342
rect 26700 7278 26752 7284
rect 26528 7002 26556 7278
rect 26606 7168 26662 7177
rect 26606 7103 26662 7112
rect 26620 7002 26648 7103
rect 26516 6996 26568 7002
rect 26516 6938 26568 6944
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 26528 6866 26556 6938
rect 26804 6866 26832 9658
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 26988 8838 27016 9522
rect 27172 9432 27200 9998
rect 27356 9586 27384 11630
rect 27540 11558 27568 12038
rect 27436 11552 27488 11558
rect 27436 11494 27488 11500
rect 27528 11552 27580 11558
rect 27528 11494 27580 11500
rect 27448 11082 27476 11494
rect 27436 11076 27488 11082
rect 27436 11018 27488 11024
rect 27540 11070 27844 11098
rect 27540 11014 27568 11070
rect 27528 11008 27580 11014
rect 27528 10950 27580 10956
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27436 10668 27488 10674
rect 27632 10656 27660 10950
rect 27488 10628 27660 10656
rect 27436 10610 27488 10616
rect 27436 10464 27488 10470
rect 27436 10406 27488 10412
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 27448 9586 27476 10406
rect 27540 9994 27568 10406
rect 27632 10130 27660 10628
rect 27816 10606 27844 11070
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27804 10464 27856 10470
rect 27710 10432 27766 10441
rect 27804 10406 27856 10412
rect 27710 10367 27766 10376
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27724 9994 27752 10367
rect 27816 10062 27844 10406
rect 27908 10198 27936 12038
rect 28000 11354 28028 12200
rect 28368 11626 28396 12200
rect 28722 12200 28778 13000
rect 29000 12436 29052 12442
rect 29000 12378 29052 12384
rect 28448 12174 28500 12180
rect 28460 11626 28488 12174
rect 28736 11642 28764 12200
rect 29012 11762 29040 12378
rect 29090 12200 29146 13000
rect 29184 12232 29236 12238
rect 29104 11898 29132 12200
rect 29458 12200 29514 13000
rect 29826 12200 29882 13000
rect 30194 12200 30250 13000
rect 30562 12200 30618 13000
rect 30654 12880 30710 12889
rect 30654 12815 30710 12824
rect 29184 12174 29236 12180
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 28356 11620 28408 11626
rect 28356 11562 28408 11568
rect 28448 11620 28500 11626
rect 28736 11614 28856 11642
rect 28448 11562 28500 11568
rect 28262 11520 28318 11529
rect 28262 11455 28318 11464
rect 28078 11384 28134 11393
rect 27988 11348 28040 11354
rect 28078 11319 28134 11328
rect 27988 11290 28040 11296
rect 27988 10464 28040 10470
rect 27988 10406 28040 10412
rect 27896 10192 27948 10198
rect 27896 10134 27948 10140
rect 27804 10056 27856 10062
rect 27804 9998 27856 10004
rect 27896 10056 27948 10062
rect 27896 9998 27948 10004
rect 27528 9988 27580 9994
rect 27528 9930 27580 9936
rect 27712 9988 27764 9994
rect 27712 9930 27764 9936
rect 27816 9722 27844 9998
rect 27620 9716 27672 9722
rect 27620 9658 27672 9664
rect 27804 9716 27856 9722
rect 27804 9658 27856 9664
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27436 9444 27488 9450
rect 27172 9404 27436 9432
rect 27436 9386 27488 9392
rect 27632 9042 27660 9658
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27620 9036 27672 9042
rect 27620 8978 27672 8984
rect 27540 8922 27568 8978
rect 27540 8894 27660 8922
rect 27632 8838 27660 8894
rect 26976 8832 27028 8838
rect 26976 8774 27028 8780
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27540 8634 27568 8774
rect 27528 8628 27580 8634
rect 27528 8570 27580 8576
rect 27618 8392 27674 8401
rect 27618 8327 27674 8336
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27540 7546 27568 7822
rect 27632 7750 27660 8327
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27632 7342 27660 7482
rect 27620 7336 27672 7342
rect 27620 7278 27672 7284
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27816 6390 27844 6598
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26528 5846 26556 6258
rect 26974 6080 27030 6089
rect 26974 6015 27030 6024
rect 26792 5908 26844 5914
rect 26792 5850 26844 5856
rect 26516 5840 26568 5846
rect 26804 5817 26832 5850
rect 26988 5817 27016 6015
rect 26516 5782 26568 5788
rect 26790 5808 26846 5817
rect 26790 5743 26846 5752
rect 26974 5808 27030 5817
rect 26974 5743 27030 5752
rect 26424 5704 26476 5710
rect 26424 5646 26476 5652
rect 26436 5302 26464 5646
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26424 5296 26476 5302
rect 26424 5238 26476 5244
rect 26424 4548 26476 4554
rect 26424 4490 26476 4496
rect 26332 4140 26384 4146
rect 26332 4082 26384 4088
rect 26344 3738 26372 4082
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 26330 3224 26386 3233
rect 26330 3159 26386 3168
rect 26240 1964 26292 1970
rect 26240 1906 26292 1912
rect 26344 1902 26372 3159
rect 26332 1896 26384 1902
rect 26332 1838 26384 1844
rect 26240 1760 26292 1766
rect 26238 1728 26240 1737
rect 26292 1728 26294 1737
rect 26238 1663 26294 1672
rect 26436 1442 26464 4490
rect 26528 2854 26556 5510
rect 27802 5400 27858 5409
rect 27802 5335 27858 5344
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26700 4004 26752 4010
rect 26700 3946 26752 3952
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 26516 2576 26568 2582
rect 26516 2518 26568 2524
rect 26528 2310 26556 2518
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 26608 1896 26660 1902
rect 26606 1864 26608 1873
rect 26660 1864 26662 1873
rect 26606 1799 26662 1808
rect 26344 1414 26464 1442
rect 26148 1352 26200 1358
rect 26148 1294 26200 1300
rect 26056 1284 26108 1290
rect 26056 1226 26108 1232
rect 26160 1018 26188 1294
rect 26148 1012 26200 1018
rect 26148 954 26200 960
rect 26344 800 26372 1414
rect 26516 1352 26568 1358
rect 26516 1294 26568 1300
rect 24582 232 24638 241
rect 24582 167 24638 176
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26528 678 26556 1294
rect 26712 800 26740 3946
rect 26988 3670 27016 4626
rect 27816 4298 27844 5335
rect 27908 4826 27936 9998
rect 28000 9926 28028 10406
rect 28092 9926 28120 11319
rect 28276 11218 28304 11455
rect 28430 11452 28726 11472
rect 28486 11450 28510 11452
rect 28566 11450 28590 11452
rect 28646 11450 28670 11452
rect 28508 11398 28510 11450
rect 28572 11398 28584 11450
rect 28646 11398 28648 11450
rect 28486 11396 28510 11398
rect 28566 11396 28590 11398
rect 28646 11396 28670 11398
rect 28430 11376 28726 11396
rect 28724 11280 28776 11286
rect 28724 11222 28776 11228
rect 28264 11212 28316 11218
rect 28264 11154 28316 11160
rect 28736 10452 28764 11222
rect 28828 10742 28856 11614
rect 29196 11354 29224 12174
rect 29368 11688 29420 11694
rect 29368 11630 29420 11636
rect 29380 11354 29408 11630
rect 29184 11348 29236 11354
rect 29184 11290 29236 11296
rect 29368 11348 29420 11354
rect 29368 11290 29420 11296
rect 29092 11076 29144 11082
rect 29092 11018 29144 11024
rect 29104 10742 29132 11018
rect 28816 10736 28868 10742
rect 28816 10678 28868 10684
rect 29092 10736 29144 10742
rect 29092 10678 29144 10684
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 28736 10424 28856 10452
rect 28430 10364 28726 10384
rect 28486 10362 28510 10364
rect 28566 10362 28590 10364
rect 28646 10362 28670 10364
rect 28508 10310 28510 10362
rect 28572 10310 28584 10362
rect 28646 10310 28648 10362
rect 28486 10308 28510 10310
rect 28566 10308 28590 10310
rect 28646 10308 28670 10310
rect 28262 10296 28318 10305
rect 28430 10288 28726 10308
rect 28318 10254 28396 10282
rect 28262 10231 28318 10240
rect 27988 9920 28040 9926
rect 27988 9862 28040 9868
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 28368 9500 28396 10254
rect 28828 9722 28856 10424
rect 29012 10198 29040 10610
rect 29472 10606 29500 12200
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29460 10600 29512 10606
rect 29460 10542 29512 10548
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29104 10266 29408 10282
rect 29092 10260 29408 10266
rect 29144 10254 29408 10260
rect 29092 10202 29144 10208
rect 29000 10192 29052 10198
rect 28998 10160 29000 10169
rect 29052 10160 29054 10169
rect 29380 10130 29408 10254
rect 28998 10095 29054 10104
rect 29368 10124 29420 10130
rect 29012 10069 29040 10095
rect 29368 10066 29420 10072
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 29012 9738 29040 9862
rect 29564 9738 29592 10542
rect 29656 9926 29684 11086
rect 29644 9920 29696 9926
rect 29644 9862 29696 9868
rect 28816 9716 28868 9722
rect 29012 9710 29592 9738
rect 28816 9658 28868 9664
rect 28368 9472 29408 9500
rect 29380 9382 29408 9472
rect 29840 9450 29868 12200
rect 30208 9586 30236 12200
rect 30576 10742 30604 12200
rect 30668 12102 30696 12815
rect 30930 12200 30986 13000
rect 31298 12200 31354 13000
rect 31666 12200 31722 13000
rect 32034 12200 32090 13000
rect 32220 12912 32272 12918
rect 32220 12854 32272 12860
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30748 12096 30800 12102
rect 30748 12038 30800 12044
rect 30760 11286 30788 12038
rect 30944 11830 30972 12200
rect 31114 12064 31170 12073
rect 31114 11999 31170 12008
rect 30932 11824 30984 11830
rect 30932 11766 30984 11772
rect 30748 11280 30800 11286
rect 30748 11222 30800 11228
rect 30760 11150 30788 11222
rect 30748 11144 30800 11150
rect 30748 11086 30800 11092
rect 30564 10736 30616 10742
rect 30564 10678 30616 10684
rect 30748 10668 30800 10674
rect 30748 10610 30800 10616
rect 30760 10266 30788 10610
rect 30748 10260 30800 10266
rect 30748 10202 30800 10208
rect 30746 10160 30802 10169
rect 30746 10095 30802 10104
rect 30760 9994 30788 10095
rect 30748 9988 30800 9994
rect 30748 9930 30800 9936
rect 30288 9920 30340 9926
rect 31128 9897 31156 11999
rect 31206 11928 31262 11937
rect 31206 11863 31262 11872
rect 31220 10169 31248 11863
rect 31312 11354 31340 12200
rect 31482 11928 31538 11937
rect 31482 11863 31538 11872
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31392 10668 31444 10674
rect 31392 10610 31444 10616
rect 31206 10160 31262 10169
rect 31206 10095 31262 10104
rect 30288 9862 30340 9868
rect 31114 9888 31170 9897
rect 30300 9586 30328 9862
rect 31114 9823 31170 9832
rect 31404 9722 31432 10610
rect 31496 10470 31524 11863
rect 31576 11688 31628 11694
rect 31576 11630 31628 11636
rect 31588 10538 31616 11630
rect 31680 10742 31708 12200
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 31850 11384 31906 11393
rect 31850 11319 31906 11328
rect 31668 10736 31720 10742
rect 31668 10678 31720 10684
rect 31576 10532 31628 10538
rect 31576 10474 31628 10480
rect 31484 10464 31536 10470
rect 31484 10406 31536 10412
rect 31864 10169 31892 11319
rect 31956 11218 31984 12038
rect 32048 11898 32076 12200
rect 32036 11892 32088 11898
rect 32036 11834 32088 11840
rect 32126 11520 32182 11529
rect 32126 11455 32182 11464
rect 31944 11212 31996 11218
rect 31944 11154 31996 11160
rect 32140 11082 32168 11455
rect 32128 11076 32180 11082
rect 32128 11018 32180 11024
rect 32232 10674 32260 12854
rect 32402 12200 32458 13000
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32508 12306 32536 12378
rect 32496 12300 32548 12306
rect 32496 12242 32548 12248
rect 32770 12200 32826 13000
rect 33138 12200 33194 13000
rect 33414 12200 33470 12209
rect 33506 12200 33562 13000
rect 41142 13016 41198 13025
rect 33690 12951 33746 12960
rect 33598 12608 33654 12617
rect 33598 12543 33654 12552
rect 32416 11218 32444 12200
rect 32496 12164 32548 12170
rect 32496 12106 32548 12112
rect 32404 11212 32456 11218
rect 32404 11154 32456 11160
rect 32508 11150 32536 12106
rect 32588 11756 32640 11762
rect 32588 11698 32640 11704
rect 32600 11218 32628 11698
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32312 11008 32364 11014
rect 32312 10950 32364 10956
rect 32496 11008 32548 11014
rect 32496 10950 32548 10956
rect 32324 10674 32352 10950
rect 32220 10668 32272 10674
rect 32220 10610 32272 10616
rect 32312 10668 32364 10674
rect 32312 10610 32364 10616
rect 31850 10160 31906 10169
rect 31850 10095 31906 10104
rect 32232 9926 32260 10610
rect 32404 10056 32456 10062
rect 32508 10044 32536 10950
rect 32784 10742 32812 12200
rect 33152 11354 33180 12200
rect 33414 12135 33470 12144
rect 33230 12064 33286 12073
rect 33230 11999 33286 12008
rect 33140 11348 33192 11354
rect 33140 11290 33192 11296
rect 32772 10736 32824 10742
rect 32772 10678 32824 10684
rect 32588 10464 32640 10470
rect 32588 10406 32640 10412
rect 32600 10062 32628 10406
rect 32456 10016 32536 10044
rect 32588 10056 32640 10062
rect 32404 9998 32456 10004
rect 32588 9998 32640 10004
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 32220 9920 32272 9926
rect 32220 9862 32272 9868
rect 32600 9722 32628 9998
rect 31392 9716 31444 9722
rect 31392 9658 31444 9664
rect 32588 9716 32640 9722
rect 32588 9658 32640 9664
rect 30196 9580 30248 9586
rect 30196 9522 30248 9528
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 31484 9580 31536 9586
rect 31944 9580 31996 9586
rect 31484 9522 31536 9528
rect 31864 9540 31944 9568
rect 29828 9444 29880 9450
rect 29828 9386 29880 9392
rect 29276 9376 29328 9382
rect 28276 9353 28856 9364
rect 28262 9344 28870 9353
rect 28318 9336 28814 9344
rect 28262 9279 28318 9288
rect 28430 9276 28726 9296
rect 29276 9318 29328 9324
rect 29368 9376 29420 9382
rect 29368 9318 29420 9324
rect 28814 9279 28870 9288
rect 28486 9274 28510 9276
rect 28566 9274 28590 9276
rect 28646 9274 28670 9276
rect 28508 9222 28510 9274
rect 28572 9222 28584 9274
rect 28646 9222 28648 9274
rect 28486 9220 28510 9222
rect 28566 9220 28590 9222
rect 28646 9220 28670 9222
rect 28262 9208 28318 9217
rect 28172 9172 28224 9178
rect 28430 9200 28726 9220
rect 28814 9208 28870 9217
rect 28262 9143 28318 9152
rect 28814 9143 28816 9152
rect 28172 9114 28224 9120
rect 28080 8968 28132 8974
rect 28184 8956 28212 9114
rect 28276 9092 28304 9143
rect 28868 9143 28870 9152
rect 28816 9114 28868 9120
rect 28276 9064 28488 9092
rect 28356 8968 28408 8974
rect 28184 8928 28356 8956
rect 28080 8910 28132 8916
rect 28356 8910 28408 8916
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 28000 6662 28028 6734
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 28092 5778 28120 8910
rect 28460 8378 28488 9064
rect 29184 8968 29236 8974
rect 29184 8910 29236 8916
rect 29196 8430 29224 8910
rect 29288 8430 29316 9318
rect 30300 9178 30328 9522
rect 31496 9382 31524 9522
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 31484 9376 31536 9382
rect 31484 9318 31536 9324
rect 31668 9376 31720 9382
rect 31668 9318 31720 9324
rect 30288 9172 30340 9178
rect 30288 9114 30340 9120
rect 29184 8424 29236 8430
rect 28998 8392 29054 8401
rect 28460 8350 28998 8378
rect 29184 8366 29236 8372
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 28998 8327 29054 8336
rect 28430 8188 28726 8208
rect 28486 8186 28510 8188
rect 28566 8186 28590 8188
rect 28646 8186 28670 8188
rect 28508 8134 28510 8186
rect 28572 8134 28584 8186
rect 28646 8134 28648 8186
rect 28486 8132 28510 8134
rect 28566 8132 28590 8134
rect 28646 8132 28670 8134
rect 28430 8112 28726 8132
rect 28908 7404 28960 7410
rect 28908 7346 28960 7352
rect 28920 7206 28948 7346
rect 28816 7200 28868 7206
rect 28814 7168 28816 7177
rect 28908 7200 28960 7206
rect 28868 7168 28870 7177
rect 28430 7100 28726 7120
rect 28908 7142 28960 7148
rect 28814 7103 28870 7112
rect 28486 7098 28510 7100
rect 28566 7098 28590 7100
rect 28646 7098 28670 7100
rect 28508 7046 28510 7098
rect 28572 7046 28584 7098
rect 28646 7046 28648 7098
rect 28486 7044 28510 7046
rect 28566 7044 28590 7046
rect 28646 7044 28670 7046
rect 28170 7032 28226 7041
rect 28430 7024 28726 7044
rect 28814 7032 28870 7041
rect 28170 6967 28226 6976
rect 28814 6967 28816 6976
rect 28184 6798 28212 6967
rect 28868 6967 28870 6976
rect 28816 6938 28868 6944
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28264 6656 28316 6662
rect 28356 6656 28408 6662
rect 28316 6616 28356 6644
rect 28264 6598 28316 6604
rect 28356 6598 28408 6604
rect 29288 6186 29316 6802
rect 30852 6322 30880 9318
rect 31680 9110 31708 9318
rect 31668 9104 31720 9110
rect 31668 9046 31720 9052
rect 31864 8974 31892 9540
rect 31944 9522 31996 9528
rect 31944 9444 31996 9450
rect 31944 9386 31996 9392
rect 31956 8974 31984 9386
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 32496 7268 32548 7274
rect 32496 7210 32548 7216
rect 31758 7168 31814 7177
rect 31758 7103 31814 7112
rect 31772 7018 31800 7103
rect 32034 7032 32090 7041
rect 31772 6990 32034 7018
rect 32034 6967 32090 6976
rect 31116 6452 31168 6458
rect 31116 6394 31168 6400
rect 29828 6316 29880 6322
rect 29828 6258 29880 6264
rect 30380 6316 30432 6322
rect 30380 6258 30432 6264
rect 30840 6316 30892 6322
rect 30840 6258 30892 6264
rect 29276 6180 29328 6186
rect 29276 6122 29328 6128
rect 29092 6112 29144 6118
rect 28814 6080 28870 6089
rect 28430 6012 28726 6032
rect 29092 6054 29144 6060
rect 28814 6015 28870 6024
rect 28486 6010 28510 6012
rect 28566 6010 28590 6012
rect 28646 6010 28670 6012
rect 28508 5958 28510 6010
rect 28572 5958 28584 6010
rect 28646 5958 28648 6010
rect 28486 5956 28510 5958
rect 28566 5956 28590 5958
rect 28646 5956 28670 5958
rect 28262 5944 28318 5953
rect 28430 5936 28726 5956
rect 28828 5914 28856 6015
rect 28262 5879 28318 5888
rect 28816 5908 28868 5914
rect 28276 5794 28304 5879
rect 28816 5850 28868 5856
rect 28998 5808 29054 5817
rect 28080 5772 28132 5778
rect 28276 5766 28998 5794
rect 28998 5743 29054 5752
rect 28080 5714 28132 5720
rect 27988 5704 28040 5710
rect 27988 5646 28040 5652
rect 27896 4820 27948 4826
rect 27896 4762 27948 4768
rect 27816 4270 27936 4298
rect 27804 4140 27856 4146
rect 27804 4082 27856 4088
rect 26976 3664 27028 3670
rect 26976 3606 27028 3612
rect 27252 3664 27304 3670
rect 27252 3606 27304 3612
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 26792 1964 26844 1970
rect 26792 1906 26844 1912
rect 26804 1562 26832 1906
rect 26792 1556 26844 1562
rect 26792 1498 26844 1504
rect 27080 800 27108 3402
rect 27264 3369 27292 3606
rect 27250 3360 27306 3369
rect 27250 3295 27306 3304
rect 27434 3360 27490 3369
rect 27434 3295 27490 3304
rect 27448 3058 27476 3295
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27344 2916 27396 2922
rect 27344 2858 27396 2864
rect 27356 2446 27384 2858
rect 27448 2650 27476 2994
rect 27620 2848 27672 2854
rect 27540 2796 27620 2802
rect 27540 2790 27672 2796
rect 27540 2774 27660 2790
rect 27436 2644 27488 2650
rect 27436 2586 27488 2592
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 27356 1358 27384 2382
rect 27540 1442 27568 2774
rect 27448 1414 27568 1442
rect 27344 1352 27396 1358
rect 27344 1294 27396 1300
rect 27448 800 27476 1414
rect 27712 1352 27764 1358
rect 27712 1294 27764 1300
rect 27528 808 27580 814
rect 26516 672 26568 678
rect 26516 614 26568 620
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27528 750 27580 756
rect 27540 474 27568 750
rect 27724 513 27752 1294
rect 27816 800 27844 4082
rect 27908 882 27936 4270
rect 28000 3738 28028 5646
rect 29104 5409 29132 6054
rect 28906 5400 28962 5409
rect 28906 5335 28962 5344
rect 29090 5400 29146 5409
rect 29090 5335 29146 5344
rect 28920 5114 28948 5335
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 28998 5128 29054 5137
rect 28920 5086 28998 5114
rect 28998 5063 29054 5072
rect 28430 4924 28726 4944
rect 28486 4922 28510 4924
rect 28566 4922 28590 4924
rect 28646 4922 28670 4924
rect 28508 4870 28510 4922
rect 28572 4870 28584 4922
rect 28646 4870 28648 4922
rect 28486 4868 28510 4870
rect 28566 4868 28590 4870
rect 28646 4868 28670 4870
rect 28430 4848 28726 4868
rect 29196 4865 29224 5170
rect 29182 4856 29238 4865
rect 29182 4791 29238 4800
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28078 3768 28134 3777
rect 27988 3732 28040 3738
rect 28184 3754 28212 4558
rect 28998 4040 29054 4049
rect 28276 3998 28998 4026
rect 28276 3913 28304 3998
rect 28998 3975 29054 3984
rect 28262 3904 28318 3913
rect 28814 3904 28870 3913
rect 28262 3839 28318 3848
rect 28430 3836 28726 3856
rect 28814 3839 28870 3848
rect 28486 3834 28510 3836
rect 28566 3834 28590 3836
rect 28646 3834 28670 3836
rect 28508 3782 28510 3834
rect 28572 3782 28584 3834
rect 28646 3782 28648 3834
rect 28486 3780 28510 3782
rect 28566 3780 28590 3782
rect 28646 3780 28670 3782
rect 28430 3760 28726 3780
rect 28184 3726 28396 3754
rect 28078 3703 28080 3712
rect 27988 3674 28040 3680
rect 28132 3703 28134 3712
rect 28080 3674 28132 3680
rect 28000 3534 28028 3674
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 28172 2984 28224 2990
rect 28172 2926 28224 2932
rect 28080 1420 28132 1426
rect 28080 1362 28132 1368
rect 27988 1012 28040 1018
rect 27988 954 28040 960
rect 27896 876 27948 882
rect 27896 818 27948 824
rect 27710 504 27766 513
rect 27528 468 27580 474
rect 27710 439 27766 448
rect 27528 410 27580 416
rect 27802 0 27858 800
rect 28000 746 28028 954
rect 28092 746 28120 1362
rect 28184 800 28212 2926
rect 28262 2680 28318 2689
rect 28262 2615 28264 2624
rect 28316 2615 28318 2624
rect 28264 2586 28316 2592
rect 28264 1896 28316 1902
rect 28264 1838 28316 1844
rect 28276 1562 28304 1838
rect 28264 1556 28316 1562
rect 28264 1498 28316 1504
rect 28276 1340 28304 1498
rect 28368 1442 28396 3726
rect 28828 2825 28856 3839
rect 28906 3768 28962 3777
rect 28906 3703 28908 3712
rect 28960 3703 28962 3712
rect 28908 3674 28960 3680
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 28814 2816 28870 2825
rect 28430 2748 28726 2768
rect 28814 2751 28870 2760
rect 28486 2746 28510 2748
rect 28566 2746 28590 2748
rect 28646 2746 28670 2748
rect 28508 2694 28510 2746
rect 28572 2694 28584 2746
rect 28646 2694 28648 2746
rect 28486 2692 28510 2694
rect 28566 2692 28590 2694
rect 28646 2692 28670 2694
rect 28430 2672 28726 2692
rect 28814 2680 28870 2689
rect 28814 2615 28816 2624
rect 28868 2615 28870 2624
rect 28816 2586 28868 2592
rect 28816 1964 28868 1970
rect 28816 1906 28868 1912
rect 28430 1660 28726 1680
rect 28486 1658 28510 1660
rect 28566 1658 28590 1660
rect 28646 1658 28670 1660
rect 28508 1606 28510 1658
rect 28572 1606 28584 1658
rect 28646 1606 28648 1658
rect 28486 1604 28510 1606
rect 28566 1604 28590 1606
rect 28646 1604 28670 1606
rect 28430 1584 28726 1604
rect 28828 1601 28856 1906
rect 28814 1592 28870 1601
rect 28814 1527 28870 1536
rect 28368 1414 28580 1442
rect 28356 1352 28408 1358
rect 28276 1312 28356 1340
rect 28356 1294 28408 1300
rect 28552 800 28580 1414
rect 28632 1420 28684 1426
rect 28632 1362 28684 1368
rect 28644 1290 28672 1362
rect 28632 1284 28684 1290
rect 28632 1226 28684 1232
rect 28920 800 28948 3130
rect 28998 1864 29054 1873
rect 28998 1799 29054 1808
rect 29012 1766 29040 1799
rect 29000 1760 29052 1766
rect 29000 1702 29052 1708
rect 29000 808 29052 814
rect 27988 740 28040 746
rect 27988 682 28040 688
rect 28080 740 28132 746
rect 28080 682 28132 688
rect 28170 0 28226 800
rect 28538 592 28594 800
rect 28816 672 28868 678
rect 28816 614 28868 620
rect 28430 572 28726 592
rect 28486 570 28510 572
rect 28566 570 28590 572
rect 28646 570 28670 572
rect 28508 518 28510 570
rect 28572 518 28584 570
rect 28646 518 28648 570
rect 28486 516 28510 518
rect 28566 516 28590 518
rect 28646 516 28670 518
rect 28430 496 28726 516
rect 28538 0 28594 496
rect 28828 474 28856 614
rect 28816 468 28868 474
rect 28816 410 28868 416
rect 28906 0 28962 800
rect 29288 800 29316 5170
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 29656 3738 29684 5102
rect 29736 4820 29788 4826
rect 29736 4762 29788 4768
rect 29644 3732 29696 3738
rect 29644 3674 29696 3680
rect 29552 3460 29604 3466
rect 29552 3402 29604 3408
rect 29564 3194 29592 3402
rect 29644 3392 29696 3398
rect 29644 3334 29696 3340
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29656 3058 29684 3334
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29656 2650 29684 2994
rect 29644 2644 29696 2650
rect 29644 2586 29696 2592
rect 29748 1442 29776 4762
rect 29840 4214 29868 6258
rect 30392 5914 30420 6258
rect 31128 6254 31156 6394
rect 31116 6248 31168 6254
rect 31116 6190 31168 6196
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30392 4758 30420 5510
rect 31758 5264 31814 5273
rect 31758 5199 31814 5208
rect 31496 5086 31708 5114
rect 30838 4856 30894 4865
rect 30838 4791 30894 4800
rect 31390 4856 31446 4865
rect 31390 4791 31446 4800
rect 30380 4752 30432 4758
rect 30380 4694 30432 4700
rect 30472 4684 30524 4690
rect 30472 4626 30524 4632
rect 30484 4570 30512 4626
rect 30748 4616 30800 4622
rect 30484 4564 30748 4570
rect 30484 4558 30800 4564
rect 30484 4542 30788 4558
rect 30852 4554 30880 4791
rect 30840 4548 30892 4554
rect 30840 4490 30892 4496
rect 29828 4208 29880 4214
rect 29828 4150 29880 4156
rect 31116 4208 31168 4214
rect 31116 4150 31168 4156
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 29656 1414 29776 1442
rect 29656 800 29684 1414
rect 30024 800 30052 3674
rect 30380 3188 30432 3194
rect 30380 3130 30432 3136
rect 30288 2916 30340 2922
rect 30288 2858 30340 2864
rect 30104 1964 30156 1970
rect 30104 1906 30156 1912
rect 30116 882 30144 1906
rect 30300 1494 30328 2858
rect 30288 1488 30340 1494
rect 30288 1430 30340 1436
rect 30288 1216 30340 1222
rect 30288 1158 30340 1164
rect 30300 1018 30328 1158
rect 30196 1012 30248 1018
rect 30196 954 30248 960
rect 30288 1012 30340 1018
rect 30288 954 30340 960
rect 30104 876 30156 882
rect 30104 818 30156 824
rect 29052 768 29132 796
rect 29000 750 29052 756
rect 29104 513 29132 768
rect 29090 504 29146 513
rect 29090 439 29146 448
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30208 678 30236 954
rect 30392 800 30420 3130
rect 30760 3126 30788 3878
rect 30748 3120 30800 3126
rect 30748 3062 30800 3068
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 30944 2650 30972 2994
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 30840 2304 30892 2310
rect 30840 2246 30892 2252
rect 30472 1964 30524 1970
rect 30472 1906 30524 1912
rect 30484 1562 30512 1906
rect 30472 1556 30524 1562
rect 30472 1498 30524 1504
rect 30748 1556 30800 1562
rect 30748 1498 30800 1504
rect 30760 800 30788 1498
rect 30852 1358 30880 2246
rect 30840 1352 30892 1358
rect 30840 1294 30892 1300
rect 30840 1216 30892 1222
rect 30840 1158 30892 1164
rect 30196 672 30248 678
rect 30196 614 30248 620
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 30852 202 30880 1158
rect 31128 800 31156 4150
rect 31300 4004 31352 4010
rect 31300 3946 31352 3952
rect 31206 3360 31262 3369
rect 31206 3295 31262 3304
rect 31220 3058 31248 3295
rect 31208 3052 31260 3058
rect 31208 2994 31260 3000
rect 31312 2020 31340 3946
rect 31404 3097 31432 4791
rect 31496 4622 31524 5086
rect 31680 5030 31708 5086
rect 31576 5024 31628 5030
rect 31576 4966 31628 4972
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 31772 4978 31800 5199
rect 32218 4992 32274 5001
rect 31588 4842 31616 4966
rect 31772 4950 32218 4978
rect 32218 4927 32274 4936
rect 31588 4814 31708 4842
rect 31484 4616 31536 4622
rect 31484 4558 31536 4564
rect 31680 4282 31708 4814
rect 31852 4548 31904 4554
rect 31852 4490 31904 4496
rect 31864 4282 31892 4490
rect 32508 4486 32536 7210
rect 32496 4480 32548 4486
rect 32496 4422 32548 4428
rect 31576 4276 31628 4282
rect 31576 4218 31628 4224
rect 31668 4276 31720 4282
rect 31668 4218 31720 4224
rect 31852 4276 31904 4282
rect 31852 4218 31904 4224
rect 32220 4276 32272 4282
rect 32220 4218 32272 4224
rect 31588 4162 31616 4218
rect 31588 4134 31708 4162
rect 31390 3088 31446 3097
rect 31390 3023 31446 3032
rect 31680 2990 31708 4134
rect 31942 3224 31998 3233
rect 31942 3159 31998 3168
rect 31956 3058 31984 3159
rect 31944 3052 31996 3058
rect 31944 2994 31996 3000
rect 31668 2984 31720 2990
rect 31668 2926 31720 2932
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 31864 2825 31892 2926
rect 31850 2816 31906 2825
rect 31850 2751 31906 2760
rect 31852 2304 31904 2310
rect 31852 2246 31904 2252
rect 31312 1992 31524 2020
rect 31496 800 31524 1992
rect 31864 800 31892 2246
rect 31944 1012 31996 1018
rect 31944 954 31996 960
rect 30840 196 30892 202
rect 30840 138 30892 144
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 31956 785 31984 954
rect 32232 800 32260 4218
rect 32692 4146 32720 9998
rect 33244 8566 33272 11999
rect 33428 11286 33456 12135
rect 33520 11830 33548 12200
rect 33508 11824 33560 11830
rect 33508 11766 33560 11772
rect 33416 11280 33468 11286
rect 33416 11222 33468 11228
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33428 9926 33456 9998
rect 33416 9920 33468 9926
rect 33416 9862 33468 9868
rect 33428 9722 33456 9862
rect 33416 9716 33468 9722
rect 33416 9658 33468 9664
rect 33324 9648 33376 9654
rect 33324 9590 33376 9596
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 33232 8560 33284 8566
rect 33232 8502 33284 8508
rect 33336 8265 33364 9590
rect 33520 8838 33548 9590
rect 33508 8832 33560 8838
rect 33508 8774 33560 8780
rect 33612 8634 33640 12543
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33322 8256 33378 8265
rect 33322 8191 33378 8200
rect 33704 7206 33732 12951
rect 33782 12336 33838 12345
rect 33782 12271 33838 12280
rect 33796 8362 33824 12271
rect 33874 12200 33930 13000
rect 33966 12744 34022 12753
rect 33966 12679 34022 12688
rect 33888 10742 33916 12200
rect 33876 10736 33928 10742
rect 33876 10678 33928 10684
rect 33876 10260 33928 10266
rect 33876 10202 33928 10208
rect 33888 9994 33916 10202
rect 33876 9988 33928 9994
rect 33876 9930 33928 9936
rect 33784 8356 33836 8362
rect 33784 8298 33836 8304
rect 33784 7812 33836 7818
rect 33784 7754 33836 7760
rect 33876 7812 33928 7818
rect 33876 7754 33928 7760
rect 33692 7200 33744 7206
rect 33692 7142 33744 7148
rect 33796 7002 33824 7754
rect 33784 6996 33836 7002
rect 33784 6938 33836 6944
rect 33784 6792 33836 6798
rect 33888 6780 33916 7754
rect 33980 7546 34008 12679
rect 34242 12200 34298 13000
rect 34428 12436 34480 12442
rect 34428 12378 34480 12384
rect 34440 12209 34468 12378
rect 34426 12200 34482 12209
rect 34610 12200 34666 13000
rect 34978 12200 35034 13000
rect 35346 12200 35402 13000
rect 35622 12880 35678 12889
rect 35622 12815 35678 12824
rect 35636 12442 35664 12815
rect 35624 12436 35676 12442
rect 35624 12378 35676 12384
rect 35714 12200 35770 13000
rect 35900 12912 35952 12918
rect 35898 12880 35900 12889
rect 35992 12912 36044 12918
rect 35952 12880 35954 12889
rect 35992 12854 36044 12860
rect 35898 12815 35954 12824
rect 34060 12164 34112 12170
rect 34060 12106 34112 12112
rect 34072 11354 34100 12106
rect 34256 11694 34284 12200
rect 34426 12135 34482 12144
rect 34244 11688 34296 11694
rect 34244 11630 34296 11636
rect 34060 11348 34112 11354
rect 34060 11290 34112 11296
rect 34624 11234 34652 12200
rect 34992 11354 35020 12200
rect 35256 11756 35308 11762
rect 35256 11698 35308 11704
rect 34980 11348 35032 11354
rect 34980 11290 35032 11296
rect 34624 11206 34928 11234
rect 34612 11076 34664 11082
rect 34612 11018 34664 11024
rect 34336 10192 34388 10198
rect 34336 10134 34388 10140
rect 34520 10192 34572 10198
rect 34520 10134 34572 10140
rect 34348 9178 34376 10134
rect 34428 9648 34480 9654
rect 34428 9590 34480 9596
rect 34440 9382 34468 9590
rect 34428 9376 34480 9382
rect 34428 9318 34480 9324
rect 34336 9172 34388 9178
rect 34336 9114 34388 9120
rect 34152 9036 34204 9042
rect 34152 8978 34204 8984
rect 34164 8566 34192 8978
rect 34428 8628 34480 8634
rect 34428 8570 34480 8576
rect 34152 8560 34204 8566
rect 34152 8502 34204 8508
rect 34440 8498 34468 8570
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34336 8424 34388 8430
rect 34336 8366 34388 8372
rect 33968 7540 34020 7546
rect 33968 7482 34020 7488
rect 34152 7472 34204 7478
rect 34152 7414 34204 7420
rect 34244 7472 34296 7478
rect 34244 7414 34296 7420
rect 33968 7200 34020 7206
rect 33968 7142 34020 7148
rect 33980 6798 34008 7142
rect 33836 6752 33916 6780
rect 33968 6792 34020 6798
rect 33784 6734 33836 6740
rect 33968 6734 34020 6740
rect 33692 6248 33744 6254
rect 33692 6190 33744 6196
rect 33704 5914 33732 6190
rect 33692 5908 33744 5914
rect 33692 5850 33744 5856
rect 34164 5710 34192 7414
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 34256 5642 34284 7414
rect 34244 5636 34296 5642
rect 34244 5578 34296 5584
rect 34348 5250 34376 8366
rect 34428 7812 34480 7818
rect 34428 7754 34480 7760
rect 34440 7342 34468 7754
rect 34428 7336 34480 7342
rect 34428 7278 34480 7284
rect 34072 5222 34376 5250
rect 34428 5296 34480 5302
rect 34428 5238 34480 5244
rect 34072 5166 34100 5222
rect 34060 5160 34112 5166
rect 34060 5102 34112 5108
rect 34440 4706 34468 5238
rect 34532 4758 34560 10134
rect 34624 9654 34652 11018
rect 34612 9648 34664 9654
rect 34612 9590 34664 9596
rect 34900 9568 34928 11206
rect 35164 10668 35216 10674
rect 35164 10610 35216 10616
rect 35072 10464 35124 10470
rect 35072 10406 35124 10412
rect 35084 10062 35112 10406
rect 35176 10305 35204 10610
rect 35162 10296 35218 10305
rect 35162 10231 35164 10240
rect 35216 10231 35218 10240
rect 35164 10202 35216 10208
rect 35176 10171 35204 10202
rect 35072 10056 35124 10062
rect 35072 9998 35124 10004
rect 34980 9580 35032 9586
rect 34900 9540 34980 9568
rect 34980 9522 35032 9528
rect 34612 9512 34664 9518
rect 34612 9454 34664 9460
rect 34624 9110 34652 9454
rect 34612 9104 34664 9110
rect 34612 9046 34664 9052
rect 35084 9042 35112 9998
rect 34888 9036 34940 9042
rect 34888 8978 34940 8984
rect 35072 9036 35124 9042
rect 35072 8978 35124 8984
rect 34900 8838 34928 8978
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34888 8832 34940 8838
rect 34888 8774 34940 8780
rect 34808 8498 34836 8774
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 34888 8492 34940 8498
rect 34888 8434 34940 8440
rect 34808 8090 34836 8434
rect 34612 8084 34664 8090
rect 34612 8026 34664 8032
rect 34796 8084 34848 8090
rect 34796 8026 34848 8032
rect 34624 7546 34652 8026
rect 34612 7540 34664 7546
rect 34612 7482 34664 7488
rect 34796 7336 34848 7342
rect 34796 7278 34848 7284
rect 34612 7200 34664 7206
rect 34612 7142 34664 7148
rect 34256 4678 34468 4706
rect 34520 4752 34572 4758
rect 34520 4694 34572 4700
rect 34256 4570 34284 4678
rect 33980 4542 34284 4570
rect 34428 4616 34480 4622
rect 34428 4558 34480 4564
rect 33980 4486 34008 4542
rect 33968 4480 34020 4486
rect 33968 4422 34020 4428
rect 34060 4480 34112 4486
rect 34060 4422 34112 4428
rect 32680 4140 32732 4146
rect 32680 4082 32732 4088
rect 33232 4140 33284 4146
rect 33232 4082 33284 4088
rect 32494 3904 32550 3913
rect 32494 3839 32550 3848
rect 32508 3670 32536 3839
rect 32692 3670 32720 4082
rect 32496 3664 32548 3670
rect 32496 3606 32548 3612
rect 32680 3664 32732 3670
rect 32680 3606 32732 3612
rect 32956 3664 33008 3670
rect 32956 3606 33008 3612
rect 32588 2984 32640 2990
rect 32588 2926 32640 2932
rect 32496 2032 32548 2038
rect 32496 1974 32548 1980
rect 32508 1426 32536 1974
rect 32496 1420 32548 1426
rect 32496 1362 32548 1368
rect 32600 800 32628 2926
rect 32680 2440 32732 2446
rect 32680 2382 32732 2388
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 32692 2038 32720 2382
rect 32680 2032 32732 2038
rect 32680 1974 32732 1980
rect 32784 1562 32812 2382
rect 32772 1556 32824 1562
rect 32772 1498 32824 1504
rect 32770 1320 32826 1329
rect 32770 1255 32826 1264
rect 31942 776 31998 785
rect 31942 711 31998 720
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32784 474 32812 1255
rect 32968 800 32996 3606
rect 33244 3194 33272 4082
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 33324 3188 33376 3194
rect 33324 3130 33376 3136
rect 33140 1284 33192 1290
rect 33140 1226 33192 1232
rect 32862 504 32918 513
rect 32772 468 32824 474
rect 32862 439 32864 448
rect 32772 410 32824 416
rect 32916 439 32918 448
rect 32864 410 32916 416
rect 32954 0 33010 800
rect 33152 513 33180 1226
rect 33336 800 33364 3130
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 33600 1896 33652 1902
rect 33600 1838 33652 1844
rect 33508 1828 33560 1834
rect 33508 1770 33560 1776
rect 33416 1556 33468 1562
rect 33416 1498 33468 1504
rect 33428 882 33456 1498
rect 33520 1494 33548 1770
rect 33508 1488 33560 1494
rect 33508 1430 33560 1436
rect 33612 1358 33640 1838
rect 33600 1352 33652 1358
rect 33600 1294 33652 1300
rect 33416 876 33468 882
rect 33416 818 33468 824
rect 33704 800 33732 2994
rect 33876 1488 33928 1494
rect 33876 1430 33928 1436
rect 33888 882 33916 1430
rect 33876 876 33928 882
rect 33876 818 33928 824
rect 34072 800 34100 4422
rect 34336 1488 34388 1494
rect 34336 1430 34388 1436
rect 33138 504 33194 513
rect 33138 439 33194 448
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34348 66 34376 1430
rect 34440 800 34468 4558
rect 34624 3398 34652 7142
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 34716 6322 34744 6734
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 34808 5642 34836 7278
rect 34796 5636 34848 5642
rect 34796 5578 34848 5584
rect 34900 5234 34928 8434
rect 35164 7744 35216 7750
rect 35164 7686 35216 7692
rect 35176 6882 35204 7686
rect 35268 7342 35296 11698
rect 35360 11642 35388 12200
rect 35360 11614 35664 11642
rect 35636 11558 35664 11614
rect 35532 11552 35584 11558
rect 35532 11494 35584 11500
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35544 11218 35572 11494
rect 35532 11212 35584 11218
rect 35532 11154 35584 11160
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 35360 9926 35388 10610
rect 35624 10600 35676 10606
rect 35624 10542 35676 10548
rect 35636 10470 35664 10542
rect 35624 10464 35676 10470
rect 35624 10406 35676 10412
rect 35440 10192 35492 10198
rect 35440 10134 35492 10140
rect 35348 9920 35400 9926
rect 35348 9862 35400 9868
rect 35256 7336 35308 7342
rect 35256 7278 35308 7284
rect 35084 6854 35204 6882
rect 35452 6866 35480 10134
rect 35728 9654 35756 12200
rect 36004 11937 36032 12854
rect 36082 12200 36138 13000
rect 36450 12200 36506 13000
rect 36726 12472 36782 12481
rect 36726 12407 36782 12416
rect 35990 11928 36046 11937
rect 35990 11863 36046 11872
rect 36096 11132 36124 12200
rect 36266 11928 36322 11937
rect 36266 11863 36322 11872
rect 36176 11144 36228 11150
rect 36096 11104 36176 11132
rect 36176 11086 36228 11092
rect 36084 10600 36136 10606
rect 36084 10542 36136 10548
rect 36096 9926 36124 10542
rect 36084 9920 36136 9926
rect 36084 9862 36136 9868
rect 35624 9648 35676 9654
rect 35624 9590 35676 9596
rect 35716 9648 35768 9654
rect 35716 9590 35768 9596
rect 35532 9512 35584 9518
rect 35532 9454 35584 9460
rect 35636 9466 35664 9590
rect 36280 9466 36308 11863
rect 36358 11520 36414 11529
rect 36358 11455 36414 11464
rect 36372 10606 36400 11455
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 35544 8498 35572 9454
rect 35636 9438 36308 9466
rect 36266 9072 36322 9081
rect 36266 9007 36322 9016
rect 35532 8492 35584 8498
rect 35532 8434 35584 8440
rect 35544 8090 35572 8434
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35900 8084 35952 8090
rect 35900 8026 35952 8032
rect 35532 7880 35584 7886
rect 35532 7822 35584 7828
rect 35544 6866 35572 7822
rect 35912 7410 35940 8026
rect 36280 7750 36308 9007
rect 36464 8974 36492 12200
rect 36634 11520 36690 11529
rect 36634 11455 36690 11464
rect 36542 9072 36598 9081
rect 36648 9042 36676 11455
rect 36740 11218 36768 12407
rect 36818 12200 36874 13000
rect 37186 12200 37242 13000
rect 37554 12200 37610 13000
rect 37922 12200 37978 13000
rect 38016 12572 38068 12578
rect 38016 12514 38068 12520
rect 36728 11212 36780 11218
rect 36728 11154 36780 11160
rect 36832 10266 36860 12200
rect 37200 12102 37228 12200
rect 37096 12096 37148 12102
rect 37096 12038 37148 12044
rect 37188 12096 37240 12102
rect 37188 12038 37240 12044
rect 37004 11688 37056 11694
rect 37004 11630 37056 11636
rect 37016 11218 37044 11630
rect 37108 11218 37136 12038
rect 37188 11824 37240 11830
rect 37188 11766 37240 11772
rect 37568 11778 37596 12200
rect 37200 11694 37228 11766
rect 37568 11750 37688 11778
rect 37660 11694 37688 11750
rect 37188 11688 37240 11694
rect 37188 11630 37240 11636
rect 37648 11688 37700 11694
rect 37648 11630 37700 11636
rect 37740 11280 37792 11286
rect 37740 11222 37792 11228
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 37096 11212 37148 11218
rect 37096 11154 37148 11160
rect 37648 11144 37700 11150
rect 37648 11086 37700 11092
rect 37660 11014 37688 11086
rect 37556 11008 37608 11014
rect 37556 10950 37608 10956
rect 37648 11008 37700 11014
rect 37648 10950 37700 10956
rect 37568 10674 37596 10950
rect 37464 10668 37516 10674
rect 37464 10610 37516 10616
rect 37556 10668 37608 10674
rect 37556 10610 37608 10616
rect 37004 10600 37056 10606
rect 37056 10548 37228 10554
rect 37004 10542 37228 10548
rect 37016 10526 37228 10542
rect 36820 10260 36872 10266
rect 36820 10202 36872 10208
rect 37096 10124 37148 10130
rect 37096 10066 37148 10072
rect 37108 9926 37136 10066
rect 37004 9920 37056 9926
rect 37004 9862 37056 9868
rect 37096 9920 37148 9926
rect 37096 9862 37148 9868
rect 36820 9580 36872 9586
rect 36820 9522 36872 9528
rect 36912 9580 36964 9586
rect 36912 9522 36964 9528
rect 36832 9042 36860 9522
rect 36542 9007 36598 9016
rect 36636 9036 36688 9042
rect 36452 8968 36504 8974
rect 36452 8910 36504 8916
rect 36556 8401 36584 9007
rect 36636 8978 36688 8984
rect 36820 9036 36872 9042
rect 36820 8978 36872 8984
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36542 8392 36598 8401
rect 36542 8327 36598 8336
rect 36740 7886 36768 8434
rect 36832 8401 36860 8978
rect 36924 8566 36952 9522
rect 37016 9042 37044 9862
rect 37004 9036 37056 9042
rect 37004 8978 37056 8984
rect 37200 8650 37228 10526
rect 37476 10169 37504 10610
rect 37648 10600 37700 10606
rect 37648 10542 37700 10548
rect 37278 10160 37334 10169
rect 37278 10095 37334 10104
rect 37462 10160 37518 10169
rect 37660 10130 37688 10542
rect 37752 10130 37780 11222
rect 37462 10095 37464 10104
rect 37292 9042 37320 10095
rect 37516 10095 37518 10104
rect 37648 10124 37700 10130
rect 37464 10066 37516 10072
rect 37648 10066 37700 10072
rect 37740 10124 37792 10130
rect 37740 10066 37792 10072
rect 37936 9382 37964 12200
rect 38028 11218 38056 12514
rect 38290 12200 38346 13000
rect 38384 12300 38436 12306
rect 38384 12242 38436 12248
rect 38568 12300 38620 12306
rect 38568 12242 38620 12248
rect 38016 11212 38068 11218
rect 38016 11154 38068 11160
rect 38304 10996 38332 12200
rect 38120 10968 38332 10996
rect 37924 9376 37976 9382
rect 37924 9318 37976 9324
rect 38120 9110 38148 10968
rect 38396 10554 38424 12242
rect 38580 11762 38608 12242
rect 38658 12200 38714 13000
rect 38936 12572 38988 12578
rect 38936 12514 38988 12520
rect 38568 11756 38620 11762
rect 38568 11698 38620 11704
rect 38672 11098 38700 12200
rect 38672 11070 38884 11098
rect 38948 11082 38976 12514
rect 39026 12200 39082 13000
rect 39394 12200 39450 13000
rect 39762 12200 39818 13000
rect 40130 12200 40186 13000
rect 40406 12880 40462 12889
rect 40406 12815 40462 12824
rect 40420 12782 40448 12815
rect 40408 12776 40460 12782
rect 40408 12718 40460 12724
rect 40406 12336 40462 12345
rect 40406 12271 40462 12280
rect 40314 12200 40370 12209
rect 38752 11008 38804 11014
rect 38752 10950 38804 10956
rect 38396 10538 38700 10554
rect 38396 10532 38712 10538
rect 38396 10526 38660 10532
rect 38660 10474 38712 10480
rect 38764 10282 38792 10950
rect 38672 10254 38792 10282
rect 38476 9580 38528 9586
rect 38672 9568 38700 10254
rect 38856 10248 38884 11070
rect 38936 11076 38988 11082
rect 38936 11018 38988 11024
rect 38856 10220 38976 10248
rect 38844 10124 38896 10130
rect 38844 10066 38896 10072
rect 38856 9874 38884 10066
rect 38528 9540 38700 9568
rect 38764 9846 38884 9874
rect 38476 9522 38528 9528
rect 38566 9344 38622 9353
rect 38566 9279 38622 9288
rect 38292 9172 38344 9178
rect 38292 9114 38344 9120
rect 38108 9104 38160 9110
rect 38108 9046 38160 9052
rect 37280 9036 37332 9042
rect 37280 8978 37332 8984
rect 37200 8622 37504 8650
rect 36912 8560 36964 8566
rect 36912 8502 36964 8508
rect 37188 8424 37240 8430
rect 36818 8392 36874 8401
rect 37188 8366 37240 8372
rect 36818 8327 36874 8336
rect 37200 7970 37228 8366
rect 37200 7942 37412 7970
rect 36728 7880 36780 7886
rect 37188 7880 37240 7886
rect 36728 7822 36780 7828
rect 36832 7840 37188 7868
rect 36268 7744 36320 7750
rect 36268 7686 36320 7692
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 36268 7404 36320 7410
rect 36268 7346 36320 7352
rect 35440 6860 35492 6866
rect 35084 6848 35112 6854
rect 34992 6820 35112 6848
rect 34992 5778 35020 6820
rect 35440 6802 35492 6808
rect 35532 6860 35584 6866
rect 35532 6802 35584 6808
rect 36280 6798 36308 7346
rect 36832 7324 36860 7840
rect 37188 7822 37240 7828
rect 37188 7404 37240 7410
rect 37188 7346 37240 7352
rect 36372 7296 36860 7324
rect 36372 7206 36400 7296
rect 37004 7268 37056 7274
rect 36464 7228 36952 7256
rect 36360 7200 36412 7206
rect 36360 7142 36412 7148
rect 36464 7002 36492 7228
rect 36924 7002 36952 7228
rect 37004 7210 37056 7216
rect 36452 6996 36504 7002
rect 36452 6938 36504 6944
rect 36912 6996 36964 7002
rect 36912 6938 36964 6944
rect 36360 6860 36412 6866
rect 36360 6802 36412 6808
rect 36464 6854 36676 6882
rect 36084 6792 36136 6798
rect 36084 6734 36136 6740
rect 36268 6792 36320 6798
rect 36268 6734 36320 6740
rect 35440 6656 35492 6662
rect 35440 6598 35492 6604
rect 35072 6316 35124 6322
rect 35072 6258 35124 6264
rect 35084 5846 35112 6258
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 35072 5840 35124 5846
rect 35072 5782 35124 5788
rect 35256 5840 35308 5846
rect 35256 5782 35308 5788
rect 34980 5772 35032 5778
rect 34980 5714 35032 5720
rect 34888 5228 34940 5234
rect 34888 5170 34940 5176
rect 34980 5228 35032 5234
rect 34980 5170 35032 5176
rect 34900 4758 34928 5170
rect 34888 4752 34940 4758
rect 34888 4694 34940 4700
rect 34992 4282 35020 5170
rect 35072 5024 35124 5030
rect 35072 4966 35124 4972
rect 34980 4276 35032 4282
rect 34980 4218 35032 4224
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 34716 2854 34744 3334
rect 34704 2848 34756 2854
rect 34704 2790 34756 2796
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 34704 876 34756 882
rect 34704 818 34756 824
rect 34336 60 34388 66
rect 34336 2 34388 8
rect 34426 0 34482 800
rect 34716 746 34744 818
rect 34808 800 34836 2790
rect 35084 2650 35112 4966
rect 35162 4856 35218 4865
rect 35162 4791 35218 4800
rect 35176 4758 35204 4791
rect 35164 4752 35216 4758
rect 35164 4694 35216 4700
rect 35164 4276 35216 4282
rect 35164 4218 35216 4224
rect 35176 3913 35204 4218
rect 35162 3904 35218 3913
rect 35162 3839 35218 3848
rect 35072 2644 35124 2650
rect 35072 2586 35124 2592
rect 35268 2446 35296 5782
rect 35360 5778 35388 5850
rect 35348 5772 35400 5778
rect 35348 5714 35400 5720
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 35360 2310 35388 2586
rect 35348 2304 35400 2310
rect 35452 2292 35480 6598
rect 36096 6322 36124 6734
rect 36280 6458 36308 6734
rect 36176 6452 36228 6458
rect 36176 6394 36228 6400
rect 36268 6452 36320 6458
rect 36268 6394 36320 6400
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 36004 6100 36032 6258
rect 36188 6118 36216 6394
rect 36084 6112 36136 6118
rect 36004 6072 36084 6100
rect 36084 6054 36136 6060
rect 36176 6112 36228 6118
rect 36176 6054 36228 6060
rect 36096 5914 36124 6054
rect 36084 5908 36136 5914
rect 36084 5850 36136 5856
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 35900 5636 35952 5642
rect 35900 5578 35952 5584
rect 35714 3904 35770 3913
rect 35714 3839 35770 3848
rect 35624 2848 35676 2854
rect 35624 2790 35676 2796
rect 35532 2440 35584 2446
rect 35530 2408 35532 2417
rect 35584 2408 35586 2417
rect 35530 2343 35586 2352
rect 35636 2310 35664 2790
rect 35728 2514 35756 3839
rect 35912 3602 35940 5578
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 35820 3482 35848 3538
rect 35820 3454 36124 3482
rect 35806 2952 35862 2961
rect 35806 2887 35862 2896
rect 35990 2952 36046 2961
rect 35990 2887 36046 2896
rect 35820 2514 35848 2887
rect 35898 2680 35954 2689
rect 35898 2615 35954 2624
rect 35716 2508 35768 2514
rect 35716 2450 35768 2456
rect 35808 2508 35860 2514
rect 35808 2450 35860 2456
rect 35912 2417 35940 2615
rect 35898 2408 35954 2417
rect 35898 2343 35954 2352
rect 35624 2304 35676 2310
rect 35452 2264 35572 2292
rect 35348 2246 35400 2252
rect 35348 1896 35400 1902
rect 35348 1838 35400 1844
rect 35360 1358 35388 1838
rect 35348 1352 35400 1358
rect 35348 1294 35400 1300
rect 35440 1352 35492 1358
rect 35440 1294 35492 1300
rect 34888 1284 34940 1290
rect 34888 1226 34940 1232
rect 35072 1284 35124 1290
rect 35072 1226 35124 1232
rect 34704 740 34756 746
rect 34704 682 34756 688
rect 34518 504 34574 513
rect 34518 439 34574 448
rect 34532 66 34560 439
rect 34520 60 34572 66
rect 34520 2 34572 8
rect 34794 0 34850 800
rect 34900 746 34928 1226
rect 35084 950 35112 1226
rect 35072 944 35124 950
rect 35072 886 35124 892
rect 35452 882 35480 1294
rect 35440 876 35492 882
rect 35176 836 35296 864
rect 35176 800 35204 836
rect 34888 740 34940 746
rect 34888 682 34940 688
rect 35162 0 35218 800
rect 35268 513 35296 836
rect 35440 818 35492 824
rect 35544 800 35572 2264
rect 35624 2246 35676 2252
rect 36004 1442 36032 2887
rect 36096 2689 36124 3454
rect 36082 2680 36138 2689
rect 36082 2615 36138 2624
rect 36280 2446 36308 5646
rect 36372 5250 36400 6802
rect 36464 5574 36492 6854
rect 36648 6848 36676 6854
rect 36728 6860 36780 6866
rect 36648 6820 36728 6848
rect 37016 6848 37044 7210
rect 37200 7206 37228 7346
rect 37280 7336 37332 7342
rect 37280 7278 37332 7284
rect 37188 7200 37240 7206
rect 37188 7142 37240 7148
rect 36728 6802 36780 6808
rect 36924 6820 37044 6848
rect 36924 6730 36952 6820
rect 37292 6798 37320 7278
rect 37280 6792 37332 6798
rect 37108 6752 37280 6780
rect 36636 6724 36688 6730
rect 36636 6666 36688 6672
rect 36912 6724 36964 6730
rect 36912 6666 36964 6672
rect 37004 6724 37056 6730
rect 37004 6666 37056 6672
rect 36648 6610 36676 6666
rect 37016 6610 37044 6666
rect 36648 6582 37044 6610
rect 36636 6452 36688 6458
rect 36636 6394 36688 6400
rect 36648 5778 36676 6394
rect 37108 5778 37136 6752
rect 37280 6734 37332 6740
rect 37280 6316 37332 6322
rect 37280 6258 37332 6264
rect 37292 5778 37320 6258
rect 36636 5772 36688 5778
rect 36636 5714 36688 5720
rect 37096 5772 37148 5778
rect 37096 5714 37148 5720
rect 37280 5772 37332 5778
rect 37280 5714 37332 5720
rect 36452 5568 36504 5574
rect 36452 5510 36504 5516
rect 36372 5222 37044 5250
rect 36464 5086 36676 5114
rect 36464 5030 36492 5086
rect 36452 5024 36504 5030
rect 36452 4966 36504 4972
rect 36544 5024 36596 5030
rect 36544 4966 36596 4972
rect 36358 4856 36414 4865
rect 36556 4826 36584 4966
rect 36648 4842 36676 5086
rect 37016 5001 37044 5222
rect 37002 4992 37058 5001
rect 37002 4927 37058 4936
rect 36358 4791 36414 4800
rect 36544 4820 36596 4826
rect 36372 4321 36400 4791
rect 36648 4814 36952 4842
rect 36544 4762 36596 4768
rect 36452 4752 36504 4758
rect 36820 4752 36872 4758
rect 36504 4700 36768 4706
rect 36452 4694 36768 4700
rect 36820 4694 36872 4700
rect 36464 4678 36768 4694
rect 36740 4554 36768 4678
rect 36832 4622 36860 4694
rect 36924 4622 36952 4814
rect 37004 4752 37056 4758
rect 37004 4694 37056 4700
rect 36820 4616 36872 4622
rect 36820 4558 36872 4564
rect 36912 4616 36964 4622
rect 36912 4558 36964 4564
rect 36636 4548 36688 4554
rect 36636 4490 36688 4496
rect 36728 4548 36780 4554
rect 36728 4490 36780 4496
rect 36648 4434 36676 4490
rect 36648 4406 36860 4434
rect 36358 4312 36414 4321
rect 36636 4276 36688 4282
rect 36358 4247 36414 4256
rect 36464 4236 36636 4264
rect 36360 4208 36412 4214
rect 36464 4162 36492 4236
rect 36636 4218 36688 4224
rect 36832 4214 36860 4406
rect 36412 4156 36492 4162
rect 36360 4150 36492 4156
rect 36728 4208 36780 4214
rect 36728 4150 36780 4156
rect 36820 4208 36872 4214
rect 36820 4150 36872 4156
rect 36372 4134 36492 4150
rect 36634 4040 36690 4049
rect 36372 3998 36634 4026
rect 36372 3913 36400 3998
rect 36740 4026 36768 4150
rect 37016 4026 37044 4694
rect 37384 4604 37412 7942
rect 37476 7750 37504 8622
rect 38304 8498 38332 9114
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 37464 7744 37516 7750
rect 37464 7686 37516 7692
rect 38476 7404 38528 7410
rect 38476 7346 38528 7352
rect 37464 7336 37516 7342
rect 37464 7278 37516 7284
rect 37476 6390 37504 7278
rect 38488 7002 38516 7346
rect 38580 7206 38608 9279
rect 38764 9081 38792 9846
rect 38948 9704 38976 10220
rect 38856 9676 38976 9704
rect 38856 9178 38884 9676
rect 39040 9466 39068 12200
rect 39212 11756 39264 11762
rect 39212 11698 39264 11704
rect 39120 10056 39172 10062
rect 39120 9998 39172 10004
rect 39132 9654 39160 9998
rect 39224 9926 39252 11698
rect 39408 11014 39436 12200
rect 39776 12152 39804 12200
rect 39684 12124 39804 12152
rect 39580 12096 39632 12102
rect 39684 12073 39712 12124
rect 39580 12038 39632 12044
rect 39670 12064 39726 12073
rect 39592 11336 39620 12038
rect 39670 11999 39726 12008
rect 39854 12064 39910 12073
rect 39854 11999 39910 12008
rect 39868 11762 39896 11999
rect 39856 11756 39908 11762
rect 39856 11698 39908 11704
rect 39764 11348 39816 11354
rect 39592 11308 39764 11336
rect 39764 11290 39816 11296
rect 39396 11008 39448 11014
rect 39396 10950 39448 10956
rect 40144 10282 40172 12200
rect 40314 12135 40370 12144
rect 40420 12152 40448 12271
rect 40498 12200 40554 13000
rect 40590 12880 40646 12889
rect 40590 12815 40646 12824
rect 40512 12152 40540 12200
rect 40144 10254 40264 10282
rect 40130 10160 40186 10169
rect 40130 10095 40186 10104
rect 39212 9920 39264 9926
rect 39212 9862 39264 9868
rect 40040 9920 40092 9926
rect 40040 9862 40092 9868
rect 39120 9648 39172 9654
rect 39120 9590 39172 9596
rect 39212 9580 39264 9586
rect 39212 9522 39264 9528
rect 39304 9580 39356 9586
rect 39304 9522 39356 9528
rect 38948 9438 39068 9466
rect 38844 9172 38896 9178
rect 38844 9114 38896 9120
rect 38750 9072 38806 9081
rect 38750 9007 38806 9016
rect 38948 8838 38976 9438
rect 39028 9376 39080 9382
rect 39224 9353 39252 9522
rect 39028 9318 39080 9324
rect 39210 9344 39266 9353
rect 39040 9081 39068 9318
rect 39210 9279 39266 9288
rect 39224 9178 39252 9279
rect 39212 9172 39264 9178
rect 39212 9114 39264 9120
rect 39026 9072 39082 9081
rect 39026 9007 39082 9016
rect 39040 8974 39068 9007
rect 39028 8968 39080 8974
rect 39028 8910 39080 8916
rect 38936 8832 38988 8838
rect 38936 8774 38988 8780
rect 39212 8424 39264 8430
rect 39212 8366 39264 8372
rect 39224 8090 39252 8366
rect 39212 8084 39264 8090
rect 39212 8026 39264 8032
rect 38936 7948 38988 7954
rect 38856 7908 38936 7936
rect 38752 7880 38804 7886
rect 38856 7834 38884 7908
rect 38936 7890 38988 7896
rect 38804 7828 38884 7834
rect 38752 7822 38884 7828
rect 38764 7806 38884 7822
rect 39316 7342 39344 9522
rect 39946 9480 40002 9489
rect 39946 9415 40002 9424
rect 39580 9172 39632 9178
rect 39580 9114 39632 9120
rect 39396 8492 39448 8498
rect 39396 8434 39448 8440
rect 39408 8090 39436 8434
rect 39396 8084 39448 8090
rect 39396 8026 39448 8032
rect 39592 7750 39620 9114
rect 39960 9110 39988 9415
rect 39856 9104 39908 9110
rect 39856 9046 39908 9052
rect 39948 9104 40000 9110
rect 39948 9046 40000 9052
rect 39868 8786 39896 9046
rect 39868 8758 39988 8786
rect 39856 8492 39908 8498
rect 39856 8434 39908 8440
rect 39868 8378 39896 8434
rect 39776 8362 39896 8378
rect 39764 8356 39896 8362
rect 39816 8350 39896 8356
rect 39764 8298 39816 8304
rect 39672 7948 39724 7954
rect 39672 7890 39724 7896
rect 39764 7948 39816 7954
rect 39764 7890 39816 7896
rect 39580 7744 39632 7750
rect 39580 7686 39632 7692
rect 39684 7478 39712 7890
rect 39672 7472 39724 7478
rect 39672 7414 39724 7420
rect 39488 7404 39540 7410
rect 39488 7346 39540 7352
rect 38660 7336 38712 7342
rect 38660 7278 38712 7284
rect 39304 7336 39356 7342
rect 39304 7278 39356 7284
rect 39396 7336 39448 7342
rect 39396 7278 39448 7284
rect 38568 7200 38620 7206
rect 38568 7142 38620 7148
rect 38292 6996 38344 7002
rect 38292 6938 38344 6944
rect 38476 6996 38528 7002
rect 38476 6938 38528 6944
rect 38304 6882 38332 6938
rect 38672 6882 38700 7278
rect 39408 7002 39436 7278
rect 39500 7002 39528 7346
rect 38844 6996 38896 7002
rect 38844 6938 38896 6944
rect 39396 6996 39448 7002
rect 39396 6938 39448 6944
rect 39488 6996 39540 7002
rect 39488 6938 39540 6944
rect 38304 6854 38700 6882
rect 38016 6792 38068 6798
rect 38016 6734 38068 6740
rect 38028 6662 38056 6734
rect 38856 6662 38884 6938
rect 39776 6882 39804 7890
rect 39960 7274 39988 8758
rect 40052 8362 40080 9862
rect 40144 9489 40172 10095
rect 40236 9586 40264 10254
rect 40328 10169 40356 12135
rect 40420 12124 40540 12152
rect 40604 11082 40632 12815
rect 40774 12744 40830 12753
rect 40774 12679 40830 12688
rect 40682 12608 40738 12617
rect 40682 12543 40738 12552
rect 40696 12345 40724 12543
rect 40682 12336 40738 12345
rect 40682 12271 40738 12280
rect 40788 12152 40816 12679
rect 40866 12200 40922 13000
rect 50894 13016 50950 13025
rect 41142 12951 41198 12960
rect 40958 12608 41014 12617
rect 40958 12543 40960 12552
rect 41012 12543 41014 12552
rect 41052 12572 41104 12578
rect 40960 12514 41012 12520
rect 41052 12514 41104 12520
rect 40880 12152 40908 12200
rect 40788 12124 40908 12152
rect 40682 12064 40738 12073
rect 40682 11999 40738 12008
rect 40592 11076 40644 11082
rect 40592 11018 40644 11024
rect 40314 10160 40370 10169
rect 40314 10095 40370 10104
rect 40408 9920 40460 9926
rect 40408 9862 40460 9868
rect 40224 9580 40276 9586
rect 40224 9522 40276 9528
rect 40130 9480 40186 9489
rect 40130 9415 40186 9424
rect 40224 9376 40276 9382
rect 40224 9318 40276 9324
rect 40316 9376 40368 9382
rect 40316 9318 40368 9324
rect 40132 9036 40184 9042
rect 40132 8978 40184 8984
rect 40040 8356 40092 8362
rect 40040 8298 40092 8304
rect 40040 8084 40092 8090
rect 40040 8026 40092 8032
rect 39948 7268 40000 7274
rect 39948 7210 40000 7216
rect 39592 6854 39804 6882
rect 38016 6656 38068 6662
rect 38016 6598 38068 6604
rect 38844 6656 38896 6662
rect 38844 6598 38896 6604
rect 38936 6656 38988 6662
rect 38936 6598 38988 6604
rect 37464 6384 37516 6390
rect 37464 6326 37516 6332
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 37844 5778 37872 6258
rect 38028 5914 38056 6598
rect 38948 6322 38976 6598
rect 39592 6458 39620 6854
rect 39764 6792 39816 6798
rect 39764 6734 39816 6740
rect 39948 6792 40000 6798
rect 39948 6734 40000 6740
rect 39776 6458 39804 6734
rect 39580 6452 39632 6458
rect 39580 6394 39632 6400
rect 39764 6452 39816 6458
rect 39764 6394 39816 6400
rect 39856 6452 39908 6458
rect 39856 6394 39908 6400
rect 38936 6316 38988 6322
rect 38936 6258 38988 6264
rect 39488 6248 39540 6254
rect 39040 6208 39488 6236
rect 37924 5908 37976 5914
rect 37924 5850 37976 5856
rect 38016 5908 38068 5914
rect 38016 5850 38068 5856
rect 37936 5778 37964 5850
rect 37832 5772 37884 5778
rect 37832 5714 37884 5720
rect 37924 5772 37976 5778
rect 37924 5714 37976 5720
rect 38200 5568 38252 5574
rect 38200 5510 38252 5516
rect 37384 4576 37504 4604
rect 36740 3998 37044 4026
rect 36634 3975 36690 3984
rect 36358 3904 36414 3913
rect 36358 3839 36414 3848
rect 36360 3596 36412 3602
rect 36360 3538 36412 3544
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 36372 2990 36400 3538
rect 36544 3120 36596 3126
rect 36544 3062 36596 3068
rect 37004 3120 37056 3126
rect 37004 3062 37056 3068
rect 36360 2984 36412 2990
rect 36360 2926 36412 2932
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 36372 2446 36400 2790
rect 36556 2666 36584 3062
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 36740 2854 36768 2994
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 36556 2638 36768 2666
rect 36268 2440 36320 2446
rect 36268 2382 36320 2388
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 36636 2440 36688 2446
rect 36636 2382 36688 2388
rect 36648 1970 36676 2382
rect 36740 1970 36768 2638
rect 37016 2514 37044 3062
rect 37004 2508 37056 2514
rect 37004 2450 37056 2456
rect 36636 1964 36688 1970
rect 36636 1906 36688 1912
rect 36728 1964 36780 1970
rect 36728 1906 36780 1912
rect 37004 1896 37056 1902
rect 37280 1896 37332 1902
rect 37004 1838 37056 1844
rect 37108 1856 37280 1884
rect 36452 1828 36504 1834
rect 36452 1770 36504 1776
rect 35820 1414 36032 1442
rect 36464 1426 36492 1770
rect 36820 1760 36872 1766
rect 36820 1702 36872 1708
rect 36452 1420 36504 1426
rect 35820 1034 35848 1414
rect 36452 1362 36504 1368
rect 36832 1358 36860 1702
rect 37016 1358 37044 1838
rect 37108 1766 37136 1856
rect 37280 1838 37332 1844
rect 37096 1760 37148 1766
rect 37096 1702 37148 1708
rect 35900 1352 35952 1358
rect 36820 1352 36872 1358
rect 35900 1294 35952 1300
rect 36542 1320 36598 1329
rect 35912 1170 35940 1294
rect 35992 1284 36044 1290
rect 36044 1244 36492 1272
rect 36820 1294 36872 1300
rect 37004 1352 37056 1358
rect 37004 1294 37056 1300
rect 36542 1255 36598 1264
rect 35992 1226 36044 1232
rect 35912 1142 36400 1170
rect 35716 1012 35768 1018
rect 35820 1006 35940 1034
rect 36372 1018 36400 1142
rect 36464 1018 36492 1244
rect 35716 954 35768 960
rect 35254 504 35310 513
rect 35254 439 35310 448
rect 35530 0 35586 800
rect 35728 762 35756 954
rect 35912 800 35940 1006
rect 36360 1012 36412 1018
rect 36360 954 36412 960
rect 36452 1012 36504 1018
rect 36452 954 36504 960
rect 36556 898 36584 1255
rect 36280 870 36584 898
rect 36280 800 36308 870
rect 36648 836 36768 864
rect 36648 800 36676 836
rect 35806 776 35862 785
rect 35728 734 35806 762
rect 35806 711 35862 720
rect 35806 640 35862 649
rect 35806 575 35862 584
rect 35820 66 35848 575
rect 35808 60 35860 66
rect 35808 2 35860 8
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36544 740 36596 746
rect 36544 682 36596 688
rect 36452 672 36504 678
rect 36452 614 36504 620
rect 36464 134 36492 614
rect 36556 134 36584 682
rect 36452 128 36504 134
rect 36452 70 36504 76
rect 36544 128 36596 134
rect 36544 70 36596 76
rect 36634 0 36690 800
rect 36740 134 36768 836
rect 37016 836 37136 864
rect 37016 800 37044 836
rect 36728 128 36780 134
rect 36728 70 36780 76
rect 37002 0 37058 800
rect 37108 513 37136 836
rect 37384 800 37412 3538
rect 37476 3534 37504 4576
rect 37464 3528 37516 3534
rect 38108 3528 38160 3534
rect 37464 3470 37516 3476
rect 37844 3488 38108 3516
rect 37844 3058 37872 3488
rect 38108 3470 38160 3476
rect 37832 3052 37884 3058
rect 37832 2994 37884 3000
rect 38016 2984 38068 2990
rect 38016 2926 38068 2932
rect 37462 2816 37518 2825
rect 37462 2751 37518 2760
rect 37476 950 37504 2751
rect 38028 2650 38056 2926
rect 38212 2854 38240 5510
rect 39040 5114 39068 6208
rect 39488 6190 39540 6196
rect 39868 5710 39896 6394
rect 39856 5704 39908 5710
rect 39856 5646 39908 5652
rect 38948 5086 39068 5114
rect 38948 4758 38976 5086
rect 39960 4978 39988 6734
rect 39040 4950 39988 4978
rect 38936 4752 38988 4758
rect 38936 4694 38988 4700
rect 39040 3516 39068 4950
rect 39212 4752 39264 4758
rect 40052 4706 40080 8026
rect 39212 4694 39264 4700
rect 38764 3488 39068 3516
rect 38764 2990 38792 3488
rect 39224 3448 39252 4694
rect 39856 4684 39908 4690
rect 39040 3420 39252 3448
rect 39316 4644 39856 4672
rect 39040 3210 39068 3420
rect 38948 3182 39068 3210
rect 38948 3074 38976 3182
rect 39316 3176 39344 4644
rect 39856 4626 39908 4632
rect 39960 4678 40080 4706
rect 39960 4298 39988 4678
rect 40040 4616 40092 4622
rect 40144 4604 40172 8978
rect 40236 4622 40264 9318
rect 40328 8838 40356 9318
rect 40316 8832 40368 8838
rect 40316 8774 40368 8780
rect 40316 6860 40368 6866
rect 40316 6802 40368 6808
rect 40328 5710 40356 6802
rect 40316 5704 40368 5710
rect 40316 5646 40368 5652
rect 40092 4576 40172 4604
rect 40224 4616 40276 4622
rect 40040 4558 40092 4564
rect 40224 4558 40276 4564
rect 39684 4270 39988 4298
rect 39684 4214 39712 4270
rect 39672 4208 39724 4214
rect 40040 4208 40092 4214
rect 39672 4150 39724 4156
rect 39776 4168 40040 4196
rect 39500 3318 39712 3346
rect 39500 3194 39528 3318
rect 39224 3148 39344 3176
rect 39488 3188 39540 3194
rect 38856 3046 38976 3074
rect 39028 3120 39080 3126
rect 39028 3062 39080 3068
rect 38752 2984 38804 2990
rect 38752 2926 38804 2932
rect 38200 2848 38252 2854
rect 38200 2790 38252 2796
rect 38292 2848 38344 2854
rect 38292 2790 38344 2796
rect 38474 2816 38530 2825
rect 38016 2644 38068 2650
rect 38016 2586 38068 2592
rect 38108 1760 38160 1766
rect 38108 1702 38160 1708
rect 37556 1352 37608 1358
rect 37556 1294 37608 1300
rect 37464 944 37516 950
rect 37464 886 37516 892
rect 37568 882 37596 1294
rect 37556 876 37608 882
rect 37832 876 37884 882
rect 37556 818 37608 824
rect 37752 836 37832 864
rect 37752 800 37780 836
rect 37832 818 37884 824
rect 38120 800 38148 1702
rect 38304 814 38332 2790
rect 38474 2751 38530 2760
rect 38384 2644 38436 2650
rect 38384 2586 38436 2592
rect 38396 1000 38424 2586
rect 38488 2038 38516 2751
rect 38752 2508 38804 2514
rect 38752 2450 38804 2456
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38476 2032 38528 2038
rect 38476 1974 38528 1980
rect 38568 2032 38620 2038
rect 38568 1974 38620 1980
rect 38580 1766 38608 1974
rect 38672 1766 38700 2382
rect 38568 1760 38620 1766
rect 38568 1702 38620 1708
rect 38660 1760 38712 1766
rect 38660 1702 38712 1708
rect 38764 1329 38792 2450
rect 38750 1320 38806 1329
rect 38750 1255 38806 1264
rect 38396 972 38516 1000
rect 38292 808 38344 814
rect 37094 504 37150 513
rect 37094 439 37150 448
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38488 800 38516 972
rect 38856 800 38884 3046
rect 39040 2990 39068 3062
rect 38936 2984 38988 2990
rect 38936 2926 38988 2932
rect 39028 2984 39080 2990
rect 39224 2961 39252 3148
rect 39488 3130 39540 3136
rect 39580 3188 39632 3194
rect 39580 3130 39632 3136
rect 39592 3074 39620 3130
rect 39500 3046 39620 3074
rect 39684 3058 39712 3318
rect 39672 3052 39724 3058
rect 39028 2926 39080 2932
rect 39210 2952 39266 2961
rect 38948 2446 38976 2926
rect 39394 2952 39450 2961
rect 39210 2887 39266 2896
rect 39316 2910 39394 2938
rect 39316 2530 39344 2910
rect 39394 2887 39450 2896
rect 39040 2502 39344 2530
rect 38936 2440 38988 2446
rect 38936 2382 38988 2388
rect 38948 882 38976 2382
rect 39040 1766 39068 2502
rect 39120 2440 39172 2446
rect 39120 2382 39172 2388
rect 39396 2440 39448 2446
rect 39500 2428 39528 3046
rect 39672 2994 39724 3000
rect 39580 2984 39632 2990
rect 39580 2926 39632 2932
rect 39592 2632 39620 2926
rect 39672 2644 39724 2650
rect 39592 2604 39672 2632
rect 39672 2586 39724 2592
rect 39448 2400 39528 2428
rect 39396 2382 39448 2388
rect 39028 1760 39080 1766
rect 39028 1702 39080 1708
rect 39132 1358 39160 2382
rect 39776 2292 39804 4168
rect 40040 4150 40092 4156
rect 39868 3998 40080 4026
rect 39868 3534 39896 3998
rect 40052 3942 40080 3998
rect 39948 3936 40000 3942
rect 39948 3878 40000 3884
rect 40040 3936 40092 3942
rect 40040 3878 40092 3884
rect 39960 3754 39988 3878
rect 39960 3726 40080 3754
rect 39856 3528 39908 3534
rect 39856 3470 39908 3476
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 39960 3126 39988 3470
rect 40052 3126 40080 3726
rect 40420 3448 40448 9862
rect 40592 9512 40644 9518
rect 40592 9454 40644 9460
rect 40500 9172 40552 9178
rect 40500 9114 40552 9120
rect 40512 6338 40540 9114
rect 40604 9042 40632 9454
rect 40592 9036 40644 9042
rect 40592 8978 40644 8984
rect 40592 8900 40644 8906
rect 40592 8842 40644 8848
rect 40604 8276 40632 8842
rect 40696 8430 40724 11999
rect 41064 11762 41092 12514
rect 41156 12152 41184 12951
rect 41234 12200 41290 13000
rect 41328 12844 41380 12850
rect 41328 12786 41380 12792
rect 41248 12152 41276 12200
rect 41156 12124 41276 12152
rect 41144 11892 41196 11898
rect 41144 11834 41196 11840
rect 41236 11892 41288 11898
rect 41236 11834 41288 11840
rect 41156 11762 41184 11834
rect 40776 11756 40828 11762
rect 40776 11698 40828 11704
rect 41052 11756 41104 11762
rect 41052 11698 41104 11704
rect 41144 11756 41196 11762
rect 41144 11698 41196 11704
rect 40788 11014 40816 11698
rect 41052 11144 41104 11150
rect 41052 11086 41104 11092
rect 40776 11008 40828 11014
rect 40776 10950 40828 10956
rect 40960 11008 41012 11014
rect 40960 10950 41012 10956
rect 40868 9172 40920 9178
rect 40868 9114 40920 9120
rect 40684 8424 40736 8430
rect 40684 8366 40736 8372
rect 40776 8424 40828 8430
rect 40776 8366 40828 8372
rect 40788 8276 40816 8366
rect 40604 8248 40816 8276
rect 40776 8084 40828 8090
rect 40880 8072 40908 9114
rect 40972 8634 41000 10950
rect 41064 10674 41092 11086
rect 41052 10668 41104 10674
rect 41052 10610 41104 10616
rect 41248 9704 41276 11834
rect 41340 11558 41368 12786
rect 41418 12744 41474 12753
rect 41418 12679 41474 12688
rect 41432 12209 41460 12679
rect 41510 12608 41566 12617
rect 41510 12543 41512 12552
rect 41564 12543 41566 12552
rect 41512 12514 41564 12520
rect 41418 12200 41474 12209
rect 41602 12200 41658 13000
rect 41696 12640 41748 12646
rect 41694 12608 41696 12617
rect 41788 12640 41840 12646
rect 41748 12608 41750 12617
rect 41788 12582 41840 12588
rect 41694 12543 41750 12552
rect 41418 12135 41474 12144
rect 41616 12073 41644 12200
rect 41602 12064 41658 12073
rect 41602 11999 41658 12008
rect 41800 11762 41828 12582
rect 41970 12200 42026 13000
rect 42154 12200 42210 12209
rect 42338 12200 42394 13000
rect 42522 12744 42578 12753
rect 42522 12679 42578 12688
rect 41788 11756 41840 11762
rect 41788 11698 41840 11704
rect 41328 11552 41380 11558
rect 41328 11494 41380 11500
rect 41984 11200 42012 12200
rect 42154 12135 42210 12144
rect 42064 11688 42116 11694
rect 42064 11630 42116 11636
rect 41800 11172 42012 11200
rect 41800 11014 41828 11172
rect 42076 11098 42104 11630
rect 41892 11070 42104 11098
rect 41788 11008 41840 11014
rect 41788 10950 41840 10956
rect 41604 10668 41656 10674
rect 41604 10610 41656 10616
rect 41696 10668 41748 10674
rect 41696 10610 41748 10616
rect 41616 10266 41644 10610
rect 41708 10538 41736 10610
rect 41696 10532 41748 10538
rect 41696 10474 41748 10480
rect 41788 10532 41840 10538
rect 41788 10474 41840 10480
rect 41604 10260 41656 10266
rect 41604 10202 41656 10208
rect 41800 9874 41828 10474
rect 41892 10266 41920 11070
rect 42064 11008 42116 11014
rect 42064 10950 42116 10956
rect 42076 10826 42104 10950
rect 41984 10798 42104 10826
rect 41984 10742 42012 10798
rect 41972 10736 42024 10742
rect 41972 10678 42024 10684
rect 42064 10736 42116 10742
rect 42064 10678 42116 10684
rect 42076 10554 42104 10678
rect 41984 10538 42104 10554
rect 41972 10532 42104 10538
rect 42024 10526 42104 10532
rect 41972 10474 42024 10480
rect 42064 10464 42116 10470
rect 42064 10406 42116 10412
rect 42076 10266 42104 10406
rect 41880 10260 41932 10266
rect 41880 10202 41932 10208
rect 42064 10260 42116 10266
rect 42064 10202 42116 10208
rect 41972 10192 42024 10198
rect 41972 10134 42024 10140
rect 41064 9676 41276 9704
rect 41524 9846 41828 9874
rect 41064 9586 41092 9676
rect 41328 9648 41380 9654
rect 41328 9590 41380 9596
rect 41052 9580 41104 9586
rect 41052 9522 41104 9528
rect 41340 9518 41368 9590
rect 41328 9512 41380 9518
rect 41328 9454 41380 9460
rect 41524 9382 41552 9846
rect 41984 9722 42012 10134
rect 41788 9716 41840 9722
rect 41788 9658 41840 9664
rect 41972 9716 42024 9722
rect 41972 9658 42024 9664
rect 41800 9518 41828 9658
rect 41880 9580 41932 9586
rect 41880 9522 41932 9528
rect 41972 9580 42024 9586
rect 41972 9522 42024 9528
rect 41788 9512 41840 9518
rect 41788 9454 41840 9460
rect 41512 9376 41564 9382
rect 41512 9318 41564 9324
rect 41248 9132 41736 9160
rect 41248 9042 41276 9132
rect 41236 9036 41288 9042
rect 41236 8978 41288 8984
rect 41512 9036 41564 9042
rect 41512 8978 41564 8984
rect 41236 8900 41288 8906
rect 41236 8842 41288 8848
rect 40960 8628 41012 8634
rect 40960 8570 41012 8576
rect 41248 8548 41276 8842
rect 41524 8634 41552 8978
rect 41604 8968 41656 8974
rect 41604 8910 41656 8916
rect 41512 8628 41564 8634
rect 41512 8570 41564 8576
rect 41248 8520 41368 8548
rect 40960 8492 41012 8498
rect 40960 8434 41012 8440
rect 40972 8276 41000 8434
rect 40972 8248 41276 8276
rect 40828 8044 40908 8072
rect 40776 8026 40828 8032
rect 41248 8022 41276 8248
rect 41236 8016 41288 8022
rect 41236 7958 41288 7964
rect 41340 7954 41368 8520
rect 41616 8498 41644 8910
rect 41708 8498 41736 9132
rect 41892 9042 41920 9522
rect 41984 9178 42012 9522
rect 41972 9172 42024 9178
rect 42168 9160 42196 12135
rect 42246 12064 42302 12073
rect 42246 11999 42302 12008
rect 42260 11898 42288 11999
rect 42352 11937 42380 12200
rect 42536 12152 42564 12679
rect 42706 12200 42762 13000
rect 43074 12200 43130 13000
rect 43166 12744 43222 12753
rect 43166 12679 43222 12688
rect 42720 12152 42748 12200
rect 42536 12124 42748 12152
rect 42338 11928 42394 11937
rect 42248 11892 42300 11898
rect 42338 11863 42394 11872
rect 42432 11892 42484 11898
rect 42248 11834 42300 11840
rect 42432 11834 42484 11840
rect 41972 9114 42024 9120
rect 42076 9132 42196 9160
rect 41880 9036 41932 9042
rect 41880 8978 41932 8984
rect 41972 9036 42024 9042
rect 41972 8978 42024 8984
rect 41604 8492 41656 8498
rect 41604 8434 41656 8440
rect 41696 8492 41748 8498
rect 41696 8434 41748 8440
rect 41604 8084 41656 8090
rect 41524 8044 41604 8072
rect 41328 7948 41380 7954
rect 41328 7890 41380 7896
rect 41144 7880 41196 7886
rect 40604 7806 41000 7834
rect 41420 7880 41472 7886
rect 41196 7828 41420 7834
rect 41144 7822 41472 7828
rect 41156 7806 41460 7822
rect 40604 7546 40632 7806
rect 40972 7750 41000 7806
rect 40868 7744 40920 7750
rect 40868 7686 40920 7692
rect 40960 7744 41012 7750
rect 40960 7686 41012 7692
rect 41144 7744 41196 7750
rect 41524 7732 41552 8044
rect 41604 8026 41656 8032
rect 41196 7704 41552 7732
rect 41604 7744 41656 7750
rect 41144 7686 41196 7692
rect 41604 7686 41656 7692
rect 40880 7562 40908 7686
rect 41616 7562 41644 7686
rect 40592 7540 40644 7546
rect 40592 7482 40644 7488
rect 40684 7540 40736 7546
rect 40880 7534 41644 7562
rect 40684 7482 40736 7488
rect 40592 7404 40644 7410
rect 40592 7346 40644 7352
rect 40604 6866 40632 7346
rect 40696 7342 40724 7482
rect 41340 7410 41828 7426
rect 41340 7404 41840 7410
rect 41340 7398 41788 7404
rect 40684 7336 40736 7342
rect 40684 7278 40736 7284
rect 40868 7268 40920 7274
rect 40868 7210 40920 7216
rect 40592 6860 40644 6866
rect 40592 6802 40644 6808
rect 40880 6458 40908 7210
rect 41236 6792 41288 6798
rect 41340 6780 41368 7398
rect 41788 7346 41840 7352
rect 41420 7336 41472 7342
rect 41604 7336 41656 7342
rect 41472 7296 41552 7324
rect 41420 7278 41472 7284
rect 41420 6996 41472 7002
rect 41420 6938 41472 6944
rect 41432 6866 41460 6938
rect 41420 6860 41472 6866
rect 41420 6802 41472 6808
rect 41288 6752 41368 6780
rect 41236 6734 41288 6740
rect 41524 6662 41552 7296
rect 41604 7278 41656 7284
rect 41696 7336 41748 7342
rect 41696 7278 41748 7284
rect 41984 7290 42012 8978
rect 42076 8906 42104 9132
rect 42260 9092 42288 11834
rect 42444 10826 42472 11834
rect 42800 11144 42852 11150
rect 42800 11086 42852 11092
rect 42352 10798 42472 10826
rect 42352 10742 42380 10798
rect 42340 10736 42392 10742
rect 42340 10678 42392 10684
rect 42432 10736 42484 10742
rect 42432 10678 42484 10684
rect 42444 10266 42472 10678
rect 42812 10266 42840 11086
rect 42432 10260 42484 10266
rect 42432 10202 42484 10208
rect 42800 10260 42852 10266
rect 42800 10202 42852 10208
rect 42616 9920 42668 9926
rect 42616 9862 42668 9868
rect 42628 9654 42656 9862
rect 42616 9648 42668 9654
rect 42616 9590 42668 9596
rect 42984 9648 43036 9654
rect 42984 9590 43036 9596
rect 42432 9580 42484 9586
rect 42432 9522 42484 9528
rect 42444 9178 42472 9522
rect 42536 9438 42932 9466
rect 42432 9172 42484 9178
rect 42432 9114 42484 9120
rect 42168 9064 42288 9092
rect 42064 8900 42116 8906
rect 42064 8842 42116 8848
rect 42168 8838 42196 9064
rect 42536 9024 42564 9438
rect 42616 9376 42668 9382
rect 42800 9376 42852 9382
rect 42616 9318 42668 9324
rect 42706 9344 42762 9353
rect 42628 9178 42656 9318
rect 42904 9353 42932 9438
rect 42800 9318 42852 9324
rect 42890 9344 42946 9353
rect 42706 9279 42762 9288
rect 42616 9172 42668 9178
rect 42616 9114 42668 9120
rect 42720 9081 42748 9279
rect 42260 8996 42564 9024
rect 42706 9072 42762 9081
rect 42706 9007 42762 9016
rect 42156 8832 42208 8838
rect 42156 8774 42208 8780
rect 42260 8401 42288 8996
rect 42812 8974 42840 9318
rect 42890 9279 42946 9288
rect 42996 9110 43024 9590
rect 42984 9104 43036 9110
rect 42984 9046 43036 9052
rect 42800 8968 42852 8974
rect 42800 8910 42852 8916
rect 42892 8968 42944 8974
rect 42892 8910 42944 8916
rect 42432 8900 42484 8906
rect 42432 8842 42484 8848
rect 42444 8566 42472 8842
rect 42536 8622 42840 8650
rect 42432 8560 42484 8566
rect 42432 8502 42484 8508
rect 42246 8392 42302 8401
rect 42246 8327 42302 8336
rect 42536 8242 42564 8622
rect 42616 8560 42668 8566
rect 42616 8502 42668 8508
rect 42076 8214 42564 8242
rect 42076 7886 42104 8214
rect 42628 8004 42656 8502
rect 42260 7976 42656 8004
rect 42064 7880 42116 7886
rect 42064 7822 42116 7828
rect 42260 7546 42288 7976
rect 42708 7948 42760 7954
rect 42444 7908 42708 7936
rect 42340 7744 42392 7750
rect 42340 7686 42392 7692
rect 42248 7540 42300 7546
rect 42248 7482 42300 7488
rect 42248 7404 42300 7410
rect 42352 7392 42380 7686
rect 42300 7364 42380 7392
rect 42248 7346 42300 7352
rect 42156 7336 42208 7342
rect 41616 6798 41644 7278
rect 41708 7041 41736 7278
rect 41984 7262 42104 7290
rect 42208 7284 42288 7290
rect 42156 7278 42288 7284
rect 42168 7262 42288 7278
rect 42444 7274 42472 7908
rect 42708 7890 42760 7896
rect 42616 7540 42668 7546
rect 42536 7500 42616 7528
rect 41694 7032 41750 7041
rect 41878 7032 41934 7041
rect 41800 7002 41878 7018
rect 41694 6967 41750 6976
rect 41788 6996 41878 7002
rect 41840 6990 41878 6996
rect 41878 6967 41934 6976
rect 41788 6938 41840 6944
rect 41696 6928 41748 6934
rect 41696 6870 41748 6876
rect 41604 6792 41656 6798
rect 41604 6734 41656 6740
rect 41420 6656 41472 6662
rect 41420 6598 41472 6604
rect 41512 6656 41564 6662
rect 41512 6598 41564 6604
rect 40868 6452 40920 6458
rect 40868 6394 40920 6400
rect 41144 6452 41196 6458
rect 41144 6394 41196 6400
rect 40512 6310 40724 6338
rect 41156 6322 41184 6394
rect 41432 6390 41460 6598
rect 41708 6440 41736 6870
rect 41972 6792 42024 6798
rect 41972 6734 42024 6740
rect 41616 6412 41736 6440
rect 41328 6384 41380 6390
rect 41328 6326 41380 6332
rect 41420 6384 41472 6390
rect 41420 6326 41472 6332
rect 40500 5772 40552 5778
rect 40500 5714 40552 5720
rect 40328 3420 40448 3448
rect 40222 3360 40278 3369
rect 40222 3295 40278 3304
rect 39948 3120 40000 3126
rect 39948 3062 40000 3068
rect 40040 3120 40092 3126
rect 40040 3062 40092 3068
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 39948 2984 40000 2990
rect 39946 2952 39948 2961
rect 40000 2952 40002 2961
rect 39946 2887 40002 2896
rect 39856 2848 39908 2854
rect 39856 2790 39908 2796
rect 39224 2264 39804 2292
rect 39868 2292 39896 2790
rect 40144 2666 40172 2994
rect 40236 2961 40264 3295
rect 40328 3058 40356 3420
rect 40406 3360 40462 3369
rect 40406 3295 40462 3304
rect 40316 3052 40368 3058
rect 40316 2994 40368 3000
rect 40222 2952 40278 2961
rect 40222 2887 40278 2896
rect 40420 2825 40448 3295
rect 40512 2854 40540 5714
rect 40696 5386 40724 6310
rect 41144 6316 41196 6322
rect 41144 6258 41196 6264
rect 41340 6254 41368 6326
rect 41616 6322 41644 6412
rect 41604 6316 41656 6322
rect 41604 6258 41656 6264
rect 41696 6316 41748 6322
rect 41696 6258 41748 6264
rect 41880 6316 41932 6322
rect 41880 6258 41932 6264
rect 41328 6248 41380 6254
rect 41328 6190 41380 6196
rect 41708 5778 41736 6258
rect 41696 5772 41748 5778
rect 41696 5714 41748 5720
rect 41892 5574 41920 6258
rect 41984 5574 42012 6734
rect 41880 5568 41932 5574
rect 41880 5510 41932 5516
rect 41972 5568 42024 5574
rect 41972 5510 42024 5516
rect 42076 5386 42104 7262
rect 42156 6928 42208 6934
rect 42156 6870 42208 6876
rect 42168 6322 42196 6870
rect 42260 6798 42288 7262
rect 42432 7268 42484 7274
rect 42432 7210 42484 7216
rect 42536 6866 42564 7500
rect 42616 7482 42668 7488
rect 42616 7336 42668 7342
rect 42616 7278 42668 7284
rect 42628 6866 42656 7278
rect 42812 7274 42840 8622
rect 42800 7268 42852 7274
rect 42800 7210 42852 7216
rect 42524 6860 42576 6866
rect 42524 6802 42576 6808
rect 42616 6860 42668 6866
rect 42904 6848 42932 8910
rect 43088 8566 43116 12200
rect 43180 10606 43208 12679
rect 43442 12200 43498 13000
rect 43810 12200 43866 13000
rect 44178 12200 44234 13000
rect 44546 12200 44602 13000
rect 44914 12200 44970 13000
rect 45098 12336 45154 12345
rect 45098 12271 45154 12280
rect 43352 10668 43404 10674
rect 43352 10610 43404 10616
rect 43168 10600 43220 10606
rect 43168 10542 43220 10548
rect 43180 9926 43208 10542
rect 43364 10470 43392 10610
rect 43352 10464 43404 10470
rect 43352 10406 43404 10412
rect 43168 9920 43220 9926
rect 43168 9862 43220 9868
rect 43352 9172 43404 9178
rect 43352 9114 43404 9120
rect 43364 8974 43392 9114
rect 43352 8968 43404 8974
rect 43352 8910 43404 8916
rect 43076 8560 43128 8566
rect 43076 8502 43128 8508
rect 42904 6820 43024 6848
rect 42616 6802 42668 6808
rect 42248 6792 42300 6798
rect 42248 6734 42300 6740
rect 42524 6724 42576 6730
rect 42892 6724 42944 6730
rect 42576 6684 42892 6712
rect 42524 6666 42576 6672
rect 42892 6666 42944 6672
rect 42996 6474 43024 6820
rect 43456 6474 43484 12200
rect 43718 11928 43774 11937
rect 43824 11898 43852 12200
rect 43718 11863 43774 11872
rect 43812 11892 43864 11898
rect 43732 11354 43760 11863
rect 43812 11834 43864 11840
rect 44086 11792 44142 11801
rect 44086 11727 44142 11736
rect 43720 11348 43772 11354
rect 43720 11290 43772 11296
rect 44100 9926 44128 11727
rect 44088 9920 44140 9926
rect 44088 9862 44140 9868
rect 43904 9648 43956 9654
rect 43904 9590 43956 9596
rect 43916 8906 43944 9590
rect 43904 8900 43956 8906
rect 43904 8842 43956 8848
rect 43536 8832 43588 8838
rect 43536 8774 43588 8780
rect 43548 8498 43576 8774
rect 43536 8492 43588 8498
rect 43536 8434 43588 8440
rect 44192 7206 44220 12200
rect 44560 10198 44588 12200
rect 44548 10192 44600 10198
rect 44548 10134 44600 10140
rect 44928 9738 44956 12200
rect 45112 12152 45140 12271
rect 45282 12200 45338 13000
rect 45650 12200 45706 13000
rect 45928 12776 45980 12782
rect 45928 12718 45980 12724
rect 45296 12152 45324 12200
rect 45112 12124 45324 12152
rect 45558 11520 45614 11529
rect 45558 11455 45614 11464
rect 45572 10470 45600 11455
rect 45664 11150 45692 12200
rect 45742 11792 45798 11801
rect 45742 11727 45798 11736
rect 45652 11144 45704 11150
rect 45652 11086 45704 11092
rect 45756 10985 45784 11727
rect 45836 11348 45888 11354
rect 45836 11290 45888 11296
rect 45848 11150 45876 11290
rect 45940 11150 45968 12718
rect 46018 12200 46074 13000
rect 46296 12912 46348 12918
rect 46294 12880 46296 12889
rect 46348 12880 46350 12889
rect 46294 12815 46350 12824
rect 46386 12200 46442 13000
rect 46480 12776 46532 12782
rect 46478 12744 46480 12753
rect 46532 12744 46534 12753
rect 46478 12679 46534 12688
rect 46478 12608 46534 12617
rect 46478 12543 46534 12552
rect 45836 11144 45888 11150
rect 45836 11086 45888 11092
rect 45928 11144 45980 11150
rect 45928 11086 45980 11092
rect 45742 10976 45798 10985
rect 45742 10911 45798 10920
rect 45848 10742 45876 11086
rect 45836 10736 45888 10742
rect 45836 10678 45888 10684
rect 45836 10600 45888 10606
rect 45836 10542 45888 10548
rect 45560 10464 45612 10470
rect 45560 10406 45612 10412
rect 45112 10130 45324 10146
rect 45100 10124 45336 10130
rect 45152 10118 45284 10124
rect 45100 10066 45152 10072
rect 45284 10066 45336 10072
rect 45848 10062 45876 10542
rect 45836 10056 45888 10062
rect 45836 9998 45888 10004
rect 44744 9710 44956 9738
rect 44456 9376 44508 9382
rect 44456 9318 44508 9324
rect 44272 7336 44324 7342
rect 44272 7278 44324 7284
rect 44284 7206 44312 7278
rect 43536 7200 43588 7206
rect 43536 7142 43588 7148
rect 44180 7200 44232 7206
rect 44180 7142 44232 7148
rect 44272 7200 44324 7206
rect 44272 7142 44324 7148
rect 42536 6446 43024 6474
rect 43180 6446 43484 6474
rect 43548 6458 43576 7142
rect 43628 6860 43680 6866
rect 43628 6802 43680 6808
rect 43536 6452 43588 6458
rect 42156 6316 42208 6322
rect 42156 6258 42208 6264
rect 42156 5704 42208 5710
rect 42156 5646 42208 5652
rect 40696 5358 41000 5386
rect 40776 5228 40828 5234
rect 40776 5170 40828 5176
rect 40868 5228 40920 5234
rect 40868 5170 40920 5176
rect 40788 4604 40816 5170
rect 40880 4865 40908 5170
rect 40866 4856 40922 4865
rect 40972 4842 41000 5358
rect 41340 5358 42104 5386
rect 41340 5234 41368 5358
rect 41328 5228 41380 5234
rect 41328 5170 41380 5176
rect 41420 5228 41472 5234
rect 41420 5170 41472 5176
rect 41050 4856 41106 4865
rect 40972 4814 41050 4842
rect 40866 4791 40922 4800
rect 41050 4791 41106 4800
rect 40868 4616 40920 4622
rect 40788 4576 40868 4604
rect 40868 4558 40920 4564
rect 41432 4554 41460 5170
rect 41510 5128 41566 5137
rect 41566 5086 41644 5114
rect 41510 5063 41566 5072
rect 41616 4690 41644 5086
rect 41512 4684 41564 4690
rect 41512 4626 41564 4632
rect 41604 4684 41656 4690
rect 41604 4626 41656 4632
rect 41524 4554 41552 4626
rect 41420 4548 41472 4554
rect 41420 4490 41472 4496
rect 41512 4548 41564 4554
rect 42168 4536 42196 5646
rect 42340 5568 42392 5574
rect 42340 5510 42392 5516
rect 42432 5568 42484 5574
rect 42432 5510 42484 5516
rect 41512 4490 41564 4496
rect 41616 4508 42196 4536
rect 41512 4208 41564 4214
rect 41616 4196 41644 4508
rect 41878 4448 41934 4457
rect 41878 4383 41934 4392
rect 41892 4264 41920 4383
rect 41564 4168 41644 4196
rect 41708 4236 41920 4264
rect 41708 4185 41736 4236
rect 41694 4176 41750 4185
rect 41512 4150 41564 4156
rect 41694 4111 41750 4120
rect 41878 4176 41934 4185
rect 41878 4111 41934 4120
rect 41972 4140 42024 4146
rect 40776 4072 40828 4078
rect 40776 4014 40828 4020
rect 41052 4072 41104 4078
rect 41052 4014 41104 4020
rect 40788 3058 40816 4014
rect 41064 3466 41092 4014
rect 41512 4004 41564 4010
rect 41432 3964 41512 3992
rect 41236 3664 41288 3670
rect 41236 3606 41288 3612
rect 41052 3460 41104 3466
rect 41052 3402 41104 3408
rect 41248 3398 41276 3606
rect 41432 3466 41460 3964
rect 41512 3946 41564 3952
rect 41786 3768 41842 3777
rect 41524 3726 41786 3754
rect 41524 3641 41552 3726
rect 41786 3703 41842 3712
rect 41510 3632 41566 3641
rect 41510 3567 41566 3576
rect 41604 3528 41656 3534
rect 41524 3488 41604 3516
rect 41420 3460 41472 3466
rect 41420 3402 41472 3408
rect 41236 3392 41288 3398
rect 41236 3334 41288 3340
rect 41524 3194 41552 3488
rect 41604 3470 41656 3476
rect 41892 3466 41920 4111
rect 41972 4082 42024 4088
rect 41984 3602 42012 4082
rect 41972 3596 42024 3602
rect 41972 3538 42024 3544
rect 42064 3596 42116 3602
rect 42352 3584 42380 5510
rect 42444 4457 42472 5510
rect 42430 4448 42486 4457
rect 42430 4383 42486 4392
rect 42536 4146 42564 6446
rect 43180 6390 43208 6446
rect 43536 6394 43588 6400
rect 42984 6384 43036 6390
rect 42984 6326 43036 6332
rect 43168 6384 43220 6390
rect 43168 6326 43220 6332
rect 43444 6384 43496 6390
rect 43444 6326 43496 6332
rect 42800 6316 42852 6322
rect 42800 6258 42852 6264
rect 42812 5930 42840 6258
rect 42996 6066 43024 6326
rect 43352 6180 43404 6186
rect 43352 6122 43404 6128
rect 43364 6066 43392 6122
rect 42996 6038 43392 6066
rect 42720 5914 42840 5930
rect 42708 5908 42840 5914
rect 42760 5902 42840 5908
rect 42708 5850 42760 5856
rect 42984 5840 43036 5846
rect 43456 5794 43484 6326
rect 43536 6248 43588 6254
rect 43536 6190 43588 6196
rect 43036 5788 43484 5794
rect 42984 5782 43484 5788
rect 42996 5766 43484 5782
rect 43548 5624 43576 6190
rect 43088 5596 43576 5624
rect 43088 5234 43116 5596
rect 43640 5522 43668 6802
rect 43720 6792 43772 6798
rect 43720 6734 43772 6740
rect 43732 6458 43760 6734
rect 43720 6452 43772 6458
rect 43720 6394 43772 6400
rect 44364 5908 44416 5914
rect 44364 5850 44416 5856
rect 43180 5494 43668 5522
rect 43076 5228 43128 5234
rect 43076 5170 43128 5176
rect 42800 4208 42852 4214
rect 42800 4150 42852 4156
rect 42524 4140 42576 4146
rect 42524 4082 42576 4088
rect 42616 4140 42668 4146
rect 42616 4082 42668 4088
rect 42352 3556 42472 3584
rect 42064 3538 42116 3544
rect 41880 3460 41932 3466
rect 41880 3402 41932 3408
rect 41512 3188 41564 3194
rect 41512 3130 41564 3136
rect 41604 3188 41656 3194
rect 41604 3130 41656 3136
rect 41052 3120 41104 3126
rect 41616 3074 41644 3130
rect 41104 3068 41644 3074
rect 41052 3062 41644 3068
rect 40776 3052 40828 3058
rect 41064 3046 41644 3062
rect 41696 3052 41748 3058
rect 40776 2994 40828 3000
rect 42076 3040 42104 3538
rect 42340 3460 42392 3466
rect 42340 3402 42392 3408
rect 42352 3058 42380 3402
rect 41696 2994 41748 3000
rect 41800 3012 42104 3040
rect 42340 3052 42392 3058
rect 41708 2922 41736 2994
rect 41696 2916 41748 2922
rect 40788 2876 41092 2904
rect 40500 2848 40552 2854
rect 40406 2816 40462 2825
rect 40788 2825 40816 2876
rect 40500 2790 40552 2796
rect 40774 2816 40830 2825
rect 40406 2751 40462 2760
rect 40774 2751 40830 2760
rect 40958 2816 41014 2825
rect 40958 2751 41014 2760
rect 40144 2650 40264 2666
rect 40144 2644 40276 2650
rect 40144 2638 40224 2644
rect 40224 2586 40276 2592
rect 39948 2576 40000 2582
rect 40500 2576 40552 2582
rect 40420 2536 40500 2564
rect 40420 2530 40448 2536
rect 40000 2524 40448 2530
rect 39948 2518 40448 2524
rect 40500 2518 40552 2524
rect 39960 2502 40448 2518
rect 40868 2508 40920 2514
rect 40868 2450 40920 2456
rect 40500 2440 40552 2446
rect 40880 2394 40908 2450
rect 40552 2388 40908 2394
rect 40500 2382 40908 2388
rect 40512 2366 40908 2382
rect 39868 2264 40724 2292
rect 39028 1352 39080 1358
rect 39028 1294 39080 1300
rect 39120 1352 39172 1358
rect 39120 1294 39172 1300
rect 38936 876 38988 882
rect 38936 818 38988 824
rect 39040 814 39068 1294
rect 39028 808 39080 814
rect 38292 750 38344 756
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39224 800 39252 2264
rect 39500 1686 40632 1714
rect 39500 1290 39528 1686
rect 39592 1550 40448 1578
rect 39592 1426 39620 1550
rect 40132 1488 40184 1494
rect 40184 1436 40356 1442
rect 40132 1430 40356 1436
rect 39580 1420 39632 1426
rect 39580 1362 39632 1368
rect 39672 1420 39724 1426
rect 40144 1414 40356 1430
rect 39672 1362 39724 1368
rect 39488 1284 39540 1290
rect 39488 1226 39540 1232
rect 39684 864 39712 1362
rect 40224 1352 40276 1358
rect 40052 1312 40224 1340
rect 40052 1204 40080 1312
rect 40224 1294 40276 1300
rect 39592 836 39712 864
rect 39960 1176 40080 1204
rect 39304 808 39356 814
rect 39028 750 39080 756
rect 39210 0 39266 800
rect 39592 800 39620 836
rect 39960 800 39988 1176
rect 40328 800 40356 1414
rect 40420 1358 40448 1550
rect 40500 1556 40552 1562
rect 40500 1498 40552 1504
rect 40408 1352 40460 1358
rect 40408 1294 40460 1300
rect 40408 1216 40460 1222
rect 40408 1158 40460 1164
rect 40512 1170 40540 1498
rect 40604 1290 40632 1686
rect 40696 1562 40724 2264
rect 40684 1556 40736 1562
rect 40972 1544 41000 2751
rect 41064 2530 41092 2876
rect 41696 2858 41748 2864
rect 41328 2644 41380 2650
rect 41800 2632 41828 3012
rect 42340 2994 42392 3000
rect 41880 2916 41932 2922
rect 41880 2858 41932 2864
rect 41972 2916 42024 2922
rect 41972 2858 42024 2864
rect 41892 2650 41920 2858
rect 41380 2604 41828 2632
rect 41880 2644 41932 2650
rect 41328 2586 41380 2592
rect 41880 2586 41932 2592
rect 41064 2502 41552 2530
rect 41984 2514 42012 2858
rect 42444 2650 42472 3556
rect 42432 2644 42484 2650
rect 42432 2586 42484 2592
rect 41144 2440 41196 2446
rect 41144 2382 41196 2388
rect 41156 2122 41184 2382
rect 41156 2094 41460 2122
rect 41432 2038 41460 2094
rect 41328 2032 41380 2038
rect 41328 1974 41380 1980
rect 41420 2032 41472 2038
rect 41420 1974 41472 1980
rect 41052 1896 41104 1902
rect 41052 1838 41104 1844
rect 41144 1896 41196 1902
rect 41144 1838 41196 1844
rect 40684 1498 40736 1504
rect 40880 1516 41000 1544
rect 40880 1426 40908 1516
rect 40868 1420 40920 1426
rect 40868 1362 40920 1368
rect 40960 1420 41012 1426
rect 40960 1362 41012 1368
rect 40866 1320 40922 1329
rect 40592 1284 40644 1290
rect 40972 1306 41000 1362
rect 41064 1329 41092 1838
rect 40922 1278 41000 1306
rect 41050 1320 41106 1329
rect 40866 1255 40922 1264
rect 41050 1255 41106 1264
rect 40592 1226 40644 1232
rect 41156 1170 41184 1838
rect 41340 1766 41368 1974
rect 41328 1760 41380 1766
rect 41524 1748 41552 2502
rect 41972 2508 42024 2514
rect 41972 2450 42024 2456
rect 42628 2394 42656 4082
rect 42708 2984 42760 2990
rect 42708 2926 42760 2932
rect 42352 2366 42656 2394
rect 41604 1964 41656 1970
rect 41604 1906 41656 1912
rect 41616 1816 41644 1906
rect 41616 1788 42288 1816
rect 41524 1720 42196 1748
rect 41328 1702 41380 1708
rect 41972 1556 42024 1562
rect 41972 1498 42024 1504
rect 41328 1420 41380 1426
rect 41512 1420 41564 1426
rect 41380 1380 41460 1408
rect 41328 1362 41380 1368
rect 39304 750 39356 756
rect 39316 678 39344 750
rect 39304 672 39356 678
rect 39304 614 39356 620
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40420 746 40448 1158
rect 40512 1142 40632 1170
rect 40604 814 40632 1142
rect 40788 1142 41184 1170
rect 40788 1018 40816 1142
rect 40776 1012 40828 1018
rect 40776 954 40828 960
rect 40960 1012 41012 1018
rect 40960 954 41012 960
rect 40684 944 40736 950
rect 40684 886 40736 892
rect 40868 944 40920 950
rect 40868 886 40920 892
rect 40500 808 40552 814
rect 40500 750 40552 756
rect 40592 808 40644 814
rect 40696 800 40724 886
rect 40592 750 40644 756
rect 40408 740 40460 746
rect 40408 682 40460 688
rect 40512 513 40540 750
rect 40498 504 40554 513
rect 40498 439 40554 448
rect 40682 0 40738 800
rect 40880 746 40908 886
rect 40868 740 40920 746
rect 40868 682 40920 688
rect 40972 134 41000 954
rect 41064 836 41184 864
rect 41064 800 41092 836
rect 40960 128 41012 134
rect 40960 70 41012 76
rect 41050 0 41106 800
rect 41156 66 41184 836
rect 41432 800 41460 1380
rect 41512 1362 41564 1368
rect 41524 882 41552 1362
rect 41696 1352 41748 1358
rect 41616 1312 41696 1340
rect 41512 876 41564 882
rect 41512 818 41564 824
rect 41326 504 41382 513
rect 41326 439 41382 448
rect 41340 134 41368 439
rect 41328 128 41380 134
rect 41328 70 41380 76
rect 41144 60 41196 66
rect 41144 2 41196 8
rect 41418 0 41474 800
rect 41616 678 41644 1312
rect 41696 1294 41748 1300
rect 41984 950 42012 1498
rect 41972 944 42024 950
rect 41972 886 42024 892
rect 41708 836 41828 864
rect 41708 746 41736 836
rect 41800 800 41828 836
rect 42168 800 42196 1720
rect 42260 1562 42288 1788
rect 42248 1556 42300 1562
rect 42248 1498 42300 1504
rect 42352 1170 42380 2366
rect 42616 2304 42668 2310
rect 42616 2246 42668 2252
rect 42628 2106 42656 2246
rect 42616 2100 42668 2106
rect 42616 2042 42668 2048
rect 42720 2088 42748 2926
rect 42812 2836 42840 4150
rect 43180 3720 43208 5494
rect 43536 5364 43588 5370
rect 43536 5306 43588 5312
rect 43628 5364 43680 5370
rect 43628 5306 43680 5312
rect 43352 5160 43404 5166
rect 43352 5102 43404 5108
rect 43364 5030 43392 5102
rect 43548 5030 43576 5306
rect 43352 5024 43404 5030
rect 43352 4966 43404 4972
rect 43536 5024 43588 5030
rect 43536 4966 43588 4972
rect 43258 4448 43314 4457
rect 43258 4383 43314 4392
rect 42996 3692 43208 3720
rect 42996 3602 43024 3692
rect 42984 3596 43036 3602
rect 42984 3538 43036 3544
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 43088 3126 43116 3538
rect 43076 3120 43128 3126
rect 43076 3062 43128 3068
rect 43272 2961 43300 4383
rect 43352 4140 43404 4146
rect 43352 4082 43404 4088
rect 43364 3058 43392 4082
rect 43536 3528 43588 3534
rect 43536 3470 43588 3476
rect 43548 3398 43576 3470
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 43536 3392 43588 3398
rect 43536 3334 43588 3340
rect 43456 3126 43484 3334
rect 43444 3120 43496 3126
rect 43444 3062 43496 3068
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 43536 3052 43588 3058
rect 43536 2994 43588 3000
rect 43258 2952 43314 2961
rect 43258 2887 43314 2896
rect 42984 2848 43036 2854
rect 42812 2808 42984 2836
rect 42984 2790 43036 2796
rect 43548 2106 43576 2994
rect 42800 2100 42852 2106
rect 42720 2060 42800 2088
rect 42524 1352 42576 1358
rect 42524 1294 42576 1300
rect 42616 1352 42668 1358
rect 42720 1340 42748 2060
rect 42800 2042 42852 2048
rect 43536 2100 43588 2106
rect 43536 2042 43588 2048
rect 43548 1850 43576 2042
rect 43640 1970 43668 5306
rect 44088 3460 44140 3466
rect 44088 3402 44140 3408
rect 44100 3194 44128 3402
rect 44088 3188 44140 3194
rect 44088 3130 44140 3136
rect 43812 3052 43864 3058
rect 43812 2994 43864 3000
rect 43628 1964 43680 1970
rect 43628 1906 43680 1912
rect 43548 1822 43760 1850
rect 43732 1766 43760 1822
rect 43628 1760 43680 1766
rect 43628 1702 43680 1708
rect 43720 1760 43772 1766
rect 43720 1702 43772 1708
rect 42668 1312 42748 1340
rect 42616 1294 42668 1300
rect 42536 1204 42564 1294
rect 43260 1216 43312 1222
rect 42536 1176 43116 1204
rect 42260 1142 42380 1170
rect 42260 1018 42288 1142
rect 42248 1012 42300 1018
rect 42248 954 42300 960
rect 42340 1012 42392 1018
rect 42340 954 42392 960
rect 41696 740 41748 746
rect 41696 682 41748 688
rect 41604 672 41656 678
rect 41604 614 41656 620
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42352 474 42380 954
rect 43088 950 43116 1176
rect 43260 1158 43312 1164
rect 42524 944 42576 950
rect 42524 886 42576 892
rect 43076 944 43128 950
rect 43076 886 43128 892
rect 42536 800 42564 886
rect 42984 876 43036 882
rect 42812 836 42932 864
rect 42340 468 42392 474
rect 42340 410 42392 416
rect 42522 0 42578 800
rect 42812 474 42840 836
rect 42904 800 42932 836
rect 42984 818 43036 824
rect 42800 468 42852 474
rect 42800 410 42852 416
rect 42890 0 42946 800
rect 42996 474 43024 818
rect 43272 800 43300 1158
rect 43640 800 43668 1702
rect 43824 1426 43852 2994
rect 44086 2952 44142 2961
rect 44086 2887 44142 2896
rect 44100 2650 44128 2887
rect 44088 2644 44140 2650
rect 44088 2586 44140 2592
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 44192 2530 44220 2586
rect 43916 2514 44220 2530
rect 43904 2508 44220 2514
rect 43956 2502 44220 2508
rect 44272 2508 44324 2514
rect 43904 2450 43956 2456
rect 44272 2450 44324 2456
rect 44180 2440 44232 2446
rect 44180 2382 44232 2388
rect 44192 2106 44220 2382
rect 44284 2106 44312 2450
rect 44180 2100 44232 2106
rect 44180 2042 44232 2048
rect 44272 2100 44324 2106
rect 44272 2042 44324 2048
rect 44192 1970 44220 2042
rect 44180 1964 44232 1970
rect 44180 1906 44232 1912
rect 43996 1488 44048 1494
rect 44376 1476 44404 5850
rect 44468 3602 44496 9318
rect 44744 8090 44772 9710
rect 46032 9625 46060 12200
rect 46204 12164 46256 12170
rect 46204 12106 46256 12112
rect 46216 11898 46244 12106
rect 46204 11892 46256 11898
rect 46204 11834 46256 11840
rect 46296 11688 46348 11694
rect 46296 11630 46348 11636
rect 46202 11520 46258 11529
rect 46202 11455 46258 11464
rect 46110 10976 46166 10985
rect 46110 10911 46166 10920
rect 46124 10577 46152 10911
rect 46110 10568 46166 10577
rect 46110 10503 46166 10512
rect 46216 9897 46244 11455
rect 46308 11354 46336 11630
rect 46296 11348 46348 11354
rect 46296 11290 46348 11296
rect 46400 11200 46428 12200
rect 46492 11694 46520 12543
rect 46754 12200 46810 13000
rect 47122 12200 47178 13000
rect 47490 12200 47546 13000
rect 47858 12200 47914 13000
rect 48226 12200 48282 13000
rect 48502 12608 48558 12617
rect 48502 12543 48558 12552
rect 48516 12209 48544 12543
rect 48502 12200 48558 12209
rect 48594 12200 48650 13000
rect 48962 12200 49018 13000
rect 49330 12200 49386 13000
rect 49698 12200 49754 13000
rect 50066 12200 50122 13000
rect 50434 12200 50490 13000
rect 50712 12504 50764 12510
rect 50712 12446 50764 12452
rect 50618 12200 50674 12209
rect 46570 11928 46626 11937
rect 46570 11863 46626 11872
rect 46480 11688 46532 11694
rect 46480 11630 46532 11636
rect 46584 11354 46612 11863
rect 46572 11348 46624 11354
rect 46572 11290 46624 11296
rect 46308 11172 46428 11200
rect 46202 9888 46258 9897
rect 46202 9823 46258 9832
rect 46018 9616 46074 9625
rect 46018 9551 46074 9560
rect 46202 9616 46258 9625
rect 46202 9551 46258 9560
rect 46216 9042 46244 9551
rect 46308 9518 46336 11172
rect 46664 11144 46716 11150
rect 46664 11086 46716 11092
rect 46388 11076 46440 11082
rect 46388 11018 46440 11024
rect 46400 10674 46428 11018
rect 46676 11014 46704 11086
rect 46664 11008 46716 11014
rect 46664 10950 46716 10956
rect 46388 10668 46440 10674
rect 46388 10610 46440 10616
rect 46572 10532 46624 10538
rect 46572 10474 46624 10480
rect 46584 10266 46612 10474
rect 46572 10260 46624 10266
rect 46572 10202 46624 10208
rect 46386 9888 46442 9897
rect 46386 9823 46442 9832
rect 46296 9512 46348 9518
rect 46296 9454 46348 9460
rect 46204 9036 46256 9042
rect 46204 8978 46256 8984
rect 45928 8628 45980 8634
rect 45928 8570 45980 8576
rect 46112 8628 46164 8634
rect 46112 8570 46164 8576
rect 45560 8424 45612 8430
rect 45560 8366 45612 8372
rect 44732 8084 44784 8090
rect 44732 8026 44784 8032
rect 44824 8084 44876 8090
rect 44824 8026 44876 8032
rect 44836 7954 44864 8026
rect 44824 7948 44876 7954
rect 44824 7890 44876 7896
rect 45572 7546 45600 8366
rect 45940 8362 45968 8570
rect 46124 8537 46152 8570
rect 46110 8528 46166 8537
rect 46110 8463 46166 8472
rect 45928 8356 45980 8362
rect 45928 8298 45980 8304
rect 45744 8288 45796 8294
rect 45744 8230 45796 8236
rect 45756 7954 45784 8230
rect 45744 7948 45796 7954
rect 45744 7890 45796 7896
rect 45836 7948 45888 7954
rect 45836 7890 45888 7896
rect 45756 7546 45784 7890
rect 45560 7540 45612 7546
rect 45560 7482 45612 7488
rect 45744 7540 45796 7546
rect 45744 7482 45796 7488
rect 44548 7404 44600 7410
rect 44548 7346 44600 7352
rect 44560 5710 44588 7346
rect 45100 7268 45152 7274
rect 45100 7210 45152 7216
rect 44916 7200 44968 7206
rect 44916 7142 44968 7148
rect 44928 6798 44956 7142
rect 45112 7002 45140 7210
rect 45100 6996 45152 7002
rect 45100 6938 45152 6944
rect 45468 6996 45520 7002
rect 45468 6938 45520 6944
rect 44916 6792 44968 6798
rect 44916 6734 44968 6740
rect 45376 6792 45428 6798
rect 45376 6734 45428 6740
rect 44548 5704 44600 5710
rect 44548 5646 44600 5652
rect 45284 5636 45336 5642
rect 45284 5578 45336 5584
rect 44916 4548 44968 4554
rect 44916 4490 44968 4496
rect 45192 4548 45244 4554
rect 45192 4490 45244 4496
rect 44548 4140 44600 4146
rect 44548 4082 44600 4088
rect 44824 4140 44876 4146
rect 44824 4082 44876 4088
rect 44560 3602 44588 4082
rect 44456 3596 44508 3602
rect 44456 3538 44508 3544
rect 44548 3596 44600 3602
rect 44548 3538 44600 3544
rect 44836 3194 44864 4082
rect 44928 3194 44956 4490
rect 44824 3188 44876 3194
rect 44824 3130 44876 3136
rect 44916 3188 44968 3194
rect 44916 3130 44968 3136
rect 44836 3058 44864 3130
rect 44824 3052 44876 3058
rect 44824 2994 44876 3000
rect 44916 3052 44968 3058
rect 44916 2994 44968 3000
rect 44928 2496 44956 2994
rect 44048 1448 44404 1476
rect 44560 2468 44956 2496
rect 43996 1430 44048 1436
rect 43812 1420 43864 1426
rect 43812 1362 43864 1368
rect 44364 1352 44416 1358
rect 44364 1294 44416 1300
rect 43902 1184 43958 1193
rect 43958 1142 44128 1170
rect 43902 1119 43958 1128
rect 44100 882 44128 1142
rect 43904 876 43956 882
rect 44088 876 44140 882
rect 43956 836 44036 864
rect 43904 818 43956 824
rect 44008 800 44036 836
rect 44088 818 44140 824
rect 44376 800 44404 1294
rect 44560 1018 44588 2468
rect 44824 2372 44876 2378
rect 44824 2314 44876 2320
rect 44732 1284 44784 1290
rect 44732 1226 44784 1232
rect 44640 1216 44692 1222
rect 44640 1158 44692 1164
rect 44548 1012 44600 1018
rect 44548 954 44600 960
rect 44652 814 44680 1158
rect 44640 808 44692 814
rect 42984 468 43036 474
rect 42984 410 43036 416
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44744 800 44772 1226
rect 44836 1018 44864 2314
rect 45100 1964 45152 1970
rect 45100 1906 45152 1912
rect 44916 1420 44968 1426
rect 44916 1362 44968 1368
rect 44928 1222 44956 1362
rect 44916 1216 44968 1222
rect 44916 1158 44968 1164
rect 44824 1012 44876 1018
rect 44824 954 44876 960
rect 44916 1012 44968 1018
rect 44916 954 44968 960
rect 44928 882 44956 954
rect 44916 876 44968 882
rect 44916 818 44968 824
rect 45112 800 45140 1906
rect 44640 750 44692 756
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45204 513 45232 4490
rect 45296 4010 45324 5578
rect 45388 5352 45416 6734
rect 45480 6254 45508 6938
rect 45560 6860 45612 6866
rect 45848 6848 45876 7890
rect 46400 7886 46428 9823
rect 46768 9722 46796 12200
rect 47136 11914 47164 12200
rect 46952 11886 47164 11914
rect 46756 9716 46808 9722
rect 46756 9658 46808 9664
rect 46572 9580 46624 9586
rect 46572 9522 46624 9528
rect 46584 9042 46612 9522
rect 46664 9376 46716 9382
rect 46664 9318 46716 9324
rect 46572 9036 46624 9042
rect 46572 8978 46624 8984
rect 46676 8974 46704 9318
rect 46952 9110 46980 11886
rect 47124 11756 47176 11762
rect 47124 11698 47176 11704
rect 47136 11150 47164 11698
rect 47124 11144 47176 11150
rect 47124 11086 47176 11092
rect 47032 11008 47084 11014
rect 47032 10950 47084 10956
rect 46940 9104 46992 9110
rect 46940 9046 46992 9052
rect 47044 8974 47072 10950
rect 47124 10668 47176 10674
rect 47124 10610 47176 10616
rect 47136 9994 47164 10610
rect 47124 9988 47176 9994
rect 47124 9930 47176 9936
rect 47124 9580 47176 9586
rect 47124 9522 47176 9528
rect 47136 9110 47164 9522
rect 47308 9444 47360 9450
rect 47308 9386 47360 9392
rect 47320 9110 47348 9386
rect 47124 9104 47176 9110
rect 47124 9046 47176 9052
rect 47308 9104 47360 9110
rect 47308 9046 47360 9052
rect 46664 8968 46716 8974
rect 46570 8936 46626 8945
rect 46492 8894 46570 8922
rect 46492 8498 46520 8894
rect 46664 8910 46716 8916
rect 47032 8968 47084 8974
rect 47032 8910 47084 8916
rect 46570 8871 46626 8880
rect 47504 8634 47532 12200
rect 47492 8628 47544 8634
rect 47492 8570 47544 8576
rect 47584 8628 47636 8634
rect 47584 8570 47636 8576
rect 47596 8514 47624 8570
rect 46480 8492 46532 8498
rect 46480 8434 46532 8440
rect 46676 8486 47624 8514
rect 46388 7880 46440 7886
rect 46110 7848 46166 7857
rect 46388 7822 46440 7828
rect 46110 7783 46166 7792
rect 46124 7698 46152 7783
rect 46386 7712 46442 7721
rect 46124 7670 46386 7698
rect 46386 7647 46442 7656
rect 46676 7002 46704 8486
rect 46756 8424 46808 8430
rect 46756 8366 46808 8372
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 46768 7410 46796 8366
rect 46756 7404 46808 7410
rect 46756 7346 46808 7352
rect 46768 7002 46796 7346
rect 46664 6996 46716 7002
rect 46664 6938 46716 6944
rect 46756 6996 46808 7002
rect 46756 6938 46808 6944
rect 45612 6820 45876 6848
rect 45560 6802 45612 6808
rect 45836 6656 45888 6662
rect 46480 6656 46532 6662
rect 45836 6598 45888 6604
rect 46110 6624 46166 6633
rect 45848 6254 45876 6598
rect 46480 6598 46532 6604
rect 46110 6559 46166 6568
rect 46124 6474 46152 6559
rect 46386 6488 46442 6497
rect 46124 6446 46386 6474
rect 46386 6423 46442 6432
rect 46492 6254 46520 6598
rect 46860 6338 46888 8366
rect 47872 8362 47900 12200
rect 48240 12050 48268 12200
rect 48502 12135 48558 12144
rect 48056 12022 48268 12050
rect 47952 9036 48004 9042
rect 47952 8978 48004 8984
rect 47860 8356 47912 8362
rect 47860 8298 47912 8304
rect 47492 8016 47544 8022
rect 47492 7958 47544 7964
rect 46940 7948 46992 7954
rect 46940 7890 46992 7896
rect 46952 7818 46980 7890
rect 46940 7812 46992 7818
rect 46940 7754 46992 7760
rect 47308 7744 47360 7750
rect 47308 7686 47360 7692
rect 46940 7404 46992 7410
rect 46940 7346 46992 7352
rect 46952 7206 46980 7346
rect 46940 7200 46992 7206
rect 46940 7142 46992 7148
rect 47032 7200 47084 7206
rect 47032 7142 47084 7148
rect 47044 6882 47072 7142
rect 47124 6996 47176 7002
rect 47124 6938 47176 6944
rect 46952 6854 47072 6882
rect 46952 6798 46980 6854
rect 46940 6792 46992 6798
rect 46940 6734 46992 6740
rect 46860 6310 46980 6338
rect 45468 6248 45520 6254
rect 45468 6190 45520 6196
rect 45652 6248 45704 6254
rect 45652 6190 45704 6196
rect 45836 6248 45888 6254
rect 45836 6190 45888 6196
rect 45928 6248 45980 6254
rect 45928 6190 45980 6196
rect 46480 6248 46532 6254
rect 46480 6190 46532 6196
rect 46848 6248 46900 6254
rect 46848 6190 46900 6196
rect 45664 5658 45692 6190
rect 45940 5914 45968 6190
rect 46032 6140 46336 6168
rect 46032 6089 46060 6140
rect 46018 6080 46074 6089
rect 46018 6015 46074 6024
rect 46202 6080 46258 6089
rect 46202 6015 46258 6024
rect 45928 5908 45980 5914
rect 45928 5850 45980 5856
rect 46216 5817 46244 6015
rect 46202 5808 46258 5817
rect 46308 5794 46336 6140
rect 46386 5808 46442 5817
rect 46308 5766 46386 5794
rect 46202 5743 46258 5752
rect 46386 5743 46442 5752
rect 46296 5704 46348 5710
rect 45940 5664 46296 5692
rect 45664 5630 45876 5658
rect 45848 5370 45876 5630
rect 45652 5364 45704 5370
rect 45388 5324 45508 5352
rect 45480 4128 45508 5324
rect 45652 5306 45704 5312
rect 45836 5364 45888 5370
rect 45836 5306 45888 5312
rect 45664 5250 45692 5306
rect 45940 5250 45968 5664
rect 46296 5646 46348 5652
rect 46860 5574 46888 6190
rect 46952 5692 46980 6310
rect 46952 5664 47072 5692
rect 46848 5568 46900 5574
rect 46032 5494 46520 5522
rect 46848 5510 46900 5516
rect 46032 5302 46060 5494
rect 46112 5364 46164 5370
rect 46112 5306 46164 5312
rect 45664 5222 45968 5250
rect 46020 5296 46072 5302
rect 46020 5238 46072 5244
rect 46124 4978 46152 5306
rect 46492 5284 46520 5494
rect 46664 5296 46716 5302
rect 46492 5256 46664 5284
rect 46664 5238 46716 5244
rect 46388 5228 46440 5234
rect 46440 5188 46612 5216
rect 46388 5170 46440 5176
rect 46204 5160 46256 5166
rect 46204 5102 46256 5108
rect 45664 4950 46152 4978
rect 45664 4690 45692 4950
rect 46216 4842 46244 5102
rect 45848 4814 46244 4842
rect 46388 4820 46440 4826
rect 45652 4684 45704 4690
rect 45652 4626 45704 4632
rect 45560 4616 45612 4622
rect 45848 4570 45876 4814
rect 46388 4762 46440 4768
rect 46584 4808 46612 5188
rect 47044 4808 47072 5664
rect 46584 4780 47072 4808
rect 46204 4752 46256 4758
rect 46256 4712 46336 4740
rect 46204 4694 46256 4700
rect 46112 4684 46164 4690
rect 45612 4564 45876 4570
rect 45560 4558 45876 4564
rect 45572 4542 45876 4558
rect 45940 4644 46112 4672
rect 45744 4480 45796 4486
rect 45796 4440 45876 4468
rect 45744 4422 45796 4428
rect 45388 4100 45508 4128
rect 45284 4004 45336 4010
rect 45284 3946 45336 3952
rect 45388 3346 45416 4100
rect 45848 4060 45876 4440
rect 45940 4214 45968 4644
rect 46112 4626 46164 4632
rect 46204 4548 46256 4554
rect 46204 4490 46256 4496
rect 46018 4448 46074 4457
rect 46018 4383 46074 4392
rect 46032 4214 46060 4383
rect 45928 4208 45980 4214
rect 45928 4150 45980 4156
rect 46020 4208 46072 4214
rect 46020 4150 46072 4156
rect 46216 4060 46244 4490
rect 45848 4032 46244 4060
rect 46308 4060 46336 4712
rect 46400 4690 46428 4762
rect 46584 4690 46612 4780
rect 46388 4684 46440 4690
rect 46388 4626 46440 4632
rect 46572 4684 46624 4690
rect 46572 4626 46624 4632
rect 46848 4684 46900 4690
rect 46848 4626 46900 4632
rect 46480 4616 46532 4622
rect 46386 4584 46442 4593
rect 46480 4558 46532 4564
rect 46386 4519 46442 4528
rect 46400 4185 46428 4519
rect 46492 4486 46520 4558
rect 46664 4548 46716 4554
rect 46584 4508 46664 4536
rect 46480 4480 46532 4486
rect 46480 4422 46532 4428
rect 46386 4176 46442 4185
rect 46386 4111 46442 4120
rect 46584 4060 46612 4508
rect 46664 4490 46716 4496
rect 46860 4185 46888 4626
rect 46846 4176 46902 4185
rect 46846 4111 46902 4120
rect 47030 4176 47086 4185
rect 47030 4111 47086 4120
rect 46308 4032 46612 4060
rect 45480 3998 45784 4026
rect 45480 3602 45508 3998
rect 45756 3992 45784 3998
rect 45756 3964 46796 3992
rect 45652 3936 45704 3942
rect 45652 3878 45704 3884
rect 45664 3754 45692 3878
rect 45664 3726 45876 3754
rect 45652 3664 45704 3670
rect 45652 3606 45704 3612
rect 45468 3596 45520 3602
rect 45468 3538 45520 3544
rect 45468 3460 45520 3466
rect 45664 3448 45692 3606
rect 45848 3534 45876 3726
rect 46296 3664 46348 3670
rect 46296 3606 46348 3612
rect 45836 3528 45888 3534
rect 45836 3470 45888 3476
rect 46112 3528 46164 3534
rect 46112 3470 46164 3476
rect 45520 3420 45692 3448
rect 45468 3402 45520 3408
rect 45388 3318 45600 3346
rect 45572 3058 45600 3318
rect 45560 3052 45612 3058
rect 45560 2994 45612 3000
rect 45744 3052 45796 3058
rect 45744 2994 45796 3000
rect 45374 2816 45430 2825
rect 45374 2751 45430 2760
rect 45388 2378 45416 2751
rect 45572 2650 45600 2994
rect 45652 2916 45704 2922
rect 45652 2858 45704 2864
rect 45560 2644 45612 2650
rect 45560 2586 45612 2592
rect 45376 2372 45428 2378
rect 45376 2314 45428 2320
rect 45468 1760 45520 1766
rect 45468 1702 45520 1708
rect 45376 1420 45428 1426
rect 45376 1362 45428 1368
rect 45388 746 45416 1362
rect 45480 800 45508 1702
rect 45664 1494 45692 2858
rect 45756 2446 45784 2994
rect 45836 2916 45888 2922
rect 45836 2858 45888 2864
rect 45848 2582 45876 2858
rect 45836 2576 45888 2582
rect 45836 2518 45888 2524
rect 45744 2440 45796 2446
rect 45744 2382 45796 2388
rect 46124 1970 46152 3470
rect 46308 3466 46336 3606
rect 46768 3534 46796 3964
rect 46756 3528 46808 3534
rect 46756 3470 46808 3476
rect 46204 3460 46256 3466
rect 46204 3402 46256 3408
rect 46296 3460 46348 3466
rect 46296 3402 46348 3408
rect 46216 3074 46244 3402
rect 46400 3318 46796 3346
rect 46296 3188 46348 3194
rect 46400 3176 46428 3318
rect 46348 3148 46428 3176
rect 46480 3188 46532 3194
rect 46296 3130 46348 3136
rect 46480 3130 46532 3136
rect 46664 3188 46716 3194
rect 46664 3130 46716 3136
rect 46216 3046 46428 3074
rect 46204 2644 46256 2650
rect 46204 2586 46256 2592
rect 46216 2446 46244 2586
rect 46296 2508 46348 2514
rect 46296 2450 46348 2456
rect 46204 2440 46256 2446
rect 46204 2382 46256 2388
rect 46112 1964 46164 1970
rect 46112 1906 46164 1912
rect 45652 1488 45704 1494
rect 45652 1430 45704 1436
rect 45652 1284 45704 1290
rect 45652 1226 45704 1232
rect 45836 1284 45888 1290
rect 45836 1226 45888 1232
rect 45664 882 45692 1226
rect 45652 876 45704 882
rect 45652 818 45704 824
rect 45848 800 45876 1226
rect 46308 882 46336 2450
rect 46400 2428 46428 3046
rect 46492 2650 46520 3130
rect 46572 2984 46624 2990
rect 46572 2926 46624 2932
rect 46584 2650 46612 2926
rect 46480 2644 46532 2650
rect 46480 2586 46532 2592
rect 46572 2644 46624 2650
rect 46572 2586 46624 2592
rect 46492 2530 46520 2586
rect 46492 2502 46612 2530
rect 46480 2440 46532 2446
rect 46400 2400 46480 2428
rect 46480 2382 46532 2388
rect 46480 1964 46532 1970
rect 46480 1906 46532 1912
rect 46492 1562 46520 1906
rect 46480 1556 46532 1562
rect 46480 1498 46532 1504
rect 46584 1426 46612 2502
rect 46480 1420 46532 1426
rect 46480 1362 46532 1368
rect 46572 1420 46624 1426
rect 46572 1362 46624 1368
rect 46492 1306 46520 1362
rect 46676 1306 46704 3130
rect 46768 1494 46796 3318
rect 46846 3224 46902 3233
rect 46846 3159 46902 3168
rect 46860 2378 46888 3159
rect 47044 2825 47072 4111
rect 47136 3194 47164 6938
rect 47320 6322 47348 7686
rect 47400 6792 47452 6798
rect 47400 6734 47452 6740
rect 47216 6316 47268 6322
rect 47216 6258 47268 6264
rect 47308 6316 47360 6322
rect 47308 6258 47360 6264
rect 47228 5574 47256 6258
rect 47412 5642 47440 6734
rect 47504 5778 47532 7958
rect 47584 7880 47636 7886
rect 47584 7822 47636 7828
rect 47596 7750 47624 7822
rect 47768 7812 47820 7818
rect 47768 7754 47820 7760
rect 47584 7744 47636 7750
rect 47584 7686 47636 7692
rect 47676 7744 47728 7750
rect 47676 7686 47728 7692
rect 47492 5772 47544 5778
rect 47492 5714 47544 5720
rect 47400 5636 47452 5642
rect 47400 5578 47452 5584
rect 47492 5636 47544 5642
rect 47492 5578 47544 5584
rect 47216 5568 47268 5574
rect 47216 5510 47268 5516
rect 47504 4146 47532 5578
rect 47492 4140 47544 4146
rect 47492 4082 47544 4088
rect 47596 3194 47624 7686
rect 47688 6458 47716 7686
rect 47780 7410 47808 7754
rect 47860 7472 47912 7478
rect 47860 7414 47912 7420
rect 47768 7404 47820 7410
rect 47768 7346 47820 7352
rect 47676 6452 47728 6458
rect 47676 6394 47728 6400
rect 47768 6452 47820 6458
rect 47768 6394 47820 6400
rect 47676 4684 47728 4690
rect 47780 4672 47808 6394
rect 47872 5778 47900 7414
rect 47860 5772 47912 5778
rect 47860 5714 47912 5720
rect 47728 4644 47808 4672
rect 47676 4626 47728 4632
rect 47964 4146 47992 8978
rect 48056 8838 48084 12022
rect 48228 11008 48280 11014
rect 48228 10950 48280 10956
rect 48240 10674 48268 10950
rect 48228 10668 48280 10674
rect 48228 10610 48280 10616
rect 48240 10266 48268 10610
rect 48608 10418 48636 12200
rect 48780 11280 48832 11286
rect 48780 11222 48832 11228
rect 48792 11150 48820 11222
rect 48688 11144 48740 11150
rect 48688 11086 48740 11092
rect 48780 11144 48832 11150
rect 48780 11086 48832 11092
rect 48332 10390 48636 10418
rect 48228 10260 48280 10266
rect 48228 10202 48280 10208
rect 48332 10146 48360 10390
rect 48596 10260 48648 10266
rect 48596 10202 48648 10208
rect 48240 10118 48360 10146
rect 48240 10062 48268 10118
rect 48228 10056 48280 10062
rect 48228 9998 48280 10004
rect 48412 10056 48464 10062
rect 48412 9998 48464 10004
rect 48320 9716 48372 9722
rect 48320 9658 48372 9664
rect 48332 9625 48360 9658
rect 48424 9654 48452 9998
rect 48412 9648 48464 9654
rect 48318 9616 48374 9625
rect 48412 9590 48464 9596
rect 48318 9551 48374 9560
rect 48320 9444 48372 9450
rect 48320 9386 48372 9392
rect 48136 8900 48188 8906
rect 48136 8842 48188 8848
rect 48228 8900 48280 8906
rect 48228 8842 48280 8848
rect 48044 8832 48096 8838
rect 48044 8774 48096 8780
rect 48148 7342 48176 8842
rect 48240 8634 48268 8842
rect 48228 8628 48280 8634
rect 48228 8570 48280 8576
rect 48332 8566 48360 9386
rect 48412 8832 48464 8838
rect 48412 8774 48464 8780
rect 48424 8566 48452 8774
rect 48504 8628 48556 8634
rect 48504 8570 48556 8576
rect 48320 8560 48372 8566
rect 48320 8502 48372 8508
rect 48412 8560 48464 8566
rect 48412 8502 48464 8508
rect 48412 8356 48464 8362
rect 48412 8298 48464 8304
rect 48136 7336 48188 7342
rect 48136 7278 48188 7284
rect 48136 6792 48188 6798
rect 48136 6734 48188 6740
rect 48148 6186 48176 6734
rect 48424 6304 48452 8298
rect 48516 7818 48544 8570
rect 48504 7812 48556 7818
rect 48504 7754 48556 7760
rect 48504 7472 48556 7478
rect 48504 7414 48556 7420
rect 48516 6662 48544 7414
rect 48504 6656 48556 6662
rect 48504 6598 48556 6604
rect 48424 6276 48544 6304
rect 48044 6180 48096 6186
rect 48044 6122 48096 6128
rect 48136 6180 48188 6186
rect 48136 6122 48188 6128
rect 48056 6066 48084 6122
rect 48056 6038 48360 6066
rect 48044 5228 48096 5234
rect 48044 5170 48096 5176
rect 48056 4554 48084 5170
rect 48044 4548 48096 4554
rect 48044 4490 48096 4496
rect 48228 4548 48280 4554
rect 48228 4490 48280 4496
rect 48240 4282 48268 4490
rect 48228 4276 48280 4282
rect 48228 4218 48280 4224
rect 47952 4140 48004 4146
rect 48228 4140 48280 4146
rect 48004 4100 48084 4128
rect 47952 4082 48004 4088
rect 47688 3998 47992 4026
rect 47688 3738 47716 3998
rect 47964 3942 47992 3998
rect 47768 3936 47820 3942
rect 47952 3936 48004 3942
rect 47820 3896 47900 3924
rect 47768 3878 47820 3884
rect 47676 3732 47728 3738
rect 47676 3674 47728 3680
rect 47124 3188 47176 3194
rect 47124 3130 47176 3136
rect 47584 3188 47636 3194
rect 47584 3130 47636 3136
rect 47216 3052 47268 3058
rect 47216 2994 47268 3000
rect 47584 3052 47636 3058
rect 47584 2994 47636 3000
rect 47228 2825 47256 2994
rect 47030 2816 47086 2825
rect 47030 2751 47086 2760
rect 47214 2816 47270 2825
rect 47214 2751 47270 2760
rect 47228 2650 47256 2751
rect 47032 2644 47084 2650
rect 47032 2586 47084 2592
rect 47216 2644 47268 2650
rect 47216 2586 47268 2592
rect 46848 2372 46900 2378
rect 46848 2314 46900 2320
rect 46848 1964 46900 1970
rect 46848 1906 46900 1912
rect 46756 1488 46808 1494
rect 46756 1430 46808 1436
rect 46492 1278 46704 1306
rect 46860 1034 46888 1906
rect 46940 1352 46992 1358
rect 46940 1294 46992 1300
rect 46584 1006 46888 1034
rect 46386 912 46442 921
rect 46296 876 46348 882
rect 46124 836 46244 864
rect 45376 740 45428 746
rect 45376 682 45428 688
rect 45190 504 45246 513
rect 45190 439 45246 448
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46124 746 46152 836
rect 46216 800 46244 836
rect 46386 847 46442 856
rect 46296 818 46348 824
rect 46112 740 46164 746
rect 46112 682 46164 688
rect 46202 0 46258 800
rect 46400 649 46428 847
rect 46584 800 46612 1006
rect 46952 800 46980 1294
rect 47044 921 47072 2586
rect 47596 2378 47624 2994
rect 47768 2644 47820 2650
rect 47768 2586 47820 2592
rect 47124 2372 47176 2378
rect 47124 2314 47176 2320
rect 47584 2372 47636 2378
rect 47584 2314 47636 2320
rect 47136 1193 47164 2314
rect 47308 2100 47360 2106
rect 47308 2042 47360 2048
rect 47584 2100 47636 2106
rect 47584 2042 47636 2048
rect 47216 2032 47268 2038
rect 47216 1974 47268 1980
rect 47228 1578 47256 1974
rect 47320 1748 47348 2042
rect 47596 1970 47624 2042
rect 47676 2032 47728 2038
rect 47676 1974 47728 1980
rect 47584 1964 47636 1970
rect 47584 1906 47636 1912
rect 47492 1760 47544 1766
rect 47320 1720 47492 1748
rect 47492 1702 47544 1708
rect 47688 1578 47716 1974
rect 47228 1550 47716 1578
rect 47780 1408 47808 2586
rect 47228 1380 47808 1408
rect 47122 1184 47178 1193
rect 47122 1119 47178 1128
rect 47228 1018 47256 1380
rect 47320 1290 47716 1306
rect 47308 1284 47716 1290
rect 47360 1278 47716 1284
rect 47688 1272 47716 1278
rect 47768 1284 47820 1290
rect 47688 1244 47768 1272
rect 47308 1226 47360 1232
rect 47768 1226 47820 1232
rect 47584 1216 47636 1222
rect 47306 1184 47362 1193
rect 47584 1158 47636 1164
rect 47306 1119 47362 1128
rect 47216 1012 47268 1018
rect 47216 954 47268 960
rect 47030 912 47086 921
rect 47030 847 47086 856
rect 47320 800 47348 1119
rect 47400 808 47452 814
rect 46386 640 46442 649
rect 46386 575 46442 584
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47400 750 47452 756
rect 47412 134 47440 750
rect 47596 134 47624 1158
rect 47872 1018 47900 3896
rect 47952 3878 48004 3884
rect 48056 3738 48084 4100
rect 48228 4082 48280 4088
rect 48044 3732 48096 3738
rect 48044 3674 48096 3680
rect 48136 3732 48188 3738
rect 48136 3674 48188 3680
rect 48148 3210 48176 3674
rect 47964 3182 48176 3210
rect 47860 1012 47912 1018
rect 47860 954 47912 960
rect 47964 898 47992 3182
rect 48044 3120 48096 3126
rect 48044 3062 48096 3068
rect 47688 870 47992 898
rect 47688 800 47716 870
rect 48056 800 48084 3062
rect 48240 3058 48268 4082
rect 48228 3052 48280 3058
rect 48228 2994 48280 3000
rect 48136 1964 48188 1970
rect 48136 1906 48188 1912
rect 47400 128 47452 134
rect 47400 70 47452 76
rect 47584 128 47636 134
rect 47584 70 47636 76
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48148 134 48176 1906
rect 48332 513 48360 6038
rect 48516 5234 48544 6276
rect 48608 5914 48636 10202
rect 48700 9625 48728 11086
rect 48976 10690 49004 12200
rect 49148 11756 49200 11762
rect 49148 11698 49200 11704
rect 49160 11286 49188 11698
rect 49240 11688 49292 11694
rect 49240 11630 49292 11636
rect 49252 11286 49280 11630
rect 49148 11280 49200 11286
rect 49148 11222 49200 11228
rect 49240 11280 49292 11286
rect 49240 11222 49292 11228
rect 48792 10662 49004 10690
rect 49238 10704 49294 10713
rect 48686 9616 48742 9625
rect 48686 9551 48742 9560
rect 48688 8900 48740 8906
rect 48688 8842 48740 8848
rect 48700 6882 48728 8842
rect 48792 8498 48820 10662
rect 49238 10639 49294 10648
rect 48964 10600 49016 10606
rect 48964 10542 49016 10548
rect 49056 10600 49108 10606
rect 49056 10542 49108 10548
rect 48976 10198 49004 10542
rect 48964 10192 49016 10198
rect 48964 10134 49016 10140
rect 49068 9042 49096 10542
rect 49056 9036 49108 9042
rect 49056 8978 49108 8984
rect 48780 8492 48832 8498
rect 48780 8434 48832 8440
rect 48872 8016 48924 8022
rect 48924 7976 49004 8004
rect 48872 7958 48924 7964
rect 48780 7880 48832 7886
rect 48832 7840 48912 7868
rect 48780 7822 48832 7828
rect 48884 7478 48912 7840
rect 48872 7472 48924 7478
rect 48872 7414 48924 7420
rect 48872 7336 48924 7342
rect 48872 7278 48924 7284
rect 48884 7002 48912 7278
rect 48976 7002 49004 7976
rect 49056 7948 49108 7954
rect 49056 7890 49108 7896
rect 48872 6996 48924 7002
rect 48872 6938 48924 6944
rect 48964 6996 49016 7002
rect 48964 6938 49016 6944
rect 48700 6854 48820 6882
rect 48596 5908 48648 5914
rect 48596 5850 48648 5856
rect 48504 5228 48556 5234
rect 48504 5170 48556 5176
rect 48596 4208 48648 4214
rect 48596 4150 48648 4156
rect 48504 3936 48556 3942
rect 48504 3878 48556 3884
rect 48412 3392 48464 3398
rect 48412 3334 48464 3340
rect 48424 2514 48452 3334
rect 48412 2508 48464 2514
rect 48412 2450 48464 2456
rect 48516 1748 48544 3878
rect 48608 3466 48636 4150
rect 48596 3460 48648 3466
rect 48596 3402 48648 3408
rect 48792 3058 48820 6854
rect 49068 4978 49096 7890
rect 48884 4950 49096 4978
rect 48884 3534 48912 4950
rect 48964 4616 49016 4622
rect 49252 4604 49280 10639
rect 49344 8634 49372 12200
rect 49712 11880 49740 12200
rect 49528 11852 49740 11880
rect 49424 11688 49476 11694
rect 49424 11630 49476 11636
rect 49436 11150 49464 11630
rect 49424 11144 49476 11150
rect 49424 11086 49476 11092
rect 49528 9518 49556 11852
rect 49608 11756 49660 11762
rect 49608 11698 49660 11704
rect 49792 11756 49844 11762
rect 49792 11698 49844 11704
rect 49620 11082 49648 11698
rect 49700 11688 49752 11694
rect 49700 11630 49752 11636
rect 49712 11150 49740 11630
rect 49700 11144 49752 11150
rect 49700 11086 49752 11092
rect 49608 11076 49660 11082
rect 49608 11018 49660 11024
rect 49700 10668 49752 10674
rect 49700 10610 49752 10616
rect 49712 10198 49740 10610
rect 49804 10470 49832 11698
rect 49792 10464 49844 10470
rect 49792 10406 49844 10412
rect 49976 10464 50028 10470
rect 49976 10406 50028 10412
rect 49700 10192 49752 10198
rect 49700 10134 49752 10140
rect 49884 10192 49936 10198
rect 49884 10134 49936 10140
rect 49516 9512 49568 9518
rect 49516 9454 49568 9460
rect 49790 8800 49846 8809
rect 49790 8735 49846 8744
rect 49804 8634 49832 8735
rect 49332 8628 49384 8634
rect 49332 8570 49384 8576
rect 49792 8628 49844 8634
rect 49792 8570 49844 8576
rect 49896 8430 49924 10134
rect 49988 10062 50016 10406
rect 49976 10056 50028 10062
rect 49976 9998 50028 10004
rect 49988 9722 50016 9998
rect 49976 9716 50028 9722
rect 49976 9658 50028 9664
rect 49976 8560 50028 8566
rect 49976 8502 50028 8508
rect 49884 8424 49936 8430
rect 49884 8366 49936 8372
rect 49988 8090 50016 8502
rect 49792 8084 49844 8090
rect 49792 8026 49844 8032
rect 49976 8084 50028 8090
rect 49976 8026 50028 8032
rect 49516 7948 49568 7954
rect 49516 7890 49568 7896
rect 49528 7818 49556 7890
rect 49516 7812 49568 7818
rect 49516 7754 49568 7760
rect 49608 7812 49660 7818
rect 49608 7754 49660 7760
rect 49332 5160 49384 5166
rect 49332 5102 49384 5108
rect 49344 4758 49372 5102
rect 49332 4752 49384 4758
rect 49332 4694 49384 4700
rect 49016 4576 49280 4604
rect 48964 4558 49016 4564
rect 49252 4486 49280 4576
rect 49240 4480 49292 4486
rect 49240 4422 49292 4428
rect 49620 4146 49648 7754
rect 49804 7478 49832 8026
rect 50080 8022 50108 12200
rect 50160 11552 50212 11558
rect 50160 11494 50212 11500
rect 50252 11552 50304 11558
rect 50252 11494 50304 11500
rect 50172 11082 50200 11494
rect 50264 11150 50292 11494
rect 50252 11144 50304 11150
rect 50252 11086 50304 11092
rect 50160 11076 50212 11082
rect 50160 11018 50212 11024
rect 50342 10704 50398 10713
rect 50342 10639 50398 10648
rect 50160 10464 50212 10470
rect 50160 10406 50212 10412
rect 50172 9654 50200 10406
rect 50356 9994 50384 10639
rect 50252 9988 50304 9994
rect 50252 9930 50304 9936
rect 50344 9988 50396 9994
rect 50344 9930 50396 9936
rect 50264 9722 50292 9930
rect 50252 9716 50304 9722
rect 50252 9658 50304 9664
rect 50160 9648 50212 9654
rect 50160 9590 50212 9596
rect 50448 9382 50476 12200
rect 50618 12135 50674 12144
rect 50528 11144 50580 11150
rect 50528 11086 50580 11092
rect 50540 9586 50568 11086
rect 50632 10674 50660 12135
rect 50724 11937 50752 12446
rect 50802 12200 50858 13000
rect 50894 12951 50896 12960
rect 50948 12951 50950 12960
rect 50896 12922 50948 12928
rect 50894 12472 50950 12481
rect 50894 12407 50950 12416
rect 50710 11928 50766 11937
rect 50710 11863 50766 11872
rect 50712 11688 50764 11694
rect 50712 11630 50764 11636
rect 50724 11150 50752 11630
rect 50712 11144 50764 11150
rect 50712 11086 50764 11092
rect 50620 10668 50672 10674
rect 50620 10610 50672 10616
rect 50712 10668 50764 10674
rect 50712 10610 50764 10616
rect 50724 9926 50752 10610
rect 50816 10266 50844 12200
rect 50804 10260 50856 10266
rect 50804 10202 50856 10208
rect 50908 10146 50936 12407
rect 51170 12200 51226 13000
rect 51354 12608 51410 12617
rect 51354 12543 51410 12552
rect 51262 12200 51318 12209
rect 51184 11694 51212 12200
rect 51262 12135 51318 12144
rect 51368 12152 51396 12543
rect 51538 12200 51594 13000
rect 51906 12200 51962 13000
rect 52274 12200 52330 13000
rect 52642 12200 52698 13000
rect 53010 12200 53066 13000
rect 53104 12232 53156 12238
rect 51552 12152 51580 12200
rect 51172 11688 51224 11694
rect 51172 11630 51224 11636
rect 51080 11280 51132 11286
rect 51080 11222 51132 11228
rect 50988 11144 51040 11150
rect 51092 11132 51120 11222
rect 51040 11104 51120 11132
rect 50988 11086 51040 11092
rect 51276 10810 51304 12135
rect 51368 12124 51580 12152
rect 51920 12073 51948 12200
rect 51906 12064 51962 12073
rect 51906 11999 51962 12008
rect 51816 11688 51868 11694
rect 51816 11630 51868 11636
rect 51448 11008 51500 11014
rect 51448 10950 51500 10956
rect 51540 11008 51592 11014
rect 51540 10950 51592 10956
rect 51172 10804 51224 10810
rect 51172 10746 51224 10752
rect 51264 10804 51316 10810
rect 51264 10746 51316 10752
rect 50988 10260 51040 10266
rect 50988 10202 51040 10208
rect 50816 10118 50936 10146
rect 50620 9920 50672 9926
rect 50620 9862 50672 9868
rect 50712 9920 50764 9926
rect 50712 9862 50764 9868
rect 50528 9580 50580 9586
rect 50528 9522 50580 9528
rect 50632 9518 50660 9862
rect 50620 9512 50672 9518
rect 50620 9454 50672 9460
rect 50436 9376 50488 9382
rect 50436 9318 50488 9324
rect 50618 9208 50674 9217
rect 50618 9143 50674 9152
rect 50632 8888 50660 9143
rect 50724 9042 50752 9862
rect 50816 9217 50844 10118
rect 50896 10056 50948 10062
rect 51000 10044 51028 10202
rect 50948 10016 51028 10044
rect 50896 9998 50948 10004
rect 51184 9654 51212 10746
rect 51460 10742 51488 10950
rect 51448 10736 51500 10742
rect 51448 10678 51500 10684
rect 51448 10464 51500 10470
rect 51448 10406 51500 10412
rect 51264 10192 51316 10198
rect 51264 10134 51316 10140
rect 51172 9648 51224 9654
rect 51172 9590 51224 9596
rect 51276 9586 51304 10134
rect 51460 10112 51488 10406
rect 51552 10266 51580 10950
rect 51828 10674 51856 11630
rect 52184 11552 52236 11558
rect 52184 11494 52236 11500
rect 51724 10668 51776 10674
rect 51724 10610 51776 10616
rect 51816 10668 51868 10674
rect 51816 10610 51868 10616
rect 51632 10464 51684 10470
rect 51632 10406 51684 10412
rect 51540 10260 51592 10266
rect 51540 10202 51592 10208
rect 51460 10084 51580 10112
rect 51552 9908 51580 10084
rect 51644 10062 51672 10406
rect 51736 10266 51764 10610
rect 51724 10260 51776 10266
rect 51724 10202 51776 10208
rect 51632 10056 51684 10062
rect 51684 10016 51764 10044
rect 51632 9998 51684 10004
rect 51552 9880 51672 9908
rect 51356 9716 51408 9722
rect 51356 9658 51408 9664
rect 51368 9602 51396 9658
rect 51080 9580 51132 9586
rect 51080 9522 51132 9528
rect 51264 9580 51316 9586
rect 51368 9574 51580 9602
rect 51264 9522 51316 9528
rect 50802 9208 50858 9217
rect 50802 9143 50858 9152
rect 50712 9036 50764 9042
rect 50712 8978 50764 8984
rect 50632 8860 50936 8888
rect 50160 8832 50212 8838
rect 50160 8774 50212 8780
rect 50528 8832 50580 8838
rect 50528 8774 50580 8780
rect 50172 8430 50200 8774
rect 50252 8628 50304 8634
rect 50252 8570 50304 8576
rect 50160 8424 50212 8430
rect 50160 8366 50212 8372
rect 50160 8084 50212 8090
rect 50160 8026 50212 8032
rect 50068 8016 50120 8022
rect 50068 7958 50120 7964
rect 49976 7880 50028 7886
rect 49976 7822 50028 7828
rect 49988 7562 50016 7822
rect 50172 7750 50200 8026
rect 50264 8022 50292 8570
rect 50540 8294 50568 8774
rect 50908 8378 50936 8860
rect 50986 8392 51042 8401
rect 50712 8356 50764 8362
rect 50908 8350 50986 8378
rect 50986 8327 51042 8336
rect 50712 8298 50764 8304
rect 50528 8288 50580 8294
rect 50528 8230 50580 8236
rect 50252 8016 50304 8022
rect 50252 7958 50304 7964
rect 50540 7886 50568 8230
rect 50528 7880 50580 7886
rect 50528 7822 50580 7828
rect 50160 7744 50212 7750
rect 50160 7686 50212 7692
rect 50252 7744 50304 7750
rect 50252 7686 50304 7692
rect 50264 7562 50292 7686
rect 49988 7534 50292 7562
rect 49792 7472 49844 7478
rect 49792 7414 49844 7420
rect 50264 7126 50660 7154
rect 50264 7002 50292 7126
rect 50252 6996 50304 7002
rect 50252 6938 50304 6944
rect 50344 6996 50396 7002
rect 50344 6938 50396 6944
rect 49792 6792 49844 6798
rect 49792 6734 49844 6740
rect 49804 5914 49832 6734
rect 50160 6316 50212 6322
rect 50160 6258 50212 6264
rect 49792 5908 49844 5914
rect 49792 5850 49844 5856
rect 50068 5704 50120 5710
rect 50068 5646 50120 5652
rect 49700 5228 49752 5234
rect 49700 5170 49752 5176
rect 49712 4826 49740 5170
rect 50080 4826 50108 5646
rect 49700 4820 49752 4826
rect 49700 4762 49752 4768
rect 50068 4820 50120 4826
rect 50068 4762 50120 4768
rect 49976 4480 50028 4486
rect 49976 4422 50028 4428
rect 49988 4282 50016 4422
rect 49976 4276 50028 4282
rect 49976 4218 50028 4224
rect 49792 4208 49844 4214
rect 49844 4168 49924 4196
rect 49792 4150 49844 4156
rect 49608 4140 49660 4146
rect 49608 4082 49660 4088
rect 49700 4140 49752 4146
rect 49700 4082 49752 4088
rect 49424 4004 49476 4010
rect 49424 3946 49476 3952
rect 49436 3670 49464 3946
rect 49620 3738 49648 4082
rect 49608 3732 49660 3738
rect 49608 3674 49660 3680
rect 49424 3664 49476 3670
rect 49424 3606 49476 3612
rect 48872 3528 48924 3534
rect 48872 3470 48924 3476
rect 48964 3460 49016 3466
rect 49016 3420 49188 3448
rect 48964 3402 49016 3408
rect 49160 3058 49188 3420
rect 49332 3188 49384 3194
rect 49332 3130 49384 3136
rect 49516 3188 49568 3194
rect 49516 3130 49568 3136
rect 48780 3052 48832 3058
rect 48780 2994 48832 3000
rect 49056 3052 49108 3058
rect 49056 2994 49108 3000
rect 49148 3052 49200 3058
rect 49148 2994 49200 3000
rect 48964 2848 49016 2854
rect 48964 2790 49016 2796
rect 48872 2644 48924 2650
rect 48976 2632 49004 2790
rect 49068 2650 49096 2994
rect 49344 2990 49372 3130
rect 49332 2984 49384 2990
rect 49332 2926 49384 2932
rect 49148 2916 49200 2922
rect 49148 2858 49200 2864
rect 49160 2650 49188 2858
rect 48924 2604 49004 2632
rect 49056 2644 49108 2650
rect 48872 2586 48924 2592
rect 49056 2586 49108 2592
rect 49148 2644 49200 2650
rect 49148 2586 49200 2592
rect 48596 2440 48648 2446
rect 48596 2382 48648 2388
rect 48424 1720 48544 1748
rect 48424 800 48452 1720
rect 48608 1562 48636 2382
rect 49056 2100 49108 2106
rect 49056 2042 49108 2048
rect 48688 1964 48740 1970
rect 48688 1906 48740 1912
rect 48700 1562 48728 1906
rect 49068 1766 49096 2042
rect 49424 2032 49476 2038
rect 49424 1974 49476 1980
rect 49056 1760 49108 1766
rect 49056 1702 49108 1708
rect 49148 1760 49200 1766
rect 49148 1702 49200 1708
rect 48596 1556 48648 1562
rect 48596 1498 48648 1504
rect 48688 1556 48740 1562
rect 48688 1498 48740 1504
rect 48780 1352 48832 1358
rect 49056 1352 49108 1358
rect 48832 1312 49056 1340
rect 48780 1294 48832 1300
rect 49056 1294 49108 1300
rect 48792 836 48912 864
rect 48792 800 48820 836
rect 48318 504 48374 513
rect 48318 439 48374 448
rect 48136 128 48188 134
rect 48136 70 48188 76
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 48884 728 48912 836
rect 49160 800 49188 1702
rect 49436 882 49464 1974
rect 49424 876 49476 882
rect 49424 818 49476 824
rect 49528 800 49556 3130
rect 49608 1012 49660 1018
rect 49608 954 49660 960
rect 49056 740 49108 746
rect 48884 700 49056 728
rect 49056 682 49108 688
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49620 626 49648 954
rect 49712 746 49740 4082
rect 49896 3992 49924 4168
rect 50068 4004 50120 4010
rect 49896 3964 50068 3992
rect 50068 3946 50120 3952
rect 50172 3738 50200 6258
rect 50356 4842 50384 6938
rect 50632 6730 50660 7126
rect 50724 6934 50752 8298
rect 51092 8294 51120 9522
rect 51356 9444 51408 9450
rect 51276 9404 51356 9432
rect 51080 8288 51132 8294
rect 51080 8230 51132 8236
rect 50908 7772 51212 7800
rect 50804 7744 50856 7750
rect 50804 7686 50856 7692
rect 50816 7478 50844 7686
rect 50908 7585 50936 7772
rect 51184 7721 51212 7772
rect 51170 7712 51226 7721
rect 51170 7647 51226 7656
rect 50894 7576 50950 7585
rect 50894 7511 50950 7520
rect 50804 7472 50856 7478
rect 50804 7414 50856 7420
rect 51276 7256 51304 9404
rect 51356 9386 51408 9392
rect 51552 8906 51580 9574
rect 51644 9518 51672 9880
rect 51632 9512 51684 9518
rect 51632 9454 51684 9460
rect 51632 9376 51684 9382
rect 51632 9318 51684 9324
rect 51644 9178 51672 9318
rect 51632 9172 51684 9178
rect 51632 9114 51684 9120
rect 51540 8900 51592 8906
rect 51540 8842 51592 8848
rect 51736 8786 51764 10016
rect 52196 9654 52224 11494
rect 52092 9648 52144 9654
rect 52092 9590 52144 9596
rect 52184 9648 52236 9654
rect 52184 9590 52236 9596
rect 52104 8974 52132 9590
rect 52288 9382 52316 12200
rect 52460 11552 52512 11558
rect 52460 11494 52512 11500
rect 52472 11150 52500 11494
rect 52460 11144 52512 11150
rect 52460 11086 52512 11092
rect 52368 10668 52420 10674
rect 52368 10610 52420 10616
rect 52380 10266 52408 10610
rect 52368 10260 52420 10266
rect 52368 10202 52420 10208
rect 52472 9636 52500 11086
rect 52472 9608 52592 9636
rect 52276 9376 52328 9382
rect 52276 9318 52328 9324
rect 52460 9376 52512 9382
rect 52460 9318 52512 9324
rect 52472 9217 52500 9318
rect 52458 9208 52514 9217
rect 52458 9143 52514 9152
rect 52092 8968 52144 8974
rect 52092 8910 52144 8916
rect 51552 8758 51764 8786
rect 52368 8832 52420 8838
rect 52368 8774 52420 8780
rect 51552 8634 51580 8758
rect 51540 8628 51592 8634
rect 51540 8570 51592 8576
rect 51724 8628 51776 8634
rect 51724 8570 51776 8576
rect 51368 8362 51672 8378
rect 51368 8356 51684 8362
rect 51368 8350 51632 8356
rect 51368 7886 51396 8350
rect 51632 8298 51684 8304
rect 51736 7970 51764 8570
rect 52380 8566 52408 8774
rect 52368 8560 52420 8566
rect 52368 8502 52420 8508
rect 52000 8492 52052 8498
rect 52000 8434 52052 8440
rect 51816 8288 51868 8294
rect 51816 8230 51868 8236
rect 51908 8288 51960 8294
rect 51908 8230 51960 8236
rect 51552 7942 51764 7970
rect 51552 7886 51580 7942
rect 51356 7880 51408 7886
rect 51356 7822 51408 7828
rect 51540 7880 51592 7886
rect 51540 7822 51592 7828
rect 51724 7880 51776 7886
rect 51724 7822 51776 7828
rect 51448 7472 51500 7478
rect 51552 7460 51580 7822
rect 51500 7432 51580 7460
rect 51632 7472 51684 7478
rect 51448 7414 51500 7420
rect 51632 7414 51684 7420
rect 51092 7228 51304 7256
rect 50712 6928 50764 6934
rect 50712 6870 50764 6876
rect 50896 6928 50948 6934
rect 50896 6870 50948 6876
rect 50528 6724 50580 6730
rect 50528 6666 50580 6672
rect 50620 6724 50672 6730
rect 50620 6666 50672 6672
rect 50264 4814 50384 4842
rect 50540 4826 50568 6666
rect 50712 6452 50764 6458
rect 50712 6394 50764 6400
rect 50804 6452 50856 6458
rect 50804 6394 50856 6400
rect 50724 6322 50752 6394
rect 50712 6316 50764 6322
rect 50712 6258 50764 6264
rect 50712 6180 50764 6186
rect 50816 6168 50844 6394
rect 50764 6140 50844 6168
rect 50712 6122 50764 6128
rect 50908 5817 50936 6870
rect 51092 5914 51120 7228
rect 51644 7154 51672 7414
rect 51276 7126 51672 7154
rect 51276 6798 51304 7126
rect 51448 6996 51500 7002
rect 51448 6938 51500 6944
rect 51460 6905 51488 6938
rect 51446 6896 51502 6905
rect 51446 6831 51502 6840
rect 51264 6792 51316 6798
rect 51264 6734 51316 6740
rect 51448 6724 51500 6730
rect 51500 6684 51672 6712
rect 51448 6666 51500 6672
rect 51276 6582 51580 6610
rect 51276 6458 51304 6582
rect 51264 6452 51316 6458
rect 51264 6394 51316 6400
rect 51448 6452 51500 6458
rect 51448 6394 51500 6400
rect 51172 6316 51224 6322
rect 51172 6258 51224 6264
rect 51080 5908 51132 5914
rect 51080 5850 51132 5856
rect 50894 5808 50950 5817
rect 50894 5743 50950 5752
rect 51078 5808 51134 5817
rect 51184 5778 51212 6258
rect 51460 6186 51488 6394
rect 51448 6180 51500 6186
rect 51448 6122 51500 6128
rect 51264 6112 51316 6118
rect 51264 6054 51316 6060
rect 51356 6112 51408 6118
rect 51356 6054 51408 6060
rect 51276 5914 51304 6054
rect 51264 5908 51316 5914
rect 51264 5850 51316 5856
rect 51078 5743 51134 5752
rect 51172 5772 51224 5778
rect 51092 5370 51120 5743
rect 51172 5714 51224 5720
rect 51368 5556 51396 6054
rect 51184 5528 51396 5556
rect 51080 5364 51132 5370
rect 51080 5306 51132 5312
rect 51184 5250 51212 5528
rect 51356 5364 51408 5370
rect 51356 5306 51408 5312
rect 51000 5222 51212 5250
rect 51000 5030 51028 5222
rect 51368 5137 51396 5306
rect 51354 5128 51410 5137
rect 51354 5063 51410 5072
rect 50988 5024 51040 5030
rect 51264 5024 51316 5030
rect 50988 4966 51040 4972
rect 51184 4972 51264 4978
rect 51184 4966 51316 4972
rect 51184 4950 51304 4966
rect 50528 4820 50580 4826
rect 50160 3732 50212 3738
rect 50160 3674 50212 3680
rect 50264 2446 50292 4814
rect 50528 4762 50580 4768
rect 51184 4536 51212 4950
rect 51000 4508 51212 4536
rect 50620 4480 50672 4486
rect 50620 4422 50672 4428
rect 50632 2514 50660 4422
rect 51000 3890 51028 4508
rect 51552 4214 51580 6582
rect 51644 6322 51672 6684
rect 51632 6316 51684 6322
rect 51632 6258 51684 6264
rect 51632 4480 51684 4486
rect 51632 4422 51684 4428
rect 51264 4208 51316 4214
rect 51262 4176 51264 4185
rect 51540 4208 51592 4214
rect 51316 4176 51318 4185
rect 51540 4150 51592 4156
rect 51644 4146 51672 4422
rect 51262 4111 51318 4120
rect 51632 4140 51684 4146
rect 51632 4082 51684 4088
rect 51448 4072 51500 4078
rect 51500 4032 51580 4060
rect 51448 4014 51500 4020
rect 50816 3862 51028 3890
rect 50816 3233 50844 3862
rect 50894 3768 50950 3777
rect 50894 3703 50950 3712
rect 50802 3224 50858 3233
rect 50802 3159 50858 3168
rect 50712 3052 50764 3058
rect 50712 2994 50764 3000
rect 50804 3052 50856 3058
rect 50804 2994 50856 3000
rect 50724 2514 50752 2994
rect 50816 2650 50844 2994
rect 50908 2650 50936 3703
rect 51080 3596 51132 3602
rect 51080 3538 51132 3544
rect 51092 3482 51120 3538
rect 51552 3516 51580 4032
rect 51736 3738 51764 7822
rect 51828 5137 51856 8230
rect 51920 8090 51948 8230
rect 51908 8084 51960 8090
rect 51908 8026 51960 8032
rect 52012 7478 52040 8434
rect 52368 8424 52420 8430
rect 52368 8366 52420 8372
rect 52184 8356 52236 8362
rect 52184 8298 52236 8304
rect 52092 7880 52144 7886
rect 52092 7822 52144 7828
rect 52000 7472 52052 7478
rect 52000 7414 52052 7420
rect 52104 7206 52132 7822
rect 51908 7200 51960 7206
rect 51908 7142 51960 7148
rect 52092 7200 52144 7206
rect 52092 7142 52144 7148
rect 51920 6746 51948 7142
rect 52196 6866 52224 8298
rect 52276 7880 52328 7886
rect 52276 7822 52328 7828
rect 52288 7750 52316 7822
rect 52380 7750 52408 8366
rect 52276 7744 52328 7750
rect 52276 7686 52328 7692
rect 52368 7744 52420 7750
rect 52368 7686 52420 7692
rect 52460 6996 52512 7002
rect 52460 6938 52512 6944
rect 52184 6860 52236 6866
rect 52184 6802 52236 6808
rect 52276 6860 52328 6866
rect 52276 6802 52328 6808
rect 52288 6746 52316 6802
rect 51920 6718 52316 6746
rect 52368 6656 52420 6662
rect 51906 6624 51962 6633
rect 52472 6633 52500 6938
rect 52368 6598 52420 6604
rect 52458 6624 52514 6633
rect 51906 6559 51962 6568
rect 51920 6254 51948 6559
rect 52380 6458 52408 6598
rect 52458 6559 52514 6568
rect 52564 6474 52592 9608
rect 52656 8634 52684 12200
rect 52736 11756 52788 11762
rect 52736 11698 52788 11704
rect 52748 10985 52776 11698
rect 53024 11014 53052 12200
rect 53378 12200 53434 13000
rect 53746 12200 53802 13000
rect 54114 12200 54170 13000
rect 54482 12200 54538 13000
rect 54574 12200 54630 12209
rect 54850 12200 54906 13000
rect 55218 12200 55274 13000
rect 55404 12232 55456 12238
rect 53104 12174 53156 12180
rect 53116 11558 53144 12174
rect 53194 11928 53250 11937
rect 53194 11863 53250 11872
rect 53208 11558 53236 11863
rect 53104 11552 53156 11558
rect 53104 11494 53156 11500
rect 53196 11552 53248 11558
rect 53196 11494 53248 11500
rect 53012 11008 53064 11014
rect 52734 10976 52790 10985
rect 53012 10950 53064 10956
rect 52734 10911 52790 10920
rect 52828 10464 52880 10470
rect 52828 10406 52880 10412
rect 52644 8628 52696 8634
rect 52644 8570 52696 8576
rect 52736 8492 52788 8498
rect 52736 8434 52788 8440
rect 52748 8090 52776 8434
rect 52736 8084 52788 8090
rect 52736 8026 52788 8032
rect 52736 7472 52788 7478
rect 52736 7414 52788 7420
rect 52748 7002 52776 7414
rect 52736 6996 52788 7002
rect 52736 6938 52788 6944
rect 52564 6458 52776 6474
rect 52368 6452 52420 6458
rect 52564 6452 52788 6458
rect 52564 6446 52736 6452
rect 52368 6394 52420 6400
rect 52736 6394 52788 6400
rect 52276 6384 52328 6390
rect 52276 6326 52328 6332
rect 51908 6248 51960 6254
rect 52288 6236 52316 6326
rect 52460 6316 52512 6322
rect 52644 6316 52696 6322
rect 52512 6276 52592 6304
rect 52460 6258 52512 6264
rect 52368 6248 52420 6254
rect 52288 6208 52368 6236
rect 51908 6190 51960 6196
rect 52368 6190 52420 6196
rect 52274 6080 52330 6089
rect 52274 6015 52330 6024
rect 52458 6080 52514 6089
rect 52458 6015 52514 6024
rect 52288 5817 52316 6015
rect 52274 5808 52330 5817
rect 52274 5743 52330 5752
rect 52472 5409 52500 6015
rect 52564 5658 52592 6276
rect 52644 6258 52696 6264
rect 52656 5778 52684 6258
rect 52644 5772 52696 5778
rect 52644 5714 52696 5720
rect 52736 5772 52788 5778
rect 52736 5714 52788 5720
rect 52748 5658 52776 5714
rect 52564 5630 52776 5658
rect 52458 5400 52514 5409
rect 52458 5335 52514 5344
rect 52840 5234 52868 10406
rect 53392 10062 53420 12200
rect 53472 11756 53524 11762
rect 53472 11698 53524 11704
rect 53484 11642 53512 11698
rect 53484 11614 53604 11642
rect 53576 11082 53604 11614
rect 53564 11076 53616 11082
rect 53564 11018 53616 11024
rect 53472 10668 53524 10674
rect 53472 10610 53524 10616
rect 53380 10056 53432 10062
rect 53380 9998 53432 10004
rect 53484 9994 53512 10610
rect 53472 9988 53524 9994
rect 53472 9930 53524 9936
rect 53286 9616 53342 9625
rect 53196 9580 53248 9586
rect 53286 9551 53342 9560
rect 53196 9522 53248 9528
rect 53102 9344 53158 9353
rect 53102 9279 53158 9288
rect 53116 8673 53144 9279
rect 53208 9042 53236 9522
rect 53300 9353 53328 9551
rect 53484 9518 53512 9930
rect 53472 9512 53524 9518
rect 53472 9454 53524 9460
rect 53286 9344 53342 9353
rect 53286 9279 53342 9288
rect 53196 9036 53248 9042
rect 53196 8978 53248 8984
rect 53288 8900 53340 8906
rect 53288 8842 53340 8848
rect 52918 8664 52974 8673
rect 52918 8599 52974 8608
rect 53102 8664 53158 8673
rect 53102 8599 53158 8608
rect 53196 8628 53248 8634
rect 52932 8514 52960 8599
rect 53196 8570 53248 8576
rect 52932 8486 53144 8514
rect 53012 8424 53064 8430
rect 53012 8366 53064 8372
rect 53024 8090 53052 8366
rect 53012 8084 53064 8090
rect 53012 8026 53064 8032
rect 53116 5409 53144 8486
rect 53208 6866 53236 8570
rect 53300 8362 53328 8842
rect 53288 8356 53340 8362
rect 53288 8298 53340 8304
rect 53576 7478 53604 11018
rect 53760 9738 53788 12200
rect 54022 11928 54078 11937
rect 54022 11863 54078 11872
rect 53668 9710 53788 9738
rect 53668 9178 53696 9710
rect 53746 9616 53802 9625
rect 53746 9551 53802 9560
rect 53840 9580 53892 9586
rect 53760 9450 53788 9551
rect 53840 9522 53892 9528
rect 53748 9444 53800 9450
rect 53748 9386 53800 9392
rect 53852 9353 53880 9522
rect 53838 9344 53894 9353
rect 53838 9279 53894 9288
rect 53656 9172 53708 9178
rect 53656 9114 53708 9120
rect 54036 8634 54064 11863
rect 54128 8974 54156 12200
rect 54496 9994 54524 12200
rect 54574 12135 54630 12144
rect 54588 11762 54616 12135
rect 54864 11778 54892 12200
rect 55232 12073 55260 12200
rect 55586 12200 55642 13000
rect 55678 12608 55734 12617
rect 55678 12543 55680 12552
rect 55732 12543 55734 12552
rect 55680 12514 55732 12520
rect 55770 12472 55826 12481
rect 55770 12407 55826 12416
rect 55678 12336 55734 12345
rect 55678 12271 55734 12280
rect 55404 12174 55456 12180
rect 55218 12064 55274 12073
rect 55218 11999 55274 12008
rect 55416 11801 55444 12174
rect 54576 11756 54628 11762
rect 54576 11698 54628 11704
rect 54772 11750 54892 11778
rect 55402 11792 55458 11801
rect 54588 11014 54616 11698
rect 54668 11076 54720 11082
rect 54668 11018 54720 11024
rect 54576 11008 54628 11014
rect 54576 10950 54628 10956
rect 54484 9988 54536 9994
rect 54484 9930 54536 9936
rect 54576 9988 54628 9994
rect 54576 9930 54628 9936
rect 54588 9897 54616 9930
rect 54574 9888 54630 9897
rect 54574 9823 54630 9832
rect 54680 9654 54708 11018
rect 54668 9648 54720 9654
rect 54668 9590 54720 9596
rect 54300 9444 54352 9450
rect 54300 9386 54352 9392
rect 54116 8968 54168 8974
rect 54116 8910 54168 8916
rect 54024 8628 54076 8634
rect 54024 8570 54076 8576
rect 54024 7880 54076 7886
rect 54024 7822 54076 7828
rect 53564 7472 53616 7478
rect 53564 7414 53616 7420
rect 53196 6860 53248 6866
rect 53196 6802 53248 6808
rect 54036 6458 54064 7822
rect 54116 6996 54168 7002
rect 54116 6938 54168 6944
rect 54024 6452 54076 6458
rect 54024 6394 54076 6400
rect 53746 5808 53802 5817
rect 53746 5743 53802 5752
rect 53102 5400 53158 5409
rect 53102 5335 53158 5344
rect 52828 5228 52880 5234
rect 52828 5170 52880 5176
rect 53656 5228 53708 5234
rect 53656 5170 53708 5176
rect 51814 5128 51870 5137
rect 51814 5063 51870 5072
rect 53668 4826 53696 5170
rect 53760 5030 53788 5743
rect 53748 5024 53800 5030
rect 53748 4966 53800 4972
rect 52828 4820 52880 4826
rect 52828 4762 52880 4768
rect 53656 4820 53708 4826
rect 53656 4762 53708 4768
rect 52092 4480 52144 4486
rect 52092 4422 52144 4428
rect 51816 4072 51868 4078
rect 51816 4014 51868 4020
rect 52000 4072 52052 4078
rect 52000 4014 52052 4020
rect 51724 3732 51776 3738
rect 51828 3720 51856 4014
rect 51908 3732 51960 3738
rect 51828 3692 51908 3720
rect 51724 3674 51776 3680
rect 51908 3674 51960 3680
rect 52012 3670 52040 4014
rect 52000 3664 52052 3670
rect 52000 3606 52052 3612
rect 51816 3528 51868 3534
rect 51552 3488 51816 3516
rect 51092 3454 51304 3482
rect 51816 3470 51868 3476
rect 51276 2990 51304 3454
rect 52104 3074 52132 4422
rect 52368 4140 52420 4146
rect 52368 4082 52420 4088
rect 52380 3602 52408 4082
rect 52642 3632 52698 3641
rect 52368 3596 52420 3602
rect 52642 3567 52698 3576
rect 52368 3538 52420 3544
rect 52184 3392 52236 3398
rect 52184 3334 52236 3340
rect 51736 3046 52132 3074
rect 51264 2984 51316 2990
rect 51264 2926 51316 2932
rect 51736 2922 51764 3046
rect 52196 2922 52224 3334
rect 51080 2916 51132 2922
rect 51080 2858 51132 2864
rect 51724 2916 51776 2922
rect 51724 2858 51776 2864
rect 52184 2916 52236 2922
rect 52184 2858 52236 2864
rect 51092 2666 51120 2858
rect 50804 2644 50856 2650
rect 50804 2586 50856 2592
rect 50896 2644 50948 2650
rect 51092 2638 51580 2666
rect 50896 2586 50948 2592
rect 50620 2508 50672 2514
rect 50620 2450 50672 2456
rect 50712 2508 50764 2514
rect 50712 2450 50764 2456
rect 50816 2502 51396 2530
rect 50252 2440 50304 2446
rect 50252 2382 50304 2388
rect 50252 2032 50304 2038
rect 50816 1986 50844 2502
rect 51368 2446 51396 2502
rect 51552 2446 51580 2638
rect 51724 2644 51776 2650
rect 51724 2586 51776 2592
rect 51172 2440 51224 2446
rect 50252 1974 50304 1980
rect 50068 1352 50120 1358
rect 50068 1294 50120 1300
rect 50080 1222 50108 1294
rect 50068 1216 50120 1222
rect 50068 1158 50120 1164
rect 50160 1216 50212 1222
rect 50160 1158 50212 1164
rect 50172 1018 50200 1158
rect 50160 1012 50212 1018
rect 50264 1000 50292 1974
rect 50356 1958 50844 1986
rect 50908 2400 51172 2428
rect 50356 1494 50384 1958
rect 50712 1896 50764 1902
rect 50712 1838 50764 1844
rect 50724 1766 50752 1838
rect 50620 1760 50672 1766
rect 50620 1702 50672 1708
rect 50712 1760 50764 1766
rect 50712 1702 50764 1708
rect 50344 1488 50396 1494
rect 50344 1430 50396 1436
rect 50528 1420 50580 1426
rect 50448 1380 50528 1408
rect 50344 1352 50396 1358
rect 50448 1306 50476 1380
rect 50528 1362 50580 1368
rect 50396 1300 50476 1306
rect 50344 1294 50476 1300
rect 50356 1278 50476 1294
rect 50632 1170 50660 1702
rect 50802 1184 50858 1193
rect 50632 1142 50802 1170
rect 50802 1119 50858 1128
rect 50908 1034 50936 2400
rect 51172 2382 51224 2388
rect 51356 2440 51408 2446
rect 51356 2382 51408 2388
rect 51540 2440 51592 2446
rect 51540 2382 51592 2388
rect 51264 2372 51316 2378
rect 51264 2314 51316 2320
rect 51276 2106 51304 2314
rect 51356 2304 51408 2310
rect 51356 2246 51408 2252
rect 51448 2304 51500 2310
rect 51448 2246 51500 2252
rect 51080 2100 51132 2106
rect 51080 2042 51132 2048
rect 51264 2100 51316 2106
rect 51264 2042 51316 2048
rect 51092 1850 51120 2042
rect 51092 1822 51304 1850
rect 51276 1766 51304 1822
rect 51264 1760 51316 1766
rect 51000 1686 51120 1714
rect 51264 1702 51316 1708
rect 51000 1562 51028 1686
rect 51092 1562 51120 1686
rect 50988 1556 51040 1562
rect 50988 1498 51040 1504
rect 51080 1556 51132 1562
rect 51080 1498 51132 1504
rect 50436 1012 50488 1018
rect 50264 972 50436 1000
rect 50160 954 50212 960
rect 50436 954 50488 960
rect 50632 1006 50936 1034
rect 50172 882 50200 954
rect 50160 876 50212 882
rect 49896 836 50016 864
rect 49896 800 49924 836
rect 49700 740 49752 746
rect 49700 682 49752 688
rect 49792 740 49844 746
rect 49792 682 49844 688
rect 49804 626 49832 682
rect 49620 598 49832 626
rect 49882 0 49938 800
rect 49988 66 50016 836
rect 50160 818 50212 824
rect 50264 836 50384 864
rect 50264 800 50292 836
rect 50160 740 50212 746
rect 50160 682 50212 688
rect 50172 134 50200 682
rect 50160 128 50212 134
rect 50160 70 50212 76
rect 49976 60 50028 66
rect 49976 2 50028 8
rect 50250 0 50306 800
rect 50356 134 50384 836
rect 50632 800 50660 1006
rect 50816 870 51028 898
rect 50816 814 50844 870
rect 50804 808 50856 814
rect 50344 128 50396 134
rect 50344 70 50396 76
rect 50618 0 50674 800
rect 50804 750 50856 756
rect 50896 808 50948 814
rect 51000 800 51028 870
rect 51368 800 51396 2246
rect 51460 1902 51488 2246
rect 51448 1896 51500 1902
rect 51448 1838 51500 1844
rect 51736 800 51764 2586
rect 52656 2514 52684 3567
rect 52840 2650 52868 4762
rect 53196 4276 53248 4282
rect 53196 4218 53248 4224
rect 53208 3126 53236 4218
rect 54024 3528 54076 3534
rect 54024 3470 54076 3476
rect 53288 3392 53340 3398
rect 53288 3334 53340 3340
rect 53104 3120 53156 3126
rect 53104 3062 53156 3068
rect 53196 3120 53248 3126
rect 53196 3062 53248 3068
rect 52828 2644 52880 2650
rect 52828 2586 52880 2592
rect 52644 2508 52696 2514
rect 52644 2450 52696 2456
rect 52092 2440 52144 2446
rect 52092 2382 52144 2388
rect 51816 2304 51868 2310
rect 51816 2246 51868 2252
rect 51908 2304 51960 2310
rect 51908 2246 51960 2252
rect 51828 1834 51856 2246
rect 51920 1970 51948 2246
rect 51908 1964 51960 1970
rect 51908 1906 51960 1912
rect 51816 1828 51868 1834
rect 51816 1770 51868 1776
rect 51908 1352 51960 1358
rect 51960 1312 52040 1340
rect 51908 1294 51960 1300
rect 50896 750 50948 756
rect 50908 474 50936 750
rect 50896 468 50948 474
rect 50896 410 50948 416
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51722 0 51778 800
rect 52012 746 52040 1312
rect 52104 800 52132 2382
rect 53116 2106 53144 3062
rect 53300 2650 53328 3334
rect 53472 3052 53524 3058
rect 53472 2994 53524 3000
rect 53656 3052 53708 3058
rect 53656 2994 53708 3000
rect 53288 2644 53340 2650
rect 53288 2586 53340 2592
rect 53300 2446 53328 2586
rect 53288 2440 53340 2446
rect 53288 2382 53340 2388
rect 52460 2100 52512 2106
rect 52460 2042 52512 2048
rect 53104 2100 53156 2106
rect 53104 2042 53156 2048
rect 52184 1896 52236 1902
rect 52184 1838 52236 1844
rect 52196 1358 52224 1838
rect 52184 1352 52236 1358
rect 52184 1294 52236 1300
rect 52472 800 52500 2042
rect 53484 1426 53512 2994
rect 53668 2650 53696 2994
rect 53656 2644 53708 2650
rect 53656 2586 53708 2592
rect 54036 2514 54064 3470
rect 54024 2508 54076 2514
rect 54024 2450 54076 2456
rect 54128 2038 54156 6938
rect 54312 4146 54340 9386
rect 54680 9042 54708 9590
rect 54668 9036 54720 9042
rect 54668 8978 54720 8984
rect 54772 8498 54800 11750
rect 55402 11727 55458 11736
rect 54944 11688 54996 11694
rect 54944 11630 54996 11636
rect 55128 11688 55180 11694
rect 55128 11630 55180 11636
rect 54956 10674 54984 11630
rect 55140 11150 55168 11630
rect 55128 11144 55180 11150
rect 55128 11086 55180 11092
rect 55312 11144 55364 11150
rect 55312 11086 55364 11092
rect 55496 11144 55548 11150
rect 55496 11086 55548 11092
rect 55128 11008 55180 11014
rect 55128 10950 55180 10956
rect 54944 10668 54996 10674
rect 54944 10610 54996 10616
rect 54956 10266 54984 10610
rect 55140 10441 55168 10950
rect 55324 10742 55352 11086
rect 55312 10736 55364 10742
rect 55312 10678 55364 10684
rect 55508 10470 55536 11086
rect 55220 10464 55272 10470
rect 55126 10432 55182 10441
rect 55220 10406 55272 10412
rect 55496 10464 55548 10470
rect 55496 10406 55548 10412
rect 55126 10367 55182 10376
rect 54944 10260 54996 10266
rect 54944 10202 54996 10208
rect 55128 9920 55180 9926
rect 55128 9862 55180 9868
rect 54852 9648 54904 9654
rect 54852 9590 54904 9596
rect 54864 9110 54892 9590
rect 55140 9586 55168 9862
rect 54944 9580 54996 9586
rect 54944 9522 54996 9528
rect 55128 9580 55180 9586
rect 55128 9522 55180 9528
rect 54956 9432 54984 9522
rect 55036 9444 55088 9450
rect 54956 9404 55036 9432
rect 55036 9386 55088 9392
rect 55140 9178 55168 9522
rect 55128 9172 55180 9178
rect 55128 9114 55180 9120
rect 54852 9104 54904 9110
rect 54852 9046 54904 9052
rect 54760 8492 54812 8498
rect 54760 8434 54812 8440
rect 54852 8424 54904 8430
rect 54852 8366 54904 8372
rect 54392 8288 54444 8294
rect 54392 8230 54444 8236
rect 54404 7886 54432 8230
rect 54392 7880 54444 7886
rect 54392 7822 54444 7828
rect 54576 7880 54628 7886
rect 54576 7822 54628 7828
rect 54404 7478 54432 7822
rect 54392 7472 54444 7478
rect 54392 7414 54444 7420
rect 54482 5128 54538 5137
rect 54482 5063 54538 5072
rect 54300 4140 54352 4146
rect 54300 4082 54352 4088
rect 54496 3466 54524 5063
rect 54484 3460 54536 3466
rect 54484 3402 54536 3408
rect 54588 2854 54616 7822
rect 54864 7478 54892 8366
rect 54944 8356 54996 8362
rect 54944 8298 54996 8304
rect 54852 7472 54904 7478
rect 54852 7414 54904 7420
rect 54852 7336 54904 7342
rect 54852 7278 54904 7284
rect 54760 6792 54812 6798
rect 54760 6734 54812 6740
rect 54668 6384 54720 6390
rect 54668 6326 54720 6332
rect 54680 5778 54708 6326
rect 54668 5772 54720 5778
rect 54668 5714 54720 5720
rect 54772 4622 54800 6734
rect 54864 5817 54892 7278
rect 54850 5808 54906 5817
rect 54850 5743 54906 5752
rect 54852 5636 54904 5642
rect 54852 5578 54904 5584
rect 54760 4616 54812 4622
rect 54760 4558 54812 4564
rect 54760 4072 54812 4078
rect 54760 4014 54812 4020
rect 54772 3670 54800 4014
rect 54760 3664 54812 3670
rect 54760 3606 54812 3612
rect 54864 2938 54892 5578
rect 54956 3058 54984 8298
rect 55126 7712 55182 7721
rect 55126 7647 55182 7656
rect 55140 7002 55168 7647
rect 55128 6996 55180 7002
rect 55128 6938 55180 6944
rect 55036 6248 55088 6254
rect 55036 6190 55088 6196
rect 55048 5574 55076 6190
rect 55128 5704 55180 5710
rect 55128 5646 55180 5652
rect 55140 5574 55168 5646
rect 55036 5568 55088 5574
rect 55036 5510 55088 5516
rect 55128 5568 55180 5574
rect 55128 5510 55180 5516
rect 55034 5128 55090 5137
rect 55034 5063 55090 5072
rect 55048 4282 55076 5063
rect 55232 4826 55260 10406
rect 55404 10260 55456 10266
rect 55404 10202 55456 10208
rect 55496 10260 55548 10266
rect 55496 10202 55548 10208
rect 55312 8356 55364 8362
rect 55312 8298 55364 8304
rect 55220 4820 55272 4826
rect 55220 4762 55272 4768
rect 55128 4480 55180 4486
rect 55128 4422 55180 4428
rect 55140 4282 55168 4422
rect 55036 4276 55088 4282
rect 55036 4218 55088 4224
rect 55128 4276 55180 4282
rect 55128 4218 55180 4224
rect 55324 4146 55352 8298
rect 55416 5234 55444 10202
rect 55508 10130 55536 10202
rect 55496 10124 55548 10130
rect 55496 10066 55548 10072
rect 55600 9518 55628 12200
rect 55692 9654 55720 12271
rect 55680 9648 55732 9654
rect 55680 9590 55732 9596
rect 55588 9512 55640 9518
rect 55588 9454 55640 9460
rect 55496 8968 55548 8974
rect 55496 8910 55548 8916
rect 55508 7970 55536 8910
rect 55784 8906 55812 12407
rect 55954 12200 56010 13000
rect 56140 12504 56192 12510
rect 56140 12446 56192 12452
rect 55864 12096 55916 12102
rect 55864 12038 55916 12044
rect 55876 11898 55904 12038
rect 55864 11892 55916 11898
rect 55864 11834 55916 11840
rect 55864 10736 55916 10742
rect 55864 10678 55916 10684
rect 55876 10062 55904 10678
rect 55864 10056 55916 10062
rect 55864 9998 55916 10004
rect 55864 9920 55916 9926
rect 55968 9897 55996 12200
rect 56152 11558 56180 12446
rect 56322 12200 56378 13000
rect 56508 12980 56560 12986
rect 56508 12922 56560 12928
rect 56336 11937 56364 12200
rect 56322 11928 56378 11937
rect 56322 11863 56378 11872
rect 56322 11792 56378 11801
rect 56520 11762 56548 12922
rect 56690 12200 56746 13000
rect 56968 12504 57020 12510
rect 56782 12472 56838 12481
rect 56968 12446 57020 12452
rect 56782 12407 56838 12416
rect 56704 12152 56732 12200
rect 56796 12152 56824 12407
rect 56704 12124 56824 12152
rect 56641 11996 56937 12016
rect 56697 11994 56721 11996
rect 56777 11994 56801 11996
rect 56857 11994 56881 11996
rect 56719 11942 56721 11994
rect 56783 11942 56795 11994
rect 56857 11942 56859 11994
rect 56697 11940 56721 11942
rect 56777 11940 56801 11942
rect 56857 11940 56881 11942
rect 56641 11920 56937 11940
rect 56322 11727 56324 11736
rect 56376 11727 56378 11736
rect 56508 11756 56560 11762
rect 56324 11698 56376 11704
rect 56508 11698 56560 11704
rect 56876 11756 56928 11762
rect 56876 11698 56928 11704
rect 56140 11552 56192 11558
rect 56140 11494 56192 11500
rect 56048 11144 56100 11150
rect 56048 11086 56100 11092
rect 56060 10470 56088 11086
rect 56138 10840 56194 10849
rect 56138 10775 56194 10784
rect 56048 10464 56100 10470
rect 56048 10406 56100 10412
rect 55864 9862 55916 9868
rect 55954 9888 56010 9897
rect 55876 9738 55904 9862
rect 55954 9823 56010 9832
rect 55954 9752 56010 9761
rect 55876 9710 55954 9738
rect 55954 9687 56010 9696
rect 55864 9580 55916 9586
rect 55864 9522 55916 9528
rect 55876 9042 55904 9522
rect 55956 9172 56008 9178
rect 55956 9114 56008 9120
rect 55864 9036 55916 9042
rect 55864 8978 55916 8984
rect 55772 8900 55824 8906
rect 55772 8842 55824 8848
rect 55864 8900 55916 8906
rect 55864 8842 55916 8848
rect 55772 8628 55824 8634
rect 55772 8570 55824 8576
rect 55680 8492 55732 8498
rect 55680 8434 55732 8440
rect 55692 8090 55720 8434
rect 55680 8084 55732 8090
rect 55680 8026 55732 8032
rect 55508 7942 55720 7970
rect 55588 7812 55640 7818
rect 55588 7754 55640 7760
rect 55494 7712 55550 7721
rect 55494 7647 55550 7656
rect 55508 7206 55536 7647
rect 55600 7410 55628 7754
rect 55588 7404 55640 7410
rect 55588 7346 55640 7352
rect 55496 7200 55548 7206
rect 55496 7142 55548 7148
rect 55692 7018 55720 7942
rect 55784 7750 55812 8570
rect 55876 8294 55904 8842
rect 55968 8498 55996 9114
rect 56060 8498 56088 10406
rect 56152 10130 56180 10775
rect 56232 10668 56284 10674
rect 56232 10610 56284 10616
rect 56140 10124 56192 10130
rect 56140 10066 56192 10072
rect 56244 10010 56272 10610
rect 56336 10470 56364 11698
rect 56520 11150 56548 11698
rect 56784 11688 56836 11694
rect 56784 11630 56836 11636
rect 56796 11150 56824 11630
rect 56508 11144 56560 11150
rect 56508 11086 56560 11092
rect 56784 11144 56836 11150
rect 56784 11086 56836 11092
rect 56888 10996 56916 11698
rect 56980 11286 57008 12446
rect 57058 12200 57114 13000
rect 57426 12200 57482 13000
rect 57610 12200 57666 12209
rect 57794 12200 57850 13000
rect 58162 12200 58218 13000
rect 58256 12300 58308 12306
rect 58256 12242 58308 12248
rect 56968 11280 57020 11286
rect 56968 11222 57020 11228
rect 56414 10976 56470 10985
rect 56888 10968 57008 10996
rect 56414 10911 56470 10920
rect 56428 10792 56456 10911
rect 56641 10908 56937 10928
rect 56697 10906 56721 10908
rect 56777 10906 56801 10908
rect 56857 10906 56881 10908
rect 56719 10854 56721 10906
rect 56783 10854 56795 10906
rect 56857 10854 56859 10906
rect 56697 10852 56721 10854
rect 56777 10852 56801 10854
rect 56857 10852 56881 10854
rect 56641 10832 56937 10852
rect 56428 10764 56640 10792
rect 56416 10668 56468 10674
rect 56416 10610 56468 10616
rect 56324 10464 56376 10470
rect 56324 10406 56376 10412
rect 56152 9982 56272 10010
rect 56152 9654 56180 9982
rect 56322 9888 56378 9897
rect 56322 9823 56378 9832
rect 56140 9648 56192 9654
rect 56140 9590 56192 9596
rect 56140 9444 56192 9450
rect 56140 9386 56192 9392
rect 56152 9042 56180 9386
rect 56140 9036 56192 9042
rect 56140 8978 56192 8984
rect 56336 8906 56364 9823
rect 56428 9761 56456 10610
rect 56508 10532 56560 10538
rect 56508 10474 56560 10480
rect 56520 10130 56548 10474
rect 56508 10124 56560 10130
rect 56508 10066 56560 10072
rect 56612 9994 56640 10764
rect 56980 10606 57008 10968
rect 56968 10600 57020 10606
rect 56968 10542 57020 10548
rect 56980 10282 57008 10542
rect 56796 10254 57008 10282
rect 56796 10062 56824 10254
rect 57072 10180 57100 12200
rect 57440 11762 57468 12200
rect 57610 12135 57666 12144
rect 57428 11756 57480 11762
rect 57428 11698 57480 11704
rect 57152 11144 57204 11150
rect 57204 11104 57284 11132
rect 57152 11086 57204 11092
rect 57152 11008 57204 11014
rect 57150 10976 57152 10985
rect 57204 10976 57206 10985
rect 57150 10911 57206 10920
rect 56888 10152 57100 10180
rect 56784 10056 56836 10062
rect 56784 9998 56836 10004
rect 56888 10010 56916 10152
rect 56600 9988 56652 9994
rect 56888 9982 57008 10010
rect 56600 9930 56652 9936
rect 56641 9820 56937 9840
rect 56697 9818 56721 9820
rect 56777 9818 56801 9820
rect 56857 9818 56881 9820
rect 56719 9766 56721 9818
rect 56783 9766 56795 9818
rect 56857 9766 56859 9818
rect 56697 9764 56721 9766
rect 56777 9764 56801 9766
rect 56857 9764 56881 9766
rect 56414 9752 56470 9761
rect 56641 9744 56937 9764
rect 56414 9687 56470 9696
rect 56980 9602 57008 9982
rect 57060 9988 57112 9994
rect 57060 9930 57112 9936
rect 56796 9586 57008 9602
rect 56784 9580 57008 9586
rect 56836 9574 57008 9580
rect 56784 9522 56836 9528
rect 56508 9376 56560 9382
rect 56876 9376 56928 9382
rect 56508 9318 56560 9324
rect 56612 9336 56876 9364
rect 56520 8974 56548 9318
rect 56508 8968 56560 8974
rect 56508 8910 56560 8916
rect 56324 8900 56376 8906
rect 56324 8842 56376 8848
rect 56612 8820 56640 9336
rect 56876 9318 56928 9324
rect 56784 8968 56836 8974
rect 56836 8928 57008 8956
rect 56784 8910 56836 8916
rect 56520 8809 56640 8820
rect 56322 8800 56378 8809
rect 56322 8735 56378 8744
rect 56506 8800 56640 8809
rect 56562 8792 56640 8800
rect 56506 8735 56562 8744
rect 55956 8492 56008 8498
rect 55956 8434 56008 8440
rect 56048 8492 56100 8498
rect 56048 8434 56100 8440
rect 56232 8492 56284 8498
rect 56232 8434 56284 8440
rect 55864 8288 55916 8294
rect 55864 8230 55916 8236
rect 56140 8288 56192 8294
rect 56140 8230 56192 8236
rect 56048 7948 56100 7954
rect 56048 7890 56100 7896
rect 55864 7812 55916 7818
rect 56060 7800 56088 7890
rect 55916 7772 56088 7800
rect 55864 7754 55916 7760
rect 55772 7744 55824 7750
rect 55772 7686 55824 7692
rect 56152 7562 56180 8230
rect 56244 7750 56272 8434
rect 56232 7744 56284 7750
rect 56232 7686 56284 7692
rect 55508 6990 55720 7018
rect 55968 7534 56180 7562
rect 55508 6390 55536 6990
rect 55680 6928 55732 6934
rect 55680 6870 55732 6876
rect 55586 6488 55642 6497
rect 55586 6423 55642 6432
rect 55496 6384 55548 6390
rect 55496 6326 55548 6332
rect 55494 5808 55550 5817
rect 55494 5743 55550 5752
rect 55508 5642 55536 5743
rect 55496 5636 55548 5642
rect 55496 5578 55548 5584
rect 55404 5228 55456 5234
rect 55404 5170 55456 5176
rect 55600 5114 55628 6423
rect 55692 5386 55720 6870
rect 55864 6180 55916 6186
rect 55864 6122 55916 6128
rect 55876 5817 55904 6122
rect 55862 5808 55918 5817
rect 55862 5743 55918 5752
rect 55968 5574 55996 7534
rect 56140 7404 56192 7410
rect 56140 7346 56192 7352
rect 56048 7268 56100 7274
rect 56048 7210 56100 7216
rect 56060 6497 56088 7210
rect 56152 6866 56180 7346
rect 56140 6860 56192 6866
rect 56140 6802 56192 6808
rect 56244 6798 56272 7686
rect 56336 6916 56364 8735
rect 56641 8732 56937 8752
rect 56697 8730 56721 8732
rect 56777 8730 56801 8732
rect 56857 8730 56881 8732
rect 56719 8678 56721 8730
rect 56783 8678 56795 8730
rect 56857 8678 56859 8730
rect 56697 8676 56721 8678
rect 56777 8676 56801 8678
rect 56857 8676 56881 8678
rect 56641 8656 56937 8676
rect 56784 8560 56836 8566
rect 56784 8502 56836 8508
rect 56796 8362 56824 8502
rect 56784 8356 56836 8362
rect 56784 8298 56836 8304
rect 56876 8084 56928 8090
rect 56876 8026 56928 8032
rect 56888 7800 56916 8026
rect 56980 7936 57008 8928
rect 57072 8090 57100 9930
rect 57150 9344 57206 9353
rect 57150 9279 57206 9288
rect 57164 8809 57192 9279
rect 57150 8800 57206 8809
rect 57150 8735 57206 8744
rect 57256 8294 57284 11104
rect 57426 10568 57482 10577
rect 57426 10503 57428 10512
rect 57480 10503 57482 10512
rect 57428 10474 57480 10480
rect 57428 9988 57480 9994
rect 57480 9948 57560 9976
rect 57428 9930 57480 9936
rect 57532 9636 57560 9948
rect 57624 9897 57652 12135
rect 57808 11880 57836 12200
rect 58070 12064 58126 12073
rect 58070 11999 58126 12008
rect 57716 11852 57836 11880
rect 57716 10130 57744 11852
rect 58084 11762 58112 11999
rect 57796 11756 57848 11762
rect 57796 11698 57848 11704
rect 58072 11756 58124 11762
rect 58072 11698 58124 11704
rect 57808 11082 57836 11698
rect 57796 11076 57848 11082
rect 57796 11018 57848 11024
rect 58072 11008 58124 11014
rect 58072 10950 58124 10956
rect 58084 10742 58112 10950
rect 58072 10736 58124 10742
rect 58072 10678 58124 10684
rect 57888 10668 57940 10674
rect 57888 10610 57940 10616
rect 57900 10130 57928 10610
rect 57980 10600 58032 10606
rect 57980 10542 58032 10548
rect 57704 10124 57756 10130
rect 57704 10066 57756 10072
rect 57888 10124 57940 10130
rect 57888 10066 57940 10072
rect 57796 10056 57848 10062
rect 57796 9998 57848 10004
rect 57610 9888 57666 9897
rect 57808 9874 57836 9998
rect 57610 9823 57666 9832
rect 57716 9846 57836 9874
rect 57716 9654 57744 9846
rect 57888 9716 57940 9722
rect 57888 9658 57940 9664
rect 57440 9608 57560 9636
rect 57704 9648 57756 9654
rect 57336 9376 57388 9382
rect 57336 9318 57388 9324
rect 57348 8673 57376 9318
rect 57334 8664 57390 8673
rect 57334 8599 57390 8608
rect 57440 8498 57468 9608
rect 57704 9590 57756 9596
rect 57900 9586 57928 9658
rect 57888 9580 57940 9586
rect 57888 9522 57940 9528
rect 57796 9444 57848 9450
rect 57796 9386 57848 9392
rect 57520 9376 57572 9382
rect 57520 9318 57572 9324
rect 57610 9344 57666 9353
rect 57428 8492 57480 8498
rect 57428 8434 57480 8440
rect 57244 8288 57296 8294
rect 57244 8230 57296 8236
rect 57428 8288 57480 8294
rect 57428 8230 57480 8236
rect 57060 8084 57112 8090
rect 57060 8026 57112 8032
rect 57336 7948 57388 7954
rect 56980 7908 57192 7936
rect 57060 7812 57112 7818
rect 56888 7772 57060 7800
rect 57060 7754 57112 7760
rect 56508 7744 56560 7750
rect 56506 7712 56508 7721
rect 56560 7712 56562 7721
rect 56506 7647 56562 7656
rect 56641 7644 56937 7664
rect 56697 7642 56721 7644
rect 56777 7642 56801 7644
rect 56857 7642 56881 7644
rect 56719 7590 56721 7642
rect 56783 7590 56795 7642
rect 56857 7590 56859 7642
rect 56697 7588 56721 7590
rect 56777 7588 56801 7590
rect 56857 7588 56881 7590
rect 56506 7576 56562 7585
rect 56641 7568 56937 7588
rect 57058 7576 57114 7585
rect 56506 7511 56562 7520
rect 57058 7511 57114 7520
rect 56520 7290 56548 7511
rect 56784 7404 56836 7410
rect 56968 7404 57020 7410
rect 56836 7364 56968 7392
rect 56784 7346 56836 7352
rect 56968 7346 57020 7352
rect 56520 7274 57008 7290
rect 56520 7268 57020 7274
rect 56520 7262 56968 7268
rect 56968 7210 57020 7216
rect 56600 7200 56652 7206
rect 57072 7154 57100 7511
rect 56652 7148 57100 7154
rect 56600 7142 57100 7148
rect 56612 7126 57100 7142
rect 56508 6928 56560 6934
rect 56336 6888 56508 6916
rect 56508 6870 56560 6876
rect 56232 6792 56284 6798
rect 56232 6734 56284 6740
rect 56324 6792 56376 6798
rect 56324 6734 56376 6740
rect 56336 6662 56364 6734
rect 56324 6656 56376 6662
rect 56230 6624 56286 6633
rect 56324 6598 56376 6604
rect 56416 6656 56468 6662
rect 56416 6598 56468 6604
rect 56968 6656 57020 6662
rect 56968 6598 57020 6604
rect 56230 6559 56286 6568
rect 56046 6488 56102 6497
rect 56046 6423 56102 6432
rect 55956 5568 56008 5574
rect 55956 5510 56008 5516
rect 56140 5568 56192 5574
rect 56140 5510 56192 5516
rect 55692 5358 55812 5386
rect 55678 5264 55734 5273
rect 55784 5234 55812 5358
rect 56152 5273 56180 5510
rect 56138 5264 56194 5273
rect 55678 5199 55734 5208
rect 55772 5228 55824 5234
rect 55416 5086 55628 5114
rect 55312 4140 55364 4146
rect 55312 4082 55364 4088
rect 55324 3738 55352 4082
rect 55312 3732 55364 3738
rect 55312 3674 55364 3680
rect 55220 3188 55272 3194
rect 55220 3130 55272 3136
rect 54944 3052 54996 3058
rect 54944 2994 54996 3000
rect 55128 3052 55180 3058
rect 55232 3040 55260 3130
rect 55180 3012 55260 3040
rect 55128 2994 55180 3000
rect 54864 2910 55076 2938
rect 54208 2848 54260 2854
rect 54208 2790 54260 2796
rect 54576 2848 54628 2854
rect 54576 2790 54628 2796
rect 54220 2514 54248 2790
rect 54208 2508 54260 2514
rect 54208 2450 54260 2456
rect 54588 2446 54616 2790
rect 54576 2440 54628 2446
rect 54576 2382 54628 2388
rect 53840 2032 53892 2038
rect 53840 1974 53892 1980
rect 54116 2032 54168 2038
rect 54116 1974 54168 1980
rect 53656 1964 53708 1970
rect 53656 1906 53708 1912
rect 53668 1766 53696 1906
rect 53656 1760 53708 1766
rect 53656 1702 53708 1708
rect 53196 1420 53248 1426
rect 53196 1362 53248 1368
rect 53472 1420 53524 1426
rect 53472 1362 53524 1368
rect 52564 972 52960 1000
rect 52564 882 52592 972
rect 52552 876 52604 882
rect 52552 818 52604 824
rect 52748 836 52868 864
rect 52000 740 52052 746
rect 52000 682 52052 688
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52748 474 52776 836
rect 52840 800 52868 836
rect 52736 468 52788 474
rect 52736 410 52788 416
rect 52826 0 52882 800
rect 52932 746 52960 972
rect 53012 876 53064 882
rect 53012 818 53064 824
rect 52920 740 52972 746
rect 52920 682 52972 688
rect 53024 474 53052 818
rect 53208 800 53236 1362
rect 53668 1358 53696 1702
rect 53852 1358 53880 1974
rect 54944 1896 54996 1902
rect 54944 1838 54996 1844
rect 54956 1737 54984 1838
rect 54942 1728 54998 1737
rect 54942 1663 54998 1672
rect 54300 1420 54352 1426
rect 54300 1362 54352 1368
rect 53656 1352 53708 1358
rect 53656 1294 53708 1300
rect 53840 1352 53892 1358
rect 53840 1294 53892 1300
rect 53484 836 53604 864
rect 53012 468 53064 474
rect 53012 410 53064 416
rect 53194 0 53250 800
rect 53484 678 53512 836
rect 53576 800 53604 836
rect 53852 836 53972 864
rect 53472 672 53524 678
rect 53472 614 53524 620
rect 53562 0 53618 800
rect 53656 672 53708 678
rect 53852 649 53880 836
rect 53944 800 53972 836
rect 54312 800 54340 1362
rect 54496 870 54708 898
rect 54496 814 54524 870
rect 54484 808 54536 814
rect 53656 614 53708 620
rect 53838 640 53894 649
rect 53668 513 53696 614
rect 53838 575 53894 584
rect 53654 504 53710 513
rect 53654 439 53710 448
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54680 800 54708 870
rect 55048 800 55076 2910
rect 55232 2650 55260 3012
rect 55312 2916 55364 2922
rect 55312 2858 55364 2864
rect 55220 2644 55272 2650
rect 55220 2586 55272 2592
rect 55126 2408 55182 2417
rect 55126 2343 55182 2352
rect 55140 1737 55168 2343
rect 55220 1964 55272 1970
rect 55220 1906 55272 1912
rect 55126 1728 55182 1737
rect 55126 1663 55182 1672
rect 55232 1494 55260 1906
rect 55324 1578 55352 2858
rect 55416 2854 55444 5086
rect 55692 5001 55720 5199
rect 56138 5199 56194 5208
rect 55772 5170 55824 5176
rect 56048 5024 56100 5030
rect 55678 4992 55734 5001
rect 56244 5012 56272 6559
rect 56428 6322 56456 6598
rect 56641 6556 56937 6576
rect 56697 6554 56721 6556
rect 56777 6554 56801 6556
rect 56857 6554 56881 6556
rect 56719 6502 56721 6554
rect 56783 6502 56795 6554
rect 56857 6502 56859 6554
rect 56697 6500 56721 6502
rect 56777 6500 56801 6502
rect 56857 6500 56881 6502
rect 56641 6480 56937 6500
rect 56416 6316 56468 6322
rect 56416 6258 56468 6264
rect 56980 6066 57008 6598
rect 56704 6038 57008 6066
rect 56600 5704 56652 5710
rect 56704 5692 56732 6038
rect 56968 5908 57020 5914
rect 56968 5850 57020 5856
rect 56652 5664 56732 5692
rect 56600 5646 56652 5652
rect 56322 5536 56378 5545
rect 56322 5471 56378 5480
rect 56336 5273 56364 5471
rect 56641 5468 56937 5488
rect 56697 5466 56721 5468
rect 56777 5466 56801 5468
rect 56857 5466 56881 5468
rect 56719 5414 56721 5466
rect 56783 5414 56795 5466
rect 56857 5414 56859 5466
rect 56697 5412 56721 5414
rect 56777 5412 56801 5414
rect 56857 5412 56881 5414
rect 56506 5400 56562 5409
rect 56641 5392 56937 5412
rect 56506 5335 56562 5344
rect 56322 5264 56378 5273
rect 56322 5199 56378 5208
rect 56048 4966 56100 4972
rect 56152 4984 56272 5012
rect 56324 5024 56376 5030
rect 55678 4927 55734 4936
rect 55496 4820 55548 4826
rect 55496 4762 55548 4768
rect 55508 4729 55536 4762
rect 55494 4720 55550 4729
rect 55494 4655 55550 4664
rect 55588 4616 55640 4622
rect 55494 4584 55550 4593
rect 55772 4616 55824 4622
rect 55640 4564 55720 4570
rect 55588 4558 55720 4564
rect 55772 4558 55824 4564
rect 55600 4542 55720 4558
rect 55494 4519 55550 4528
rect 55508 4486 55536 4519
rect 55496 4480 55548 4486
rect 55496 4422 55548 4428
rect 55588 4208 55640 4214
rect 55588 4150 55640 4156
rect 55496 4140 55548 4146
rect 55496 4082 55548 4088
rect 55508 3942 55536 4082
rect 55496 3936 55548 3942
rect 55496 3878 55548 3884
rect 55496 2984 55548 2990
rect 55494 2952 55496 2961
rect 55548 2952 55550 2961
rect 55494 2887 55550 2896
rect 55404 2848 55456 2854
rect 55404 2790 55456 2796
rect 55496 2848 55548 2854
rect 55496 2790 55548 2796
rect 55402 2408 55458 2417
rect 55402 2343 55458 2352
rect 55416 2145 55444 2343
rect 55402 2136 55458 2145
rect 55508 2106 55536 2790
rect 55402 2071 55458 2080
rect 55496 2100 55548 2106
rect 55496 2042 55548 2048
rect 55600 1766 55628 4150
rect 55692 3670 55720 4542
rect 55784 4282 55812 4558
rect 56060 4486 56088 4966
rect 56048 4480 56100 4486
rect 56048 4422 56100 4428
rect 55772 4276 55824 4282
rect 55772 4218 55824 4224
rect 55772 4072 55824 4078
rect 55772 4014 55824 4020
rect 55784 3942 55812 4014
rect 56048 4004 56100 4010
rect 56048 3946 56100 3952
rect 55772 3936 55824 3942
rect 55772 3878 55824 3884
rect 55680 3664 55732 3670
rect 55680 3606 55732 3612
rect 55864 3460 55916 3466
rect 55864 3402 55916 3408
rect 55680 3120 55732 3126
rect 55680 3062 55732 3068
rect 55692 2650 55720 3062
rect 55876 3058 55904 3402
rect 55956 3392 56008 3398
rect 55956 3334 56008 3340
rect 55864 3052 55916 3058
rect 55864 2994 55916 3000
rect 55968 2938 55996 3334
rect 56060 3233 56088 3946
rect 56046 3224 56102 3233
rect 56152 3194 56180 4984
rect 56324 4966 56376 4972
rect 56336 4690 56364 4966
rect 56324 4684 56376 4690
rect 56324 4626 56376 4632
rect 56520 4264 56548 5335
rect 56980 4758 57008 5850
rect 57060 5228 57112 5234
rect 57060 5170 57112 5176
rect 57072 5098 57100 5170
rect 57060 5092 57112 5098
rect 57060 5034 57112 5040
rect 56968 4752 57020 4758
rect 56968 4694 57020 4700
rect 56641 4380 56937 4400
rect 56697 4378 56721 4380
rect 56777 4378 56801 4380
rect 56857 4378 56881 4380
rect 56719 4326 56721 4378
rect 56783 4326 56795 4378
rect 56857 4326 56859 4378
rect 56697 4324 56721 4326
rect 56777 4324 56801 4326
rect 56857 4324 56881 4326
rect 56641 4304 56937 4324
rect 56980 4282 57008 4694
rect 56968 4276 57020 4282
rect 56244 4236 56456 4264
rect 56520 4236 56640 4264
rect 56244 4146 56272 4236
rect 56428 4162 56456 4236
rect 56612 4162 56640 4236
rect 56968 4218 57020 4224
rect 57060 4276 57112 4282
rect 57060 4218 57112 4224
rect 57072 4162 57100 4218
rect 56232 4140 56284 4146
rect 56232 4082 56284 4088
rect 56324 4140 56376 4146
rect 56428 4134 56548 4162
rect 56612 4134 57100 4162
rect 56324 4082 56376 4088
rect 56336 3534 56364 4082
rect 56416 3664 56468 3670
rect 56416 3606 56468 3612
rect 56324 3528 56376 3534
rect 56324 3470 56376 3476
rect 56046 3159 56102 3168
rect 56140 3188 56192 3194
rect 56140 3130 56192 3136
rect 56324 3052 56376 3058
rect 56324 2994 56376 3000
rect 55772 2916 55824 2922
rect 55772 2858 55824 2864
rect 55876 2910 55996 2938
rect 56140 2916 56192 2922
rect 55680 2644 55732 2650
rect 55680 2586 55732 2592
rect 55680 2508 55732 2514
rect 55680 2450 55732 2456
rect 55692 2281 55720 2450
rect 55678 2272 55734 2281
rect 55678 2207 55734 2216
rect 55404 1760 55456 1766
rect 55588 1760 55640 1766
rect 55456 1708 55536 1714
rect 55404 1702 55536 1708
rect 55588 1702 55640 1708
rect 55416 1686 55536 1702
rect 55324 1550 55444 1578
rect 55220 1488 55272 1494
rect 55220 1430 55272 1436
rect 55220 1352 55272 1358
rect 55220 1294 55272 1300
rect 54484 750 54536 756
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55232 746 55260 1294
rect 55312 1216 55364 1222
rect 55312 1158 55364 1164
rect 55324 882 55352 1158
rect 55312 876 55364 882
rect 55312 818 55364 824
rect 55416 800 55444 1550
rect 55508 1494 55536 1686
rect 55496 1488 55548 1494
rect 55496 1430 55548 1436
rect 55600 1358 55628 1702
rect 55588 1352 55640 1358
rect 55588 1294 55640 1300
rect 55678 912 55734 921
rect 55496 876 55548 882
rect 55678 847 55734 856
rect 55496 818 55548 824
rect 55220 740 55272 746
rect 55220 682 55272 688
rect 55402 0 55458 800
rect 55508 649 55536 818
rect 55692 649 55720 847
rect 55784 800 55812 2858
rect 55876 2038 55904 2910
rect 56140 2858 56192 2864
rect 56048 2440 56100 2446
rect 56048 2382 56100 2388
rect 56060 2310 56088 2382
rect 56048 2304 56100 2310
rect 56048 2246 56100 2252
rect 55954 2136 56010 2145
rect 55954 2071 56010 2080
rect 55864 2032 55916 2038
rect 55864 1974 55916 1980
rect 55968 1970 55996 2071
rect 55956 1964 56008 1970
rect 55956 1906 56008 1912
rect 56152 1766 56180 2858
rect 56232 2644 56284 2650
rect 56232 2586 56284 2592
rect 56140 1760 56192 1766
rect 56140 1702 56192 1708
rect 56244 1358 56272 2586
rect 56336 2038 56364 2994
rect 56324 2032 56376 2038
rect 56324 1974 56376 1980
rect 56232 1352 56284 1358
rect 56232 1294 56284 1300
rect 56048 1216 56100 1222
rect 56428 1204 56456 3606
rect 56520 3448 56548 4134
rect 57164 3602 57192 7908
rect 57336 7890 57388 7896
rect 57244 7744 57296 7750
rect 57242 7712 57244 7721
rect 57296 7712 57298 7721
rect 57242 7647 57298 7656
rect 57348 7562 57376 7890
rect 57256 7534 57376 7562
rect 57256 5914 57284 7534
rect 57440 7410 57468 8230
rect 57532 7954 57560 9318
rect 57610 9279 57666 9288
rect 57624 8974 57652 9279
rect 57808 9178 57836 9386
rect 57796 9172 57848 9178
rect 57796 9114 57848 9120
rect 57612 8968 57664 8974
rect 57612 8910 57664 8916
rect 57900 8634 57928 9522
rect 57992 9518 58020 10542
rect 58176 9738 58204 12200
rect 58268 11830 58296 12242
rect 58530 12200 58586 13000
rect 58898 12200 58954 13000
rect 59266 12200 59322 13000
rect 59452 12504 59504 12510
rect 59452 12446 59504 12452
rect 58438 12064 58494 12073
rect 58438 11999 58494 12008
rect 58256 11824 58308 11830
rect 58256 11766 58308 11772
rect 58452 11014 58480 11999
rect 58440 11008 58492 11014
rect 58440 10950 58492 10956
rect 58176 9710 58296 9738
rect 58268 9602 58296 9710
rect 58176 9574 58296 9602
rect 57980 9512 58032 9518
rect 57980 9454 58032 9460
rect 57980 9172 58032 9178
rect 57980 9114 58032 9120
rect 57796 8628 57848 8634
rect 57796 8570 57848 8576
rect 57888 8628 57940 8634
rect 57888 8570 57940 8576
rect 57612 8492 57664 8498
rect 57664 8452 57744 8480
rect 57612 8434 57664 8440
rect 57520 7948 57572 7954
rect 57520 7890 57572 7896
rect 57428 7404 57480 7410
rect 57428 7346 57480 7352
rect 57440 7290 57468 7346
rect 57348 7262 57468 7290
rect 57348 7002 57376 7262
rect 57612 7200 57664 7206
rect 57612 7142 57664 7148
rect 57336 6996 57388 7002
rect 57336 6938 57388 6944
rect 57520 6996 57572 7002
rect 57520 6938 57572 6944
rect 57428 6928 57480 6934
rect 57426 6896 57428 6905
rect 57480 6896 57482 6905
rect 57336 6860 57388 6866
rect 57426 6831 57482 6840
rect 57336 6802 57388 6808
rect 57348 6633 57376 6802
rect 57334 6624 57390 6633
rect 57334 6559 57390 6568
rect 57428 6316 57480 6322
rect 57428 6258 57480 6264
rect 57440 5914 57468 6258
rect 57244 5908 57296 5914
rect 57244 5850 57296 5856
rect 57428 5908 57480 5914
rect 57428 5850 57480 5856
rect 57532 5710 57560 6938
rect 57624 6798 57652 7142
rect 57716 7002 57744 8452
rect 57704 6996 57756 7002
rect 57704 6938 57756 6944
rect 57612 6792 57664 6798
rect 57612 6734 57664 6740
rect 57624 6458 57652 6734
rect 57612 6452 57664 6458
rect 57612 6394 57664 6400
rect 57808 6186 57836 8570
rect 57992 8242 58020 9114
rect 57992 8214 58112 8242
rect 57978 8120 58034 8129
rect 57978 8055 58034 8064
rect 57992 7954 58020 8055
rect 57980 7948 58032 7954
rect 57980 7890 58032 7896
rect 57980 7336 58032 7342
rect 57980 7278 58032 7284
rect 57992 6934 58020 7278
rect 57980 6928 58032 6934
rect 57980 6870 58032 6876
rect 57888 6792 57940 6798
rect 57888 6734 57940 6740
rect 57612 6180 57664 6186
rect 57612 6122 57664 6128
rect 57796 6180 57848 6186
rect 57796 6122 57848 6128
rect 57520 5704 57572 5710
rect 57520 5646 57572 5652
rect 57244 5364 57296 5370
rect 57244 5306 57296 5312
rect 57256 4457 57284 5306
rect 57426 5264 57482 5273
rect 57336 5228 57388 5234
rect 57426 5199 57482 5208
rect 57336 5170 57388 5176
rect 57348 4758 57376 5170
rect 57440 4826 57468 5199
rect 57518 5128 57574 5137
rect 57518 5063 57574 5072
rect 57428 4820 57480 4826
rect 57428 4762 57480 4768
rect 57336 4752 57388 4758
rect 57336 4694 57388 4700
rect 57532 4554 57560 5063
rect 57624 4826 57652 6122
rect 57612 4820 57664 4826
rect 57612 4762 57664 4768
rect 57612 4684 57664 4690
rect 57612 4626 57664 4632
rect 57520 4548 57572 4554
rect 57520 4490 57572 4496
rect 57624 4486 57652 4626
rect 57612 4480 57664 4486
rect 57242 4448 57298 4457
rect 57612 4422 57664 4428
rect 57704 4480 57756 4486
rect 57704 4422 57756 4428
rect 57242 4383 57298 4392
rect 57716 4214 57744 4422
rect 57704 4208 57756 4214
rect 57704 4150 57756 4156
rect 57244 3732 57296 3738
rect 57244 3674 57296 3680
rect 57152 3596 57204 3602
rect 57152 3538 57204 3544
rect 56692 3460 56744 3466
rect 56520 3420 56692 3448
rect 56692 3402 56744 3408
rect 56968 3392 57020 3398
rect 56968 3334 57020 3340
rect 57060 3392 57112 3398
rect 57060 3334 57112 3340
rect 56641 3292 56937 3312
rect 56697 3290 56721 3292
rect 56777 3290 56801 3292
rect 56857 3290 56881 3292
rect 56719 3238 56721 3290
rect 56783 3238 56795 3290
rect 56857 3238 56859 3290
rect 56697 3236 56721 3238
rect 56777 3236 56801 3238
rect 56857 3236 56881 3238
rect 56641 3216 56937 3236
rect 56980 3194 57008 3334
rect 56968 3188 57020 3194
rect 56968 3130 57020 3136
rect 56980 2446 57008 3130
rect 57072 3058 57100 3334
rect 57256 3058 57284 3674
rect 57426 3088 57482 3097
rect 57060 3052 57112 3058
rect 57060 2994 57112 3000
rect 57244 3052 57296 3058
rect 57426 3023 57482 3032
rect 57244 2994 57296 3000
rect 57072 2650 57100 2994
rect 57440 2990 57468 3023
rect 57428 2984 57480 2990
rect 57428 2926 57480 2932
rect 57336 2848 57388 2854
rect 57336 2790 57388 2796
rect 57704 2848 57756 2854
rect 57704 2790 57756 2796
rect 57060 2644 57112 2650
rect 57060 2586 57112 2592
rect 57152 2644 57204 2650
rect 57152 2586 57204 2592
rect 56508 2440 56560 2446
rect 56508 2382 56560 2388
rect 56968 2440 57020 2446
rect 56968 2382 57020 2388
rect 56520 1766 56548 2382
rect 56641 2204 56937 2224
rect 56697 2202 56721 2204
rect 56777 2202 56801 2204
rect 56857 2202 56881 2204
rect 56719 2150 56721 2202
rect 56783 2150 56795 2202
rect 56857 2150 56859 2202
rect 56697 2148 56721 2150
rect 56777 2148 56801 2150
rect 56857 2148 56881 2150
rect 56641 2128 56937 2148
rect 56508 1760 56560 1766
rect 56508 1702 56560 1708
rect 56968 1760 57020 1766
rect 56968 1702 57020 1708
rect 56980 1358 57008 1702
rect 56968 1352 57020 1358
rect 56968 1294 57020 1300
rect 56100 1176 56456 1204
rect 56508 1216 56560 1222
rect 56048 1158 56100 1164
rect 56508 1158 56560 1164
rect 56230 1048 56286 1057
rect 56230 983 56286 992
rect 56520 1000 56548 1158
rect 56641 1116 56937 1136
rect 56697 1114 56721 1116
rect 56777 1114 56801 1116
rect 56857 1114 56881 1116
rect 56719 1062 56721 1114
rect 56783 1062 56795 1114
rect 56857 1062 56859 1114
rect 56697 1060 56721 1062
rect 56777 1060 56801 1062
rect 56857 1060 56881 1062
rect 56641 1040 56937 1060
rect 56060 836 56180 864
rect 55494 640 55550 649
rect 55494 575 55550 584
rect 55678 640 55734 649
rect 55678 575 55734 584
rect 55770 0 55826 800
rect 56060 678 56088 836
rect 56152 800 56180 836
rect 56048 672 56100 678
rect 56048 614 56100 620
rect 56138 0 56194 800
rect 56244 678 56272 983
rect 56520 972 56916 1000
rect 56428 836 56548 864
rect 56428 746 56456 836
rect 56520 800 56548 836
rect 56888 800 56916 972
rect 56980 814 57008 1294
rect 56968 808 57020 814
rect 56416 740 56468 746
rect 56416 682 56468 688
rect 56232 672 56284 678
rect 56232 614 56284 620
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 56968 750 57020 756
rect 57164 474 57192 2586
rect 57348 2514 57376 2790
rect 57244 2508 57296 2514
rect 57244 2450 57296 2456
rect 57336 2508 57388 2514
rect 57336 2450 57388 2456
rect 57256 2417 57284 2450
rect 57612 2440 57664 2446
rect 57242 2408 57298 2417
rect 57612 2382 57664 2388
rect 57242 2343 57298 2352
rect 57242 2272 57298 2281
rect 57242 2207 57298 2216
rect 57256 1737 57284 2207
rect 57336 1896 57388 1902
rect 57336 1838 57388 1844
rect 57242 1728 57298 1737
rect 57348 1714 57376 1838
rect 57426 1728 57482 1737
rect 57348 1686 57426 1714
rect 57242 1663 57298 1672
rect 57426 1663 57482 1672
rect 57244 1284 57296 1290
rect 57244 1226 57296 1232
rect 57256 800 57284 1226
rect 57334 912 57390 921
rect 57334 847 57390 856
rect 57152 468 57204 474
rect 57152 410 57204 416
rect 57242 0 57298 800
rect 57348 649 57376 847
rect 57624 800 57652 2382
rect 57716 1970 57744 2790
rect 57900 1970 57928 6734
rect 57980 5092 58032 5098
rect 57980 5034 58032 5040
rect 57992 3126 58020 5034
rect 57980 3120 58032 3126
rect 57980 3062 58032 3068
rect 58084 2922 58112 8214
rect 58176 6798 58204 9574
rect 58348 9172 58400 9178
rect 58348 9114 58400 9120
rect 58360 8974 58388 9114
rect 58348 8968 58400 8974
rect 58348 8910 58400 8916
rect 58544 8820 58572 12200
rect 58806 11928 58862 11937
rect 58806 11863 58862 11872
rect 58624 10464 58676 10470
rect 58624 10406 58676 10412
rect 58636 10062 58664 10406
rect 58624 10056 58676 10062
rect 58624 9998 58676 10004
rect 58820 9586 58848 11863
rect 58912 11286 58940 12200
rect 59280 12050 59308 12200
rect 59004 12022 59308 12050
rect 58900 11280 58952 11286
rect 58900 11222 58952 11228
rect 58808 9580 58860 9586
rect 58808 9522 58860 9528
rect 58544 8792 58664 8820
rect 58532 8628 58584 8634
rect 58532 8570 58584 8576
rect 58256 8560 58308 8566
rect 58544 8514 58572 8570
rect 58308 8508 58572 8514
rect 58256 8502 58572 8508
rect 58268 8486 58572 8502
rect 58348 8424 58400 8430
rect 58348 8366 58400 8372
rect 58360 8129 58388 8366
rect 58346 8120 58402 8129
rect 58346 8055 58402 8064
rect 58440 7948 58492 7954
rect 58636 7936 58664 8792
rect 59004 8498 59032 12022
rect 59084 11280 59136 11286
rect 59084 11222 59136 11228
rect 59096 9654 59124 11222
rect 59464 10674 59492 12446
rect 59634 12200 59690 13000
rect 60002 12200 60058 13000
rect 60370 12200 60426 13000
rect 60554 12200 60610 12209
rect 60738 12200 60794 13000
rect 61106 12200 61162 13000
rect 61292 12572 61344 12578
rect 61292 12514 61344 12520
rect 59544 11144 59596 11150
rect 59544 11086 59596 11092
rect 59452 10668 59504 10674
rect 59452 10610 59504 10616
rect 59464 10130 59492 10610
rect 59556 10305 59584 11086
rect 59542 10296 59598 10305
rect 59542 10231 59598 10240
rect 59452 10124 59504 10130
rect 59452 10066 59504 10072
rect 59360 9716 59412 9722
rect 59648 9704 59676 12200
rect 59728 11552 59780 11558
rect 59728 11494 59780 11500
rect 59740 11150 59768 11494
rect 59728 11144 59780 11150
rect 59728 11086 59780 11092
rect 59820 10056 59872 10062
rect 59360 9658 59412 9664
rect 59464 9676 59676 9704
rect 59740 10016 59820 10044
rect 59084 9648 59136 9654
rect 59084 9590 59136 9596
rect 59372 9586 59400 9658
rect 59360 9580 59412 9586
rect 59360 9522 59412 9528
rect 59084 9376 59136 9382
rect 59084 9318 59136 9324
rect 59096 8498 59124 9318
rect 59372 9178 59400 9522
rect 59360 9172 59412 9178
rect 59360 9114 59412 9120
rect 59464 9024 59492 9676
rect 59544 9376 59596 9382
rect 59544 9318 59596 9324
rect 59280 8996 59492 9024
rect 59176 8832 59228 8838
rect 59176 8774 59228 8780
rect 59188 8514 59216 8774
rect 59280 8634 59308 8996
rect 59452 8832 59504 8838
rect 59452 8774 59504 8780
rect 59464 8634 59492 8774
rect 59268 8628 59320 8634
rect 59268 8570 59320 8576
rect 59452 8628 59504 8634
rect 59452 8570 59504 8576
rect 58992 8492 59044 8498
rect 58992 8434 59044 8440
rect 59084 8492 59136 8498
rect 59188 8486 59400 8514
rect 59084 8434 59136 8440
rect 59004 8090 59032 8434
rect 59176 8424 59228 8430
rect 59176 8366 59228 8372
rect 58992 8084 59044 8090
rect 58992 8026 59044 8032
rect 58492 7908 58664 7936
rect 58440 7890 58492 7896
rect 58348 7880 58400 7886
rect 58348 7822 58400 7828
rect 58360 7206 58388 7822
rect 59084 7744 59136 7750
rect 59084 7686 59136 7692
rect 59096 7342 59124 7686
rect 59084 7336 59136 7342
rect 59084 7278 59136 7284
rect 58348 7200 58400 7206
rect 58348 7142 58400 7148
rect 58256 6860 58308 6866
rect 58256 6802 58308 6808
rect 58164 6792 58216 6798
rect 58164 6734 58216 6740
rect 58268 3738 58296 6802
rect 58360 5642 58388 7142
rect 59096 7002 59124 7278
rect 59084 6996 59136 7002
rect 59084 6938 59136 6944
rect 58532 6792 58584 6798
rect 58532 6734 58584 6740
rect 58544 6390 58572 6734
rect 58532 6384 58584 6390
rect 58532 6326 58584 6332
rect 58348 5636 58400 5642
rect 58348 5578 58400 5584
rect 58992 5568 59044 5574
rect 58992 5510 59044 5516
rect 59004 5098 59032 5510
rect 59188 5386 59216 8366
rect 59372 7886 59400 8486
rect 59360 7880 59412 7886
rect 59360 7822 59412 7828
rect 59452 6656 59504 6662
rect 59452 6598 59504 6604
rect 59464 6390 59492 6598
rect 59452 6384 59504 6390
rect 59452 6326 59504 6332
rect 59268 6316 59320 6322
rect 59268 6258 59320 6264
rect 59280 5574 59308 6258
rect 59268 5568 59320 5574
rect 59268 5510 59320 5516
rect 59188 5358 59400 5386
rect 58992 5092 59044 5098
rect 58992 5034 59044 5040
rect 58532 3936 58584 3942
rect 58532 3878 58584 3884
rect 58716 3936 58768 3942
rect 58716 3878 58768 3884
rect 58256 3732 58308 3738
rect 58256 3674 58308 3680
rect 58440 2984 58492 2990
rect 58346 2952 58402 2961
rect 58072 2916 58124 2922
rect 58440 2926 58492 2932
rect 58346 2887 58402 2896
rect 58072 2858 58124 2864
rect 57704 1964 57756 1970
rect 57704 1906 57756 1912
rect 57888 1964 57940 1970
rect 57888 1906 57940 1912
rect 57704 1828 57756 1834
rect 57704 1770 57756 1776
rect 57716 1426 57744 1770
rect 57796 1760 57848 1766
rect 57796 1702 57848 1708
rect 57704 1420 57756 1426
rect 57704 1362 57756 1368
rect 57808 882 57836 1702
rect 57900 1358 57928 1906
rect 57980 1896 58032 1902
rect 57980 1838 58032 1844
rect 57888 1352 57940 1358
rect 57888 1294 57940 1300
rect 57796 876 57848 882
rect 57796 818 57848 824
rect 57992 800 58020 1838
rect 58360 800 58388 2887
rect 58452 1970 58480 2926
rect 58440 1964 58492 1970
rect 58440 1906 58492 1912
rect 58544 882 58572 3878
rect 58728 3738 58756 3878
rect 58716 3732 58768 3738
rect 58716 3674 58768 3680
rect 58992 3120 59044 3126
rect 58992 3062 59044 3068
rect 58808 3052 58860 3058
rect 58808 2994 58860 3000
rect 58900 3052 58952 3058
rect 58900 2994 58952 3000
rect 58820 2854 58848 2994
rect 58808 2848 58860 2854
rect 58808 2790 58860 2796
rect 58820 2650 58848 2790
rect 58808 2644 58860 2650
rect 58808 2586 58860 2592
rect 58912 2530 58940 2994
rect 59004 2922 59032 3062
rect 58992 2916 59044 2922
rect 58992 2858 59044 2864
rect 58728 2502 58940 2530
rect 58532 876 58584 882
rect 58532 818 58584 824
rect 58728 800 58756 2502
rect 59372 2446 59400 5358
rect 59556 5234 59584 9318
rect 59740 5914 59768 10016
rect 59820 9998 59872 10004
rect 59912 9580 59964 9586
rect 59912 9522 59964 9528
rect 59818 9344 59874 9353
rect 59818 9279 59874 9288
rect 59832 8430 59860 9279
rect 59924 9178 59952 9522
rect 59912 9172 59964 9178
rect 59912 9114 59964 9120
rect 60016 8566 60044 12200
rect 60384 10656 60412 12200
rect 60554 12135 60610 12144
rect 60462 11792 60518 11801
rect 60462 11727 60518 11736
rect 60476 11014 60504 11727
rect 60464 11008 60516 11014
rect 60464 10950 60516 10956
rect 60568 10826 60596 12135
rect 60752 12050 60780 12200
rect 60752 12022 61056 12050
rect 60832 11892 60884 11898
rect 60832 11834 60884 11840
rect 60646 11792 60702 11801
rect 60646 11727 60702 11736
rect 60660 11642 60688 11727
rect 60660 11614 60780 11642
rect 60648 11552 60700 11558
rect 60648 11494 60700 11500
rect 60476 10810 60596 10826
rect 60464 10804 60596 10810
rect 60516 10798 60596 10804
rect 60464 10746 60516 10752
rect 60660 10674 60688 11494
rect 60752 10810 60780 11614
rect 60740 10804 60792 10810
rect 60740 10746 60792 10752
rect 60648 10668 60700 10674
rect 60384 10628 60504 10656
rect 60372 10532 60424 10538
rect 60372 10474 60424 10480
rect 60188 10464 60240 10470
rect 60384 10418 60412 10474
rect 60240 10412 60412 10418
rect 60188 10406 60412 10412
rect 60200 10390 60412 10406
rect 60476 10146 60504 10628
rect 60648 10610 60700 10616
rect 60740 10600 60792 10606
rect 60740 10542 60792 10548
rect 60752 10266 60780 10542
rect 60740 10260 60792 10266
rect 60740 10202 60792 10208
rect 60384 10118 60504 10146
rect 60740 10124 60792 10130
rect 60280 9988 60332 9994
rect 60280 9930 60332 9936
rect 60292 9897 60320 9930
rect 60094 9888 60150 9897
rect 60094 9823 60150 9832
rect 60278 9888 60334 9897
rect 60278 9823 60334 9832
rect 60108 9178 60136 9823
rect 60384 9450 60412 10118
rect 60740 10066 60792 10072
rect 60464 10056 60516 10062
rect 60464 9998 60516 10004
rect 60556 10056 60608 10062
rect 60556 9998 60608 10004
rect 60372 9444 60424 9450
rect 60372 9386 60424 9392
rect 60476 9382 60504 9998
rect 60568 9722 60596 9998
rect 60752 9722 60780 10066
rect 60556 9716 60608 9722
rect 60556 9658 60608 9664
rect 60740 9716 60792 9722
rect 60740 9658 60792 9664
rect 60844 9586 60872 11834
rect 60924 11688 60976 11694
rect 60924 11630 60976 11636
rect 60936 11286 60964 11630
rect 60924 11280 60976 11286
rect 60924 11222 60976 11228
rect 60924 10804 60976 10810
rect 60924 10746 60976 10752
rect 60936 10606 60964 10746
rect 60924 10600 60976 10606
rect 60924 10542 60976 10548
rect 60924 10260 60976 10266
rect 60924 10202 60976 10208
rect 60936 9926 60964 10202
rect 60924 9920 60976 9926
rect 60924 9862 60976 9868
rect 61028 9738 61056 12022
rect 61120 10826 61148 12200
rect 61200 12164 61252 12170
rect 61200 12106 61252 12112
rect 61212 11558 61240 12106
rect 61200 11552 61252 11558
rect 61200 11494 61252 11500
rect 61304 11286 61332 12514
rect 61474 12200 61530 13000
rect 61842 12200 61898 13000
rect 62210 12200 62266 13000
rect 62302 12200 62358 12209
rect 62578 12200 62634 13000
rect 62762 12608 62818 12617
rect 62762 12543 62818 12552
rect 61384 11756 61436 11762
rect 61384 11698 61436 11704
rect 61396 11286 61424 11698
rect 61292 11280 61344 11286
rect 61292 11222 61344 11228
rect 61384 11280 61436 11286
rect 61384 11222 61436 11228
rect 61292 11144 61344 11150
rect 61292 11086 61344 11092
rect 61120 10798 61240 10826
rect 60936 9710 61056 9738
rect 60832 9580 60884 9586
rect 60832 9522 60884 9528
rect 60464 9376 60516 9382
rect 60464 9318 60516 9324
rect 60096 9172 60148 9178
rect 60096 9114 60148 9120
rect 60740 9104 60792 9110
rect 60740 9046 60792 9052
rect 60188 8832 60240 8838
rect 60188 8774 60240 8780
rect 60648 8832 60700 8838
rect 60648 8774 60700 8780
rect 60004 8560 60056 8566
rect 60004 8502 60056 8508
rect 60200 8498 60228 8774
rect 60188 8492 60240 8498
rect 60188 8434 60240 8440
rect 60372 8492 60424 8498
rect 60372 8434 60424 8440
rect 60556 8492 60608 8498
rect 60556 8434 60608 8440
rect 59820 8424 59872 8430
rect 59820 8366 59872 8372
rect 60200 8090 60228 8434
rect 60188 8084 60240 8090
rect 60188 8026 60240 8032
rect 59820 7404 59872 7410
rect 59820 7346 59872 7352
rect 59832 6662 59860 7346
rect 60280 7200 60332 7206
rect 60280 7142 60332 7148
rect 60292 6866 60320 7142
rect 60280 6860 60332 6866
rect 60280 6802 60332 6808
rect 59820 6656 59872 6662
rect 59820 6598 59872 6604
rect 59728 5908 59780 5914
rect 59728 5850 59780 5856
rect 59832 5778 59860 6598
rect 60292 6458 60320 6802
rect 60280 6452 60332 6458
rect 60280 6394 60332 6400
rect 59820 5772 59872 5778
rect 59820 5714 59872 5720
rect 59544 5228 59596 5234
rect 59544 5170 59596 5176
rect 59910 3632 59966 3641
rect 59910 3567 59966 3576
rect 60186 3632 60242 3641
rect 60186 3567 60242 3576
rect 59636 2984 59688 2990
rect 59636 2926 59688 2932
rect 59452 2916 59504 2922
rect 59452 2858 59504 2864
rect 59360 2440 59412 2446
rect 59360 2382 59412 2388
rect 58808 1964 58860 1970
rect 58808 1906 58860 1912
rect 58820 1562 58848 1906
rect 58808 1556 58860 1562
rect 58808 1498 58860 1504
rect 59084 1556 59136 1562
rect 59084 1498 59136 1504
rect 58992 1216 59044 1222
rect 58992 1158 59044 1164
rect 59004 814 59032 1158
rect 58992 808 59044 814
rect 57428 672 57480 678
rect 57334 640 57390 649
rect 57428 614 57480 620
rect 57334 575 57390 584
rect 57440 474 57468 614
rect 57428 468 57480 474
rect 57428 410 57480 416
rect 57610 0 57666 800
rect 57978 0 58034 800
rect 58346 0 58402 800
rect 58714 0 58770 800
rect 59096 800 59124 1498
rect 59464 800 59492 2858
rect 58992 750 59044 756
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59648 678 59676 2926
rect 59728 2508 59780 2514
rect 59728 2450 59780 2456
rect 59820 2508 59872 2514
rect 59820 2450 59872 2456
rect 59740 882 59768 2450
rect 59728 876 59780 882
rect 59728 818 59780 824
rect 59832 800 59860 2450
rect 59924 1902 59952 3567
rect 60096 3528 60148 3534
rect 60096 3470 60148 3476
rect 60004 2372 60056 2378
rect 60004 2314 60056 2320
rect 60016 2106 60044 2314
rect 60004 2100 60056 2106
rect 60004 2042 60056 2048
rect 59912 1896 59964 1902
rect 59912 1838 59964 1844
rect 60108 1766 60136 3470
rect 60096 1760 60148 1766
rect 60096 1702 60148 1708
rect 59912 1420 59964 1426
rect 59912 1362 59964 1368
rect 59924 814 59952 1362
rect 59912 808 59964 814
rect 59636 672 59688 678
rect 59636 614 59688 620
rect 59818 0 59874 800
rect 60200 800 60228 3567
rect 60384 3482 60412 8434
rect 60568 8090 60596 8434
rect 60556 8084 60608 8090
rect 60556 8026 60608 8032
rect 60660 7886 60688 8774
rect 60752 8480 60780 9046
rect 60936 8974 60964 9710
rect 60924 8968 60976 8974
rect 60924 8910 60976 8916
rect 60832 8492 60884 8498
rect 60752 8452 60832 8480
rect 60832 8434 60884 8440
rect 61212 8378 61240 10798
rect 61304 9926 61332 11086
rect 61488 10554 61516 12200
rect 61856 11937 61884 12200
rect 61842 11928 61898 11937
rect 61842 11863 61898 11872
rect 61660 11756 61712 11762
rect 61660 11698 61712 11704
rect 61488 10526 61608 10554
rect 61292 9920 61344 9926
rect 61292 9862 61344 9868
rect 61384 9172 61436 9178
rect 61384 9114 61436 9120
rect 61396 8974 61424 9114
rect 61580 9042 61608 10526
rect 61672 10470 61700 11698
rect 61936 11008 61988 11014
rect 61936 10950 61988 10956
rect 61752 10804 61804 10810
rect 61752 10746 61804 10752
rect 61660 10464 61712 10470
rect 61660 10406 61712 10412
rect 61672 9654 61700 10406
rect 61660 9648 61712 9654
rect 61660 9590 61712 9596
rect 61764 9364 61792 10746
rect 61948 10606 61976 10950
rect 61936 10600 61988 10606
rect 61936 10542 61988 10548
rect 62028 10056 62080 10062
rect 62028 9998 62080 10004
rect 62040 9722 62068 9998
rect 62028 9716 62080 9722
rect 62028 9658 62080 9664
rect 61936 9512 61988 9518
rect 61936 9454 61988 9460
rect 61948 9364 61976 9454
rect 62224 9450 62252 12200
rect 62302 12135 62358 12144
rect 62316 10674 62344 12135
rect 62488 11756 62540 11762
rect 62488 11698 62540 11704
rect 62500 11014 62528 11698
rect 62488 11008 62540 11014
rect 62488 10950 62540 10956
rect 62304 10668 62356 10674
rect 62304 10610 62356 10616
rect 62500 9586 62528 10950
rect 62592 9897 62620 12200
rect 62776 10062 62804 12543
rect 62946 12200 63002 13000
rect 63222 12336 63278 12345
rect 63222 12271 63278 12280
rect 62764 10056 62816 10062
rect 62764 9998 62816 10004
rect 62578 9888 62634 9897
rect 62578 9823 62634 9832
rect 62488 9580 62540 9586
rect 62488 9522 62540 9528
rect 62212 9444 62264 9450
rect 62212 9386 62264 9392
rect 62960 9382 62988 12200
rect 63236 11898 63264 12271
rect 63314 12200 63370 13000
rect 63682 12200 63738 13000
rect 64050 12200 64106 13000
rect 64418 12200 64474 13000
rect 64786 12200 64842 13000
rect 65154 12200 65210 13000
rect 65522 12200 65578 13000
rect 65616 12232 65668 12238
rect 63224 11892 63276 11898
rect 63224 11834 63276 11840
rect 63038 11520 63094 11529
rect 63038 11455 63094 11464
rect 63052 9897 63080 11455
rect 63038 9888 63094 9897
rect 63038 9823 63094 9832
rect 61764 9336 61976 9364
rect 62948 9376 63000 9382
rect 62948 9318 63000 9324
rect 63040 9376 63092 9382
rect 63040 9318 63092 9324
rect 62764 9104 62816 9110
rect 62764 9046 62816 9052
rect 61568 9036 61620 9042
rect 61568 8978 61620 8984
rect 61384 8968 61436 8974
rect 61384 8910 61436 8916
rect 60844 8350 61240 8378
rect 60844 8294 60872 8350
rect 60832 8288 60884 8294
rect 60832 8230 60884 8236
rect 61016 8288 61068 8294
rect 61016 8230 61068 8236
rect 61028 7954 61056 8230
rect 61016 7948 61068 7954
rect 61016 7890 61068 7896
rect 62120 7948 62172 7954
rect 62120 7890 62172 7896
rect 60648 7880 60700 7886
rect 60648 7822 60700 7828
rect 60922 7576 60978 7585
rect 60922 7511 60978 7520
rect 60936 7177 60964 7511
rect 61028 7478 61056 7890
rect 61016 7472 61068 7478
rect 61016 7414 61068 7420
rect 60922 7168 60978 7177
rect 60922 7103 60978 7112
rect 60462 7032 60518 7041
rect 60462 6967 60518 6976
rect 60476 6866 60504 6967
rect 61474 6896 61530 6905
rect 60464 6860 60516 6866
rect 61474 6831 61530 6840
rect 60464 6802 60516 6808
rect 60462 6760 60518 6769
rect 60462 6695 60518 6704
rect 60830 6760 60886 6769
rect 60830 6695 60886 6704
rect 60476 4758 60504 6695
rect 60844 5953 60872 6695
rect 60830 5944 60886 5953
rect 60830 5879 60886 5888
rect 60464 4752 60516 4758
rect 60464 4694 60516 4700
rect 60740 4752 60792 4758
rect 60740 4694 60792 4700
rect 60648 4548 60700 4554
rect 60648 4490 60700 4496
rect 60556 4140 60608 4146
rect 60556 4082 60608 4088
rect 60568 3602 60596 4082
rect 60660 3738 60688 4490
rect 60752 3738 60780 4694
rect 61292 4616 61344 4622
rect 61292 4558 61344 4564
rect 61108 4140 61160 4146
rect 61108 4082 61160 4088
rect 60648 3732 60700 3738
rect 60648 3674 60700 3680
rect 60740 3732 60792 3738
rect 60740 3674 60792 3680
rect 61120 3670 61148 4082
rect 61108 3664 61160 3670
rect 61108 3606 61160 3612
rect 60556 3596 60608 3602
rect 60556 3538 60608 3544
rect 60384 3454 60596 3482
rect 60372 3392 60424 3398
rect 60372 3334 60424 3340
rect 60464 3392 60516 3398
rect 60464 3334 60516 3340
rect 60384 2106 60412 3334
rect 60476 3194 60504 3334
rect 60568 3194 60596 3454
rect 60464 3188 60516 3194
rect 60464 3130 60516 3136
rect 60556 3188 60608 3194
rect 60556 3130 60608 3136
rect 61108 3188 61160 3194
rect 61108 3130 61160 3136
rect 60464 3052 60516 3058
rect 60464 2994 60516 3000
rect 60556 3052 60608 3058
rect 60556 2994 60608 3000
rect 60372 2100 60424 2106
rect 60372 2042 60424 2048
rect 60384 1970 60412 2042
rect 60372 1964 60424 1970
rect 60372 1906 60424 1912
rect 60476 1850 60504 2994
rect 60568 2632 60596 2994
rect 60648 2984 60700 2990
rect 60924 2984 60976 2990
rect 60700 2944 60924 2972
rect 60648 2926 60700 2932
rect 60924 2926 60976 2932
rect 60936 2650 60964 2926
rect 60740 2644 60792 2650
rect 60568 2604 60688 2632
rect 60556 2508 60608 2514
rect 60556 2450 60608 2456
rect 60568 2310 60596 2450
rect 60556 2304 60608 2310
rect 60556 2246 60608 2252
rect 60660 1850 60688 2604
rect 60740 2586 60792 2592
rect 60924 2644 60976 2650
rect 60924 2586 60976 2592
rect 60752 2496 60780 2586
rect 61016 2508 61068 2514
rect 60752 2468 61016 2496
rect 61016 2450 61068 2456
rect 61120 2446 61148 3130
rect 61304 2650 61332 4558
rect 61384 4548 61436 4554
rect 61384 4490 61436 4496
rect 61396 4010 61424 4490
rect 61488 4282 61516 6831
rect 62132 5545 62160 7890
rect 62118 5536 62174 5545
rect 62118 5471 62174 5480
rect 62302 5264 62358 5273
rect 62302 5199 62358 5208
rect 61476 4276 61528 4282
rect 61476 4218 61528 4224
rect 62212 4140 62264 4146
rect 62212 4082 62264 4088
rect 61384 4004 61436 4010
rect 61384 3946 61436 3952
rect 62224 3466 62252 4082
rect 62028 3460 62080 3466
rect 62028 3402 62080 3408
rect 62212 3460 62264 3466
rect 62212 3402 62264 3408
rect 61566 2952 61622 2961
rect 61566 2887 61622 2896
rect 61292 2644 61344 2650
rect 61292 2586 61344 2592
rect 61476 2576 61528 2582
rect 61396 2524 61476 2530
rect 61396 2518 61528 2524
rect 61396 2514 61516 2518
rect 61384 2508 61516 2514
rect 61436 2502 61516 2508
rect 61384 2450 61436 2456
rect 61108 2440 61160 2446
rect 61108 2382 61160 2388
rect 60832 2100 60884 2106
rect 60832 2042 60884 2048
rect 60740 1964 60792 1970
rect 60740 1906 60792 1912
rect 60384 1822 60504 1850
rect 60568 1822 60688 1850
rect 60280 1284 60332 1290
rect 60280 1226 60332 1232
rect 60292 1193 60320 1226
rect 60278 1184 60334 1193
rect 60278 1119 60334 1128
rect 59912 750 59964 756
rect 60186 0 60242 800
rect 60384 746 60412 1822
rect 60568 1748 60596 1822
rect 60476 1720 60596 1748
rect 60646 1728 60702 1737
rect 60476 882 60504 1720
rect 60646 1663 60702 1672
rect 60660 1290 60688 1663
rect 60648 1284 60700 1290
rect 60648 1226 60700 1232
rect 60752 1222 60780 1906
rect 60844 1426 60872 2042
rect 61580 1970 61608 2887
rect 61752 2508 61804 2514
rect 61752 2450 61804 2456
rect 61660 2440 61712 2446
rect 61660 2382 61712 2388
rect 61568 1964 61620 1970
rect 61568 1906 61620 1912
rect 61016 1896 61068 1902
rect 61016 1838 61068 1844
rect 60922 1728 60978 1737
rect 60922 1663 60978 1672
rect 60832 1420 60884 1426
rect 60832 1362 60884 1368
rect 60740 1216 60792 1222
rect 60740 1158 60792 1164
rect 60464 876 60516 882
rect 60464 818 60516 824
rect 60568 836 60688 864
rect 60568 800 60596 836
rect 60372 740 60424 746
rect 60372 682 60424 688
rect 60464 672 60516 678
rect 60462 640 60464 649
rect 60516 640 60518 649
rect 60462 575 60518 584
rect 60554 0 60610 800
rect 60660 678 60688 836
rect 60936 800 60964 1663
rect 61028 1358 61056 1838
rect 61580 1562 61608 1906
rect 61568 1556 61620 1562
rect 61568 1498 61620 1504
rect 61016 1352 61068 1358
rect 61016 1294 61068 1300
rect 61200 1284 61252 1290
rect 61200 1226 61252 1232
rect 61212 1193 61240 1226
rect 61476 1216 61528 1222
rect 61198 1184 61254 1193
rect 61382 1184 61438 1193
rect 61198 1119 61254 1128
rect 61304 1142 61382 1170
rect 61304 800 61332 1142
rect 61476 1158 61528 1164
rect 61382 1119 61438 1128
rect 61488 882 61516 1158
rect 61476 876 61528 882
rect 61476 818 61528 824
rect 61672 800 61700 2382
rect 61764 2038 61792 2450
rect 61752 2032 61804 2038
rect 61752 1974 61804 1980
rect 62040 800 62068 3402
rect 62316 3194 62344 5199
rect 62672 5160 62724 5166
rect 62672 5102 62724 5108
rect 62488 5024 62540 5030
rect 62488 4966 62540 4972
rect 62500 3398 62528 4966
rect 62488 3392 62540 3398
rect 62488 3334 62540 3340
rect 62684 3194 62712 5102
rect 62776 4146 62804 9046
rect 63052 8634 63080 9318
rect 63328 9042 63356 12200
rect 63590 11792 63646 11801
rect 63590 11727 63646 11736
rect 63604 11150 63632 11727
rect 63408 11144 63460 11150
rect 63408 11086 63460 11092
rect 63592 11144 63644 11150
rect 63592 11086 63644 11092
rect 63420 10996 63448 11086
rect 63420 10968 63540 10996
rect 63512 9654 63540 10968
rect 63500 9648 63552 9654
rect 63696 9625 63724 12200
rect 63776 10804 63828 10810
rect 63776 10746 63828 10752
rect 63788 10305 63816 10746
rect 63774 10296 63830 10305
rect 63774 10231 63830 10240
rect 63500 9590 63552 9596
rect 63682 9616 63738 9625
rect 63682 9551 63738 9560
rect 63316 9036 63368 9042
rect 63316 8978 63368 8984
rect 63408 8968 63460 8974
rect 63408 8910 63460 8916
rect 63420 8634 63448 8910
rect 63040 8628 63092 8634
rect 63040 8570 63092 8576
rect 63408 8628 63460 8634
rect 63408 8570 63460 8576
rect 64064 8537 64092 12200
rect 64236 10260 64288 10266
rect 64236 10202 64288 10208
rect 64248 9722 64276 10202
rect 64236 9716 64288 9722
rect 64432 9704 64460 12200
rect 64512 12096 64564 12102
rect 64512 12038 64564 12044
rect 64524 11558 64552 12038
rect 64696 11756 64748 11762
rect 64696 11698 64748 11704
rect 64512 11552 64564 11558
rect 64512 11494 64564 11500
rect 64708 11150 64736 11698
rect 64696 11144 64748 11150
rect 64696 11086 64748 11092
rect 64236 9658 64288 9664
rect 64340 9676 64460 9704
rect 64050 8528 64106 8537
rect 64050 8463 64106 8472
rect 62856 8424 62908 8430
rect 62856 8366 62908 8372
rect 63868 8424 63920 8430
rect 63868 8366 63920 8372
rect 62868 8090 62896 8366
rect 62856 8084 62908 8090
rect 62856 8026 62908 8032
rect 63880 7410 63908 8366
rect 64340 8362 64368 9676
rect 64800 8838 64828 12200
rect 65168 11914 65196 12200
rect 65536 12073 65564 12200
rect 65890 12200 65946 13000
rect 66076 12980 66128 12986
rect 66076 12922 66128 12928
rect 65616 12174 65668 12180
rect 65522 12064 65578 12073
rect 65522 11999 65578 12008
rect 65076 11886 65196 11914
rect 64788 8832 64840 8838
rect 64788 8774 64840 8780
rect 65076 8566 65104 11886
rect 65628 11830 65656 12174
rect 65616 11824 65668 11830
rect 65616 11766 65668 11772
rect 65156 11756 65208 11762
rect 65156 11698 65208 11704
rect 65168 11082 65196 11698
rect 65904 11694 65932 12200
rect 66088 12152 66116 12922
rect 66258 12200 66314 13000
rect 66352 12640 66404 12646
rect 66352 12582 66404 12588
rect 66272 12152 66300 12200
rect 66088 12124 66300 12152
rect 65892 11688 65944 11694
rect 65892 11630 65944 11636
rect 65156 11076 65208 11082
rect 65156 11018 65208 11024
rect 65248 11008 65300 11014
rect 65248 10950 65300 10956
rect 65340 11008 65392 11014
rect 65340 10950 65392 10956
rect 66166 10976 66222 10985
rect 65260 10606 65288 10950
rect 65352 10674 65380 10950
rect 66166 10911 66222 10920
rect 65340 10668 65392 10674
rect 65340 10610 65392 10616
rect 65248 10600 65300 10606
rect 65248 10542 65300 10548
rect 65260 10266 65288 10542
rect 66180 10538 66208 10911
rect 66260 10668 66312 10674
rect 66260 10610 66312 10616
rect 66168 10532 66220 10538
rect 66168 10474 66220 10480
rect 65248 10260 65300 10266
rect 65248 10202 65300 10208
rect 66272 9926 66300 10610
rect 66364 10538 66392 12582
rect 66626 12200 66682 13000
rect 66994 12200 67050 13000
rect 67362 12200 67418 13000
rect 67730 12200 67786 13000
rect 67824 12300 67876 12306
rect 67824 12242 67876 12248
rect 66352 10532 66404 10538
rect 66352 10474 66404 10480
rect 66260 9920 66312 9926
rect 66260 9862 66312 9868
rect 66272 8566 66300 9862
rect 65064 8560 65116 8566
rect 65064 8502 65116 8508
rect 66260 8560 66312 8566
rect 66260 8502 66312 8508
rect 64420 8492 64472 8498
rect 64420 8434 64472 8440
rect 64328 8356 64380 8362
rect 64328 8298 64380 8304
rect 64432 7818 64460 8434
rect 66640 8129 66668 12200
rect 67008 9518 67036 12200
rect 66996 9512 67048 9518
rect 66996 9454 67048 9460
rect 67376 8906 67404 12200
rect 67744 12152 67772 12200
rect 67836 12152 67864 12242
rect 68098 12200 68154 13000
rect 68466 12200 68522 13000
rect 68834 12200 68890 13000
rect 69202 12200 69258 13000
rect 69570 12200 69626 13000
rect 69938 12200 69994 13000
rect 70306 12200 70362 13000
rect 70674 12200 70730 13000
rect 70860 12912 70912 12918
rect 70860 12854 70912 12860
rect 67744 12124 67864 12152
rect 68008 12164 68060 12170
rect 68008 12106 68060 12112
rect 67824 11688 67876 11694
rect 67824 11630 67876 11636
rect 67916 11688 67968 11694
rect 67916 11630 67968 11636
rect 67836 10674 67864 11630
rect 67928 11150 67956 11630
rect 67916 11144 67968 11150
rect 67916 11086 67968 11092
rect 67824 10668 67876 10674
rect 67824 10610 67876 10616
rect 67364 8900 67416 8906
rect 67364 8842 67416 8848
rect 66626 8120 66682 8129
rect 66626 8055 66682 8064
rect 68020 7954 68048 12106
rect 68112 8430 68140 12200
rect 68480 9382 68508 12200
rect 68744 10668 68796 10674
rect 68744 10610 68796 10616
rect 68756 10266 68784 10610
rect 68744 10260 68796 10266
rect 68744 10202 68796 10208
rect 68848 9654 68876 12200
rect 69020 11552 69072 11558
rect 69020 11494 69072 11500
rect 68928 11144 68980 11150
rect 68928 11086 68980 11092
rect 68940 10130 68968 11086
rect 69032 10441 69060 11494
rect 69018 10432 69074 10441
rect 69018 10367 69074 10376
rect 68928 10124 68980 10130
rect 68928 10066 68980 10072
rect 68836 9648 68888 9654
rect 68836 9590 68888 9596
rect 69112 9580 69164 9586
rect 69216 9568 69244 12200
rect 69294 11384 69350 11393
rect 69294 11319 69350 11328
rect 69308 10441 69336 11319
rect 69584 11082 69612 12200
rect 69952 11286 69980 12200
rect 70320 11762 70348 12200
rect 70308 11756 70360 11762
rect 70308 11698 70360 11704
rect 69940 11280 69992 11286
rect 69940 11222 69992 11228
rect 70320 11150 70348 11698
rect 70492 11688 70544 11694
rect 70492 11630 70544 11636
rect 70308 11144 70360 11150
rect 70308 11086 70360 11092
rect 69572 11076 69624 11082
rect 69572 11018 69624 11024
rect 70504 10674 70532 11630
rect 70584 11552 70636 11558
rect 70584 11494 70636 11500
rect 70596 11150 70624 11494
rect 70584 11144 70636 11150
rect 70584 11086 70636 11092
rect 69388 10668 69440 10674
rect 69388 10610 69440 10616
rect 70492 10668 70544 10674
rect 70492 10610 70544 10616
rect 69294 10432 69350 10441
rect 69294 10367 69350 10376
rect 69400 10266 69428 10610
rect 70504 10266 70532 10610
rect 69388 10260 69440 10266
rect 69388 10202 69440 10208
rect 70492 10260 70544 10266
rect 70492 10202 70544 10208
rect 70596 9586 70624 11086
rect 70688 10742 70716 12200
rect 70768 11348 70820 11354
rect 70768 11290 70820 11296
rect 70676 10736 70728 10742
rect 70676 10678 70728 10684
rect 69164 9540 69244 9568
rect 70584 9580 70636 9586
rect 69112 9522 69164 9528
rect 70584 9522 70636 9528
rect 68468 9376 68520 9382
rect 68468 9318 68520 9324
rect 70780 8673 70808 11290
rect 70872 10266 70900 12854
rect 71042 12200 71098 13000
rect 71410 12200 71466 13000
rect 71778 12200 71834 13000
rect 72146 12200 72202 13000
rect 72424 12300 72476 12306
rect 72424 12242 72476 12248
rect 71056 11132 71084 12200
rect 71136 11144 71188 11150
rect 71056 11104 71136 11132
rect 71136 11086 71188 11092
rect 70860 10260 70912 10266
rect 70860 10202 70912 10208
rect 71424 10062 71452 12200
rect 71792 11778 71820 12200
rect 71792 11762 71912 11778
rect 71688 11756 71740 11762
rect 71792 11756 71924 11762
rect 71792 11750 71872 11756
rect 71688 11698 71740 11704
rect 71872 11698 71924 11704
rect 71700 11642 71728 11698
rect 71700 11614 71820 11642
rect 71792 10810 71820 11614
rect 71688 10804 71740 10810
rect 71688 10746 71740 10752
rect 71780 10804 71832 10810
rect 71780 10746 71832 10752
rect 71504 10532 71556 10538
rect 71504 10474 71556 10480
rect 70860 10056 70912 10062
rect 70860 9998 70912 10004
rect 71412 10056 71464 10062
rect 71412 9998 71464 10004
rect 70872 9654 70900 9998
rect 71516 9761 71544 10474
rect 71502 9752 71558 9761
rect 71700 9722 71728 10746
rect 71502 9687 71558 9696
rect 71688 9716 71740 9722
rect 71688 9658 71740 9664
rect 71792 9654 71820 10746
rect 72056 10532 72108 10538
rect 72056 10474 72108 10480
rect 72068 10130 72096 10474
rect 72056 10124 72108 10130
rect 72160 10112 72188 12200
rect 72332 11756 72384 11762
rect 72332 11698 72384 11704
rect 72344 11354 72372 11698
rect 72332 11348 72384 11354
rect 72332 11290 72384 11296
rect 72436 11218 72464 12242
rect 72514 12200 72570 13000
rect 72882 12200 72938 13000
rect 73250 12200 73306 13000
rect 73618 12200 73674 13000
rect 73986 12200 74042 13000
rect 74354 12200 74410 13000
rect 74722 12200 74778 13000
rect 75000 12368 75052 12374
rect 75000 12310 75052 12316
rect 72424 11212 72476 11218
rect 72424 11154 72476 11160
rect 72528 10742 72556 12200
rect 72896 11694 72924 12200
rect 72884 11688 72936 11694
rect 72884 11630 72936 11636
rect 72792 11552 72844 11558
rect 72792 11494 72844 11500
rect 72804 11218 72832 11494
rect 72792 11212 72844 11218
rect 72792 11154 72844 11160
rect 72516 10736 72568 10742
rect 72516 10678 72568 10684
rect 72424 10464 72476 10470
rect 72424 10406 72476 10412
rect 72240 10124 72292 10130
rect 72160 10084 72240 10112
rect 72056 10066 72108 10072
rect 72240 10066 72292 10072
rect 72436 10062 72464 10406
rect 72424 10056 72476 10062
rect 72424 9998 72476 10004
rect 72608 10056 72660 10062
rect 72608 9998 72660 10004
rect 70860 9648 70912 9654
rect 70860 9590 70912 9596
rect 71780 9648 71832 9654
rect 71780 9590 71832 9596
rect 72436 9042 72464 9998
rect 72620 9081 72648 9998
rect 72804 9654 72832 11154
rect 73264 10810 73292 12200
rect 73632 12102 73660 12200
rect 73620 12096 73672 12102
rect 73620 12038 73672 12044
rect 73528 11212 73580 11218
rect 73528 11154 73580 11160
rect 73252 10804 73304 10810
rect 73252 10746 73304 10752
rect 72792 9648 72844 9654
rect 72792 9590 72844 9596
rect 72606 9072 72662 9081
rect 72424 9036 72476 9042
rect 72606 9007 72662 9016
rect 72424 8978 72476 8984
rect 70766 8664 70822 8673
rect 70766 8599 70822 8608
rect 68100 8424 68152 8430
rect 68100 8366 68152 8372
rect 71780 8424 71832 8430
rect 71780 8366 71832 8372
rect 69846 8256 69902 8265
rect 69846 8191 69902 8200
rect 68008 7948 68060 7954
rect 68008 7890 68060 7896
rect 67546 7848 67602 7857
rect 64420 7812 64472 7818
rect 67546 7783 67602 7792
rect 64420 7754 64472 7760
rect 63868 7404 63920 7410
rect 63868 7346 63920 7352
rect 63408 6860 63460 6866
rect 63408 6802 63460 6808
rect 65432 6860 65484 6866
rect 65432 6802 65484 6808
rect 63316 5704 63368 5710
rect 63316 5646 63368 5652
rect 63328 5234 63356 5646
rect 63316 5228 63368 5234
rect 63316 5170 63368 5176
rect 63420 5166 63448 6802
rect 64512 6656 64564 6662
rect 64512 6598 64564 6604
rect 64524 6322 64552 6598
rect 64602 6488 64658 6497
rect 64602 6423 64658 6432
rect 63868 6316 63920 6322
rect 63868 6258 63920 6264
rect 64512 6316 64564 6322
rect 64512 6258 64564 6264
rect 63880 5370 63908 6258
rect 64524 5914 64552 6258
rect 64512 5908 64564 5914
rect 64512 5850 64564 5856
rect 64420 5568 64472 5574
rect 64420 5510 64472 5516
rect 63868 5364 63920 5370
rect 63868 5306 63920 5312
rect 63408 5160 63460 5166
rect 63408 5102 63460 5108
rect 63866 5128 63922 5137
rect 63866 5063 63922 5072
rect 63314 4856 63370 4865
rect 63314 4791 63370 4800
rect 62854 4312 62910 4321
rect 62854 4247 62910 4256
rect 62764 4140 62816 4146
rect 62764 4082 62816 4088
rect 62764 3528 62816 3534
rect 62764 3470 62816 3476
rect 62776 3398 62804 3470
rect 62764 3392 62816 3398
rect 62764 3334 62816 3340
rect 62304 3188 62356 3194
rect 62304 3130 62356 3136
rect 62672 3188 62724 3194
rect 62672 3130 62724 3136
rect 62396 3052 62448 3058
rect 62396 2994 62448 3000
rect 62408 2310 62436 2994
rect 62578 2952 62634 2961
rect 62578 2887 62634 2896
rect 62764 2916 62816 2922
rect 62592 2650 62620 2887
rect 62764 2858 62816 2864
rect 62580 2644 62632 2650
rect 62580 2586 62632 2592
rect 62212 2304 62264 2310
rect 62212 2246 62264 2252
rect 62396 2304 62448 2310
rect 62396 2246 62448 2252
rect 62224 1834 62252 2246
rect 62212 1828 62264 1834
rect 62212 1770 62264 1776
rect 62120 1760 62172 1766
rect 62120 1702 62172 1708
rect 62132 1562 62160 1702
rect 62120 1556 62172 1562
rect 62120 1498 62172 1504
rect 62304 1352 62356 1358
rect 62304 1294 62356 1300
rect 62316 1222 62344 1294
rect 62304 1216 62356 1222
rect 62304 1158 62356 1164
rect 62408 800 62436 2246
rect 62488 1964 62540 1970
rect 62488 1906 62540 1912
rect 62500 1562 62528 1906
rect 62672 1896 62724 1902
rect 62672 1838 62724 1844
rect 62488 1556 62540 1562
rect 62488 1498 62540 1504
rect 62684 1222 62712 1838
rect 62672 1216 62724 1222
rect 62672 1158 62724 1164
rect 62776 800 62804 2858
rect 62868 2650 62896 4247
rect 63328 4146 63356 4791
rect 63684 4684 63736 4690
rect 63684 4626 63736 4632
rect 62948 4140 63000 4146
rect 62948 4082 63000 4088
rect 63224 4140 63276 4146
rect 63224 4082 63276 4088
rect 63316 4140 63368 4146
rect 63316 4082 63368 4088
rect 62960 3534 62988 4082
rect 63236 3602 63264 4082
rect 63592 3664 63644 3670
rect 63592 3606 63644 3612
rect 63040 3596 63092 3602
rect 63040 3538 63092 3544
rect 63224 3596 63276 3602
rect 63224 3538 63276 3544
rect 62948 3528 63000 3534
rect 62948 3470 63000 3476
rect 62856 2644 62908 2650
rect 62856 2586 62908 2592
rect 62856 1964 62908 1970
rect 62856 1906 62908 1912
rect 62868 1426 62896 1906
rect 63052 1902 63080 3538
rect 63500 3052 63552 3058
rect 63500 2994 63552 3000
rect 63512 2922 63540 2994
rect 63500 2916 63552 2922
rect 63500 2858 63552 2864
rect 63224 2848 63276 2854
rect 63224 2790 63276 2796
rect 63236 2514 63264 2790
rect 63512 2650 63540 2858
rect 63500 2644 63552 2650
rect 63500 2586 63552 2592
rect 63224 2508 63276 2514
rect 63224 2450 63276 2456
rect 63316 2508 63368 2514
rect 63316 2450 63368 2456
rect 63040 1896 63092 1902
rect 63040 1838 63092 1844
rect 63328 1562 63356 2450
rect 63500 2440 63552 2446
rect 63500 2382 63552 2388
rect 63512 2310 63540 2382
rect 63500 2304 63552 2310
rect 63500 2246 63552 2252
rect 63500 1964 63552 1970
rect 63420 1924 63500 1952
rect 63316 1556 63368 1562
rect 63316 1498 63368 1504
rect 63420 1442 63448 1924
rect 63500 1906 63552 1912
rect 63604 1850 63632 3606
rect 63696 2650 63724 4626
rect 63880 3670 63908 5063
rect 64432 5030 64460 5510
rect 64420 5024 64472 5030
rect 64420 4966 64472 4972
rect 64616 4282 64644 6423
rect 65444 5846 65472 6802
rect 66076 6316 66128 6322
rect 66076 6258 66128 6264
rect 65524 6248 65576 6254
rect 65522 6216 65524 6225
rect 65576 6216 65578 6225
rect 65522 6151 65578 6160
rect 65432 5840 65484 5846
rect 65432 5782 65484 5788
rect 66088 5574 66116 6258
rect 66812 5772 66864 5778
rect 66812 5714 66864 5720
rect 66076 5568 66128 5574
rect 66076 5510 66128 5516
rect 64694 5400 64750 5409
rect 64694 5335 64750 5344
rect 64604 4276 64656 4282
rect 64604 4218 64656 4224
rect 64420 4072 64472 4078
rect 64420 4014 64472 4020
rect 64052 3936 64104 3942
rect 64052 3878 64104 3884
rect 63868 3664 63920 3670
rect 63774 3632 63830 3641
rect 63868 3606 63920 3612
rect 63774 3567 63830 3576
rect 63788 3058 63816 3567
rect 63776 3052 63828 3058
rect 63776 2994 63828 3000
rect 63960 2984 64012 2990
rect 63960 2926 64012 2932
rect 63684 2644 63736 2650
rect 63684 2586 63736 2592
rect 63776 2100 63828 2106
rect 63776 2042 63828 2048
rect 63684 2032 63736 2038
rect 63684 1974 63736 1980
rect 62856 1420 62908 1426
rect 62856 1362 62908 1368
rect 63144 1414 63448 1442
rect 63512 1822 63632 1850
rect 63144 800 63172 1414
rect 63512 800 63540 1822
rect 63696 1426 63724 1974
rect 63788 1562 63816 2042
rect 63776 1556 63828 1562
rect 63776 1498 63828 1504
rect 63684 1420 63736 1426
rect 63684 1362 63736 1368
rect 63972 1358 64000 2926
rect 63776 1352 63828 1358
rect 63776 1294 63828 1300
rect 63960 1352 64012 1358
rect 63960 1294 64012 1300
rect 63788 882 63816 1294
rect 64064 1170 64092 3878
rect 64236 3460 64288 3466
rect 64236 3402 64288 3408
rect 63880 1142 64092 1170
rect 63776 876 63828 882
rect 63776 818 63828 824
rect 63880 800 63908 1142
rect 64248 800 64276 3402
rect 64432 3194 64460 4014
rect 64604 3936 64656 3942
rect 64604 3878 64656 3884
rect 64420 3188 64472 3194
rect 64420 3130 64472 3136
rect 64512 3188 64564 3194
rect 64512 3130 64564 3136
rect 64524 3058 64552 3130
rect 64512 3052 64564 3058
rect 64512 2994 64564 3000
rect 64524 2650 64552 2994
rect 64616 2854 64644 3878
rect 64604 2848 64656 2854
rect 64604 2790 64656 2796
rect 64512 2644 64564 2650
rect 64512 2586 64564 2592
rect 64708 2106 64736 5335
rect 66536 5228 66588 5234
rect 66536 5170 66588 5176
rect 65064 5092 65116 5098
rect 65064 5034 65116 5040
rect 64972 2304 65024 2310
rect 64972 2246 65024 2252
rect 64696 2100 64748 2106
rect 64696 2042 64748 2048
rect 64604 1896 64656 1902
rect 64604 1838 64656 1844
rect 64616 800 64644 1838
rect 64984 800 65012 2246
rect 65076 2106 65104 5034
rect 66444 4480 66496 4486
rect 66444 4422 66496 4428
rect 65248 3596 65300 3602
rect 65248 3538 65300 3544
rect 65064 2100 65116 2106
rect 65064 2042 65116 2048
rect 65260 1442 65288 3538
rect 66076 3392 66128 3398
rect 66076 3334 66128 3340
rect 66352 3392 66404 3398
rect 66352 3334 66404 3340
rect 65708 3120 65760 3126
rect 65708 3062 65760 3068
rect 65984 3120 66036 3126
rect 65984 3062 66036 3068
rect 65340 2984 65392 2990
rect 65340 2926 65392 2932
rect 65352 2038 65380 2926
rect 65340 2032 65392 2038
rect 65340 1974 65392 1980
rect 65432 2032 65484 2038
rect 65432 1974 65484 1980
rect 65260 1414 65380 1442
rect 65156 1216 65208 1222
rect 65156 1158 65208 1164
rect 65168 950 65196 1158
rect 65156 944 65208 950
rect 65156 886 65208 892
rect 65352 800 65380 1414
rect 60648 672 60700 678
rect 60648 614 60700 620
rect 60922 0 60978 800
rect 61200 740 61252 746
rect 61200 682 61252 688
rect 61212 649 61240 682
rect 61198 640 61254 649
rect 61198 575 61254 584
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65064 740 65116 746
rect 65064 682 65116 688
rect 65076 105 65104 682
rect 65062 96 65118 105
rect 65062 31 65118 40
rect 65338 0 65394 800
rect 65444 678 65472 1974
rect 65616 1964 65668 1970
rect 65616 1906 65668 1912
rect 65522 1728 65578 1737
rect 65522 1663 65578 1672
rect 65536 678 65564 1663
rect 65628 1426 65656 1906
rect 65616 1420 65668 1426
rect 65616 1362 65668 1368
rect 65720 800 65748 3062
rect 65996 1358 66024 3062
rect 65984 1352 66036 1358
rect 65984 1294 66036 1300
rect 66088 800 66116 3334
rect 66364 950 66392 3334
rect 66352 944 66404 950
rect 66352 886 66404 892
rect 66456 800 66484 4422
rect 66548 2650 66576 5170
rect 66720 2984 66772 2990
rect 66720 2926 66772 2932
rect 66536 2644 66588 2650
rect 66536 2586 66588 2592
rect 66732 1766 66760 2926
rect 66824 2106 66852 5714
rect 67088 5364 67140 5370
rect 67088 5306 67140 5312
rect 66902 2952 66958 2961
rect 66902 2887 66958 2896
rect 66916 2106 66944 2887
rect 66812 2100 66864 2106
rect 66812 2042 66864 2048
rect 66904 2100 66956 2106
rect 66904 2042 66956 2048
rect 66812 1896 66864 1902
rect 66812 1838 66864 1844
rect 66628 1760 66680 1766
rect 66628 1702 66680 1708
rect 66720 1760 66772 1766
rect 66720 1702 66772 1708
rect 66640 1578 66668 1702
rect 66824 1578 66852 1838
rect 66640 1550 66852 1578
rect 66812 1420 66864 1426
rect 66812 1362 66864 1368
rect 66824 800 66852 1362
rect 67100 1358 67128 5306
rect 67454 3496 67510 3505
rect 67454 3431 67456 3440
rect 67508 3431 67510 3440
rect 67456 3402 67508 3408
rect 67454 3224 67510 3233
rect 67454 3159 67510 3168
rect 67180 2916 67232 2922
rect 67180 2858 67232 2864
rect 67364 2916 67416 2922
rect 67364 2858 67416 2864
rect 67088 1352 67140 1358
rect 67088 1294 67140 1300
rect 66904 1284 66956 1290
rect 66904 1226 66956 1232
rect 66916 1170 66944 1226
rect 67088 1216 67140 1222
rect 66916 1164 67088 1170
rect 66916 1158 67140 1164
rect 66916 1142 67128 1158
rect 67192 800 67220 2858
rect 67376 1970 67404 2858
rect 67364 1964 67416 1970
rect 67364 1906 67416 1912
rect 67272 1760 67324 1766
rect 67272 1702 67324 1708
rect 67284 1358 67312 1702
rect 67376 1426 67404 1906
rect 67468 1442 67496 3159
rect 67560 2650 67588 7783
rect 67732 7744 67784 7750
rect 67732 7686 67784 7692
rect 68836 7744 68888 7750
rect 68836 7686 68888 7692
rect 67640 5296 67692 5302
rect 67640 5238 67692 5244
rect 67652 3534 67680 5238
rect 67640 3528 67692 3534
rect 67640 3470 67692 3476
rect 67744 2854 67772 7686
rect 68848 7410 68876 7686
rect 68836 7404 68888 7410
rect 68836 7346 68888 7352
rect 68848 7002 68876 7346
rect 69860 7342 69888 8191
rect 71792 8090 71820 8366
rect 71780 8084 71832 8090
rect 71780 8026 71832 8032
rect 71792 7954 71820 8026
rect 72790 7984 72846 7993
rect 71780 7948 71832 7954
rect 72790 7919 72792 7928
rect 71780 7890 71832 7896
rect 72844 7919 72846 7928
rect 72792 7890 72844 7896
rect 72884 7880 72936 7886
rect 72884 7822 72936 7828
rect 71136 7812 71188 7818
rect 71136 7754 71188 7760
rect 70124 7404 70176 7410
rect 70124 7346 70176 7352
rect 69848 7336 69900 7342
rect 69848 7278 69900 7284
rect 70136 7002 70164 7346
rect 68836 6996 68888 7002
rect 68836 6938 68888 6944
rect 70124 6996 70176 7002
rect 70124 6938 70176 6944
rect 69294 6760 69350 6769
rect 69294 6695 69350 6704
rect 69112 5636 69164 5642
rect 69112 5578 69164 5584
rect 68284 4208 68336 4214
rect 68284 4150 68336 4156
rect 67732 2848 67784 2854
rect 67732 2790 67784 2796
rect 67548 2644 67600 2650
rect 67548 2586 67600 2592
rect 67548 2304 67600 2310
rect 68008 2304 68060 2310
rect 67600 2264 67956 2292
rect 67548 2246 67600 2252
rect 67732 2100 67784 2106
rect 67732 2042 67784 2048
rect 67744 1766 67772 2042
rect 67732 1760 67784 1766
rect 67732 1702 67784 1708
rect 67364 1420 67416 1426
rect 67468 1414 67588 1442
rect 67364 1362 67416 1368
rect 67272 1352 67324 1358
rect 67272 1294 67324 1300
rect 67560 800 67588 1414
rect 67928 800 67956 2264
rect 68008 2246 68060 2252
rect 68020 1329 68048 2246
rect 68100 1964 68152 1970
rect 68100 1906 68152 1912
rect 68006 1320 68062 1329
rect 68006 1255 68062 1264
rect 65616 740 65668 746
rect 65616 682 65668 688
rect 65432 672 65484 678
rect 65432 614 65484 620
rect 65524 672 65576 678
rect 65524 614 65576 620
rect 65628 105 65656 682
rect 65614 96 65670 105
rect 65614 31 65670 40
rect 65706 0 65762 800
rect 66074 0 66130 800
rect 66442 0 66498 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68112 746 68140 1906
rect 68296 800 68324 4150
rect 68744 4140 68796 4146
rect 68744 4082 68796 4088
rect 68756 3398 68784 4082
rect 68836 3664 68888 3670
rect 68836 3606 68888 3612
rect 68744 3392 68796 3398
rect 68744 3334 68796 3340
rect 68376 3052 68428 3058
rect 68376 2994 68428 3000
rect 68388 2961 68416 2994
rect 68560 2984 68612 2990
rect 68374 2952 68430 2961
rect 68560 2926 68612 2932
rect 68374 2887 68430 2896
rect 68572 2650 68600 2926
rect 68560 2644 68612 2650
rect 68560 2586 68612 2592
rect 68756 1737 68784 3334
rect 68558 1728 68614 1737
rect 68558 1663 68614 1672
rect 68742 1728 68798 1737
rect 68742 1663 68798 1672
rect 68572 1426 68600 1663
rect 68560 1420 68612 1426
rect 68560 1362 68612 1368
rect 68744 1420 68796 1426
rect 68744 1362 68796 1368
rect 68652 1216 68704 1222
rect 68652 1158 68704 1164
rect 68664 800 68692 1158
rect 68756 950 68784 1362
rect 68848 950 68876 3606
rect 69020 3596 69072 3602
rect 69020 3538 69072 3544
rect 68744 944 68796 950
rect 68744 886 68796 892
rect 68836 944 68888 950
rect 68836 886 68888 892
rect 68928 808 68980 814
rect 68100 740 68152 746
rect 68100 682 68152 688
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69032 800 69060 3538
rect 69124 3398 69152 5578
rect 69112 3392 69164 3398
rect 69112 3334 69164 3340
rect 69308 2106 69336 6695
rect 70136 6662 70164 6938
rect 69940 6656 69992 6662
rect 69940 6598 69992 6604
rect 70124 6656 70176 6662
rect 70124 6598 70176 6604
rect 69952 6322 69980 6598
rect 70950 6352 71006 6361
rect 69940 6316 69992 6322
rect 70950 6287 71006 6296
rect 69940 6258 69992 6264
rect 69952 5914 69980 6258
rect 70964 6254 70992 6287
rect 70952 6248 71004 6254
rect 70952 6190 71004 6196
rect 69940 5908 69992 5914
rect 69940 5850 69992 5856
rect 71044 5568 71096 5574
rect 71044 5510 71096 5516
rect 70492 5160 70544 5166
rect 70492 5102 70544 5108
rect 70030 4584 70086 4593
rect 70030 4519 70086 4528
rect 70044 4146 70072 4519
rect 70032 4140 70084 4146
rect 70032 4082 70084 4088
rect 70216 4140 70268 4146
rect 70216 4082 70268 4088
rect 70124 3936 70176 3942
rect 69386 3904 69442 3913
rect 69386 3839 69442 3848
rect 70122 3904 70124 3913
rect 70176 3904 70178 3913
rect 70122 3839 70178 3848
rect 69296 2100 69348 2106
rect 69296 2042 69348 2048
rect 69204 1896 69256 1902
rect 69204 1838 69256 1844
rect 69216 882 69244 1838
rect 69204 876 69256 882
rect 69204 818 69256 824
rect 69400 800 69428 3839
rect 69570 3224 69626 3233
rect 69570 3159 69626 3168
rect 70122 3224 70178 3233
rect 70122 3159 70124 3168
rect 69584 2854 69612 3159
rect 70176 3159 70178 3168
rect 70124 3130 70176 3136
rect 70228 3058 70256 4082
rect 70400 4072 70452 4078
rect 70400 4014 70452 4020
rect 70308 3936 70360 3942
rect 70308 3878 70360 3884
rect 70216 3052 70268 3058
rect 70216 2994 70268 3000
rect 69572 2848 69624 2854
rect 69572 2790 69624 2796
rect 70228 2650 70256 2994
rect 70216 2644 70268 2650
rect 70216 2586 70268 2592
rect 69756 2508 69808 2514
rect 69756 2450 69808 2456
rect 69768 800 69796 2450
rect 70320 1970 70348 3878
rect 70412 3398 70440 4014
rect 70400 3392 70452 3398
rect 70400 3334 70452 3340
rect 70398 3224 70454 3233
rect 70398 3159 70400 3168
rect 70452 3159 70454 3168
rect 70400 3130 70452 3136
rect 70504 2922 70532 5102
rect 70676 5024 70728 5030
rect 70676 4966 70728 4972
rect 70584 4140 70636 4146
rect 70584 4082 70636 4088
rect 70596 3942 70624 4082
rect 70584 3936 70636 3942
rect 70584 3878 70636 3884
rect 70582 3768 70638 3777
rect 70582 3703 70638 3712
rect 70596 3670 70624 3703
rect 70584 3664 70636 3670
rect 70584 3606 70636 3612
rect 70582 3224 70638 3233
rect 70582 3159 70638 3168
rect 70596 3058 70624 3159
rect 70584 3052 70636 3058
rect 70584 2994 70636 3000
rect 70492 2916 70544 2922
rect 70492 2858 70544 2864
rect 70596 2650 70624 2994
rect 70584 2644 70636 2650
rect 70584 2586 70636 2592
rect 70400 2304 70452 2310
rect 70400 2246 70452 2252
rect 70308 1964 70360 1970
rect 70308 1906 70360 1912
rect 70032 1760 70084 1766
rect 70032 1702 70084 1708
rect 69848 1556 69900 1562
rect 69848 1498 69900 1504
rect 69860 814 69888 1498
rect 70044 1329 70072 1702
rect 70320 1562 70348 1906
rect 70412 1562 70440 2246
rect 70490 1728 70546 1737
rect 70490 1663 70546 1672
rect 70308 1556 70360 1562
rect 70308 1498 70360 1504
rect 70400 1556 70452 1562
rect 70400 1498 70452 1504
rect 70030 1320 70086 1329
rect 70030 1255 70086 1264
rect 70214 1184 70270 1193
rect 70214 1119 70270 1128
rect 70124 944 70176 950
rect 70124 886 70176 892
rect 69848 808 69900 814
rect 68928 750 68980 756
rect 68940 474 68968 750
rect 68928 468 68980 474
rect 68928 410 68980 416
rect 69018 0 69074 800
rect 69112 740 69164 746
rect 69112 682 69164 688
rect 69124 474 69152 682
rect 69112 468 69164 474
rect 69112 410 69164 416
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70136 800 70164 886
rect 69848 750 69900 756
rect 70122 0 70178 800
rect 70228 746 70256 1119
rect 70504 800 70532 1663
rect 70688 950 70716 4966
rect 71056 4146 71084 5510
rect 70952 4140 71004 4146
rect 70952 4082 71004 4088
rect 71044 4140 71096 4146
rect 71044 4082 71096 4088
rect 70964 3466 70992 4082
rect 71148 3534 71176 7754
rect 71688 7540 71740 7546
rect 71688 7482 71740 7488
rect 71228 4072 71280 4078
rect 71228 4014 71280 4020
rect 71320 4072 71372 4078
rect 71320 4014 71372 4020
rect 71136 3528 71188 3534
rect 71136 3470 71188 3476
rect 70952 3460 71004 3466
rect 70952 3402 71004 3408
rect 71136 3052 71188 3058
rect 71136 2994 71188 3000
rect 70952 2916 71004 2922
rect 70952 2858 71004 2864
rect 70964 1970 70992 2858
rect 71148 2650 71176 2994
rect 71136 2644 71188 2650
rect 71136 2586 71188 2592
rect 71042 2408 71098 2417
rect 71042 2343 71098 2352
rect 71056 2106 71084 2343
rect 71044 2100 71096 2106
rect 71044 2042 71096 2048
rect 70952 1964 71004 1970
rect 70952 1906 71004 1912
rect 70964 1358 70992 1906
rect 70952 1352 71004 1358
rect 70952 1294 71004 1300
rect 70676 944 70728 950
rect 70676 886 70728 892
rect 70860 944 70912 950
rect 70860 886 70912 892
rect 70872 800 70900 886
rect 71240 800 71268 4014
rect 71332 2990 71360 4014
rect 71596 3460 71648 3466
rect 71596 3402 71648 3408
rect 71320 2984 71372 2990
rect 71320 2926 71372 2932
rect 71318 2408 71374 2417
rect 71318 2343 71320 2352
rect 71372 2343 71374 2352
rect 71320 2314 71372 2320
rect 71504 1760 71556 1766
rect 71504 1702 71556 1708
rect 71516 1358 71544 1702
rect 71504 1352 71556 1358
rect 71504 1294 71556 1300
rect 71608 800 71636 3402
rect 71700 3058 71728 7482
rect 71870 7304 71926 7313
rect 71870 7239 71926 7248
rect 71780 6316 71832 6322
rect 71780 6258 71832 6264
rect 71792 5574 71820 6258
rect 71780 5568 71832 5574
rect 71780 5510 71832 5516
rect 71792 3670 71820 5510
rect 71780 3664 71832 3670
rect 71780 3606 71832 3612
rect 71780 3188 71832 3194
rect 71780 3130 71832 3136
rect 71688 3052 71740 3058
rect 71688 2994 71740 3000
rect 71688 2644 71740 2650
rect 71688 2586 71740 2592
rect 71700 1737 71728 2586
rect 71686 1728 71742 1737
rect 71686 1663 71742 1672
rect 71792 1442 71820 3130
rect 71884 2650 71912 7239
rect 72056 6724 72108 6730
rect 72056 6666 72108 6672
rect 72068 4146 72096 6666
rect 71964 4140 72016 4146
rect 71964 4082 72016 4088
rect 72056 4140 72108 4146
rect 72056 4082 72108 4088
rect 71976 3670 72004 4082
rect 72896 3670 72924 7822
rect 73540 7721 73568 11154
rect 73620 10668 73672 10674
rect 73620 10610 73672 10616
rect 73632 9926 73660 10610
rect 73896 10532 73948 10538
rect 73896 10474 73948 10480
rect 73908 10062 73936 10474
rect 73896 10056 73948 10062
rect 73896 9998 73948 10004
rect 73620 9920 73672 9926
rect 73620 9862 73672 9868
rect 73632 9042 73660 9862
rect 74000 9654 74028 12200
rect 74368 11898 74396 12200
rect 74356 11892 74408 11898
rect 74356 11834 74408 11840
rect 74448 11892 74500 11898
rect 74448 11834 74500 11840
rect 74460 11354 74488 11834
rect 74632 11552 74684 11558
rect 74632 11494 74684 11500
rect 74448 11348 74500 11354
rect 74448 11290 74500 11296
rect 74538 11248 74594 11257
rect 74538 11183 74594 11192
rect 74552 10810 74580 11183
rect 74356 10804 74408 10810
rect 74356 10746 74408 10752
rect 74540 10804 74592 10810
rect 74540 10746 74592 10752
rect 74080 10464 74132 10470
rect 74080 10406 74132 10412
rect 74092 10062 74120 10406
rect 74368 10062 74396 10746
rect 74448 10668 74500 10674
rect 74448 10610 74500 10616
rect 74460 10266 74488 10610
rect 74448 10260 74500 10266
rect 74448 10202 74500 10208
rect 74080 10056 74132 10062
rect 74080 9998 74132 10004
rect 74356 10056 74408 10062
rect 74356 9998 74408 10004
rect 73988 9648 74040 9654
rect 73988 9590 74040 9596
rect 73620 9036 73672 9042
rect 73620 8978 73672 8984
rect 74092 8634 74120 9998
rect 74448 9648 74500 9654
rect 74448 9590 74500 9596
rect 74356 9580 74408 9586
rect 74356 9522 74408 9528
rect 74368 9178 74396 9522
rect 74460 9178 74488 9590
rect 74540 9512 74592 9518
rect 74540 9454 74592 9460
rect 74552 9217 74580 9454
rect 74538 9208 74594 9217
rect 74356 9172 74408 9178
rect 74356 9114 74408 9120
rect 74448 9172 74500 9178
rect 74538 9143 74594 9152
rect 74448 9114 74500 9120
rect 74368 8634 74396 9114
rect 74080 8628 74132 8634
rect 74080 8570 74132 8576
rect 74356 8628 74408 8634
rect 74356 8570 74408 8576
rect 74644 8401 74672 11494
rect 74736 11150 74764 12200
rect 74816 11756 74868 11762
rect 74816 11698 74868 11704
rect 74724 11144 74776 11150
rect 74724 11086 74776 11092
rect 74828 11082 74856 11698
rect 75012 11354 75040 12310
rect 75090 12200 75146 13000
rect 75458 12200 75514 13000
rect 75826 12200 75882 13000
rect 76194 12200 76250 13000
rect 76562 12200 76618 13000
rect 76930 12200 76986 13000
rect 77298 12200 77354 13000
rect 77666 12200 77722 13000
rect 78034 12200 78090 13000
rect 78402 12200 78458 13000
rect 78770 12200 78826 13000
rect 79048 12232 79100 12238
rect 75000 11348 75052 11354
rect 75000 11290 75052 11296
rect 74816 11076 74868 11082
rect 74816 11018 74868 11024
rect 74828 9042 74856 11018
rect 75104 10674 75132 12200
rect 75472 11762 75500 12200
rect 75840 11830 75868 12200
rect 75828 11824 75880 11830
rect 75828 11766 75880 11772
rect 75460 11756 75512 11762
rect 75460 11698 75512 11704
rect 75368 11688 75420 11694
rect 75368 11630 75420 11636
rect 75380 11354 75408 11630
rect 75368 11348 75420 11354
rect 75368 11290 75420 11296
rect 76208 11218 76236 12200
rect 76288 11552 76340 11558
rect 76288 11494 76340 11500
rect 76196 11212 76248 11218
rect 76196 11154 76248 11160
rect 76012 11144 76064 11150
rect 76300 11121 76328 11494
rect 76012 11086 76064 11092
rect 76286 11112 76342 11121
rect 75092 10668 75144 10674
rect 75092 10610 75144 10616
rect 75104 10266 75132 10610
rect 75092 10260 75144 10266
rect 75092 10202 75144 10208
rect 76024 9042 76052 11086
rect 76286 11047 76342 11056
rect 76378 10704 76434 10713
rect 76378 10639 76434 10648
rect 76288 10600 76340 10606
rect 76288 10542 76340 10548
rect 76300 9926 76328 10542
rect 76392 10266 76420 10639
rect 76576 10266 76604 12200
rect 76840 12096 76892 12102
rect 76840 12038 76892 12044
rect 76748 11552 76800 11558
rect 76748 11494 76800 11500
rect 76760 11150 76788 11494
rect 76852 11150 76880 12038
rect 76748 11144 76800 11150
rect 76748 11086 76800 11092
rect 76840 11144 76892 11150
rect 76840 11086 76892 11092
rect 76380 10260 76432 10266
rect 76380 10202 76432 10208
rect 76564 10260 76616 10266
rect 76564 10202 76616 10208
rect 76576 10062 76604 10202
rect 76564 10056 76616 10062
rect 76564 9998 76616 10004
rect 76288 9920 76340 9926
rect 76288 9862 76340 9868
rect 76300 9042 76328 9862
rect 76944 9586 76972 12200
rect 77312 10062 77340 12200
rect 77680 11880 77708 12200
rect 77944 12096 77996 12102
rect 77944 12038 77996 12044
rect 77680 11852 77800 11880
rect 77668 11756 77720 11762
rect 77668 11698 77720 11704
rect 77576 11688 77628 11694
rect 77574 11656 77576 11665
rect 77628 11656 77630 11665
rect 77574 11591 77630 11600
rect 77680 11354 77708 11698
rect 77668 11348 77720 11354
rect 77668 11290 77720 11296
rect 77390 10840 77446 10849
rect 77390 10775 77446 10784
rect 77404 10606 77432 10775
rect 77772 10674 77800 11852
rect 77956 11354 77984 12038
rect 77944 11348 77996 11354
rect 77944 11290 77996 11296
rect 78048 10810 78076 12200
rect 78312 11008 78364 11014
rect 78312 10950 78364 10956
rect 78036 10804 78088 10810
rect 78036 10746 78088 10752
rect 77760 10668 77812 10674
rect 77760 10610 77812 10616
rect 77392 10600 77444 10606
rect 77392 10542 77444 10548
rect 78048 10062 78076 10746
rect 78220 10532 78272 10538
rect 78220 10474 78272 10480
rect 78232 10266 78260 10474
rect 78324 10266 78352 10950
rect 78220 10260 78272 10266
rect 78220 10202 78272 10208
rect 78312 10260 78364 10266
rect 78312 10202 78364 10208
rect 78416 10062 78444 12200
rect 78784 11762 78812 12200
rect 79138 12200 79194 13000
rect 79506 12200 79562 13000
rect 79874 12200 79930 13000
rect 80242 12200 80298 13000
rect 80610 12200 80666 13000
rect 80978 12200 81034 13000
rect 81346 12200 81402 13000
rect 81714 12200 81770 13000
rect 82082 12200 82138 13000
rect 82450 12200 82506 13000
rect 82818 12200 82874 13000
rect 83004 12436 83056 12442
rect 83004 12378 83056 12384
rect 79048 12174 79100 12180
rect 79060 11898 79088 12174
rect 79048 11892 79100 11898
rect 79048 11834 79100 11840
rect 78772 11756 78824 11762
rect 78772 11698 78824 11704
rect 78784 11354 78812 11698
rect 78772 11348 78824 11354
rect 78772 11290 78824 11296
rect 79152 11286 79180 12200
rect 79140 11280 79192 11286
rect 79140 11222 79192 11228
rect 79048 10668 79100 10674
rect 79048 10610 79100 10616
rect 79060 10266 79088 10610
rect 79048 10260 79100 10266
rect 79048 10202 79100 10208
rect 79416 10192 79468 10198
rect 79414 10160 79416 10169
rect 79468 10160 79470 10169
rect 79414 10095 79470 10104
rect 79520 10062 79548 12200
rect 79888 11801 79916 12200
rect 80256 12102 80284 12200
rect 80428 12164 80480 12170
rect 80428 12106 80480 12112
rect 80244 12096 80296 12102
rect 80244 12038 80296 12044
rect 79874 11792 79930 11801
rect 79874 11727 79930 11736
rect 80060 11688 80112 11694
rect 80060 11630 80112 11636
rect 80152 11688 80204 11694
rect 80152 11630 80204 11636
rect 80072 11150 80100 11630
rect 80164 11558 80192 11630
rect 80152 11552 80204 11558
rect 80152 11494 80204 11500
rect 80060 11144 80112 11150
rect 80060 11086 80112 11092
rect 77300 10056 77352 10062
rect 78036 10056 78088 10062
rect 77300 9998 77352 10004
rect 77390 10024 77446 10033
rect 78036 9998 78088 10004
rect 78404 10056 78456 10062
rect 78404 9998 78456 10004
rect 79508 10056 79560 10062
rect 79508 9998 79560 10004
rect 77390 9959 77392 9968
rect 77444 9959 77446 9968
rect 77392 9930 77444 9936
rect 78496 9920 78548 9926
rect 78496 9862 78548 9868
rect 78508 9722 78536 9862
rect 78496 9716 78548 9722
rect 78496 9658 78548 9664
rect 76932 9580 76984 9586
rect 76932 9522 76984 9528
rect 76472 9376 76524 9382
rect 76470 9344 76472 9353
rect 76564 9376 76616 9382
rect 76524 9344 76526 9353
rect 76564 9318 76616 9324
rect 76470 9279 76526 9288
rect 74816 9036 74868 9042
rect 74816 8978 74868 8984
rect 76012 9036 76064 9042
rect 76012 8978 76064 8984
rect 76288 9036 76340 9042
rect 76288 8978 76340 8984
rect 76576 8566 76604 9318
rect 76944 9178 76972 9522
rect 76932 9172 76984 9178
rect 76932 9114 76984 9120
rect 80072 9042 80100 11086
rect 80060 9036 80112 9042
rect 80060 8978 80112 8984
rect 80164 8634 80192 11494
rect 80440 11218 80468 12106
rect 80428 11212 80480 11218
rect 80428 11154 80480 11160
rect 80428 10736 80480 10742
rect 80428 10678 80480 10684
rect 80244 10600 80296 10606
rect 80244 10542 80296 10548
rect 80256 10266 80284 10542
rect 80440 10266 80468 10678
rect 80244 10260 80296 10266
rect 80244 10202 80296 10208
rect 80428 10260 80480 10266
rect 80428 10202 80480 10208
rect 80256 9654 80284 10202
rect 80244 9648 80296 9654
rect 80244 9590 80296 9596
rect 80624 9586 80652 12200
rect 80992 11914 81020 12200
rect 80992 11886 81112 11914
rect 80980 11756 81032 11762
rect 80980 11698 81032 11704
rect 80992 11354 81020 11698
rect 80980 11348 81032 11354
rect 80980 11290 81032 11296
rect 81084 10062 81112 11886
rect 81360 10690 81388 12200
rect 81728 11778 81756 12200
rect 82096 11812 82124 12200
rect 82176 11824 82228 11830
rect 82096 11784 82176 11812
rect 81728 11750 82032 11778
rect 82176 11766 82228 11772
rect 81716 11688 81768 11694
rect 81716 11630 81768 11636
rect 81728 11218 81756 11630
rect 82004 11218 82032 11750
rect 82464 11286 82492 12200
rect 82542 11792 82598 11801
rect 82542 11727 82544 11736
rect 82596 11727 82598 11736
rect 82544 11698 82596 11704
rect 82452 11280 82504 11286
rect 82452 11222 82504 11228
rect 81716 11212 81768 11218
rect 81716 11154 81768 11160
rect 81992 11212 82044 11218
rect 81992 11154 82044 11160
rect 81360 10662 81480 10690
rect 81452 10606 81480 10662
rect 81532 10668 81584 10674
rect 81532 10610 81584 10616
rect 81164 10600 81216 10606
rect 81162 10568 81164 10577
rect 81440 10600 81492 10606
rect 81216 10568 81218 10577
rect 81440 10542 81492 10548
rect 81162 10503 81218 10512
rect 81544 10266 81572 10610
rect 82728 10600 82780 10606
rect 82728 10542 82780 10548
rect 82740 10266 82768 10542
rect 81532 10260 81584 10266
rect 81532 10202 81584 10208
rect 82728 10260 82780 10266
rect 82728 10202 82780 10208
rect 81072 10056 81124 10062
rect 81072 9998 81124 10004
rect 82832 9654 82860 12200
rect 82912 12096 82964 12102
rect 82912 12038 82964 12044
rect 82924 11150 82952 12038
rect 83016 11354 83044 12378
rect 83096 12300 83148 12306
rect 83096 12242 83148 12248
rect 83004 11348 83056 11354
rect 83004 11290 83056 11296
rect 82912 11144 82964 11150
rect 82912 11086 82964 11092
rect 82912 10804 82964 10810
rect 82912 10746 82964 10752
rect 82924 10062 82952 10746
rect 82912 10056 82964 10062
rect 82912 9998 82964 10004
rect 82820 9648 82872 9654
rect 82820 9590 82872 9596
rect 80612 9580 80664 9586
rect 80612 9522 80664 9528
rect 80624 9178 80652 9522
rect 80796 9512 80848 9518
rect 80794 9480 80796 9489
rect 80848 9480 80850 9489
rect 83108 9450 83136 12242
rect 83186 12200 83242 13000
rect 83280 12708 83332 12714
rect 83280 12650 83332 12656
rect 83200 10674 83228 12200
rect 83292 11898 83320 12650
rect 83554 12200 83610 13000
rect 83922 12200 83978 13000
rect 84290 12200 84346 13000
rect 84658 12200 84714 13000
rect 85026 12200 85082 13000
rect 85394 12200 85450 13000
rect 85762 12200 85818 13000
rect 86130 12200 86186 13000
rect 86498 12200 86554 13000
rect 86866 12200 86922 13000
rect 87234 12200 87290 13000
rect 87602 12200 87658 13000
rect 87970 12200 88026 13000
rect 88338 12200 88394 13000
rect 88706 12200 88762 13000
rect 89074 12200 89130 13000
rect 89442 12200 89498 13000
rect 89810 12200 89866 13000
rect 90178 12200 90234 13000
rect 90546 12200 90602 13000
rect 90914 12200 90970 13000
rect 91282 12200 91338 13000
rect 91650 12200 91706 13000
rect 92018 12200 92074 13000
rect 92386 12200 92442 13000
rect 92754 12200 92810 13000
rect 93122 12200 93178 13000
rect 93490 12200 93546 13000
rect 93858 12200 93914 13000
rect 94226 12200 94282 13000
rect 94594 12200 94650 13000
rect 94962 12200 95018 13000
rect 95330 12200 95386 13000
rect 95698 12200 95754 13000
rect 96066 12200 96122 13000
rect 96434 12200 96490 13000
rect 96802 12200 96858 13000
rect 96896 12504 96948 12510
rect 96896 12446 96948 12452
rect 83280 11892 83332 11898
rect 83280 11834 83332 11840
rect 83372 11756 83424 11762
rect 83372 11698 83424 11704
rect 83384 11354 83412 11698
rect 83372 11348 83424 11354
rect 83372 11290 83424 11296
rect 83568 10826 83596 12200
rect 83476 10798 83596 10826
rect 83936 10810 83964 12200
rect 83924 10804 83976 10810
rect 83188 10668 83240 10674
rect 83188 10610 83240 10616
rect 83188 9580 83240 9586
rect 83188 9522 83240 9528
rect 80794 9415 80850 9424
rect 83096 9444 83148 9450
rect 83096 9386 83148 9392
rect 83200 9178 83228 9522
rect 83476 9518 83504 10798
rect 83924 10746 83976 10752
rect 83556 10668 83608 10674
rect 83556 10610 83608 10616
rect 83568 10266 83596 10610
rect 83556 10260 83608 10266
rect 83556 10202 83608 10208
rect 83464 9512 83516 9518
rect 83464 9454 83516 9460
rect 80612 9172 80664 9178
rect 80612 9114 80664 9120
rect 83188 9172 83240 9178
rect 83188 9114 83240 9120
rect 83476 9110 83504 9454
rect 83464 9104 83516 9110
rect 83464 9046 83516 9052
rect 84304 9042 84332 12200
rect 84672 10690 84700 12200
rect 84752 11756 84804 11762
rect 84752 11698 84804 11704
rect 84764 11354 84792 11698
rect 85040 11642 85068 12200
rect 85040 11614 85252 11642
rect 84852 11452 85148 11472
rect 84908 11450 84932 11452
rect 84988 11450 85012 11452
rect 85068 11450 85092 11452
rect 84930 11398 84932 11450
rect 84994 11398 85006 11450
rect 85068 11398 85070 11450
rect 84908 11396 84932 11398
rect 84988 11396 85012 11398
rect 85068 11396 85092 11398
rect 84852 11376 85148 11396
rect 84752 11348 84804 11354
rect 84752 11290 84804 11296
rect 84580 10662 84700 10690
rect 84580 9586 84608 10662
rect 84660 10600 84712 10606
rect 84660 10542 84712 10548
rect 84672 10266 84700 10542
rect 84852 10364 85148 10384
rect 84908 10362 84932 10364
rect 84988 10362 85012 10364
rect 85068 10362 85092 10364
rect 84930 10310 84932 10362
rect 84994 10310 85006 10362
rect 85068 10310 85070 10362
rect 84908 10308 84932 10310
rect 84988 10308 85012 10310
rect 85068 10308 85092 10310
rect 84852 10288 85148 10308
rect 84660 10260 84712 10266
rect 84660 10202 84712 10208
rect 85224 10198 85252 11614
rect 85212 10192 85264 10198
rect 85212 10134 85264 10140
rect 85120 10124 85172 10130
rect 85120 10066 85172 10072
rect 85132 9722 85160 10066
rect 85120 9716 85172 9722
rect 85120 9658 85172 9664
rect 84568 9580 84620 9586
rect 84568 9522 84620 9528
rect 84852 9276 85148 9296
rect 84908 9274 84932 9276
rect 84988 9274 85012 9276
rect 85068 9274 85092 9276
rect 84930 9222 84932 9274
rect 84994 9222 85006 9274
rect 85068 9222 85070 9274
rect 84908 9220 84932 9222
rect 84988 9220 85012 9222
rect 85068 9220 85092 9222
rect 84852 9200 85148 9220
rect 85408 9178 85436 12200
rect 85776 11234 85804 12200
rect 85776 11206 85896 11234
rect 85764 11076 85816 11082
rect 85764 11018 85816 11024
rect 85776 10674 85804 11018
rect 85764 10668 85816 10674
rect 85764 10610 85816 10616
rect 85672 10600 85724 10606
rect 85670 10568 85672 10577
rect 85724 10568 85726 10577
rect 85670 10503 85726 10512
rect 85396 9172 85448 9178
rect 85396 9114 85448 9120
rect 84292 9036 84344 9042
rect 84292 8978 84344 8984
rect 81990 8936 82046 8945
rect 81990 8871 81992 8880
rect 82044 8871 82046 8880
rect 81992 8842 82044 8848
rect 85578 8800 85634 8809
rect 85634 8758 85712 8786
rect 85578 8735 85634 8744
rect 80152 8628 80204 8634
rect 80152 8570 80204 8576
rect 76564 8560 76616 8566
rect 85684 8537 85712 8758
rect 85868 8634 85896 11206
rect 85948 11008 86000 11014
rect 85948 10950 86000 10956
rect 85960 10130 85988 10950
rect 85948 10124 86000 10130
rect 85948 10066 86000 10072
rect 86144 8838 86172 12200
rect 86512 9518 86540 12200
rect 86500 9512 86552 9518
rect 86500 9454 86552 9460
rect 86132 8832 86184 8838
rect 86132 8774 86184 8780
rect 85856 8628 85908 8634
rect 85856 8570 85908 8576
rect 76564 8502 76616 8508
rect 85670 8528 85726 8537
rect 83464 8492 83516 8498
rect 85670 8463 85726 8472
rect 83464 8434 83516 8440
rect 81992 8424 82044 8430
rect 74630 8392 74686 8401
rect 81992 8366 82044 8372
rect 83004 8424 83056 8430
rect 83004 8366 83056 8372
rect 74630 8327 74686 8336
rect 79416 8288 79468 8294
rect 79416 8230 79468 8236
rect 79428 7954 79456 8230
rect 82004 7954 82032 8366
rect 79416 7948 79468 7954
rect 79416 7890 79468 7896
rect 80428 7948 80480 7954
rect 80428 7890 80480 7896
rect 81992 7948 82044 7954
rect 81992 7890 82044 7896
rect 80152 7744 80204 7750
rect 73526 7712 73582 7721
rect 80152 7686 80204 7692
rect 73526 7647 73582 7656
rect 79784 7336 79836 7342
rect 79784 7278 79836 7284
rect 79796 6866 79824 7278
rect 73252 6860 73304 6866
rect 73252 6802 73304 6808
rect 79784 6860 79836 6866
rect 79784 6802 79836 6808
rect 73066 3904 73122 3913
rect 73066 3839 73122 3848
rect 71964 3664 72016 3670
rect 71964 3606 72016 3612
rect 72700 3664 72752 3670
rect 72700 3606 72752 3612
rect 72884 3664 72936 3670
rect 72884 3606 72936 3612
rect 72976 3664 73028 3670
rect 72976 3606 73028 3612
rect 72148 3596 72200 3602
rect 72148 3538 72200 3544
rect 72056 3460 72108 3466
rect 72056 3402 72108 3408
rect 72068 3126 72096 3402
rect 72056 3120 72108 3126
rect 72056 3062 72108 3068
rect 72054 2952 72110 2961
rect 72054 2887 72110 2896
rect 71872 2644 71924 2650
rect 71872 2586 71924 2592
rect 71792 1414 72004 1442
rect 71780 1352 71832 1358
rect 71780 1294 71832 1300
rect 71792 882 71820 1294
rect 71872 1216 71924 1222
rect 71872 1158 71924 1164
rect 71884 950 71912 1158
rect 71872 944 71924 950
rect 71872 886 71924 892
rect 71780 876 71832 882
rect 71780 818 71832 824
rect 71976 800 72004 1414
rect 72068 1358 72096 2887
rect 72160 2650 72188 3538
rect 72332 3528 72384 3534
rect 72332 3470 72384 3476
rect 72712 3482 72740 3606
rect 72148 2644 72200 2650
rect 72148 2586 72200 2592
rect 72056 1352 72108 1358
rect 72056 1294 72108 1300
rect 72344 800 72372 3470
rect 72424 3460 72476 3466
rect 72712 3454 72832 3482
rect 72424 3402 72476 3408
rect 72436 2854 72464 3402
rect 72424 2848 72476 2854
rect 72424 2790 72476 2796
rect 72516 1964 72568 1970
rect 72516 1906 72568 1912
rect 72424 1896 72476 1902
rect 72424 1838 72476 1844
rect 72436 1329 72464 1838
rect 72528 1358 72556 1906
rect 72608 1556 72660 1562
rect 72608 1498 72660 1504
rect 72516 1352 72568 1358
rect 72422 1320 72478 1329
rect 72516 1294 72568 1300
rect 72422 1255 72478 1264
rect 72620 1222 72648 1498
rect 72804 1442 72832 3454
rect 72988 3233 73016 3606
rect 73080 3602 73108 3839
rect 73068 3596 73120 3602
rect 73068 3538 73120 3544
rect 72974 3224 73030 3233
rect 72974 3159 73030 3168
rect 72884 2508 72936 2514
rect 72884 2450 72936 2456
rect 72896 2038 72924 2450
rect 73264 2106 73292 6802
rect 74724 6792 74776 6798
rect 74724 6734 74776 6740
rect 74354 4176 74410 4185
rect 74354 4111 74410 4120
rect 73802 3768 73858 3777
rect 73802 3703 73858 3712
rect 73344 3528 73396 3534
rect 73344 3470 73396 3476
rect 73356 3398 73384 3470
rect 73816 3398 73844 3703
rect 73344 3392 73396 3398
rect 73712 3392 73764 3398
rect 73344 3334 73396 3340
rect 73526 3360 73582 3369
rect 73712 3334 73764 3340
rect 73804 3392 73856 3398
rect 73804 3334 73856 3340
rect 73526 3295 73582 3304
rect 73540 3194 73568 3295
rect 73528 3188 73580 3194
rect 73528 3130 73580 3136
rect 73620 2984 73672 2990
rect 73620 2926 73672 2932
rect 73436 2304 73488 2310
rect 73436 2246 73488 2252
rect 73252 2100 73304 2106
rect 73252 2042 73304 2048
rect 72884 2032 72936 2038
rect 72884 1974 72936 1980
rect 72976 2032 73028 2038
rect 72976 1974 73028 1980
rect 72712 1414 72832 1442
rect 72988 1426 73016 1974
rect 72976 1420 73028 1426
rect 72608 1216 72660 1222
rect 72608 1158 72660 1164
rect 72712 800 72740 1414
rect 72976 1362 73028 1368
rect 73068 1216 73120 1222
rect 73068 1158 73120 1164
rect 72976 876 73028 882
rect 72976 818 73028 824
rect 70216 740 70268 746
rect 70216 682 70268 688
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 72988 474 73016 818
rect 73080 800 73108 1158
rect 73448 800 73476 2246
rect 73632 1766 73660 2926
rect 73724 2106 73752 3334
rect 74264 3052 74316 3058
rect 74264 2994 74316 3000
rect 74276 2854 74304 2994
rect 73804 2848 73856 2854
rect 73804 2790 73856 2796
rect 74264 2848 74316 2854
rect 74264 2790 74316 2796
rect 73712 2100 73764 2106
rect 73712 2042 73764 2048
rect 73620 1760 73672 1766
rect 73620 1702 73672 1708
rect 73816 800 73844 2790
rect 74276 2650 74304 2790
rect 74264 2644 74316 2650
rect 74264 2586 74316 2592
rect 73896 2032 73948 2038
rect 73896 1974 73948 1980
rect 73908 1290 73936 1974
rect 74172 1760 74224 1766
rect 74172 1702 74224 1708
rect 74264 1760 74316 1766
rect 74264 1702 74316 1708
rect 73896 1284 73948 1290
rect 73896 1226 73948 1232
rect 74184 800 74212 1702
rect 74276 814 74304 1702
rect 74368 1426 74396 4111
rect 74540 4004 74592 4010
rect 74540 3946 74592 3952
rect 74356 1420 74408 1426
rect 74356 1362 74408 1368
rect 74264 808 74316 814
rect 72976 468 73028 474
rect 72976 410 73028 416
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73802 0 73858 800
rect 74170 0 74226 800
rect 74552 800 74580 3946
rect 74736 2650 74764 6734
rect 79140 6656 79192 6662
rect 79140 6598 79192 6604
rect 75736 6180 75788 6186
rect 75736 6122 75788 6128
rect 75748 6066 75776 6122
rect 75828 6112 75880 6118
rect 75748 6060 75828 6066
rect 75748 6054 75880 6060
rect 75748 6038 75868 6054
rect 76012 4140 76064 4146
rect 76012 4082 76064 4088
rect 76380 4140 76432 4146
rect 76380 4082 76432 4088
rect 74908 2916 74960 2922
rect 74908 2858 74960 2864
rect 74724 2644 74776 2650
rect 74724 2586 74776 2592
rect 74632 2304 74684 2310
rect 74632 2246 74684 2252
rect 74644 1970 74672 2246
rect 74632 1964 74684 1970
rect 74632 1906 74684 1912
rect 74920 800 74948 2858
rect 75918 2680 75974 2689
rect 75918 2615 75974 2624
rect 75736 2372 75788 2378
rect 75736 2314 75788 2320
rect 75000 2304 75052 2310
rect 75000 2246 75052 2252
rect 75012 1562 75040 2246
rect 75644 1964 75696 1970
rect 75644 1906 75696 1912
rect 75092 1896 75144 1902
rect 75092 1838 75144 1844
rect 75104 1562 75132 1838
rect 75274 1728 75330 1737
rect 75274 1663 75330 1672
rect 75000 1556 75052 1562
rect 75000 1498 75052 1504
rect 75092 1556 75144 1562
rect 75092 1498 75144 1504
rect 74998 1048 75054 1057
rect 74998 983 75054 992
rect 74264 750 74316 756
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75012 785 75040 983
rect 75104 950 75132 1498
rect 75184 1216 75236 1222
rect 75184 1158 75236 1164
rect 75196 950 75224 1158
rect 75092 944 75144 950
rect 75092 886 75144 892
rect 75184 944 75236 950
rect 75184 886 75236 892
rect 75288 800 75316 1663
rect 75656 800 75684 1906
rect 74998 776 75054 785
rect 74998 711 75054 720
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 75748 746 75776 2314
rect 75932 1902 75960 2615
rect 75920 1896 75972 1902
rect 75920 1838 75972 1844
rect 75828 808 75880 814
rect 76024 800 76052 4082
rect 76104 2984 76156 2990
rect 76104 2926 76156 2932
rect 76116 1358 76144 2926
rect 76104 1352 76156 1358
rect 76104 1294 76156 1300
rect 76392 800 76420 4082
rect 77852 4072 77904 4078
rect 77852 4014 77904 4020
rect 76564 2984 76616 2990
rect 76564 2926 76616 2932
rect 76576 2446 76604 2926
rect 77300 2848 77352 2854
rect 77300 2790 77352 2796
rect 76564 2440 76616 2446
rect 76564 2382 76616 2388
rect 76656 2440 76708 2446
rect 76656 2382 76708 2388
rect 77114 2408 77170 2417
rect 76668 882 76696 2382
rect 77114 2343 77170 2352
rect 76748 1420 76800 1426
rect 76748 1362 76800 1368
rect 76656 876 76708 882
rect 76656 818 76708 824
rect 76760 800 76788 1362
rect 77128 800 77156 2343
rect 77312 1714 77340 2790
rect 77574 2136 77630 2145
rect 77574 2071 77576 2080
rect 77628 2071 77630 2080
rect 77576 2042 77628 2048
rect 77312 1686 77432 1714
rect 77298 1592 77354 1601
rect 77298 1527 77354 1536
rect 77312 1426 77340 1527
rect 77300 1420 77352 1426
rect 77300 1362 77352 1368
rect 77404 898 77432 1686
rect 77574 1184 77630 1193
rect 77574 1119 77630 1128
rect 77404 870 77524 898
rect 77496 800 77524 870
rect 77588 814 77616 1119
rect 77576 808 77628 814
rect 75828 750 75880 756
rect 75736 740 75788 746
rect 75736 682 75788 688
rect 75840 66 75868 750
rect 75828 60 75880 66
rect 75828 2 75880 8
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77482 0 77538 800
rect 77864 800 77892 4014
rect 78220 3664 78272 3670
rect 78220 3606 78272 3612
rect 78036 2100 78088 2106
rect 78036 2042 78088 2048
rect 78048 1426 78076 2042
rect 78036 1420 78088 1426
rect 78036 1362 78088 1368
rect 78232 800 78260 3606
rect 78956 3528 79008 3534
rect 78956 3470 79008 3476
rect 78588 1964 78640 1970
rect 78588 1906 78640 1912
rect 78600 1222 78628 1906
rect 78588 1216 78640 1222
rect 78588 1158 78640 1164
rect 78600 800 78628 1158
rect 78680 808 78732 814
rect 77576 750 77628 756
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78968 800 78996 3470
rect 79152 2106 79180 6598
rect 79692 2644 79744 2650
rect 79692 2586 79744 2592
rect 79324 2440 79376 2446
rect 79324 2382 79376 2388
rect 79336 2106 79364 2382
rect 79140 2100 79192 2106
rect 79140 2042 79192 2048
rect 79324 2100 79376 2106
rect 79324 2042 79376 2048
rect 79048 1964 79100 1970
rect 79048 1906 79100 1912
rect 79060 1222 79088 1906
rect 79336 1358 79364 2042
rect 79324 1352 79376 1358
rect 79324 1294 79376 1300
rect 79416 1352 79468 1358
rect 79416 1294 79468 1300
rect 79600 1352 79652 1358
rect 79600 1294 79652 1300
rect 79048 1216 79100 1222
rect 79048 1158 79100 1164
rect 79244 882 79364 898
rect 79428 882 79456 1294
rect 79232 876 79364 882
rect 79284 870 79364 876
rect 79232 818 79284 824
rect 79336 800 79364 870
rect 79416 876 79468 882
rect 79416 818 79468 824
rect 78680 750 78732 756
rect 78692 134 78720 750
rect 78680 128 78732 134
rect 78680 70 78732 76
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79612 746 79640 1294
rect 79704 800 79732 2586
rect 80164 1290 80192 7686
rect 80440 7177 80468 7890
rect 80888 7880 80940 7886
rect 80888 7822 80940 7828
rect 80794 7440 80850 7449
rect 80794 7375 80850 7384
rect 80808 7342 80836 7375
rect 80796 7336 80848 7342
rect 80796 7278 80848 7284
rect 80426 7168 80482 7177
rect 80426 7103 80482 7112
rect 80900 2650 80928 7822
rect 81348 7404 81400 7410
rect 81348 7346 81400 7352
rect 81360 6662 81388 7346
rect 81900 7200 81952 7206
rect 81900 7142 81952 7148
rect 81912 6866 81940 7142
rect 81900 6860 81952 6866
rect 81900 6802 81952 6808
rect 81348 6656 81400 6662
rect 81348 6598 81400 6604
rect 81912 6458 81940 6802
rect 82820 6792 82872 6798
rect 82820 6734 82872 6740
rect 81992 6656 82044 6662
rect 81992 6598 82044 6604
rect 81900 6452 81952 6458
rect 81900 6394 81952 6400
rect 81624 4820 81676 4826
rect 81624 4762 81676 4768
rect 80980 2984 81032 2990
rect 80980 2926 81032 2932
rect 80888 2644 80940 2650
rect 80888 2586 80940 2592
rect 80796 2508 80848 2514
rect 80796 2450 80848 2456
rect 80428 2440 80480 2446
rect 80428 2382 80480 2388
rect 80152 1284 80204 1290
rect 80152 1226 80204 1232
rect 79968 1216 80020 1222
rect 80020 1164 80100 1170
rect 79968 1158 80100 1164
rect 79980 1142 80100 1158
rect 80072 800 80100 1142
rect 80440 800 80468 2382
rect 80520 1760 80572 1766
rect 80520 1702 80572 1708
rect 80532 950 80560 1702
rect 80520 944 80572 950
rect 80520 886 80572 892
rect 80808 800 80836 2450
rect 80888 2372 80940 2378
rect 80888 2314 80940 2320
rect 80900 2106 80928 2314
rect 80888 2100 80940 2106
rect 80888 2042 80940 2048
rect 80992 1562 81020 2926
rect 81348 2100 81400 2106
rect 81348 2042 81400 2048
rect 81360 1970 81388 2042
rect 81348 1964 81400 1970
rect 81348 1906 81400 1912
rect 81072 1896 81124 1902
rect 81072 1838 81124 1844
rect 81256 1896 81308 1902
rect 81256 1838 81308 1844
rect 80980 1556 81032 1562
rect 80980 1498 81032 1504
rect 81084 882 81112 1838
rect 81268 1562 81296 1838
rect 81256 1556 81308 1562
rect 81256 1498 81308 1504
rect 81360 1290 81388 1906
rect 81348 1284 81400 1290
rect 81348 1226 81400 1232
rect 81532 1284 81584 1290
rect 81532 1226 81584 1232
rect 81164 1216 81216 1222
rect 81164 1158 81216 1164
rect 81072 876 81124 882
rect 81072 818 81124 824
rect 81176 800 81204 1158
rect 81544 800 81572 1226
rect 79600 740 79652 746
rect 79600 682 79652 688
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81636 474 81664 4762
rect 81900 3460 81952 3466
rect 81900 3402 81952 3408
rect 81912 800 81940 3402
rect 82004 2650 82032 6598
rect 82266 2816 82322 2825
rect 82266 2751 82322 2760
rect 81992 2644 82044 2650
rect 81992 2586 82044 2592
rect 82176 1964 82228 1970
rect 82176 1906 82228 1912
rect 82188 1290 82216 1906
rect 82176 1284 82228 1290
rect 82176 1226 82228 1232
rect 81992 1216 82044 1222
rect 81992 1158 82044 1164
rect 81624 468 81676 474
rect 81624 410 81676 416
rect 81898 0 81954 800
rect 82004 406 82032 1158
rect 82280 800 82308 2751
rect 82832 2106 82860 6734
rect 83016 6633 83044 8366
rect 83372 7948 83424 7954
rect 83372 7890 83424 7896
rect 83384 7546 83412 7890
rect 83476 7750 83504 8434
rect 86880 8362 86908 12200
rect 87144 11756 87196 11762
rect 87144 11698 87196 11704
rect 86960 11688 87012 11694
rect 86960 11630 87012 11636
rect 86972 10810 87000 11630
rect 87156 11354 87184 11698
rect 87144 11348 87196 11354
rect 87144 11290 87196 11296
rect 86960 10804 87012 10810
rect 86960 10746 87012 10752
rect 86960 9920 87012 9926
rect 86960 9862 87012 9868
rect 86972 9722 87000 9862
rect 86960 9716 87012 9722
rect 86960 9658 87012 9664
rect 87156 9654 87184 11290
rect 87248 10130 87276 12200
rect 87512 11076 87564 11082
rect 87512 11018 87564 11024
rect 87236 10124 87288 10130
rect 87236 10066 87288 10072
rect 87236 9920 87288 9926
rect 87236 9862 87288 9868
rect 87144 9648 87196 9654
rect 87144 9590 87196 9596
rect 86960 9580 87012 9586
rect 86960 9522 87012 9528
rect 86972 9178 87000 9522
rect 86960 9172 87012 9178
rect 86960 9114 87012 9120
rect 87248 9042 87276 9862
rect 87524 9586 87552 11018
rect 87512 9580 87564 9586
rect 87512 9522 87564 9528
rect 87236 9036 87288 9042
rect 87236 8978 87288 8984
rect 87616 8498 87644 12200
rect 87604 8492 87656 8498
rect 87604 8434 87656 8440
rect 87984 8430 88012 12200
rect 88352 11642 88380 12200
rect 88352 11614 88472 11642
rect 88340 11552 88392 11558
rect 88340 11494 88392 11500
rect 88352 10674 88380 11494
rect 88340 10668 88392 10674
rect 88340 10610 88392 10616
rect 88064 10600 88116 10606
rect 88064 10542 88116 10548
rect 88076 9897 88104 10542
rect 88062 9888 88118 9897
rect 88062 9823 88118 9832
rect 88340 8628 88392 8634
rect 88340 8570 88392 8576
rect 87236 8424 87288 8430
rect 87236 8366 87288 8372
rect 87972 8424 88024 8430
rect 87972 8366 88024 8372
rect 86868 8356 86920 8362
rect 86868 8298 86920 8304
rect 83832 8288 83884 8294
rect 83832 8230 83884 8236
rect 83844 7954 83872 8230
rect 84852 8188 85148 8208
rect 84908 8186 84932 8188
rect 84988 8186 85012 8188
rect 85068 8186 85092 8188
rect 84930 8134 84932 8186
rect 84994 8134 85006 8186
rect 85068 8134 85070 8186
rect 84908 8132 84932 8134
rect 84988 8132 85012 8134
rect 85068 8132 85092 8134
rect 84852 8112 85148 8132
rect 87248 8090 87276 8366
rect 87512 8288 87564 8294
rect 87512 8230 87564 8236
rect 87236 8084 87288 8090
rect 87236 8026 87288 8032
rect 87524 7954 87552 8230
rect 88352 7954 88380 8570
rect 83832 7948 83884 7954
rect 83832 7890 83884 7896
rect 87512 7948 87564 7954
rect 87512 7890 87564 7896
rect 88340 7948 88392 7954
rect 88340 7890 88392 7896
rect 84752 7880 84804 7886
rect 84752 7822 84804 7828
rect 83464 7744 83516 7750
rect 83464 7686 83516 7692
rect 83372 7540 83424 7546
rect 83372 7482 83424 7488
rect 83186 7032 83242 7041
rect 83186 6967 83242 6976
rect 83200 6934 83228 6967
rect 83188 6928 83240 6934
rect 83188 6870 83240 6876
rect 83002 6624 83058 6633
rect 83002 6559 83058 6568
rect 83004 3936 83056 3942
rect 83004 3878 83056 3884
rect 82820 2100 82872 2106
rect 82820 2042 82872 2048
rect 82636 1216 82688 1222
rect 82636 1158 82688 1164
rect 82648 800 82676 1158
rect 83016 800 83044 3878
rect 83096 2984 83148 2990
rect 83096 2926 83148 2932
rect 83108 2106 83136 2926
rect 83476 2650 83504 7686
rect 84660 4004 84712 4010
rect 84660 3946 84712 3952
rect 83740 3732 83792 3738
rect 83740 3674 83792 3680
rect 83464 2644 83516 2650
rect 83464 2586 83516 2592
rect 83556 2644 83608 2650
rect 83556 2586 83608 2592
rect 83096 2100 83148 2106
rect 83096 2042 83148 2048
rect 83108 1426 83136 2042
rect 83464 1896 83516 1902
rect 83462 1864 83464 1873
rect 83516 1864 83518 1873
rect 83462 1799 83518 1808
rect 83568 1766 83596 2586
rect 83556 1760 83608 1766
rect 83556 1702 83608 1708
rect 83096 1420 83148 1426
rect 83096 1362 83148 1368
rect 83384 882 83504 898
rect 83384 876 83516 882
rect 83384 870 83464 876
rect 83384 800 83412 870
rect 83464 818 83516 824
rect 83752 800 83780 3674
rect 84476 2304 84528 2310
rect 84476 2246 84528 2252
rect 84198 2000 84254 2009
rect 84198 1935 84254 1944
rect 84212 1426 84240 1935
rect 84200 1420 84252 1426
rect 84200 1362 84252 1368
rect 84028 870 84148 898
rect 84028 814 84056 870
rect 84016 808 84068 814
rect 82176 740 82228 746
rect 82176 682 82228 688
rect 81992 400 82044 406
rect 81992 342 82044 348
rect 82188 338 82216 682
rect 82176 332 82228 338
rect 82176 274 82228 280
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83280 672 83332 678
rect 83280 614 83332 620
rect 83292 270 83320 614
rect 83280 264 83332 270
rect 83280 206 83332 212
rect 83370 0 83426 800
rect 83738 0 83794 800
rect 84120 800 84148 870
rect 84488 800 84516 2246
rect 84672 1970 84700 3946
rect 84764 2106 84792 7822
rect 87604 7336 87656 7342
rect 87604 7278 87656 7284
rect 87788 7336 87840 7342
rect 87788 7278 87840 7284
rect 84852 7100 85148 7120
rect 84908 7098 84932 7100
rect 84988 7098 85012 7100
rect 85068 7098 85092 7100
rect 84930 7046 84932 7098
rect 84994 7046 85006 7098
rect 85068 7046 85070 7098
rect 84908 7044 84932 7046
rect 84988 7044 85012 7046
rect 85068 7044 85092 7046
rect 84852 7024 85148 7044
rect 87616 6866 87644 7278
rect 87800 6934 87828 7278
rect 88156 6996 88208 7002
rect 88156 6938 88208 6944
rect 87788 6928 87840 6934
rect 87788 6870 87840 6876
rect 87604 6860 87656 6866
rect 87604 6802 87656 6808
rect 87800 6458 87828 6870
rect 87788 6452 87840 6458
rect 87788 6394 87840 6400
rect 87512 6248 87564 6254
rect 87512 6190 87564 6196
rect 84852 6012 85148 6032
rect 84908 6010 84932 6012
rect 84988 6010 85012 6012
rect 85068 6010 85092 6012
rect 84930 5958 84932 6010
rect 84994 5958 85006 6010
rect 85068 5958 85070 6010
rect 84908 5956 84932 5958
rect 84988 5956 85012 5958
rect 85068 5956 85092 5958
rect 84852 5936 85148 5956
rect 87524 5778 87552 6190
rect 87512 5772 87564 5778
rect 87512 5714 87564 5720
rect 86776 5160 86828 5166
rect 86776 5102 86828 5108
rect 87788 5160 87840 5166
rect 87788 5102 87840 5108
rect 84852 4924 85148 4944
rect 84908 4922 84932 4924
rect 84988 4922 85012 4924
rect 85068 4922 85092 4924
rect 84930 4870 84932 4922
rect 84994 4870 85006 4922
rect 85068 4870 85070 4922
rect 84908 4868 84932 4870
rect 84988 4868 85012 4870
rect 85068 4868 85092 4870
rect 84852 4848 85148 4868
rect 86788 4826 86816 5102
rect 86776 4820 86828 4826
rect 86776 4762 86828 4768
rect 87800 4690 87828 5102
rect 87788 4684 87840 4690
rect 87788 4626 87840 4632
rect 84852 3836 85148 3856
rect 84908 3834 84932 3836
rect 84988 3834 85012 3836
rect 85068 3834 85092 3836
rect 84930 3782 84932 3834
rect 84994 3782 85006 3834
rect 85068 3782 85070 3834
rect 84908 3780 84932 3782
rect 84988 3780 85012 3782
rect 85068 3780 85092 3782
rect 84852 3760 85148 3780
rect 85210 3632 85266 3641
rect 85210 3567 85266 3576
rect 84852 2748 85148 2768
rect 84908 2746 84932 2748
rect 84988 2746 85012 2748
rect 85068 2746 85092 2748
rect 84930 2694 84932 2746
rect 84994 2694 85006 2746
rect 85068 2694 85070 2746
rect 84908 2692 84932 2694
rect 84988 2692 85012 2694
rect 85068 2692 85092 2694
rect 84852 2672 85148 2692
rect 84752 2100 84804 2106
rect 84752 2042 84804 2048
rect 84660 1964 84712 1970
rect 84660 1906 84712 1912
rect 84568 1896 84620 1902
rect 84568 1838 84620 1844
rect 84580 1358 84608 1838
rect 84672 1562 84700 1906
rect 84852 1660 85148 1680
rect 84908 1658 84932 1660
rect 84988 1658 85012 1660
rect 85068 1658 85092 1660
rect 84930 1606 84932 1658
rect 84994 1606 85006 1658
rect 85068 1606 85070 1658
rect 84908 1604 84932 1606
rect 84988 1604 85012 1606
rect 85068 1604 85092 1606
rect 84852 1584 85148 1604
rect 84660 1556 84712 1562
rect 84660 1498 84712 1504
rect 84568 1352 84620 1358
rect 84568 1294 84620 1300
rect 84844 944 84896 950
rect 84844 886 84896 892
rect 84856 800 84884 886
rect 85224 800 85252 3567
rect 85948 3392 86000 3398
rect 85948 3334 86000 3340
rect 85764 2576 85816 2582
rect 85764 2518 85816 2524
rect 85776 2106 85804 2518
rect 85764 2100 85816 2106
rect 85764 2042 85816 2048
rect 85672 1964 85724 1970
rect 85672 1906 85724 1912
rect 85580 1760 85632 1766
rect 85580 1702 85632 1708
rect 85488 1216 85540 1222
rect 85488 1158 85540 1164
rect 84016 750 84068 756
rect 84106 0 84162 800
rect 84292 672 84344 678
rect 84292 614 84344 620
rect 84304 377 84332 614
rect 84290 368 84346 377
rect 84290 303 84346 312
rect 84474 0 84530 800
rect 84842 592 84898 800
rect 84842 572 85148 592
rect 84842 516 84852 572
rect 84908 570 84932 572
rect 84988 570 85012 572
rect 85068 570 85092 572
rect 84930 518 84932 570
rect 84994 518 85006 570
rect 85068 518 85070 570
rect 84908 516 84932 518
rect 84988 516 85012 518
rect 85068 516 85092 518
rect 84842 496 85148 516
rect 84842 0 84898 496
rect 85210 0 85266 800
rect 85500 105 85528 1158
rect 85592 800 85620 1702
rect 85684 1426 85712 1906
rect 85672 1420 85724 1426
rect 85672 1362 85724 1368
rect 85960 800 85988 3334
rect 86684 3120 86736 3126
rect 86684 3062 86736 3068
rect 86316 2984 86368 2990
rect 86316 2926 86368 2932
rect 86328 1970 86356 2926
rect 86316 1964 86368 1970
rect 86316 1906 86368 1912
rect 86500 1216 86552 1222
rect 86500 1158 86552 1164
rect 86512 1057 86540 1158
rect 86498 1048 86554 1057
rect 86498 983 86554 992
rect 86316 944 86368 950
rect 86316 886 86368 892
rect 86328 800 86356 886
rect 86696 800 86724 3062
rect 87328 3052 87380 3058
rect 87328 2994 87380 3000
rect 86958 2952 87014 2961
rect 86958 2887 87014 2896
rect 86972 2650 87000 2887
rect 87340 2825 87368 2994
rect 88168 2990 88196 6938
rect 88444 6866 88472 11614
rect 88524 9580 88576 9586
rect 88524 9522 88576 9528
rect 88536 9382 88564 9522
rect 88524 9376 88576 9382
rect 88524 9318 88576 9324
rect 88432 6860 88484 6866
rect 88432 6802 88484 6808
rect 88536 6662 88564 9318
rect 88524 6656 88576 6662
rect 88524 6598 88576 6604
rect 88720 5778 88748 12200
rect 89088 7342 89116 12200
rect 89260 8492 89312 8498
rect 89260 8434 89312 8440
rect 89272 8022 89300 8434
rect 89260 8016 89312 8022
rect 89260 7958 89312 7964
rect 89076 7336 89128 7342
rect 89076 7278 89128 7284
rect 88708 5772 88760 5778
rect 88708 5714 88760 5720
rect 89456 5166 89484 12200
rect 89824 9110 89852 12200
rect 89904 9512 89956 9518
rect 89904 9454 89956 9460
rect 89812 9104 89864 9110
rect 89812 9046 89864 9052
rect 89916 8974 89944 9454
rect 90192 9382 90220 12200
rect 90364 11008 90416 11014
rect 90364 10950 90416 10956
rect 90376 10810 90404 10950
rect 90364 10804 90416 10810
rect 90364 10746 90416 10752
rect 90376 10130 90404 10746
rect 90364 10124 90416 10130
rect 90364 10066 90416 10072
rect 90272 9512 90324 9518
rect 90272 9454 90324 9460
rect 90180 9376 90232 9382
rect 90180 9318 90232 9324
rect 89904 8968 89956 8974
rect 89904 8910 89956 8916
rect 89536 8832 89588 8838
rect 89536 8774 89588 8780
rect 89548 6458 89576 8774
rect 90284 8634 90312 9454
rect 90272 8628 90324 8634
rect 90272 8570 90324 8576
rect 90284 7954 90312 8570
rect 90456 8560 90508 8566
rect 90456 8502 90508 8508
rect 90468 8430 90496 8502
rect 90456 8424 90508 8430
rect 90456 8366 90508 8372
rect 90272 7948 90324 7954
rect 90272 7890 90324 7896
rect 90468 7478 90496 8366
rect 90456 7472 90508 7478
rect 90456 7414 90508 7420
rect 89536 6452 89588 6458
rect 89536 6394 89588 6400
rect 89996 6384 90048 6390
rect 89996 6326 90048 6332
rect 89444 5160 89496 5166
rect 89444 5102 89496 5108
rect 88892 4208 88944 4214
rect 88892 4150 88944 4156
rect 88432 3596 88484 3602
rect 88432 3538 88484 3544
rect 88340 3392 88392 3398
rect 88340 3334 88392 3340
rect 88156 2984 88208 2990
rect 88156 2926 88208 2932
rect 87420 2848 87472 2854
rect 87326 2816 87382 2825
rect 87420 2790 87472 2796
rect 87326 2751 87382 2760
rect 87340 2650 87368 2751
rect 86960 2644 87012 2650
rect 86960 2586 87012 2592
rect 87328 2644 87380 2650
rect 87328 2586 87380 2592
rect 86972 2446 87000 2586
rect 86960 2440 87012 2446
rect 86960 2382 87012 2388
rect 87236 1964 87288 1970
rect 87236 1906 87288 1912
rect 87248 1358 87276 1906
rect 87432 1562 87460 2790
rect 87602 2680 87658 2689
rect 87602 2615 87604 2624
rect 87656 2615 87658 2624
rect 87604 2586 87656 2592
rect 88352 2582 88380 3334
rect 88444 3194 88472 3538
rect 88800 3392 88852 3398
rect 88800 3334 88852 3340
rect 88812 3194 88840 3334
rect 88432 3188 88484 3194
rect 88432 3130 88484 3136
rect 88800 3188 88852 3194
rect 88800 3130 88852 3136
rect 88432 3052 88484 3058
rect 88432 2994 88484 3000
rect 88444 2802 88472 2994
rect 88524 2848 88576 2854
rect 88444 2796 88524 2802
rect 88444 2790 88576 2796
rect 88444 2774 88564 2790
rect 88444 2650 88472 2774
rect 88432 2644 88484 2650
rect 88432 2586 88484 2592
rect 88340 2576 88392 2582
rect 88340 2518 88392 2524
rect 88800 2372 88852 2378
rect 88800 2314 88852 2320
rect 88616 2304 88668 2310
rect 88154 2272 88210 2281
rect 88616 2246 88668 2252
rect 88154 2207 88210 2216
rect 88168 1834 88196 2207
rect 88628 2038 88656 2246
rect 88616 2032 88668 2038
rect 88616 1974 88668 1980
rect 88432 1964 88484 1970
rect 88432 1906 88484 1912
rect 88156 1828 88208 1834
rect 88156 1770 88208 1776
rect 87420 1556 87472 1562
rect 87420 1498 87472 1504
rect 87420 1420 87472 1426
rect 87420 1362 87472 1368
rect 87236 1352 87288 1358
rect 87236 1294 87288 1300
rect 87052 1216 87104 1222
rect 87052 1158 87104 1164
rect 87064 800 87092 1158
rect 87432 800 87460 1362
rect 88444 1358 88472 1906
rect 88432 1352 88484 1358
rect 88432 1294 88484 1300
rect 88812 1306 88840 2314
rect 88904 2106 88932 4150
rect 89168 4140 89220 4146
rect 89168 4082 89220 4088
rect 89180 3738 89208 4082
rect 90008 4078 90036 6326
rect 90272 6248 90324 6254
rect 90272 6190 90324 6196
rect 90284 5914 90312 6190
rect 90272 5908 90324 5914
rect 90272 5850 90324 5856
rect 90364 5092 90416 5098
rect 90364 5034 90416 5040
rect 90376 4622 90404 5034
rect 90560 4758 90588 12200
rect 90928 10674 90956 12200
rect 90916 10668 90968 10674
rect 90916 10610 90968 10616
rect 91192 9376 91244 9382
rect 91192 9318 91244 9324
rect 91100 8356 91152 8362
rect 91100 8298 91152 8304
rect 91112 7954 91140 8298
rect 91100 7948 91152 7954
rect 91100 7890 91152 7896
rect 91204 6254 91232 9318
rect 91296 8276 91324 12200
rect 91664 9518 91692 12200
rect 91744 11688 91796 11694
rect 91744 11630 91796 11636
rect 91756 11082 91784 11630
rect 92032 11200 92060 12200
rect 92032 11172 92152 11200
rect 91744 11076 91796 11082
rect 91744 11018 91796 11024
rect 92020 11076 92072 11082
rect 92020 11018 92072 11024
rect 91756 10810 91784 11018
rect 91744 10804 91796 10810
rect 91744 10746 91796 10752
rect 91928 10056 91980 10062
rect 91928 9998 91980 10004
rect 91652 9512 91704 9518
rect 91652 9454 91704 9460
rect 91652 8492 91704 8498
rect 91652 8434 91704 8440
rect 91296 8248 91416 8276
rect 91284 7880 91336 7886
rect 91284 7822 91336 7828
rect 91296 7478 91324 7822
rect 91284 7472 91336 7478
rect 91284 7414 91336 7420
rect 91388 6798 91416 8248
rect 91664 7818 91692 8434
rect 91652 7812 91704 7818
rect 91652 7754 91704 7760
rect 91376 6792 91428 6798
rect 91376 6734 91428 6740
rect 91836 6316 91888 6322
rect 91836 6258 91888 6264
rect 91192 6248 91244 6254
rect 91192 6190 91244 6196
rect 91284 5636 91336 5642
rect 91284 5578 91336 5584
rect 90732 5568 90784 5574
rect 90732 5510 90784 5516
rect 90548 4752 90600 4758
rect 90548 4694 90600 4700
rect 90364 4616 90416 4622
rect 90364 4558 90416 4564
rect 89996 4072 90048 4078
rect 89442 4040 89498 4049
rect 89996 4014 90048 4020
rect 89442 3975 89498 3984
rect 89260 3936 89312 3942
rect 89260 3878 89312 3884
rect 89168 3732 89220 3738
rect 89168 3674 89220 3680
rect 88892 2100 88944 2106
rect 88892 2042 88944 2048
rect 88904 1426 88932 2042
rect 89272 1970 89300 3878
rect 89456 3670 89484 3975
rect 89444 3664 89496 3670
rect 89444 3606 89496 3612
rect 89996 3392 90048 3398
rect 89996 3334 90048 3340
rect 90456 3392 90508 3398
rect 90456 3334 90508 3340
rect 89718 2680 89774 2689
rect 89718 2615 89774 2624
rect 89260 1964 89312 1970
rect 89260 1906 89312 1912
rect 89732 1426 89760 2615
rect 89904 2304 89956 2310
rect 89904 2246 89956 2252
rect 88892 1420 88944 1426
rect 88892 1362 88944 1368
rect 89720 1420 89772 1426
rect 89720 1362 89772 1368
rect 87788 1284 87840 1290
rect 88812 1278 88932 1306
rect 87788 1226 87840 1232
rect 87604 1216 87656 1222
rect 87604 1158 87656 1164
rect 87616 921 87644 1158
rect 87602 912 87658 921
rect 87602 847 87658 856
rect 87800 800 87828 1226
rect 88156 1216 88208 1222
rect 88156 1158 88208 1164
rect 88168 800 88196 1158
rect 88536 882 88656 898
rect 88536 876 88668 882
rect 88536 870 88616 876
rect 88536 800 88564 870
rect 88616 818 88668 824
rect 88904 800 88932 1278
rect 89628 944 89680 950
rect 89272 882 89392 898
rect 89628 886 89680 892
rect 89916 898 89944 2246
rect 90008 1222 90036 3334
rect 90468 3097 90496 3334
rect 90454 3088 90510 3097
rect 90272 3052 90324 3058
rect 90744 3058 90772 5510
rect 91100 5228 91152 5234
rect 91100 5170 91152 5176
rect 90824 5160 90876 5166
rect 90822 5128 90824 5137
rect 90876 5128 90878 5137
rect 90822 5063 90878 5072
rect 91112 4554 91140 5170
rect 91100 4548 91152 4554
rect 91100 4490 91152 4496
rect 91100 4140 91152 4146
rect 91100 4082 91152 4088
rect 91112 3670 91140 4082
rect 91100 3664 91152 3670
rect 91100 3606 91152 3612
rect 90454 3023 90510 3032
rect 90732 3052 90784 3058
rect 90272 2994 90324 3000
rect 90732 2994 90784 3000
rect 90284 2650 90312 2994
rect 90364 2848 90416 2854
rect 90364 2790 90416 2796
rect 90272 2644 90324 2650
rect 90272 2586 90324 2592
rect 90180 1352 90232 1358
rect 90180 1294 90232 1300
rect 89996 1216 90048 1222
rect 89996 1158 90048 1164
rect 90192 950 90220 1294
rect 90180 944 90232 950
rect 89272 876 89404 882
rect 89272 870 89352 876
rect 89272 800 89300 870
rect 89352 818 89404 824
rect 89640 800 89668 886
rect 89916 870 90036 898
rect 90180 886 90232 892
rect 90008 800 90036 870
rect 90376 800 90404 2790
rect 91296 1902 91324 5578
rect 91848 5574 91876 6258
rect 91836 5568 91888 5574
rect 91836 5510 91888 5516
rect 91836 5024 91888 5030
rect 91836 4966 91888 4972
rect 91744 3664 91796 3670
rect 91744 3606 91796 3612
rect 91468 3392 91520 3398
rect 91468 3334 91520 3340
rect 91374 2544 91430 2553
rect 91374 2479 91376 2488
rect 91428 2479 91430 2488
rect 91376 2450 91428 2456
rect 91284 1896 91336 1902
rect 91284 1838 91336 1844
rect 91296 1562 91324 1838
rect 91284 1556 91336 1562
rect 91284 1498 91336 1504
rect 91100 1352 91152 1358
rect 90744 1300 91100 1306
rect 90744 1294 91152 1300
rect 90744 1278 91140 1294
rect 90744 800 90772 1278
rect 91100 1216 91152 1222
rect 91100 1158 91152 1164
rect 91376 1216 91428 1222
rect 91376 1158 91428 1164
rect 91112 800 91140 1158
rect 85486 96 85542 105
rect 85486 31 85542 40
rect 85578 0 85634 800
rect 85946 0 86002 800
rect 86132 672 86184 678
rect 86132 614 86184 620
rect 86144 241 86172 614
rect 86130 232 86186 241
rect 86130 167 86186 176
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87786 0 87842 800
rect 88154 0 88210 800
rect 88522 0 88578 800
rect 88890 0 88946 800
rect 88982 776 89038 785
rect 88982 711 88984 720
rect 89036 711 89038 720
rect 89076 740 89128 746
rect 88984 682 89036 688
rect 89076 682 89128 688
rect 89088 474 89116 682
rect 89076 468 89128 474
rect 89076 410 89128 416
rect 89258 0 89314 800
rect 89626 0 89682 800
rect 89994 0 90050 800
rect 90362 0 90418 800
rect 90730 0 90786 800
rect 91098 0 91154 800
rect 91388 202 91416 1158
rect 91480 800 91508 3334
rect 91756 898 91784 3606
rect 91848 3058 91876 4966
rect 91940 4078 91968 9998
rect 92032 9586 92060 11018
rect 92020 9580 92072 9586
rect 92020 9522 92072 9528
rect 92032 9178 92060 9522
rect 92020 9172 92072 9178
rect 92020 9114 92072 9120
rect 92020 8832 92072 8838
rect 92020 8774 92072 8780
rect 92032 6390 92060 8774
rect 92124 8430 92152 11172
rect 92400 10198 92428 12200
rect 92664 11756 92716 11762
rect 92664 11698 92716 11704
rect 92388 10192 92440 10198
rect 92388 10134 92440 10140
rect 92676 10062 92704 11698
rect 92768 10130 92796 12200
rect 93136 11694 93164 12200
rect 93504 11778 93532 12200
rect 93872 11914 93900 12200
rect 93872 11886 93992 11914
rect 93308 11756 93360 11762
rect 93504 11750 93900 11778
rect 93308 11698 93360 11704
rect 93124 11688 93176 11694
rect 93124 11630 93176 11636
rect 93320 11286 93348 11698
rect 93676 11688 93728 11694
rect 93676 11630 93728 11636
rect 93308 11280 93360 11286
rect 93308 11222 93360 11228
rect 93688 11218 93716 11630
rect 93872 11218 93900 11750
rect 93676 11212 93728 11218
rect 93676 11154 93728 11160
rect 93860 11212 93912 11218
rect 93860 11154 93912 11160
rect 93124 10600 93176 10606
rect 93124 10542 93176 10548
rect 92756 10124 92808 10130
rect 92756 10066 92808 10072
rect 92664 10056 92716 10062
rect 92664 9998 92716 10004
rect 93136 9926 93164 10542
rect 93492 10260 93544 10266
rect 93492 10202 93544 10208
rect 93308 10056 93360 10062
rect 93308 9998 93360 10004
rect 93124 9920 93176 9926
rect 93124 9862 93176 9868
rect 92756 9580 92808 9586
rect 92756 9522 92808 9528
rect 92768 8838 92796 9522
rect 92848 9512 92900 9518
rect 92848 9454 92900 9460
rect 92756 8832 92808 8838
rect 92756 8774 92808 8780
rect 92112 8424 92164 8430
rect 92112 8366 92164 8372
rect 92020 6384 92072 6390
rect 92020 6326 92072 6332
rect 92296 5228 92348 5234
rect 92296 5170 92348 5176
rect 92204 4548 92256 4554
rect 92204 4490 92256 4496
rect 91928 4072 91980 4078
rect 91928 4014 91980 4020
rect 91836 3052 91888 3058
rect 91836 2994 91888 3000
rect 92020 2440 92072 2446
rect 92020 2382 92072 2388
rect 91928 1964 91980 1970
rect 91928 1906 91980 1912
rect 91940 1426 91968 1906
rect 91928 1420 91980 1426
rect 91928 1362 91980 1368
rect 92032 950 92060 2382
rect 92020 944 92072 950
rect 91756 870 91876 898
rect 92020 886 92072 892
rect 91848 800 91876 870
rect 92216 800 92244 4490
rect 92308 4486 92336 5170
rect 92768 4826 92796 8774
rect 92860 8498 92888 9454
rect 93136 9042 93164 9862
rect 93320 9722 93348 9998
rect 93400 9920 93452 9926
rect 93400 9862 93452 9868
rect 93412 9722 93440 9862
rect 93504 9722 93532 10202
rect 93308 9716 93360 9722
rect 93308 9658 93360 9664
rect 93400 9716 93452 9722
rect 93400 9658 93452 9664
rect 93492 9716 93544 9722
rect 93492 9658 93544 9664
rect 93964 9178 93992 11886
rect 94240 10146 94268 12200
rect 94240 10118 94360 10146
rect 94228 10056 94280 10062
rect 94228 9998 94280 10004
rect 93952 9172 94004 9178
rect 93952 9114 94004 9120
rect 93124 9036 93176 9042
rect 93124 8978 93176 8984
rect 92848 8492 92900 8498
rect 92848 8434 92900 8440
rect 92860 8090 92888 8434
rect 92848 8084 92900 8090
rect 92848 8026 92900 8032
rect 93216 5976 93268 5982
rect 93216 5918 93268 5924
rect 92940 5364 92992 5370
rect 92940 5306 92992 5312
rect 92756 4820 92808 4826
rect 92756 4762 92808 4768
rect 92296 4480 92348 4486
rect 92296 4422 92348 4428
rect 92296 4140 92348 4146
rect 92296 4082 92348 4088
rect 92308 3398 92336 4082
rect 92572 3732 92624 3738
rect 92572 3674 92624 3680
rect 92296 3392 92348 3398
rect 92296 3334 92348 3340
rect 92308 1562 92336 3334
rect 92296 1556 92348 1562
rect 92296 1498 92348 1504
rect 92584 800 92612 3674
rect 92952 800 92980 5306
rect 93228 3738 93256 5918
rect 93216 3732 93268 3738
rect 93216 3674 93268 3680
rect 94240 3466 94268 9998
rect 94332 9586 94360 10118
rect 94320 9580 94372 9586
rect 94320 9522 94372 9528
rect 94320 9376 94372 9382
rect 94320 9318 94372 9324
rect 94332 8974 94360 9318
rect 94320 8968 94372 8974
rect 94320 8910 94372 8916
rect 94332 7478 94360 8910
rect 94608 8498 94636 12200
rect 94976 8566 95004 12200
rect 95146 8936 95202 8945
rect 95146 8871 95202 8880
rect 94964 8560 95016 8566
rect 95160 8537 95188 8871
rect 94964 8502 95016 8508
rect 95146 8528 95202 8537
rect 94596 8492 94648 8498
rect 95146 8463 95202 8472
rect 94596 8434 94648 8440
rect 94320 7472 94372 7478
rect 94320 7414 94372 7420
rect 95344 7002 95372 12200
rect 95516 11552 95568 11558
rect 95516 11494 95568 11500
rect 95528 11218 95556 11494
rect 95516 11212 95568 11218
rect 95516 11154 95568 11160
rect 95528 10810 95556 11154
rect 95516 10804 95568 10810
rect 95516 10746 95568 10752
rect 95712 9450 95740 12200
rect 96080 10674 96108 12200
rect 96068 10668 96120 10674
rect 96068 10610 96120 10616
rect 95884 10600 95936 10606
rect 95884 10542 95936 10548
rect 95896 10266 95924 10542
rect 95884 10260 95936 10266
rect 95884 10202 95936 10208
rect 95700 9444 95752 9450
rect 95700 9386 95752 9392
rect 96252 8832 96304 8838
rect 96252 8774 96304 8780
rect 95608 8356 95660 8362
rect 95608 8298 95660 8304
rect 95332 6996 95384 7002
rect 95332 6938 95384 6944
rect 95620 6866 95648 8298
rect 95608 6860 95660 6866
rect 95608 6802 95660 6808
rect 96264 6730 96292 8774
rect 96448 7682 96476 12200
rect 96620 11552 96672 11558
rect 96620 11494 96672 11500
rect 96632 11150 96660 11494
rect 96816 11370 96844 12200
rect 96908 11830 96936 12446
rect 97170 12200 97226 13000
rect 97538 12200 97594 13000
rect 97906 12200 97962 13000
rect 98184 12640 98236 12646
rect 98184 12582 98236 12588
rect 96896 11824 96948 11830
rect 96896 11766 96948 11772
rect 96816 11342 96936 11370
rect 96804 11280 96856 11286
rect 96804 11222 96856 11228
rect 96620 11144 96672 11150
rect 96620 11086 96672 11092
rect 96620 9512 96672 9518
rect 96620 9454 96672 9460
rect 96632 8838 96660 9454
rect 96816 9178 96844 11222
rect 96804 9172 96856 9178
rect 96804 9114 96856 9120
rect 96620 8832 96672 8838
rect 96620 8774 96672 8780
rect 96632 8430 96660 8774
rect 96620 8424 96672 8430
rect 96620 8366 96672 8372
rect 96436 7676 96488 7682
rect 96436 7618 96488 7624
rect 96908 7342 96936 11342
rect 97184 7750 97212 12200
rect 97552 10962 97580 12200
rect 97552 10934 97672 10962
rect 97538 10840 97594 10849
rect 97538 10775 97594 10784
rect 97552 10198 97580 10775
rect 97540 10192 97592 10198
rect 97540 10134 97592 10140
rect 97644 9654 97672 10934
rect 97920 9738 97948 12200
rect 98196 11762 98224 12582
rect 98274 12200 98330 13000
rect 98642 12200 98698 13000
rect 99010 12200 99066 13000
rect 99378 12200 99434 13000
rect 99746 12200 99802 13000
rect 100114 12200 100170 13000
rect 100482 12200 100538 13000
rect 100850 12200 100906 13000
rect 101218 12200 101274 13000
rect 101586 12200 101642 13000
rect 101954 12200 102010 13000
rect 102322 12200 102378 13000
rect 102690 12200 102746 13000
rect 103058 12200 103114 13000
rect 103426 12200 103482 13000
rect 103794 12200 103850 13000
rect 104162 12200 104218 13000
rect 104530 12200 104586 13000
rect 104898 12200 104954 13000
rect 105266 12200 105322 13000
rect 105634 12200 105690 13000
rect 106002 12200 106058 13000
rect 106370 12200 106426 13000
rect 106738 12200 106794 13000
rect 107106 12200 107162 13000
rect 107474 12200 107530 13000
rect 107842 12200 107898 13000
rect 108028 12232 108080 12238
rect 98184 11756 98236 11762
rect 98184 11698 98236 11704
rect 98196 11354 98224 11698
rect 98288 11642 98316 12200
rect 98288 11614 98500 11642
rect 98276 11552 98328 11558
rect 98276 11494 98328 11500
rect 98184 11348 98236 11354
rect 98184 11290 98236 11296
rect 98288 10266 98316 11494
rect 98368 10600 98420 10606
rect 98368 10542 98420 10548
rect 98380 10266 98408 10542
rect 98276 10260 98328 10266
rect 98276 10202 98328 10208
rect 98368 10260 98420 10266
rect 98368 10202 98420 10208
rect 98368 9920 98420 9926
rect 98366 9888 98368 9897
rect 98420 9888 98422 9897
rect 98366 9823 98422 9832
rect 97828 9710 97948 9738
rect 97632 9648 97684 9654
rect 97828 9625 97856 9710
rect 97632 9590 97684 9596
rect 97814 9616 97870 9625
rect 97814 9551 97870 9560
rect 97908 9580 97960 9586
rect 97908 9522 97960 9528
rect 97920 9042 97948 9522
rect 98184 9512 98236 9518
rect 98184 9454 98236 9460
rect 98196 9178 98224 9454
rect 98184 9172 98236 9178
rect 98184 9114 98236 9120
rect 97908 9036 97960 9042
rect 97908 8978 97960 8984
rect 97264 8832 97316 8838
rect 97264 8774 97316 8780
rect 97172 7744 97224 7750
rect 97172 7686 97224 7692
rect 96528 7336 96580 7342
rect 96528 7278 96580 7284
rect 96896 7336 96948 7342
rect 96896 7278 96948 7284
rect 96540 7188 96568 7278
rect 96540 7160 96660 7188
rect 96632 7041 96660 7160
rect 96618 7032 96674 7041
rect 96618 6967 96674 6976
rect 96252 6724 96304 6730
rect 96252 6666 96304 6672
rect 97276 6322 97304 8774
rect 98276 8628 98328 8634
rect 98276 8570 98328 8576
rect 98000 8492 98052 8498
rect 98000 8434 98052 8440
rect 98012 8294 98040 8434
rect 98000 8288 98052 8294
rect 98000 8230 98052 8236
rect 98012 6458 98040 8230
rect 98000 6452 98052 6458
rect 98000 6394 98052 6400
rect 97264 6316 97316 6322
rect 97264 6258 97316 6264
rect 98288 5953 98316 8570
rect 98472 7954 98500 11614
rect 98460 7948 98512 7954
rect 98460 7890 98512 7896
rect 98656 7478 98684 12200
rect 98920 10668 98972 10674
rect 98920 10610 98972 10616
rect 98932 10130 98960 10610
rect 98920 10124 98972 10130
rect 98920 10066 98972 10072
rect 99024 8974 99052 12200
rect 99012 8968 99064 8974
rect 99012 8910 99064 8916
rect 99392 8294 99420 12200
rect 99472 11688 99524 11694
rect 99472 11630 99524 11636
rect 99484 11218 99512 11630
rect 99472 11212 99524 11218
rect 99472 11154 99524 11160
rect 99564 10600 99616 10606
rect 99564 10542 99616 10548
rect 99576 10266 99604 10542
rect 99564 10260 99616 10266
rect 99564 10202 99616 10208
rect 99760 9602 99788 12200
rect 99760 9574 99972 9602
rect 99748 9512 99800 9518
rect 99748 9454 99800 9460
rect 99656 9376 99708 9382
rect 99656 9318 99708 9324
rect 99564 9036 99616 9042
rect 99564 8978 99616 8984
rect 99380 8288 99432 8294
rect 99380 8230 99432 8236
rect 98644 7472 98696 7478
rect 98644 7414 98696 7420
rect 99286 6488 99342 6497
rect 99286 6423 99342 6432
rect 99300 6052 99328 6423
rect 98274 5944 98330 5953
rect 98274 5879 98330 5888
rect 99104 5568 99156 5574
rect 99104 5510 99156 5516
rect 99116 5438 99144 5510
rect 99104 5432 99156 5438
rect 99104 5374 99156 5380
rect 94964 4480 95016 4486
rect 95016 4428 95280 4434
rect 94964 4422 95280 4428
rect 94976 4406 95280 4422
rect 94228 3460 94280 3466
rect 94228 3402 94280 3408
rect 93308 3188 93360 3194
rect 93308 3130 93360 3136
rect 93320 800 93348 3130
rect 95054 2952 95110 2961
rect 95054 2887 95110 2896
rect 95068 1698 95096 2887
rect 95146 2816 95202 2825
rect 95146 2751 95202 2760
rect 95160 1834 95188 2751
rect 95148 1828 95200 1834
rect 95148 1770 95200 1776
rect 95056 1692 95108 1698
rect 95056 1634 95108 1640
rect 94780 1352 94832 1358
rect 94780 1294 94832 1300
rect 94044 1216 94096 1222
rect 94044 1158 94096 1164
rect 93676 944 93728 950
rect 93676 886 93728 892
rect 93688 800 93716 886
rect 94056 800 94084 1158
rect 94412 944 94464 950
rect 94412 886 94464 892
rect 94424 800 94452 886
rect 94792 800 94820 1294
rect 95252 1034 95280 4406
rect 99576 4185 99604 8978
rect 99668 8974 99696 9318
rect 99760 9178 99788 9454
rect 99944 9178 99972 9574
rect 99748 9172 99800 9178
rect 99748 9114 99800 9120
rect 99932 9172 99984 9178
rect 99932 9114 99984 9120
rect 100128 9110 100156 12200
rect 100116 9104 100168 9110
rect 100496 9058 100524 12200
rect 100668 11076 100720 11082
rect 100668 11018 100720 11024
rect 100116 9046 100168 9052
rect 100404 9030 100524 9058
rect 100576 9104 100628 9110
rect 100576 9046 100628 9052
rect 99656 8968 99708 8974
rect 99656 8910 99708 8916
rect 100300 8492 100352 8498
rect 100300 8434 100352 8440
rect 100312 8362 100340 8434
rect 100300 8356 100352 8362
rect 100300 8298 100352 8304
rect 99562 4176 99618 4185
rect 99562 4111 99618 4120
rect 100312 4078 100340 8298
rect 100404 7954 100432 9030
rect 100588 8974 100616 9046
rect 100484 8968 100536 8974
rect 100484 8910 100536 8916
rect 100576 8968 100628 8974
rect 100576 8910 100628 8916
rect 100496 8838 100524 8910
rect 100484 8832 100536 8838
rect 100484 8774 100536 8780
rect 100392 7948 100444 7954
rect 100392 7890 100444 7896
rect 100392 7540 100444 7546
rect 100392 7482 100444 7488
rect 100404 4758 100432 7482
rect 100392 4752 100444 4758
rect 100392 4694 100444 4700
rect 100392 4480 100444 4486
rect 100392 4422 100444 4428
rect 100300 4072 100352 4078
rect 100300 4014 100352 4020
rect 100208 3936 100260 3942
rect 100208 3878 100260 3884
rect 100024 3664 100076 3670
rect 100024 3606 100076 3612
rect 100036 3482 100064 3606
rect 99944 3454 100064 3482
rect 96620 1828 96672 1834
rect 96620 1770 96672 1776
rect 97724 1828 97776 1834
rect 97724 1770 97776 1776
rect 95976 1624 96028 1630
rect 95634 1572 95976 1578
rect 95634 1566 96028 1572
rect 95634 1550 96016 1566
rect 96252 1284 96304 1290
rect 96252 1226 96304 1232
rect 95252 1006 95924 1034
rect 95068 870 95188 898
rect 91376 196 91428 202
rect 91376 138 91428 144
rect 91466 0 91522 800
rect 91834 0 91890 800
rect 92202 0 92258 800
rect 92570 0 92626 800
rect 92938 0 92994 800
rect 93306 0 93362 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95068 338 95096 870
rect 95160 800 95188 870
rect 95528 870 95648 898
rect 95528 800 95556 870
rect 95056 332 95108 338
rect 95056 274 95108 280
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95620 678 95648 870
rect 95896 800 95924 1006
rect 96264 800 96292 1226
rect 96632 800 96660 1770
rect 96988 1692 97040 1698
rect 96988 1634 97040 1640
rect 97000 800 97028 1634
rect 97356 1080 97408 1086
rect 97356 1022 97408 1028
rect 97368 800 97396 1022
rect 97736 800 97764 1770
rect 98826 1728 98882 1737
rect 98826 1663 98882 1672
rect 98090 1184 98146 1193
rect 98090 1119 98146 1128
rect 98104 800 98132 1119
rect 98472 870 98592 898
rect 98472 800 98500 870
rect 95608 672 95660 678
rect 95608 614 95660 620
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96618 0 96674 800
rect 96986 0 97042 800
rect 97354 0 97410 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98458 0 98514 800
rect 98564 406 98592 870
rect 98840 800 98868 1663
rect 99472 1624 99524 1630
rect 99472 1566 99524 1572
rect 99196 1556 99248 1562
rect 99196 1498 99248 1504
rect 99208 800 99236 1498
rect 99484 1426 99512 1566
rect 99472 1420 99524 1426
rect 99472 1362 99524 1368
rect 99564 1420 99616 1426
rect 99564 1362 99616 1368
rect 99576 800 99604 1362
rect 99944 800 99972 3454
rect 100024 3392 100076 3398
rect 100024 3334 100076 3340
rect 100036 1766 100064 3334
rect 100116 2848 100168 2854
rect 100116 2790 100168 2796
rect 100024 1760 100076 1766
rect 100024 1702 100076 1708
rect 100128 1630 100156 2790
rect 100116 1624 100168 1630
rect 100116 1566 100168 1572
rect 100220 1494 100248 3878
rect 100300 3596 100352 3602
rect 100300 3538 100352 3544
rect 100312 1698 100340 3538
rect 100404 1737 100432 4422
rect 100496 4146 100524 8774
rect 100576 6656 100628 6662
rect 100576 6598 100628 6604
rect 100588 4622 100616 6598
rect 100680 5930 100708 11018
rect 100864 10282 100892 12200
rect 100864 10254 100984 10282
rect 100852 10124 100904 10130
rect 100852 10066 100904 10072
rect 100864 9654 100892 10066
rect 100852 9648 100904 9654
rect 100852 9590 100904 9596
rect 100956 9450 100984 10254
rect 101036 9580 101088 9586
rect 101036 9522 101088 9528
rect 100944 9444 100996 9450
rect 100944 9386 100996 9392
rect 101048 8838 101076 9522
rect 101036 8832 101088 8838
rect 101036 8774 101088 8780
rect 100944 6112 100996 6118
rect 100944 6054 100996 6060
rect 100680 5902 100800 5930
rect 100666 5808 100722 5817
rect 100666 5743 100722 5752
rect 100576 4616 100628 4622
rect 100576 4558 100628 4564
rect 100484 4140 100536 4146
rect 100484 4082 100536 4088
rect 100484 4004 100536 4010
rect 100484 3946 100536 3952
rect 100390 1728 100446 1737
rect 100300 1692 100352 1698
rect 100390 1663 100446 1672
rect 100300 1634 100352 1640
rect 100208 1488 100260 1494
rect 100496 1442 100524 3946
rect 100576 3732 100628 3738
rect 100576 3674 100628 3680
rect 100208 1430 100260 1436
rect 100312 1414 100524 1442
rect 100588 1426 100616 3674
rect 100680 2038 100708 5743
rect 100772 5234 100800 5902
rect 100760 5228 100812 5234
rect 100760 5170 100812 5176
rect 100956 5137 100984 6054
rect 100942 5128 100998 5137
rect 100942 5063 100998 5072
rect 101048 4729 101076 8774
rect 101232 8362 101260 12200
rect 101404 12096 101456 12102
rect 101404 12038 101456 12044
rect 101416 11354 101444 12038
rect 101404 11348 101456 11354
rect 101404 11290 101456 11296
rect 101600 10146 101628 12200
rect 101864 11688 101916 11694
rect 101864 11630 101916 11636
rect 101876 11218 101904 11630
rect 101864 11212 101916 11218
rect 101864 11154 101916 11160
rect 101772 10668 101824 10674
rect 101772 10610 101824 10616
rect 101600 10118 101720 10146
rect 101588 10056 101640 10062
rect 101588 9998 101640 10004
rect 101220 8356 101272 8362
rect 101220 8298 101272 8304
rect 101404 5636 101456 5642
rect 101404 5578 101456 5584
rect 101416 5545 101444 5578
rect 101402 5536 101458 5545
rect 101402 5471 101458 5480
rect 101034 4720 101090 4729
rect 101034 4655 101090 4664
rect 101600 3126 101628 9998
rect 101692 6254 101720 10118
rect 101784 10062 101812 10610
rect 101772 10056 101824 10062
rect 101772 9998 101824 10004
rect 101968 9110 101996 12200
rect 102232 10600 102284 10606
rect 102232 10542 102284 10548
rect 102244 10130 102272 10542
rect 102232 10124 102284 10130
rect 102232 10066 102284 10072
rect 102140 9920 102192 9926
rect 102140 9862 102192 9868
rect 102230 9888 102286 9897
rect 101956 9104 102008 9110
rect 101956 9046 102008 9052
rect 102152 6798 102180 9862
rect 102230 9823 102286 9832
rect 102140 6792 102192 6798
rect 102140 6734 102192 6740
rect 101680 6248 101732 6254
rect 101680 6190 101732 6196
rect 102244 5574 102272 9823
rect 102336 8294 102364 12200
rect 102704 8566 102732 12200
rect 102876 8832 102928 8838
rect 102876 8774 102928 8780
rect 102692 8560 102744 8566
rect 102692 8502 102744 8508
rect 102888 8498 102916 8774
rect 102876 8492 102928 8498
rect 102876 8434 102928 8440
rect 102324 8288 102376 8294
rect 102324 8230 102376 8236
rect 102888 8090 102916 8434
rect 102876 8084 102928 8090
rect 102876 8026 102928 8032
rect 102324 7744 102376 7750
rect 102324 7686 102376 7692
rect 102336 7410 102364 7686
rect 102324 7404 102376 7410
rect 102324 7346 102376 7352
rect 102336 6934 102364 7346
rect 102324 6928 102376 6934
rect 102324 6870 102376 6876
rect 103072 6662 103100 12200
rect 103152 12164 103204 12170
rect 103152 12106 103204 12112
rect 103164 11218 103192 12106
rect 103152 11212 103204 11218
rect 103152 11154 103204 11160
rect 103244 10600 103296 10606
rect 103244 10542 103296 10548
rect 103256 9625 103284 10542
rect 103336 9920 103388 9926
rect 103336 9862 103388 9868
rect 103242 9616 103298 9625
rect 103242 9551 103298 9560
rect 103348 9518 103376 9862
rect 103336 9512 103388 9518
rect 103336 9454 103388 9460
rect 103348 8906 103376 9454
rect 103336 8900 103388 8906
rect 103336 8842 103388 8848
rect 103336 8628 103388 8634
rect 103336 8570 103388 8576
rect 103348 7954 103376 8570
rect 103336 7948 103388 7954
rect 103336 7890 103388 7896
rect 103060 6656 103112 6662
rect 103060 6598 103112 6604
rect 103336 6248 103388 6254
rect 103334 6216 103336 6225
rect 103388 6216 103390 6225
rect 103334 6151 103390 6160
rect 103440 6089 103468 12200
rect 103808 7954 103836 12200
rect 104072 11756 104124 11762
rect 104072 11698 104124 11704
rect 104084 11354 104112 11698
rect 104072 11348 104124 11354
rect 104072 11290 104124 11296
rect 103980 8968 104032 8974
rect 103980 8910 104032 8916
rect 103992 8498 104020 8910
rect 104176 8906 104204 12200
rect 104256 10668 104308 10674
rect 104256 10610 104308 10616
rect 104268 9926 104296 10610
rect 104256 9920 104308 9926
rect 104256 9862 104308 9868
rect 104164 8900 104216 8906
rect 104164 8842 104216 8848
rect 103980 8492 104032 8498
rect 103980 8434 104032 8440
rect 103796 7948 103848 7954
rect 103796 7890 103848 7896
rect 103980 7404 104032 7410
rect 103980 7346 104032 7352
rect 103992 6934 104020 7346
rect 104070 7032 104126 7041
rect 104070 6967 104126 6976
rect 104084 6934 104112 6967
rect 103980 6928 104032 6934
rect 103980 6870 104032 6876
rect 104072 6928 104124 6934
rect 104072 6870 104124 6876
rect 103992 6633 104020 6870
rect 103978 6624 104034 6633
rect 103978 6559 104034 6568
rect 103520 6180 103572 6186
rect 103520 6122 103572 6128
rect 103426 6080 103482 6089
rect 103426 6015 103482 6024
rect 103426 5944 103482 5953
rect 103532 5930 103560 6122
rect 103610 5944 103666 5953
rect 103532 5902 103610 5930
rect 103426 5879 103482 5888
rect 103610 5879 103666 5888
rect 102232 5568 102284 5574
rect 102232 5510 102284 5516
rect 102140 5364 102192 5370
rect 102140 5306 102192 5312
rect 101588 3120 101640 3126
rect 101588 3062 101640 3068
rect 102152 3058 102180 5306
rect 103060 5160 103112 5166
rect 103060 5102 103112 5108
rect 103072 4690 103100 5102
rect 103060 4684 103112 4690
rect 103060 4626 103112 4632
rect 102232 4140 102284 4146
rect 102232 4082 102284 4088
rect 102244 3466 102272 4082
rect 102324 3528 102376 3534
rect 102324 3470 102376 3476
rect 102968 3528 103020 3534
rect 102968 3470 103020 3476
rect 102232 3460 102284 3466
rect 102232 3402 102284 3408
rect 102140 3052 102192 3058
rect 102140 2994 102192 3000
rect 102140 2644 102192 2650
rect 102140 2586 102192 2592
rect 100760 2304 100812 2310
rect 100760 2246 100812 2252
rect 100668 2032 100720 2038
rect 100668 1974 100720 1980
rect 100576 1420 100628 1426
rect 100312 800 100340 1414
rect 100576 1362 100628 1368
rect 100772 1272 100800 2246
rect 101772 1556 101824 1562
rect 101772 1498 101824 1504
rect 100680 1244 100800 1272
rect 100680 800 100708 1244
rect 101402 1048 101458 1057
rect 101402 983 101458 992
rect 101048 870 101168 898
rect 101048 800 101076 870
rect 98552 400 98604 406
rect 98552 342 98604 348
rect 98826 0 98882 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100298 0 100354 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101140 474 101168 870
rect 101416 800 101444 983
rect 101784 800 101812 1498
rect 102152 800 102180 2586
rect 102336 2258 102364 3470
rect 102980 2650 103008 3470
rect 103440 3398 103468 5879
rect 104072 5636 104124 5642
rect 104072 5578 104124 5584
rect 104084 5166 104112 5578
rect 104072 5160 104124 5166
rect 104072 5102 104124 5108
rect 103796 5092 103848 5098
rect 103796 5034 103848 5040
rect 103808 4758 103836 5034
rect 103796 4752 103848 4758
rect 103796 4694 103848 4700
rect 104268 4010 104296 9862
rect 104348 7744 104400 7750
rect 104348 7686 104400 7692
rect 104360 7206 104388 7686
rect 104544 7342 104572 12200
rect 104912 11778 104940 12200
rect 104912 11750 105032 11778
rect 104900 11620 104952 11626
rect 104900 11562 104952 11568
rect 104912 11354 104940 11562
rect 104900 11348 104952 11354
rect 104900 11290 104952 11296
rect 104624 10600 104676 10606
rect 104624 10542 104676 10548
rect 104636 9926 104664 10542
rect 104624 9920 104676 9926
rect 104624 9862 104676 9868
rect 104636 9654 104664 9862
rect 105004 9654 105032 11750
rect 105280 11642 105308 12200
rect 105280 11614 105400 11642
rect 105268 11552 105320 11558
rect 105268 11494 105320 11500
rect 105280 11354 105308 11494
rect 105268 11348 105320 11354
rect 105268 11290 105320 11296
rect 104624 9648 104676 9654
rect 104624 9590 104676 9596
rect 104992 9648 105044 9654
rect 104992 9590 105044 9596
rect 104716 9580 104768 9586
rect 104716 9522 104768 9528
rect 104728 8838 104756 9522
rect 105372 9042 105400 11614
rect 105648 10538 105676 12200
rect 105636 10532 105688 10538
rect 105636 10474 105688 10480
rect 106016 9586 106044 12200
rect 106186 10840 106242 10849
rect 106186 10775 106188 10784
rect 106240 10775 106242 10784
rect 106188 10746 106240 10752
rect 106188 10668 106240 10674
rect 106188 10610 106240 10616
rect 106200 9926 106228 10610
rect 106188 9920 106240 9926
rect 106188 9862 106240 9868
rect 106188 9716 106240 9722
rect 106188 9658 106240 9664
rect 106004 9580 106056 9586
rect 106004 9522 106056 9528
rect 105360 9036 105412 9042
rect 105360 8978 105412 8984
rect 104716 8832 104768 8838
rect 104716 8774 104768 8780
rect 104624 8492 104676 8498
rect 104624 8434 104676 8440
rect 104636 7750 104664 8434
rect 104624 7744 104676 7750
rect 104624 7686 104676 7692
rect 104532 7336 104584 7342
rect 104532 7278 104584 7284
rect 104348 7200 104400 7206
rect 104348 7142 104400 7148
rect 104360 6582 104664 6610
rect 104360 6390 104388 6582
rect 104440 6452 104492 6458
rect 104440 6394 104492 6400
rect 104348 6384 104400 6390
rect 104348 6326 104400 6332
rect 104452 6100 104480 6394
rect 104636 6390 104664 6582
rect 104714 6488 104770 6497
rect 104714 6423 104716 6432
rect 104768 6423 104770 6432
rect 104716 6394 104768 6400
rect 104624 6384 104676 6390
rect 104624 6326 104676 6332
rect 104808 6248 104860 6254
rect 104808 6190 104860 6196
rect 104820 6100 104848 6190
rect 104452 6072 104572 6100
rect 104728 6089 104848 6100
rect 104440 5704 104492 5710
rect 104440 5646 104492 5652
rect 104452 5545 104480 5646
rect 104544 5574 104572 6072
rect 104714 6080 104848 6089
rect 104770 6072 104848 6080
rect 104714 6015 104770 6024
rect 104532 5568 104584 5574
rect 104438 5536 104494 5545
rect 104532 5510 104584 5516
rect 104438 5471 104494 5480
rect 105648 5324 106044 5352
rect 105648 5234 105676 5324
rect 104440 5228 104492 5234
rect 104440 5170 104492 5176
rect 105636 5228 105688 5234
rect 105636 5170 105688 5176
rect 105820 5228 105872 5234
rect 105872 5188 105952 5216
rect 105820 5170 105872 5176
rect 104452 4826 104480 5170
rect 104440 4820 104492 4826
rect 104440 4762 104492 4768
rect 105924 4486 105952 5188
rect 106016 5166 106044 5324
rect 106200 5234 106228 9658
rect 106280 8832 106332 8838
rect 106280 8774 106332 8780
rect 106292 6610 106320 8774
rect 106384 6730 106412 12200
rect 106556 11688 106608 11694
rect 106556 11630 106608 11636
rect 106568 11354 106596 11630
rect 106556 11348 106608 11354
rect 106556 11290 106608 11296
rect 106752 10198 106780 12200
rect 107120 11642 107148 12200
rect 107120 11614 107240 11642
rect 107108 11552 107160 11558
rect 107108 11494 107160 11500
rect 107120 11218 107148 11494
rect 107108 11212 107160 11218
rect 107108 11154 107160 11160
rect 107212 10305 107240 11614
rect 107198 10296 107254 10305
rect 107198 10231 107254 10240
rect 106740 10192 106792 10198
rect 106740 10134 106792 10140
rect 106556 9036 106608 9042
rect 106556 8978 106608 8984
rect 106568 8922 106596 8978
rect 106568 8906 106688 8922
rect 106568 8900 106700 8906
rect 106568 8894 106648 8900
rect 106648 8842 106700 8848
rect 106464 8832 106516 8838
rect 106464 8774 106516 8780
rect 106476 8498 106504 8774
rect 106464 8492 106516 8498
rect 106464 8434 106516 8440
rect 107108 8492 107160 8498
rect 107108 8434 107160 8440
rect 107120 8090 107148 8434
rect 107108 8084 107160 8090
rect 107108 8026 107160 8032
rect 106556 7812 106608 7818
rect 106556 7754 106608 7760
rect 106372 6724 106424 6730
rect 106372 6666 106424 6672
rect 106292 6582 106504 6610
rect 106370 6488 106426 6497
rect 106370 6423 106426 6432
rect 106280 6384 106332 6390
rect 106384 6338 106412 6423
rect 106332 6332 106412 6338
rect 106280 6326 106412 6332
rect 106292 6310 106412 6326
rect 106280 6248 106332 6254
rect 106332 6208 106412 6236
rect 106280 6190 106332 6196
rect 106384 5953 106412 6208
rect 106370 5944 106426 5953
rect 106370 5879 106426 5888
rect 106476 5370 106504 6582
rect 106464 5364 106516 5370
rect 106464 5306 106516 5312
rect 106188 5228 106240 5234
rect 106188 5170 106240 5176
rect 106004 5160 106056 5166
rect 106004 5102 106056 5108
rect 106094 5128 106150 5137
rect 106094 5063 106096 5072
rect 106148 5063 106150 5072
rect 106096 5034 106148 5040
rect 106188 5024 106240 5030
rect 106188 4966 106240 4972
rect 106200 4729 106228 4966
rect 106186 4720 106242 4729
rect 106186 4655 106242 4664
rect 105912 4480 105964 4486
rect 105912 4422 105964 4428
rect 105924 4282 105952 4422
rect 105912 4276 105964 4282
rect 105912 4218 105964 4224
rect 106464 4140 106516 4146
rect 106464 4082 106516 4088
rect 104256 4004 104308 4010
rect 104256 3946 104308 3952
rect 106476 3466 106504 4082
rect 106464 3460 106516 3466
rect 106464 3402 106516 3408
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103428 3392 103480 3398
rect 103428 3334 103480 3340
rect 103060 2984 103112 2990
rect 103060 2926 103112 2932
rect 102968 2644 103020 2650
rect 102968 2586 103020 2592
rect 102876 2508 102928 2514
rect 102876 2450 102928 2456
rect 102244 2230 102364 2258
rect 102244 1290 102272 2230
rect 102324 2100 102376 2106
rect 102324 2042 102376 2048
rect 102336 1426 102364 2042
rect 102416 1760 102468 1766
rect 102416 1702 102468 1708
rect 102508 1760 102560 1766
rect 102508 1702 102560 1708
rect 102324 1420 102376 1426
rect 102324 1362 102376 1368
rect 102232 1284 102284 1290
rect 102232 1226 102284 1232
rect 102428 1018 102456 1702
rect 102520 1562 102548 1702
rect 102508 1556 102560 1562
rect 102508 1498 102560 1504
rect 102416 1012 102468 1018
rect 102416 954 102468 960
rect 102520 870 102640 898
rect 102520 800 102548 870
rect 102612 814 102640 870
rect 102600 808 102652 814
rect 101128 468 101180 474
rect 101128 410 101180 416
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102888 800 102916 2450
rect 102600 750 102652 756
rect 102874 0 102930 800
rect 103072 678 103100 2926
rect 103244 2848 103296 2854
rect 103244 2790 103296 2796
rect 103256 2650 103284 2790
rect 103244 2644 103296 2650
rect 103244 2586 103296 2592
rect 103256 2378 103284 2586
rect 103244 2372 103296 2378
rect 103244 2314 103296 2320
rect 103348 2106 103376 3334
rect 104440 3188 104492 3194
rect 104440 3130 104492 3136
rect 103520 3120 103572 3126
rect 103440 3068 103520 3074
rect 103440 3062 103572 3068
rect 103440 3046 103560 3062
rect 103336 2100 103388 2106
rect 103336 2042 103388 2048
rect 103440 1442 103468 3046
rect 104164 2984 104216 2990
rect 104164 2926 104216 2932
rect 104348 2984 104400 2990
rect 104348 2926 104400 2932
rect 103888 2848 103940 2854
rect 103888 2790 103940 2796
rect 103900 2514 103928 2790
rect 104176 2650 104204 2926
rect 104256 2848 104308 2854
rect 104256 2790 104308 2796
rect 104164 2644 104216 2650
rect 104164 2586 104216 2592
rect 103888 2508 103940 2514
rect 103888 2450 103940 2456
rect 103256 1414 103468 1442
rect 103518 1456 103574 1465
rect 104268 1442 104296 2790
rect 104360 1970 104388 2926
rect 104348 1964 104400 1970
rect 104348 1906 104400 1912
rect 104360 1562 104388 1906
rect 104348 1556 104400 1562
rect 104348 1498 104400 1504
rect 104452 1442 104480 3130
rect 105452 2984 105504 2990
rect 105452 2926 105504 2932
rect 105268 2916 105320 2922
rect 105268 2858 105320 2864
rect 104992 2304 105044 2310
rect 104992 2246 105044 2252
rect 104900 2032 104952 2038
rect 104900 1974 104952 1980
rect 104808 1896 104860 1902
rect 104808 1838 104860 1844
rect 103256 800 103284 1414
rect 103518 1391 103520 1400
rect 103572 1391 103574 1400
rect 103992 1414 104296 1442
rect 104360 1414 104480 1442
rect 103520 1362 103572 1368
rect 103624 870 103744 898
rect 103624 800 103652 870
rect 103060 672 103112 678
rect 103060 614 103112 620
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103716 649 103744 870
rect 103992 800 104020 1414
rect 104256 876 104308 882
rect 104256 818 104308 824
rect 103702 640 103758 649
rect 103702 575 103758 584
rect 103978 0 104034 800
rect 104268 678 104296 818
rect 104360 800 104388 1414
rect 104820 1057 104848 1838
rect 104912 1193 104940 1974
rect 104898 1184 104954 1193
rect 104898 1119 104954 1128
rect 104806 1048 104862 1057
rect 105004 1018 105032 2246
rect 105280 1970 105308 2858
rect 105268 1964 105320 1970
rect 105268 1906 105320 1912
rect 105280 1562 105308 1906
rect 105268 1556 105320 1562
rect 105268 1498 105320 1504
rect 105268 1352 105320 1358
rect 105188 1300 105268 1306
rect 105188 1294 105320 1300
rect 105188 1278 105308 1294
rect 104806 983 104862 992
rect 104992 1012 105044 1018
rect 104992 954 105044 960
rect 105188 950 105216 1278
rect 105176 944 105228 950
rect 104728 870 104848 898
rect 104728 800 104756 870
rect 104256 672 104308 678
rect 104256 614 104308 620
rect 104268 134 104296 614
rect 104256 128 104308 134
rect 104256 70 104308 76
rect 104346 0 104402 800
rect 104714 0 104770 800
rect 104820 338 104848 870
rect 105004 870 105124 898
rect 105176 886 105228 892
rect 105004 814 105032 870
rect 104992 808 105044 814
rect 105096 800 105124 870
rect 105464 800 105492 2926
rect 106568 2106 106596 7754
rect 107488 6254 107516 12200
rect 107752 11756 107804 11762
rect 107752 11698 107804 11704
rect 107764 11014 107792 11698
rect 107856 11642 107884 12200
rect 108210 12200 108266 13000
rect 108488 12300 108540 12306
rect 108488 12242 108540 12248
rect 108028 12174 108080 12180
rect 107856 11614 107976 11642
rect 107844 11552 107896 11558
rect 107844 11494 107896 11500
rect 107752 11008 107804 11014
rect 107752 10950 107804 10956
rect 107856 10674 107884 11494
rect 107844 10668 107896 10674
rect 107844 10610 107896 10616
rect 107660 10600 107712 10606
rect 107660 10542 107712 10548
rect 107672 10266 107700 10542
rect 107660 10260 107712 10266
rect 107660 10202 107712 10208
rect 107672 10130 107700 10202
rect 107660 10124 107712 10130
rect 107660 10066 107712 10072
rect 107948 9450 107976 11614
rect 108040 11286 108068 12174
rect 108224 12050 108252 12200
rect 108224 12022 108436 12050
rect 108212 11892 108264 11898
rect 108212 11834 108264 11840
rect 108028 11280 108080 11286
rect 108028 11222 108080 11228
rect 108224 11150 108252 11834
rect 108212 11144 108264 11150
rect 108212 11086 108264 11092
rect 108210 9616 108266 9625
rect 108210 9551 108212 9560
rect 108264 9551 108266 9560
rect 108212 9522 108264 9528
rect 108304 9512 108356 9518
rect 108304 9454 108356 9460
rect 107936 9444 107988 9450
rect 107936 9386 107988 9392
rect 108118 9208 108174 9217
rect 108316 9178 108344 9454
rect 108118 9143 108120 9152
rect 108172 9143 108174 9152
rect 108304 9172 108356 9178
rect 108120 9114 108172 9120
rect 108304 9114 108356 9120
rect 108408 8634 108436 12022
rect 108500 11898 108528 12242
rect 108578 12200 108634 13000
rect 108946 12200 109002 13000
rect 109314 12200 109370 13000
rect 109682 12200 109738 13000
rect 109960 12572 110012 12578
rect 109960 12514 110012 12520
rect 108488 11892 108540 11898
rect 108488 11834 108540 11840
rect 108592 11234 108620 12200
rect 108960 11898 108988 12200
rect 108948 11892 109000 11898
rect 108948 11834 109000 11840
rect 109040 11688 109092 11694
rect 109040 11630 109092 11636
rect 108592 11206 108712 11234
rect 108580 11144 108632 11150
rect 108580 11086 108632 11092
rect 108592 11014 108620 11086
rect 108580 11008 108632 11014
rect 108580 10950 108632 10956
rect 108592 9722 108620 10950
rect 108580 9716 108632 9722
rect 108580 9658 108632 9664
rect 108488 9512 108540 9518
rect 108488 9454 108540 9460
rect 108500 9382 108528 9454
rect 108488 9376 108540 9382
rect 108488 9318 108540 9324
rect 108684 9081 108712 11206
rect 109052 11014 109080 11630
rect 109040 11008 109092 11014
rect 109040 10950 109092 10956
rect 108948 10668 109000 10674
rect 108948 10610 109000 10616
rect 108854 10568 108910 10577
rect 108854 10503 108856 10512
rect 108908 10503 108910 10512
rect 108856 10474 108908 10480
rect 108960 10266 108988 10610
rect 108948 10260 109000 10266
rect 108948 10202 109000 10208
rect 109052 9994 109080 10950
rect 109040 9988 109092 9994
rect 109040 9930 109092 9936
rect 108670 9072 108726 9081
rect 108670 9007 108726 9016
rect 108396 8628 108448 8634
rect 108396 8570 108448 8576
rect 108488 8492 108540 8498
rect 108488 8434 108540 8440
rect 108500 8090 108528 8434
rect 108580 8288 108632 8294
rect 108580 8230 108632 8236
rect 108488 8084 108540 8090
rect 108488 8026 108540 8032
rect 108592 7546 108620 8230
rect 108488 7540 108540 7546
rect 108488 7482 108540 7488
rect 108580 7540 108632 7546
rect 108580 7482 108632 7488
rect 107750 6624 107806 6633
rect 107750 6559 107806 6568
rect 107476 6248 107528 6254
rect 107476 6190 107528 6196
rect 107764 6118 107792 6559
rect 107842 6488 107898 6497
rect 107842 6423 107898 6432
rect 107752 6112 107804 6118
rect 107752 6054 107804 6060
rect 106738 5944 106794 5953
rect 106738 5879 106794 5888
rect 106752 5846 106780 5879
rect 106648 5840 106700 5846
rect 106648 5782 106700 5788
rect 106740 5840 106792 5846
rect 106740 5782 106792 5788
rect 106660 4146 106688 5782
rect 107660 5772 107712 5778
rect 107660 5714 107712 5720
rect 107016 4684 107068 4690
rect 107016 4626 107068 4632
rect 106648 4140 106700 4146
rect 106648 4082 106700 4088
rect 106740 3460 106792 3466
rect 106740 3402 106792 3408
rect 106646 2816 106702 2825
rect 106646 2751 106702 2760
rect 106556 2100 106608 2106
rect 106556 2042 106608 2048
rect 106370 1592 106426 1601
rect 106370 1527 106426 1536
rect 106384 1426 106412 1527
rect 106660 1442 106688 2751
rect 106372 1420 106424 1426
rect 106372 1362 106424 1368
rect 106568 1414 106688 1442
rect 105820 1284 105872 1290
rect 105820 1226 105872 1232
rect 105832 800 105860 1226
rect 106096 1216 106148 1222
rect 106096 1158 106148 1164
rect 106108 882 106136 1158
rect 106370 912 106426 921
rect 106096 876 106148 882
rect 106096 818 106148 824
rect 106200 870 106320 898
rect 106200 800 106228 870
rect 104992 750 105044 756
rect 104808 332 104860 338
rect 104808 274 104860 280
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106292 202 106320 870
rect 106370 847 106426 856
rect 106384 814 106412 847
rect 106372 808 106424 814
rect 106568 800 106596 1414
rect 106752 921 106780 3402
rect 107028 2106 107056 4626
rect 107566 4040 107622 4049
rect 107566 3975 107568 3984
rect 107620 3975 107622 3984
rect 107568 3946 107620 3952
rect 107474 3904 107530 3913
rect 107474 3839 107530 3848
rect 107488 3058 107516 3839
rect 107566 3496 107622 3505
rect 107566 3431 107622 3440
rect 107580 3398 107608 3431
rect 107568 3392 107620 3398
rect 107568 3334 107620 3340
rect 107476 3052 107528 3058
rect 107476 2994 107528 3000
rect 107672 2689 107700 5714
rect 107856 4146 107884 6423
rect 108304 6248 108356 6254
rect 108302 6216 108304 6225
rect 108356 6216 108358 6225
rect 108302 6151 108358 6160
rect 107936 5228 107988 5234
rect 107936 5170 107988 5176
rect 107752 4140 107804 4146
rect 107752 4082 107804 4088
rect 107844 4140 107896 4146
rect 107844 4082 107896 4088
rect 107764 3398 107792 4082
rect 107948 4026 107976 5170
rect 108394 4176 108450 4185
rect 108394 4111 108450 4120
rect 108408 4078 108436 4111
rect 107856 3998 107976 4026
rect 108212 4072 108264 4078
rect 108212 4014 108264 4020
rect 108396 4072 108448 4078
rect 108396 4014 108448 4020
rect 107752 3392 107804 3398
rect 107752 3334 107804 3340
rect 107856 3126 107884 3998
rect 107936 3664 107988 3670
rect 107936 3606 107988 3612
rect 108026 3632 108082 3641
rect 107948 3466 107976 3606
rect 108026 3567 108082 3576
rect 108120 3596 108172 3602
rect 108040 3534 108068 3567
rect 108120 3538 108172 3544
rect 108028 3528 108080 3534
rect 108028 3470 108080 3476
rect 107936 3460 107988 3466
rect 107936 3402 107988 3408
rect 108132 3126 108160 3538
rect 108224 3534 108252 4014
rect 108396 3732 108448 3738
rect 108396 3674 108448 3680
rect 108212 3528 108264 3534
rect 108408 3505 108436 3674
rect 108212 3470 108264 3476
rect 108394 3496 108450 3505
rect 108394 3431 108450 3440
rect 107844 3120 107896 3126
rect 107844 3062 107896 3068
rect 108120 3120 108172 3126
rect 108120 3062 108172 3068
rect 107752 3052 107804 3058
rect 107752 2994 107804 3000
rect 107658 2680 107714 2689
rect 107658 2615 107714 2624
rect 107764 2310 107792 2994
rect 108500 2650 108528 7482
rect 109328 7410 109356 12200
rect 109696 10554 109724 12200
rect 109972 11762 110000 12514
rect 110050 12200 110106 13000
rect 110418 12200 110474 13000
rect 110512 12436 110564 12442
rect 110512 12378 110564 12384
rect 109868 11756 109920 11762
rect 109868 11698 109920 11704
rect 109960 11756 110012 11762
rect 109960 11698 110012 11704
rect 109696 10526 109816 10554
rect 109684 10464 109736 10470
rect 109684 10406 109736 10412
rect 109696 10266 109724 10406
rect 109684 10260 109736 10266
rect 109684 10202 109736 10208
rect 109592 9580 109644 9586
rect 109592 9522 109644 9528
rect 109604 8838 109632 9522
rect 109592 8832 109644 8838
rect 109592 8774 109644 8780
rect 109316 7404 109368 7410
rect 109316 7346 109368 7352
rect 109500 6860 109552 6866
rect 109500 6802 109552 6808
rect 108672 6792 108724 6798
rect 108672 6734 108724 6740
rect 108946 6760 109002 6769
rect 108578 3088 108634 3097
rect 108578 3023 108634 3032
rect 108592 2990 108620 3023
rect 108580 2984 108632 2990
rect 108580 2926 108632 2932
rect 108488 2644 108540 2650
rect 108488 2586 108540 2592
rect 108580 2508 108632 2514
rect 108580 2450 108632 2456
rect 108120 2440 108172 2446
rect 108120 2382 108172 2388
rect 107844 2372 107896 2378
rect 107844 2314 107896 2320
rect 107752 2304 107804 2310
rect 107752 2246 107804 2252
rect 107016 2100 107068 2106
rect 107016 2042 107068 2048
rect 106924 1964 106976 1970
rect 106924 1906 106976 1912
rect 107752 1964 107804 1970
rect 107752 1906 107804 1912
rect 106936 1766 106964 1906
rect 106924 1760 106976 1766
rect 106924 1702 106976 1708
rect 106936 1426 106964 1702
rect 107290 1456 107346 1465
rect 106924 1420 106976 1426
rect 107764 1426 107792 1906
rect 107290 1391 107346 1400
rect 107752 1420 107804 1426
rect 106924 1362 106976 1368
rect 107016 1216 107068 1222
rect 107016 1158 107068 1164
rect 107028 1018 107056 1158
rect 107016 1012 107068 1018
rect 107016 954 107068 960
rect 106738 912 106794 921
rect 106738 847 106794 856
rect 106936 870 107056 898
rect 106936 800 106964 870
rect 106372 750 106424 756
rect 106372 672 106424 678
rect 106370 640 106372 649
rect 106424 640 106426 649
rect 106370 575 106426 584
rect 106280 196 106332 202
rect 106280 138 106332 144
rect 106554 0 106610 800
rect 106922 0 106978 800
rect 107028 785 107056 870
rect 107304 800 107332 1391
rect 107752 1362 107804 1368
rect 107856 1018 107884 2314
rect 107936 2304 107988 2310
rect 107936 2246 107988 2252
rect 107948 1562 107976 2246
rect 108132 2106 108160 2382
rect 108120 2100 108172 2106
rect 108120 2042 108172 2048
rect 108592 1902 108620 2450
rect 108684 1902 108712 6734
rect 108946 6695 109002 6704
rect 108960 6662 108988 6695
rect 108948 6656 109000 6662
rect 108948 6598 109000 6604
rect 108764 5636 108816 5642
rect 108764 5578 108816 5584
rect 108580 1896 108632 1902
rect 108580 1838 108632 1844
rect 108672 1896 108724 1902
rect 108672 1838 108724 1844
rect 107936 1556 107988 1562
rect 107936 1498 107988 1504
rect 107844 1012 107896 1018
rect 107844 954 107896 960
rect 107672 870 107792 898
rect 107672 800 107700 870
rect 107014 776 107070 785
rect 107014 711 107070 720
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 107764 66 107792 870
rect 108040 870 108160 898
rect 107936 808 107988 814
rect 108040 800 108068 870
rect 107936 750 107988 756
rect 107948 270 107976 750
rect 107936 264 107988 270
rect 107936 206 107988 212
rect 107752 60 107804 66
rect 107752 2 107804 8
rect 108026 0 108082 800
rect 108132 270 108160 870
rect 108408 836 108528 864
rect 108408 800 108436 836
rect 108120 264 108172 270
rect 108120 206 108172 212
rect 108394 0 108450 800
rect 108500 649 108528 836
rect 108776 800 108804 5578
rect 109052 4146 109448 4162
rect 109040 4140 109448 4146
rect 109092 4134 109448 4140
rect 109040 4082 109092 4088
rect 109316 4072 109368 4078
rect 109314 4040 109316 4049
rect 109368 4040 109370 4049
rect 109224 4004 109276 4010
rect 109314 3975 109370 3984
rect 109224 3946 109276 3952
rect 108856 3936 108908 3942
rect 108948 3936 109000 3942
rect 108856 3878 108908 3884
rect 108946 3904 108948 3913
rect 109000 3904 109002 3913
rect 108868 3754 108896 3878
rect 108946 3839 109002 3848
rect 108868 3726 108988 3754
rect 108960 3670 108988 3726
rect 108948 3664 109000 3670
rect 108948 3606 109000 3612
rect 109236 3534 109264 3946
rect 109420 3534 109448 4134
rect 109224 3528 109276 3534
rect 109224 3470 109276 3476
rect 109408 3528 109460 3534
rect 109408 3470 109460 3476
rect 108856 3460 108908 3466
rect 108856 3402 108908 3408
rect 108948 3460 109000 3466
rect 108948 3402 109000 3408
rect 108868 3126 108896 3402
rect 108960 3194 108988 3402
rect 108948 3188 109000 3194
rect 108948 3130 109000 3136
rect 109040 3188 109092 3194
rect 109040 3130 109092 3136
rect 108856 3120 108908 3126
rect 109052 3097 109080 3130
rect 108856 3062 108908 3068
rect 109038 3088 109094 3097
rect 109038 3023 109094 3032
rect 109408 3052 109460 3058
rect 109408 2994 109460 3000
rect 109132 2984 109184 2990
rect 108854 2952 108910 2961
rect 108854 2887 108856 2896
rect 108908 2887 108910 2896
rect 109130 2952 109132 2961
rect 109420 2961 109448 2994
rect 109184 2952 109186 2961
rect 109130 2887 109186 2896
rect 109406 2952 109462 2961
rect 109406 2887 109462 2896
rect 108856 2858 108908 2864
rect 109512 2650 109540 6802
rect 109604 4690 109632 8774
rect 109788 8294 109816 10526
rect 109880 10010 109908 11698
rect 109972 11558 110000 11698
rect 109960 11552 110012 11558
rect 109960 11494 110012 11500
rect 110064 10690 110092 12200
rect 110064 10662 110184 10690
rect 110052 10600 110104 10606
rect 110052 10542 110104 10548
rect 110064 10130 110092 10542
rect 110156 10169 110184 10662
rect 110142 10160 110198 10169
rect 110052 10124 110104 10130
rect 110142 10095 110198 10104
rect 110052 10066 110104 10072
rect 109880 9994 110092 10010
rect 109880 9988 110104 9994
rect 109880 9982 110052 9988
rect 110052 9930 110104 9936
rect 109776 8288 109828 8294
rect 109776 8230 109828 8236
rect 110432 7041 110460 12200
rect 110524 11150 110552 12378
rect 110786 12200 110842 13000
rect 111154 12200 111210 13000
rect 111522 12200 111578 13000
rect 111890 12200 111946 13000
rect 112258 12200 112314 13000
rect 112626 12200 112682 13000
rect 112994 12200 113050 13000
rect 113362 12200 113418 13000
rect 113730 12200 113786 13000
rect 114098 12200 114154 13000
rect 114466 12200 114522 13000
rect 114834 12200 114890 13000
rect 115202 12200 115258 13000
rect 115570 12200 115626 13000
rect 115938 12200 115994 13000
rect 116306 12200 116362 13000
rect 116674 12200 116730 13000
rect 117042 12200 117098 13000
rect 117410 12200 117466 13000
rect 117778 12200 117834 13000
rect 118146 12200 118202 13000
rect 118514 12200 118570 13000
rect 118882 12200 118938 13000
rect 119250 12200 119306 13000
rect 119618 12200 119674 13000
rect 119986 12200 120042 13000
rect 120354 12200 120410 13000
rect 120722 12200 120778 13000
rect 121090 12200 121146 13000
rect 121368 12504 121420 12510
rect 121368 12446 121420 12452
rect 121276 12300 121328 12306
rect 121276 12242 121328 12248
rect 110512 11144 110564 11150
rect 110512 11086 110564 11092
rect 110800 11014 110828 12200
rect 110880 11552 110932 11558
rect 111168 11506 111196 12200
rect 111536 12170 111564 12200
rect 111524 12164 111576 12170
rect 111524 12106 111576 12112
rect 111708 11688 111760 11694
rect 111708 11630 111760 11636
rect 110880 11494 110932 11500
rect 110892 11218 110920 11494
rect 111076 11478 111196 11506
rect 111248 11552 111300 11558
rect 111248 11494 111300 11500
rect 110880 11212 110932 11218
rect 110880 11154 110932 11160
rect 110972 11076 111024 11082
rect 110972 11018 111024 11024
rect 110788 11008 110840 11014
rect 110788 10950 110840 10956
rect 110880 11008 110932 11014
rect 110880 10950 110932 10956
rect 110892 10742 110920 10950
rect 110880 10736 110932 10742
rect 110880 10678 110932 10684
rect 110984 10538 111012 11018
rect 111076 10810 111104 11478
rect 111260 11218 111288 11494
rect 111248 11212 111300 11218
rect 111248 11154 111300 11160
rect 111064 10804 111116 10810
rect 111064 10746 111116 10752
rect 110972 10532 111024 10538
rect 110972 10474 111024 10480
rect 111156 10464 111208 10470
rect 111156 10406 111208 10412
rect 110972 10260 111024 10266
rect 110972 10202 111024 10208
rect 110418 7032 110474 7041
rect 110418 6967 110474 6976
rect 110880 6928 110932 6934
rect 110880 6870 110932 6876
rect 109776 5296 109828 5302
rect 109776 5238 109828 5244
rect 109592 4684 109644 4690
rect 109592 4626 109644 4632
rect 109788 3058 109816 5238
rect 110236 5228 110288 5234
rect 110236 5170 110288 5176
rect 110248 4486 110276 5170
rect 110328 5160 110380 5166
rect 110328 5102 110380 5108
rect 110340 4622 110368 5102
rect 110420 5092 110472 5098
rect 110420 5034 110472 5040
rect 110328 4616 110380 4622
rect 110328 4558 110380 4564
rect 110236 4480 110288 4486
rect 110236 4422 110288 4428
rect 109868 3392 109920 3398
rect 109868 3334 109920 3340
rect 109592 3052 109644 3058
rect 109592 2994 109644 3000
rect 109776 3052 109828 3058
rect 109776 2994 109828 3000
rect 109604 2650 109632 2994
rect 109500 2644 109552 2650
rect 109500 2586 109552 2592
rect 109592 2644 109644 2650
rect 109592 2586 109644 2592
rect 109592 2304 109644 2310
rect 109592 2246 109644 2252
rect 109604 1970 109632 2246
rect 109040 1964 109092 1970
rect 109040 1906 109092 1912
rect 109592 1964 109644 1970
rect 109592 1906 109644 1912
rect 109052 1358 109080 1906
rect 109776 1896 109828 1902
rect 109776 1838 109828 1844
rect 109236 1550 109632 1578
rect 109236 1426 109264 1550
rect 109224 1420 109276 1426
rect 109224 1362 109276 1368
rect 109040 1352 109092 1358
rect 109038 1320 109040 1329
rect 109092 1320 109094 1329
rect 109038 1255 109094 1264
rect 109224 1284 109276 1290
rect 109224 1226 109276 1232
rect 109408 1284 109460 1290
rect 109408 1226 109460 1232
rect 109040 1216 109092 1222
rect 109038 1184 109040 1193
rect 109092 1184 109094 1193
rect 109038 1119 109094 1128
rect 109236 950 109264 1226
rect 109224 944 109276 950
rect 109038 912 109094 921
rect 109224 886 109276 892
rect 109094 856 109172 864
rect 109038 847 109172 856
rect 109052 836 109172 847
rect 109144 800 109172 836
rect 109420 814 109448 1226
rect 109604 898 109632 1550
rect 109788 1358 109816 1838
rect 109776 1352 109828 1358
rect 109776 1294 109828 1300
rect 109684 1216 109736 1222
rect 109682 1184 109684 1193
rect 109736 1184 109738 1193
rect 109682 1119 109738 1128
rect 109512 870 109632 898
rect 109408 808 109460 814
rect 108486 640 108542 649
rect 108486 575 108542 584
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109512 800 109540 870
rect 109880 800 109908 3334
rect 110248 800 110276 4422
rect 110328 2916 110380 2922
rect 110328 2858 110380 2864
rect 110340 2650 110368 2858
rect 110432 2650 110460 5034
rect 110788 4752 110840 4758
rect 110788 4694 110840 4700
rect 110696 2848 110748 2854
rect 110696 2790 110748 2796
rect 110328 2644 110380 2650
rect 110328 2586 110380 2592
rect 110420 2644 110472 2650
rect 110420 2586 110472 2592
rect 110708 1902 110736 2790
rect 110800 2650 110828 4694
rect 110892 2854 110920 6870
rect 110984 5574 111012 10202
rect 111168 9654 111196 10406
rect 111260 10130 111288 11154
rect 111340 10668 111392 10674
rect 111340 10610 111392 10616
rect 111352 10538 111380 10610
rect 111340 10532 111392 10538
rect 111340 10474 111392 10480
rect 111352 10266 111380 10474
rect 111720 10470 111748 11630
rect 111904 11014 111932 12200
rect 112272 11830 112300 12200
rect 112260 11824 112312 11830
rect 112260 11766 112312 11772
rect 111892 11008 111944 11014
rect 111892 10950 111944 10956
rect 112640 10674 112668 12200
rect 113008 12152 113036 12200
rect 113376 12170 113404 12200
rect 112916 12124 113036 12152
rect 113364 12164 113416 12170
rect 112628 10668 112680 10674
rect 112628 10610 112680 10616
rect 112916 10606 112944 12124
rect 113364 12106 113416 12112
rect 113062 11996 113358 12016
rect 113118 11994 113142 11996
rect 113198 11994 113222 11996
rect 113278 11994 113302 11996
rect 113140 11942 113142 11994
rect 113204 11942 113216 11994
rect 113278 11942 113280 11994
rect 113118 11940 113142 11942
rect 113198 11940 113222 11942
rect 113278 11940 113302 11942
rect 113062 11920 113358 11940
rect 112996 11756 113048 11762
rect 112996 11698 113048 11704
rect 113008 11218 113036 11698
rect 112996 11212 113048 11218
rect 112996 11154 113048 11160
rect 113744 11082 113772 12200
rect 114112 11626 114140 12200
rect 114100 11620 114152 11626
rect 114100 11562 114152 11568
rect 114480 11286 114508 12200
rect 114652 11688 114704 11694
rect 114652 11630 114704 11636
rect 114468 11280 114520 11286
rect 114468 11222 114520 11228
rect 114664 11082 114692 11630
rect 113732 11076 113784 11082
rect 113732 11018 113784 11024
rect 114652 11076 114704 11082
rect 114652 11018 114704 11024
rect 114560 11008 114612 11014
rect 114560 10950 114612 10956
rect 113062 10908 113358 10928
rect 113118 10906 113142 10908
rect 113198 10906 113222 10908
rect 113278 10906 113302 10908
rect 113140 10854 113142 10906
rect 113204 10854 113216 10906
rect 113278 10854 113280 10906
rect 113118 10852 113142 10854
rect 113198 10852 113222 10854
rect 113278 10852 113302 10854
rect 113062 10832 113358 10852
rect 112904 10600 112956 10606
rect 113456 10600 113508 10606
rect 112904 10542 112956 10548
rect 112994 10568 113050 10577
rect 113456 10542 113508 10548
rect 112994 10503 113050 10512
rect 113008 10470 113036 10503
rect 111708 10464 111760 10470
rect 111708 10406 111760 10412
rect 112904 10464 112956 10470
rect 112904 10406 112956 10412
rect 112996 10464 113048 10470
rect 112996 10406 113048 10412
rect 111340 10260 111392 10266
rect 111340 10202 111392 10208
rect 111248 10124 111300 10130
rect 111248 10066 111300 10072
rect 112536 10124 112588 10130
rect 112536 10066 112588 10072
rect 112260 10056 112312 10062
rect 112260 9998 112312 10004
rect 111156 9648 111208 9654
rect 111156 9590 111208 9596
rect 112272 9042 112300 9998
rect 112260 9036 112312 9042
rect 112260 8978 112312 8984
rect 112260 8288 112312 8294
rect 112260 8230 112312 8236
rect 112272 7954 112300 8230
rect 112260 7948 112312 7954
rect 112260 7890 112312 7896
rect 112272 6866 112300 7890
rect 112260 6860 112312 6866
rect 112260 6802 112312 6808
rect 110972 5568 111024 5574
rect 110972 5510 111024 5516
rect 111616 4004 111668 4010
rect 111616 3946 111668 3952
rect 111524 3052 111576 3058
rect 111524 2994 111576 3000
rect 111062 2952 111118 2961
rect 111062 2887 111118 2896
rect 111432 2916 111484 2922
rect 111076 2854 111104 2887
rect 111432 2858 111484 2864
rect 110880 2848 110932 2854
rect 110880 2790 110932 2796
rect 111064 2848 111116 2854
rect 111064 2790 111116 2796
rect 110788 2644 110840 2650
rect 110788 2586 110840 2592
rect 111248 2304 111300 2310
rect 111248 2246 111300 2252
rect 111064 1964 111116 1970
rect 111064 1906 111116 1912
rect 110696 1896 110748 1902
rect 110696 1838 110748 1844
rect 110604 1760 110656 1766
rect 110604 1702 110656 1708
rect 110616 800 110644 1702
rect 110972 1556 111024 1562
rect 110972 1498 111024 1504
rect 110788 1420 110840 1426
rect 110788 1362 110840 1368
rect 110800 950 110828 1362
rect 110788 944 110840 950
rect 110788 886 110840 892
rect 110984 800 111012 1498
rect 111076 1057 111104 1906
rect 111260 1902 111288 2246
rect 111340 1964 111392 1970
rect 111340 1906 111392 1912
rect 111248 1896 111300 1902
rect 111248 1838 111300 1844
rect 111248 1352 111300 1358
rect 111248 1294 111300 1300
rect 111156 1216 111208 1222
rect 111156 1158 111208 1164
rect 111062 1048 111118 1057
rect 111062 983 111118 992
rect 111168 882 111196 1158
rect 111156 876 111208 882
rect 111156 818 111208 824
rect 109408 750 109460 756
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111260 746 111288 1294
rect 111352 1290 111380 1906
rect 111340 1284 111392 1290
rect 111340 1226 111392 1232
rect 111338 1048 111394 1057
rect 111338 983 111394 992
rect 111352 800 111380 983
rect 111444 898 111472 2858
rect 111536 2650 111564 2994
rect 111628 2922 111656 3946
rect 111616 2916 111668 2922
rect 111616 2858 111668 2864
rect 111524 2644 111576 2650
rect 111524 2586 111576 2592
rect 111524 2440 111576 2446
rect 111576 2388 111840 2394
rect 111524 2382 111840 2388
rect 111536 2366 111840 2382
rect 111616 1760 111668 1766
rect 111616 1702 111668 1708
rect 111628 1358 111656 1702
rect 111812 1426 111840 2366
rect 112260 2304 112312 2310
rect 112260 2246 112312 2252
rect 112168 1964 112220 1970
rect 112168 1906 112220 1912
rect 112076 1896 112128 1902
rect 112076 1838 112128 1844
rect 111800 1420 111852 1426
rect 111800 1362 111852 1368
rect 111616 1352 111668 1358
rect 111616 1294 111668 1300
rect 111444 870 111748 898
rect 111720 800 111748 870
rect 112088 800 112116 1838
rect 112180 1601 112208 1906
rect 112272 1902 112300 2246
rect 112260 1896 112312 1902
rect 112260 1838 112312 1844
rect 112260 1760 112312 1766
rect 112260 1702 112312 1708
rect 112166 1592 112222 1601
rect 112166 1527 112222 1536
rect 112272 1358 112300 1702
rect 112548 1562 112576 10066
rect 112916 10062 112944 10406
rect 112904 10056 112956 10062
rect 112904 9998 112956 10004
rect 113062 9820 113358 9840
rect 113118 9818 113142 9820
rect 113198 9818 113222 9820
rect 113278 9818 113302 9820
rect 113140 9766 113142 9818
rect 113204 9766 113216 9818
rect 113278 9766 113280 9818
rect 113118 9764 113142 9766
rect 113198 9764 113222 9766
rect 113278 9764 113302 9766
rect 113062 9744 113358 9764
rect 113468 9654 113496 10542
rect 114572 9926 114600 10950
rect 114848 10606 114876 12200
rect 115018 11656 115074 11665
rect 115018 11591 115074 11600
rect 115032 11218 115060 11591
rect 115216 11218 115244 12200
rect 115584 11762 115612 12200
rect 115572 11756 115624 11762
rect 115572 11698 115624 11704
rect 115020 11212 115072 11218
rect 115020 11154 115072 11160
rect 115204 11212 115256 11218
rect 115204 11154 115256 11160
rect 115572 11144 115624 11150
rect 115572 11086 115624 11092
rect 114836 10600 114888 10606
rect 114836 10542 114888 10548
rect 114652 10532 114704 10538
rect 114652 10474 114704 10480
rect 114664 10062 114692 10474
rect 115584 10130 115612 11086
rect 115848 10600 115900 10606
rect 115848 10542 115900 10548
rect 115572 10124 115624 10130
rect 115572 10066 115624 10072
rect 114652 10056 114704 10062
rect 114652 9998 114704 10004
rect 115860 9926 115888 10542
rect 115952 10062 115980 12200
rect 116320 11694 116348 12200
rect 116492 11756 116544 11762
rect 116492 11698 116544 11704
rect 116308 11688 116360 11694
rect 116308 11630 116360 11636
rect 116504 11558 116532 11698
rect 116492 11552 116544 11558
rect 116490 11520 116492 11529
rect 116544 11520 116546 11529
rect 116490 11455 116546 11464
rect 116584 11076 116636 11082
rect 116584 11018 116636 11024
rect 116596 10130 116624 11018
rect 116688 10606 116716 12200
rect 116950 11384 117006 11393
rect 116950 11319 117006 11328
rect 116676 10600 116728 10606
rect 116676 10542 116728 10548
rect 116964 10266 116992 11319
rect 117056 10713 117084 12200
rect 117042 10704 117098 10713
rect 117042 10639 117098 10648
rect 117136 10668 117188 10674
rect 117136 10610 117188 10616
rect 117148 10266 117176 10610
rect 116952 10260 117004 10266
rect 116952 10202 117004 10208
rect 117136 10260 117188 10266
rect 117136 10202 117188 10208
rect 116584 10124 116636 10130
rect 116584 10066 116636 10072
rect 115940 10056 115992 10062
rect 115940 9998 115992 10004
rect 114560 9920 114612 9926
rect 114560 9862 114612 9868
rect 115848 9920 115900 9926
rect 115848 9862 115900 9868
rect 113456 9648 113508 9654
rect 113548 9648 113600 9654
rect 113456 9590 113508 9596
rect 113546 9616 113548 9625
rect 113600 9616 113602 9625
rect 113546 9551 113602 9560
rect 115204 9580 115256 9586
rect 115204 9522 115256 9528
rect 113916 9512 113968 9518
rect 113916 9454 113968 9460
rect 113928 9042 113956 9454
rect 113916 9036 113968 9042
rect 113916 8978 113968 8984
rect 115216 8786 115244 9522
rect 115572 9512 115624 9518
rect 115572 9454 115624 9460
rect 115296 9444 115348 9450
rect 115296 9386 115348 9392
rect 115308 8974 115336 9386
rect 115584 9042 115612 9454
rect 115662 9208 115718 9217
rect 115662 9143 115718 9152
rect 115676 9042 115704 9143
rect 115572 9036 115624 9042
rect 115572 8978 115624 8984
rect 115664 9036 115716 9042
rect 115664 8978 115716 8984
rect 115296 8968 115348 8974
rect 115296 8910 115348 8916
rect 115296 8832 115348 8838
rect 115216 8780 115296 8786
rect 115216 8774 115348 8780
rect 115216 8758 115336 8774
rect 113062 8732 113358 8752
rect 113118 8730 113142 8732
rect 113198 8730 113222 8732
rect 113278 8730 113302 8732
rect 113140 8678 113142 8730
rect 113204 8678 113216 8730
rect 113278 8678 113280 8730
rect 113118 8676 113142 8678
rect 113198 8676 113222 8678
rect 113278 8676 113302 8678
rect 113062 8656 113358 8676
rect 113456 8424 113508 8430
rect 113456 8366 113508 8372
rect 112902 7712 112958 7721
rect 112902 7647 112958 7656
rect 112916 7528 112944 7647
rect 113062 7644 113358 7664
rect 113118 7642 113142 7644
rect 113198 7642 113222 7644
rect 113278 7642 113302 7644
rect 113140 7590 113142 7642
rect 113204 7590 113216 7642
rect 113278 7590 113280 7642
rect 113118 7588 113142 7590
rect 113198 7588 113222 7590
rect 113278 7588 113302 7590
rect 113062 7568 113358 7588
rect 112916 7500 113128 7528
rect 113100 7449 113128 7500
rect 113086 7440 113142 7449
rect 113086 7375 113142 7384
rect 113468 7342 113496 8366
rect 114100 7948 114152 7954
rect 114100 7890 114152 7896
rect 114112 7410 114140 7890
rect 114558 7576 114614 7585
rect 114558 7511 114614 7520
rect 114374 7440 114430 7449
rect 114100 7404 114152 7410
rect 114572 7426 114600 7511
rect 114430 7398 114600 7426
rect 114374 7375 114430 7384
rect 114100 7346 114152 7352
rect 113272 7336 113324 7342
rect 113272 7278 113324 7284
rect 113456 7336 113508 7342
rect 113456 7278 113508 7284
rect 113284 6882 113312 7278
rect 113468 7002 113496 7278
rect 113456 6996 113508 7002
rect 113456 6938 113508 6944
rect 113548 6996 113600 7002
rect 113548 6938 113600 6944
rect 113560 6882 113588 6938
rect 113284 6854 113588 6882
rect 114664 6866 114876 6882
rect 114664 6860 114888 6866
rect 114664 6854 114836 6860
rect 114664 6798 114692 6854
rect 114836 6802 114888 6808
rect 114652 6792 114704 6798
rect 113638 6760 113694 6769
rect 114652 6734 114704 6740
rect 113638 6695 113640 6704
rect 113692 6695 113694 6704
rect 113640 6666 113692 6672
rect 113456 6656 113508 6662
rect 113456 6598 113508 6604
rect 113062 6556 113358 6576
rect 113118 6554 113142 6556
rect 113198 6554 113222 6556
rect 113278 6554 113302 6556
rect 113140 6502 113142 6554
rect 113204 6502 113216 6554
rect 113278 6502 113280 6554
rect 113118 6500 113142 6502
rect 113198 6500 113222 6502
rect 113278 6500 113302 6502
rect 113062 6480 113358 6500
rect 113468 6254 113496 6598
rect 113456 6248 113508 6254
rect 113456 6190 113508 6196
rect 114836 6180 114888 6186
rect 114836 6122 114888 6128
rect 112720 5772 112772 5778
rect 112720 5714 112772 5720
rect 112732 2650 112760 5714
rect 114848 5574 114876 6122
rect 114652 5568 114704 5574
rect 114652 5510 114704 5516
rect 114836 5568 114888 5574
rect 114836 5510 114888 5516
rect 113062 5468 113358 5488
rect 113118 5466 113142 5468
rect 113198 5466 113222 5468
rect 113278 5466 113302 5468
rect 113140 5414 113142 5466
rect 113204 5414 113216 5466
rect 113278 5414 113280 5466
rect 113118 5412 113142 5414
rect 113198 5412 113222 5414
rect 113278 5412 113302 5414
rect 113062 5392 113358 5412
rect 112904 5296 112956 5302
rect 112904 5238 112956 5244
rect 112812 3052 112864 3058
rect 112812 2994 112864 3000
rect 112720 2644 112772 2650
rect 112720 2586 112772 2592
rect 112626 1728 112682 1737
rect 112626 1663 112682 1672
rect 112536 1556 112588 1562
rect 112536 1498 112588 1504
rect 112640 1426 112668 1663
rect 112444 1420 112496 1426
rect 112444 1362 112496 1368
rect 112628 1420 112680 1426
rect 112628 1362 112680 1368
rect 112260 1352 112312 1358
rect 112260 1294 112312 1300
rect 112456 800 112484 1362
rect 112824 800 112852 2994
rect 112916 1970 112944 5238
rect 113456 4548 113508 4554
rect 113456 4490 113508 4496
rect 113548 4548 113600 4554
rect 113548 4490 113600 4496
rect 113062 4380 113358 4400
rect 113118 4378 113142 4380
rect 113198 4378 113222 4380
rect 113278 4378 113302 4380
rect 113140 4326 113142 4378
rect 113204 4326 113216 4378
rect 113278 4326 113280 4378
rect 113118 4324 113142 4326
rect 113198 4324 113222 4326
rect 113278 4324 113302 4326
rect 113062 4304 113358 4324
rect 113062 3292 113358 3312
rect 113118 3290 113142 3292
rect 113198 3290 113222 3292
rect 113278 3290 113302 3292
rect 113140 3238 113142 3290
rect 113204 3238 113216 3290
rect 113278 3238 113280 3290
rect 113118 3236 113142 3238
rect 113198 3236 113222 3238
rect 113278 3236 113302 3238
rect 113062 3216 113358 3236
rect 113468 2650 113496 4490
rect 113560 4282 113588 4490
rect 113548 4276 113600 4282
rect 113548 4218 113600 4224
rect 114008 4276 114060 4282
rect 114008 4218 114060 4224
rect 113640 4140 113692 4146
rect 113640 4082 113692 4088
rect 113548 3936 113600 3942
rect 113548 3878 113600 3884
rect 113560 3738 113588 3878
rect 113652 3738 113680 4082
rect 113548 3732 113600 3738
rect 113548 3674 113600 3680
rect 113640 3732 113692 3738
rect 113640 3674 113692 3680
rect 114020 3534 114048 4218
rect 114008 3528 114060 3534
rect 114008 3470 114060 3476
rect 114560 3052 114612 3058
rect 114560 2994 114612 3000
rect 114572 2922 114600 2994
rect 114560 2916 114612 2922
rect 114560 2858 114612 2864
rect 114466 2816 114522 2825
rect 114466 2751 114522 2760
rect 113456 2644 113508 2650
rect 113456 2586 113508 2592
rect 114284 2440 114336 2446
rect 114284 2382 114336 2388
rect 114296 2310 114324 2382
rect 114480 2310 114508 2751
rect 114572 2650 114600 2858
rect 114560 2644 114612 2650
rect 114560 2586 114612 2592
rect 113916 2304 113968 2310
rect 113916 2246 113968 2252
rect 114284 2304 114336 2310
rect 114284 2246 114336 2252
rect 114468 2304 114520 2310
rect 114468 2246 114520 2252
rect 113062 2204 113358 2224
rect 113118 2202 113142 2204
rect 113198 2202 113222 2204
rect 113278 2202 113302 2204
rect 113140 2150 113142 2202
rect 113204 2150 113216 2202
rect 113278 2150 113280 2202
rect 113118 2148 113142 2150
rect 113198 2148 113222 2150
rect 113278 2148 113302 2150
rect 113062 2128 113358 2148
rect 112904 1964 112956 1970
rect 112904 1906 112956 1912
rect 113456 1896 113508 1902
rect 113456 1838 113508 1844
rect 113824 1896 113876 1902
rect 113824 1838 113876 1844
rect 113062 1116 113358 1136
rect 113118 1114 113142 1116
rect 113198 1114 113222 1116
rect 113278 1114 113302 1116
rect 113140 1062 113142 1114
rect 113204 1062 113216 1114
rect 113278 1062 113280 1114
rect 113118 1060 113142 1062
rect 113198 1060 113222 1062
rect 113278 1060 113302 1062
rect 113062 1040 113358 1060
rect 113468 898 113496 1838
rect 113836 1426 113864 1838
rect 113824 1420 113876 1426
rect 113824 1362 113876 1368
rect 113546 1320 113602 1329
rect 113546 1255 113602 1264
rect 113192 870 113496 898
rect 113192 800 113220 870
rect 113560 800 113588 1255
rect 113928 800 113956 2246
rect 114100 1284 114152 1290
rect 114100 1226 114152 1232
rect 114008 1216 114060 1222
rect 114008 1158 114060 1164
rect 114020 950 114048 1158
rect 114008 944 114060 950
rect 114008 886 114060 892
rect 111248 740 111300 746
rect 111248 682 111300 688
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113178 0 113234 800
rect 113546 0 113602 800
rect 113914 0 113970 800
rect 114112 649 114140 1226
rect 114296 800 114324 2246
rect 114466 1728 114522 1737
rect 114466 1663 114522 1672
rect 114098 640 114154 649
rect 114098 575 114154 584
rect 114282 0 114338 800
rect 114480 338 114508 1663
rect 114664 800 114692 5510
rect 115308 5098 115336 8758
rect 115860 8498 115888 9862
rect 117424 9586 117452 12200
rect 117792 11014 117820 12200
rect 117964 11552 118016 11558
rect 117964 11494 118016 11500
rect 117976 11218 118004 11494
rect 117964 11212 118016 11218
rect 117964 11154 118016 11160
rect 117780 11008 117832 11014
rect 117780 10950 117832 10956
rect 117976 10130 118004 11154
rect 117964 10124 118016 10130
rect 117964 10066 118016 10072
rect 117412 9580 117464 9586
rect 117412 9522 117464 9528
rect 118160 9353 118188 12200
rect 118332 12096 118384 12102
rect 118332 12038 118384 12044
rect 118344 11762 118372 12038
rect 118332 11756 118384 11762
rect 118332 11698 118384 11704
rect 118528 11200 118556 12200
rect 118700 12096 118752 12102
rect 118700 12038 118752 12044
rect 118712 11898 118740 12038
rect 118700 11892 118752 11898
rect 118700 11834 118752 11840
rect 118792 11892 118844 11898
rect 118792 11834 118844 11840
rect 118608 11620 118660 11626
rect 118608 11562 118660 11568
rect 118620 11354 118648 11562
rect 118804 11558 118832 11834
rect 118896 11762 118924 12200
rect 118884 11756 118936 11762
rect 118884 11698 118936 11704
rect 119264 11558 119292 12200
rect 119632 12170 119660 12200
rect 120000 12170 120028 12200
rect 119620 12164 119672 12170
rect 119620 12106 119672 12112
rect 119988 12164 120040 12170
rect 119988 12106 120040 12112
rect 120264 11688 120316 11694
rect 120264 11630 120316 11636
rect 118792 11552 118844 11558
rect 118792 11494 118844 11500
rect 119252 11552 119304 11558
rect 119252 11494 119304 11500
rect 118608 11348 118660 11354
rect 118608 11290 118660 11296
rect 118700 11212 118752 11218
rect 118528 11172 118700 11200
rect 118700 11154 118752 11160
rect 120276 11082 120304 11630
rect 120368 11098 120396 12200
rect 120264 11076 120316 11082
rect 120368 11070 120488 11098
rect 120264 11018 120316 11024
rect 119712 11008 119764 11014
rect 119712 10950 119764 10956
rect 119724 10742 119752 10950
rect 120276 10810 120304 11018
rect 120460 11014 120488 11070
rect 120448 11008 120500 11014
rect 120448 10950 120500 10956
rect 120736 10810 120764 12200
rect 121104 10826 121132 12200
rect 121288 11354 121316 12242
rect 121380 12152 121408 12446
rect 121458 12200 121514 13000
rect 121644 12640 121696 12646
rect 121644 12582 121696 12588
rect 121472 12152 121500 12200
rect 121380 12124 121500 12152
rect 121656 12152 121684 12582
rect 121826 12200 121882 13000
rect 121920 12300 121972 12306
rect 121920 12242 121972 12248
rect 121840 12152 121868 12200
rect 121656 12124 121868 12152
rect 121932 11762 121960 12242
rect 122194 12200 122250 13000
rect 122562 12200 122618 13000
rect 122930 12200 122986 13000
rect 123208 12572 123260 12578
rect 123208 12514 123260 12520
rect 122208 11830 122236 12200
rect 122196 11824 122248 11830
rect 122196 11766 122248 11772
rect 121920 11756 121972 11762
rect 121920 11698 121972 11704
rect 121736 11620 121788 11626
rect 121736 11562 121788 11568
rect 121748 11354 121776 11562
rect 121932 11354 121960 11698
rect 122576 11665 122604 12200
rect 122562 11656 122618 11665
rect 122562 11591 122618 11600
rect 122944 11393 122972 12200
rect 123220 11762 123248 12514
rect 123298 12200 123354 13000
rect 123484 12436 123536 12442
rect 123484 12378 123536 12384
rect 123116 11756 123168 11762
rect 123116 11698 123168 11704
rect 123208 11756 123260 11762
rect 123208 11698 123260 11704
rect 122930 11384 122986 11393
rect 121276 11348 121328 11354
rect 121276 11290 121328 11296
rect 121736 11348 121788 11354
rect 121736 11290 121788 11296
rect 121920 11348 121972 11354
rect 123128 11354 123156 11698
rect 122930 11319 122986 11328
rect 123116 11348 123168 11354
rect 121920 11290 121972 11296
rect 123116 11290 123168 11296
rect 122932 11212 122984 11218
rect 122932 11154 122984 11160
rect 122196 11076 122248 11082
rect 122196 11018 122248 11024
rect 120264 10804 120316 10810
rect 120264 10746 120316 10752
rect 120724 10804 120776 10810
rect 121104 10798 121224 10826
rect 120724 10746 120776 10752
rect 119620 10736 119672 10742
rect 119620 10678 119672 10684
rect 119712 10736 119764 10742
rect 119712 10678 119764 10684
rect 120538 10704 120594 10713
rect 119528 10600 119580 10606
rect 119528 10542 119580 10548
rect 119540 10266 119568 10542
rect 119632 10266 119660 10678
rect 120538 10639 120594 10648
rect 121092 10668 121144 10674
rect 120552 10606 120580 10639
rect 121092 10610 121144 10616
rect 120540 10600 120592 10606
rect 120540 10542 120592 10548
rect 119528 10260 119580 10266
rect 119528 10202 119580 10208
rect 119620 10260 119672 10266
rect 119620 10202 119672 10208
rect 120736 9994 120948 10010
rect 120736 9988 120960 9994
rect 120736 9982 120908 9988
rect 120736 9926 120764 9982
rect 120908 9930 120960 9936
rect 121104 9926 121132 10610
rect 121196 10577 121224 10798
rect 121182 10568 121238 10577
rect 121182 10503 121238 10512
rect 121184 10464 121236 10470
rect 121184 10406 121236 10412
rect 121196 10062 121224 10406
rect 122104 10260 122156 10266
rect 122104 10202 122156 10208
rect 122116 10062 122144 10202
rect 121184 10056 121236 10062
rect 121184 9998 121236 10004
rect 122104 10056 122156 10062
rect 122104 9998 122156 10004
rect 120724 9920 120776 9926
rect 120724 9862 120776 9868
rect 121092 9920 121144 9926
rect 121092 9862 121144 9868
rect 121000 9716 121052 9722
rect 121000 9658 121052 9664
rect 119252 9648 119304 9654
rect 119250 9616 119252 9625
rect 119304 9616 119306 9625
rect 119250 9551 119306 9560
rect 120448 9580 120500 9586
rect 120448 9522 120500 9528
rect 118792 9512 118844 9518
rect 118792 9454 118844 9460
rect 119896 9512 119948 9518
rect 119896 9454 119948 9460
rect 118146 9344 118202 9353
rect 118146 9279 118202 9288
rect 118804 8974 118832 9454
rect 119172 9042 119476 9058
rect 119160 9036 119488 9042
rect 119212 9030 119436 9036
rect 119160 8978 119212 8984
rect 119436 8978 119488 8984
rect 117504 8968 117556 8974
rect 117504 8910 117556 8916
rect 118792 8968 118844 8974
rect 118792 8910 118844 8916
rect 117516 8838 117544 8910
rect 118516 8900 118568 8906
rect 118516 8842 118568 8848
rect 117504 8832 117556 8838
rect 117504 8774 117556 8780
rect 115848 8492 115900 8498
rect 115848 8434 115900 8440
rect 116584 8424 116636 8430
rect 115860 8350 116532 8378
rect 116584 8366 116636 8372
rect 115860 8294 115888 8350
rect 116504 8294 116532 8350
rect 115848 8288 115900 8294
rect 115848 8230 115900 8236
rect 116492 8288 116544 8294
rect 116492 8230 116544 8236
rect 116124 7880 116176 7886
rect 116122 7848 116124 7857
rect 116176 7848 116178 7857
rect 116596 7818 116624 8366
rect 116950 7848 117006 7857
rect 116122 7783 116178 7792
rect 116216 7812 116268 7818
rect 116216 7754 116268 7760
rect 116584 7812 116636 7818
rect 116950 7783 117006 7792
rect 116584 7754 116636 7760
rect 115940 7404 115992 7410
rect 115940 7346 115992 7352
rect 115756 7336 115808 7342
rect 115756 7278 115808 7284
rect 115768 6662 115796 7278
rect 115756 6656 115808 6662
rect 115756 6598 115808 6604
rect 115768 6254 115796 6598
rect 115756 6248 115808 6254
rect 115756 6190 115808 6196
rect 115388 5228 115440 5234
rect 115388 5170 115440 5176
rect 115296 5092 115348 5098
rect 115296 5034 115348 5040
rect 115400 4486 115428 5170
rect 115388 4480 115440 4486
rect 115388 4422 115440 4428
rect 115400 4282 115428 4422
rect 115388 4276 115440 4282
rect 115388 4218 115440 4224
rect 114836 4140 114888 4146
rect 115848 4140 115900 4146
rect 114888 4100 115060 4128
rect 114836 4082 114888 4088
rect 114756 4010 114968 4026
rect 114744 4004 114980 4010
rect 114796 3998 114928 4004
rect 114744 3946 114796 3952
rect 114928 3946 114980 3952
rect 115032 3942 115060 4100
rect 115848 4082 115900 4088
rect 114836 3936 114888 3942
rect 114836 3878 114888 3884
rect 115020 3936 115072 3942
rect 115020 3878 115072 3884
rect 114848 3398 114876 3878
rect 115756 3732 115808 3738
rect 115756 3674 115808 3680
rect 115018 3632 115074 3641
rect 115018 3567 115074 3576
rect 115032 3466 115060 3567
rect 115020 3460 115072 3466
rect 115020 3402 115072 3408
rect 114836 3392 114888 3398
rect 114836 3334 114888 3340
rect 115386 2680 115442 2689
rect 115386 2615 115442 2624
rect 115112 2304 115164 2310
rect 115112 2246 115164 2252
rect 115124 1766 115152 2246
rect 115112 1760 115164 1766
rect 115112 1702 115164 1708
rect 115020 1420 115072 1426
rect 115020 1362 115072 1368
rect 114928 808 114980 814
rect 114468 332 114520 338
rect 114468 274 114520 280
rect 114650 0 114706 800
rect 115032 800 115060 1362
rect 115400 800 115428 2615
rect 115572 1964 115624 1970
rect 115572 1906 115624 1912
rect 115584 1222 115612 1906
rect 115572 1216 115624 1222
rect 115572 1158 115624 1164
rect 114928 750 114980 756
rect 114940 406 114968 750
rect 114928 400 114980 406
rect 114928 342 114980 348
rect 115018 0 115074 800
rect 115386 0 115442 800
rect 115584 678 115612 1158
rect 115768 800 115796 3674
rect 115860 3398 115888 4082
rect 115848 3392 115900 3398
rect 115848 3334 115900 3340
rect 115952 2310 115980 7346
rect 116228 5914 116256 7754
rect 116964 7478 116992 7783
rect 116952 7472 117004 7478
rect 116952 7414 117004 7420
rect 117136 7404 117188 7410
rect 117136 7346 117188 7352
rect 117148 6662 117176 7346
rect 117136 6656 117188 6662
rect 117136 6598 117188 6604
rect 116124 5908 116176 5914
rect 116124 5850 116176 5856
rect 116216 5908 116268 5914
rect 116216 5850 116268 5856
rect 116136 5624 116164 5850
rect 116136 5596 116532 5624
rect 116216 5024 116268 5030
rect 116216 4966 116268 4972
rect 116228 2854 116256 4966
rect 116124 2848 116176 2854
rect 116124 2790 116176 2796
rect 116216 2848 116268 2854
rect 116216 2790 116268 2796
rect 115940 2304 115992 2310
rect 115940 2246 115992 2252
rect 116136 800 116164 2790
rect 116216 1964 116268 1970
rect 116216 1906 116268 1912
rect 116228 1426 116256 1906
rect 116216 1420 116268 1426
rect 116216 1362 116268 1368
rect 116216 1216 116268 1222
rect 116216 1158 116268 1164
rect 116308 1216 116360 1222
rect 116308 1158 116360 1164
rect 116228 950 116256 1158
rect 116216 944 116268 950
rect 116216 886 116268 892
rect 116320 882 116348 1158
rect 116308 876 116360 882
rect 116308 818 116360 824
rect 116504 800 116532 5596
rect 116860 5568 116912 5574
rect 116860 5510 116912 5516
rect 116768 2440 116820 2446
rect 116768 2382 116820 2388
rect 116780 2310 116808 2382
rect 116768 2304 116820 2310
rect 116768 2246 116820 2252
rect 116780 1902 116808 2246
rect 116768 1896 116820 1902
rect 116768 1838 116820 1844
rect 116872 800 116900 5510
rect 117148 5234 117176 6598
rect 117136 5228 117188 5234
rect 117136 5170 117188 5176
rect 117044 4684 117096 4690
rect 117044 4626 117096 4632
rect 117056 4214 117084 4626
rect 117136 4548 117188 4554
rect 117136 4490 117188 4496
rect 117044 4208 117096 4214
rect 117044 4150 117096 4156
rect 117148 1034 117176 4490
rect 117516 3738 117544 8774
rect 118528 8498 118556 8842
rect 119908 8634 119936 9454
rect 120460 8838 120488 9522
rect 121012 9518 121040 9658
rect 122208 9586 122236 11018
rect 122944 10470 122972 11154
rect 123116 10668 123168 10674
rect 123116 10610 123168 10616
rect 122748 10464 122800 10470
rect 122748 10406 122800 10412
rect 122932 10464 122984 10470
rect 122932 10406 122984 10412
rect 122760 10062 122788 10406
rect 123128 10266 123156 10610
rect 123116 10260 123168 10266
rect 123116 10202 123168 10208
rect 122748 10056 122800 10062
rect 122748 9998 122800 10004
rect 122760 9722 122788 9998
rect 122748 9716 122800 9722
rect 122748 9658 122800 9664
rect 122470 9616 122526 9625
rect 121460 9580 121512 9586
rect 121460 9522 121512 9528
rect 122196 9580 122248 9586
rect 122470 9551 122526 9560
rect 122196 9522 122248 9528
rect 121000 9512 121052 9518
rect 121000 9454 121052 9460
rect 120724 9444 120776 9450
rect 120724 9386 120776 9392
rect 120736 9110 120764 9386
rect 121276 9376 121328 9382
rect 121276 9318 121328 9324
rect 120724 9104 120776 9110
rect 120724 9046 120776 9052
rect 121288 8974 121316 9318
rect 121472 9178 121500 9522
rect 122484 9518 122512 9551
rect 122472 9512 122524 9518
rect 122472 9454 122524 9460
rect 123312 9450 123340 12200
rect 123496 12152 123524 12378
rect 123666 12200 123722 13000
rect 124034 12200 124090 13000
rect 124402 12200 124458 13000
rect 124770 12200 124826 13000
rect 125138 12200 125194 13000
rect 125506 12200 125562 13000
rect 125600 12232 125652 12238
rect 123680 12152 123708 12200
rect 123496 12124 123708 12152
rect 124048 11898 124076 12200
rect 124036 11892 124088 11898
rect 124036 11834 124088 11840
rect 124312 11756 124364 11762
rect 124312 11698 124364 11704
rect 124324 11354 124352 11698
rect 124416 11626 124444 12200
rect 124784 11830 124812 12200
rect 124772 11824 124824 11830
rect 124772 11766 124824 11772
rect 125152 11762 125180 12200
rect 125140 11756 125192 11762
rect 125140 11698 125192 11704
rect 124404 11620 124456 11626
rect 124404 11562 124456 11568
rect 124680 11552 124732 11558
rect 124680 11494 124732 11500
rect 124770 11520 124826 11529
rect 124312 11348 124364 11354
rect 124312 11290 124364 11296
rect 123392 11280 123444 11286
rect 123392 11222 123444 11228
rect 123404 10606 123432 11222
rect 124692 11150 124720 11494
rect 124770 11455 124826 11464
rect 124680 11144 124732 11150
rect 124680 11086 124732 11092
rect 123760 10804 123812 10810
rect 123760 10746 123812 10752
rect 123392 10600 123444 10606
rect 123392 10542 123444 10548
rect 123772 10470 123800 10746
rect 123760 10464 123812 10470
rect 123760 10406 123812 10412
rect 123576 9580 123628 9586
rect 123576 9522 123628 9528
rect 123300 9444 123352 9450
rect 123300 9386 123352 9392
rect 121460 9172 121512 9178
rect 121460 9114 121512 9120
rect 121276 8968 121328 8974
rect 121276 8910 121328 8916
rect 121184 8900 121236 8906
rect 121184 8842 121236 8848
rect 120448 8832 120500 8838
rect 120448 8774 120500 8780
rect 121000 8832 121052 8838
rect 121000 8774 121052 8780
rect 119896 8628 119948 8634
rect 119896 8570 119948 8576
rect 120908 8560 120960 8566
rect 120908 8502 120960 8508
rect 118516 8492 118568 8498
rect 118516 8434 118568 8440
rect 120920 8430 120948 8502
rect 121012 8430 121040 8774
rect 121196 8498 121224 8842
rect 121288 8634 121316 8910
rect 123588 8838 123616 9522
rect 124588 9512 124640 9518
rect 124588 9454 124640 9460
rect 124600 9178 124628 9454
rect 124588 9172 124640 9178
rect 124588 9114 124640 9120
rect 124600 9042 124628 9114
rect 124588 9036 124640 9042
rect 124588 8978 124640 8984
rect 123576 8832 123628 8838
rect 123576 8774 123628 8780
rect 124692 8634 124720 11086
rect 124784 10810 124812 11455
rect 125520 11286 125548 12200
rect 125874 12200 125930 13000
rect 126242 12200 126298 13000
rect 126610 12200 126666 13000
rect 126888 12300 126940 12306
rect 126888 12242 126940 12248
rect 125600 12174 125652 12180
rect 125612 11898 125640 12174
rect 125600 11892 125652 11898
rect 125600 11834 125652 11840
rect 125508 11280 125560 11286
rect 125508 11222 125560 11228
rect 125324 11212 125376 11218
rect 125324 11154 125376 11160
rect 124772 10804 124824 10810
rect 124772 10746 124824 10752
rect 124956 10668 125008 10674
rect 124956 10610 125008 10616
rect 124968 10266 124996 10610
rect 124956 10260 125008 10266
rect 124956 10202 125008 10208
rect 125336 9654 125364 11154
rect 125600 10600 125652 10606
rect 125888 10588 125916 12200
rect 126152 11552 126204 11558
rect 126152 11494 126204 11500
rect 126164 11286 126192 11494
rect 126152 11280 126204 11286
rect 126152 11222 126204 11228
rect 126256 11150 126284 12200
rect 126244 11144 126296 11150
rect 126244 11086 126296 11092
rect 125652 10560 125916 10588
rect 126244 10600 126296 10606
rect 125600 10542 125652 10548
rect 126244 10542 126296 10548
rect 126256 9926 126284 10542
rect 126624 10266 126652 12200
rect 126612 10260 126664 10266
rect 126612 10202 126664 10208
rect 126244 9920 126296 9926
rect 126244 9862 126296 9868
rect 125324 9648 125376 9654
rect 125324 9590 125376 9596
rect 124770 9344 124826 9353
rect 124770 9279 124826 9288
rect 124784 9110 124812 9279
rect 124772 9104 124824 9110
rect 124772 9046 124824 9052
rect 125784 9036 125836 9042
rect 125784 8978 125836 8984
rect 125324 8832 125376 8838
rect 125692 8832 125744 8838
rect 125376 8780 125640 8786
rect 125324 8774 125640 8780
rect 125692 8774 125744 8780
rect 125336 8758 125640 8774
rect 121276 8628 121328 8634
rect 121276 8570 121328 8576
rect 124680 8628 124732 8634
rect 124680 8570 124732 8576
rect 121184 8492 121236 8498
rect 121184 8434 121236 8440
rect 121368 8492 121420 8498
rect 121368 8434 121420 8440
rect 119896 8424 119948 8430
rect 119896 8366 119948 8372
rect 120908 8424 120960 8430
rect 120908 8366 120960 8372
rect 121000 8424 121052 8430
rect 121000 8366 121052 8372
rect 119908 7954 119936 8366
rect 119896 7948 119948 7954
rect 119896 7890 119948 7896
rect 121380 7818 121408 8434
rect 124956 8084 125008 8090
rect 124956 8026 125008 8032
rect 120816 7812 120868 7818
rect 120816 7754 120868 7760
rect 121368 7812 121420 7818
rect 121368 7754 121420 7760
rect 122472 7812 122524 7818
rect 122472 7754 122524 7760
rect 118792 7744 118844 7750
rect 118792 7686 118844 7692
rect 118976 7744 119028 7750
rect 118976 7686 119028 7692
rect 117780 6860 117832 6866
rect 117780 6802 117832 6808
rect 117688 6112 117740 6118
rect 117688 6054 117740 6060
rect 117596 3936 117648 3942
rect 117596 3878 117648 3884
rect 117504 3732 117556 3738
rect 117504 3674 117556 3680
rect 117228 3052 117280 3058
rect 117228 2994 117280 3000
rect 117240 2650 117268 2994
rect 117228 2644 117280 2650
rect 117228 2586 117280 2592
rect 117412 2304 117464 2310
rect 117412 2246 117464 2252
rect 117424 1562 117452 2246
rect 117412 1556 117464 1562
rect 117412 1498 117464 1504
rect 117148 1006 117268 1034
rect 117240 800 117268 1006
rect 117608 800 117636 3878
rect 117700 2650 117728 6054
rect 117688 2644 117740 2650
rect 117688 2586 117740 2592
rect 117792 2038 117820 6802
rect 118608 6792 118660 6798
rect 118606 6760 118608 6769
rect 118660 6760 118662 6769
rect 118606 6695 118662 6704
rect 118332 5772 118384 5778
rect 118332 5714 118384 5720
rect 117964 3392 118016 3398
rect 117964 3334 118016 3340
rect 117780 2032 117832 2038
rect 117780 1974 117832 1980
rect 117872 2032 117924 2038
rect 117872 1974 117924 1980
rect 117688 1964 117740 1970
rect 117688 1906 117740 1912
rect 117700 1562 117728 1906
rect 117884 1850 117912 1974
rect 117792 1834 117912 1850
rect 117780 1828 117912 1834
rect 117832 1822 117912 1828
rect 117780 1770 117832 1776
rect 117688 1556 117740 1562
rect 117688 1498 117740 1504
rect 117976 800 118004 3334
rect 118056 2576 118108 2582
rect 118054 2544 118056 2553
rect 118108 2544 118110 2553
rect 118054 2479 118110 2488
rect 118240 2508 118292 2514
rect 118240 2450 118292 2456
rect 118252 1766 118280 2450
rect 118240 1760 118292 1766
rect 118240 1702 118292 1708
rect 118056 1556 118108 1562
rect 118056 1498 118108 1504
rect 118068 1057 118096 1498
rect 118148 1284 118200 1290
rect 118148 1226 118200 1232
rect 118054 1048 118110 1057
rect 118054 983 118110 992
rect 118160 882 118188 1226
rect 118148 876 118200 882
rect 118148 818 118200 824
rect 118344 800 118372 5714
rect 118700 2916 118752 2922
rect 118700 2858 118752 2864
rect 118516 2644 118568 2650
rect 118516 2586 118568 2592
rect 118528 2310 118556 2586
rect 118516 2304 118568 2310
rect 118516 2246 118568 2252
rect 118608 2304 118660 2310
rect 118608 2246 118660 2252
rect 118620 1970 118648 2246
rect 118608 1964 118660 1970
rect 118608 1906 118660 1912
rect 118424 1760 118476 1766
rect 118424 1702 118476 1708
rect 118436 1426 118464 1702
rect 118424 1420 118476 1426
rect 118424 1362 118476 1368
rect 118424 808 118476 814
rect 115572 672 115624 678
rect 115572 614 115624 620
rect 115754 0 115810 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117594 0 117650 800
rect 117962 0 118018 800
rect 118330 0 118386 800
rect 118712 800 118740 2858
rect 118804 2038 118832 7686
rect 118988 7410 119016 7686
rect 118976 7404 119028 7410
rect 118976 7346 119028 7352
rect 120632 7404 120684 7410
rect 120632 7346 120684 7352
rect 118988 7002 119016 7346
rect 118976 6996 119028 7002
rect 118976 6938 119028 6944
rect 120644 6662 120672 7346
rect 120632 6656 120684 6662
rect 120632 6598 120684 6604
rect 118884 4820 118936 4826
rect 118884 4762 118936 4768
rect 118792 2032 118844 2038
rect 118792 1974 118844 1980
rect 118790 1728 118846 1737
rect 118790 1663 118846 1672
rect 118804 1562 118832 1663
rect 118792 1556 118844 1562
rect 118792 1498 118844 1504
rect 118896 1426 118924 4762
rect 120080 4140 120132 4146
rect 120080 4082 120132 4088
rect 120092 3398 120120 4082
rect 120080 3392 120132 3398
rect 120080 3334 120132 3340
rect 119436 3052 119488 3058
rect 119436 2994 119488 3000
rect 118976 2372 119028 2378
rect 118976 2314 119028 2320
rect 118988 1766 119016 2314
rect 119160 2304 119212 2310
rect 119160 2246 119212 2252
rect 119344 2304 119396 2310
rect 119344 2246 119396 2252
rect 119172 2038 119200 2246
rect 119160 2032 119212 2038
rect 119160 1974 119212 1980
rect 118976 1760 119028 1766
rect 118976 1702 119028 1708
rect 118884 1420 118936 1426
rect 118884 1362 118936 1368
rect 119066 1048 119122 1057
rect 119066 983 119122 992
rect 119080 800 119108 983
rect 119356 882 119384 2246
rect 119344 876 119396 882
rect 119344 818 119396 824
rect 119448 800 119476 2994
rect 120080 2984 120132 2990
rect 120080 2926 120132 2932
rect 119804 2644 119856 2650
rect 119804 2586 119856 2592
rect 119712 1760 119764 1766
rect 119712 1702 119764 1708
rect 119724 1426 119752 1702
rect 119712 1420 119764 1426
rect 119712 1362 119764 1368
rect 119816 800 119844 2586
rect 119896 1760 119948 1766
rect 119896 1702 119948 1708
rect 119908 1358 119936 1702
rect 119896 1352 119948 1358
rect 119896 1294 119948 1300
rect 118424 750 118476 756
rect 118436 338 118464 750
rect 118424 332 118476 338
rect 118424 274 118476 280
rect 118698 0 118754 800
rect 119066 0 119122 800
rect 119434 0 119490 800
rect 119802 0 119858 800
rect 120092 746 120120 2926
rect 120264 2372 120316 2378
rect 120264 2314 120316 2320
rect 120172 1964 120224 1970
rect 120172 1906 120224 1912
rect 120184 1766 120212 1906
rect 120172 1760 120224 1766
rect 120172 1702 120224 1708
rect 120276 1306 120304 2314
rect 120644 2038 120672 6598
rect 120828 2650 120856 7754
rect 121460 7744 121512 7750
rect 121460 7686 121512 7692
rect 121368 7336 121420 7342
rect 121368 7278 121420 7284
rect 121380 7002 121408 7278
rect 121368 6996 121420 7002
rect 121368 6938 121420 6944
rect 121472 6254 121500 7686
rect 121828 6792 121880 6798
rect 121828 6734 121880 6740
rect 121460 6248 121512 6254
rect 121460 6190 121512 6196
rect 121472 5710 121500 6190
rect 121840 5710 121868 6734
rect 121460 5704 121512 5710
rect 121460 5646 121512 5652
rect 121828 5704 121880 5710
rect 121828 5646 121880 5652
rect 121920 5364 121972 5370
rect 121920 5306 121972 5312
rect 121932 4826 121960 5306
rect 121920 4820 121972 4826
rect 121920 4762 121972 4768
rect 121644 4140 121696 4146
rect 121644 4082 121696 4088
rect 121656 3398 121684 4082
rect 121736 4072 121788 4078
rect 121736 4014 121788 4020
rect 121748 3534 121776 4014
rect 122288 3936 122340 3942
rect 122288 3878 122340 3884
rect 121736 3528 121788 3534
rect 121736 3470 121788 3476
rect 121276 3392 121328 3398
rect 121276 3334 121328 3340
rect 121644 3392 121696 3398
rect 121644 3334 121696 3340
rect 120816 2644 120868 2650
rect 120816 2586 120868 2592
rect 120724 2576 120776 2582
rect 120722 2544 120724 2553
rect 120776 2544 120778 2553
rect 120722 2479 120778 2488
rect 120908 2440 120960 2446
rect 120908 2382 120960 2388
rect 120920 2310 120948 2382
rect 120908 2304 120960 2310
rect 120908 2246 120960 2252
rect 120540 2032 120592 2038
rect 120540 1974 120592 1980
rect 120632 2032 120684 2038
rect 120632 1974 120684 1980
rect 120356 1760 120408 1766
rect 120356 1702 120408 1708
rect 120368 1358 120396 1702
rect 120184 1278 120304 1306
rect 120356 1352 120408 1358
rect 120356 1294 120408 1300
rect 120184 800 120212 1278
rect 120552 800 120580 1974
rect 120920 800 120948 2246
rect 121184 2032 121236 2038
rect 121184 1974 121236 1980
rect 121000 1964 121052 1970
rect 121000 1906 121052 1912
rect 121012 1426 121040 1906
rect 121196 1766 121224 1974
rect 121184 1760 121236 1766
rect 121184 1702 121236 1708
rect 121000 1420 121052 1426
rect 121000 1362 121052 1368
rect 121288 800 121316 3334
rect 121656 800 121684 3334
rect 122012 1896 122064 1902
rect 122012 1838 122064 1844
rect 122024 800 122052 1838
rect 122300 1358 122328 3878
rect 122484 3058 122512 7754
rect 122746 7576 122802 7585
rect 122746 7511 122802 7520
rect 122760 7313 122788 7511
rect 122932 7404 122984 7410
rect 122932 7346 122984 7352
rect 122746 7304 122802 7313
rect 122746 7239 122802 7248
rect 122840 6248 122892 6254
rect 122840 6190 122892 6196
rect 122852 5710 122880 6190
rect 122840 5704 122892 5710
rect 122840 5646 122892 5652
rect 122748 4480 122800 4486
rect 122748 4422 122800 4428
rect 122472 3052 122524 3058
rect 122472 2994 122524 3000
rect 122380 2916 122432 2922
rect 122380 2858 122432 2864
rect 122392 2650 122420 2858
rect 122656 2848 122708 2854
rect 122656 2790 122708 2796
rect 122380 2644 122432 2650
rect 122380 2586 122432 2592
rect 122380 1964 122432 1970
rect 122380 1906 122432 1912
rect 122288 1352 122340 1358
rect 122288 1294 122340 1300
rect 122392 800 122420 1906
rect 122668 882 122696 2790
rect 122656 876 122708 882
rect 122656 818 122708 824
rect 122760 800 122788 4422
rect 122944 2038 122972 7346
rect 123022 6760 123078 6769
rect 123022 6695 123024 6704
rect 123076 6695 123078 6704
rect 123024 6666 123076 6672
rect 124220 6656 124272 6662
rect 124220 6598 124272 6604
rect 123024 6316 123076 6322
rect 123024 6258 123076 6264
rect 123036 5574 123064 6258
rect 124128 6112 124180 6118
rect 124126 6080 124128 6089
rect 124180 6080 124182 6089
rect 124126 6015 124182 6024
rect 123116 5636 123168 5642
rect 123116 5578 123168 5584
rect 123024 5568 123076 5574
rect 123024 5510 123076 5516
rect 122932 2032 122984 2038
rect 122932 1974 122984 1980
rect 122840 1964 122892 1970
rect 122840 1906 122892 1912
rect 122852 1222 122880 1906
rect 122840 1216 122892 1222
rect 122840 1158 122892 1164
rect 123128 800 123156 5578
rect 123760 5568 123812 5574
rect 123760 5510 123812 5516
rect 123484 3392 123536 3398
rect 123484 3334 123536 3340
rect 123496 800 123524 3334
rect 123772 2650 123800 5510
rect 123852 2916 123904 2922
rect 123852 2858 123904 2864
rect 123760 2644 123812 2650
rect 123760 2586 123812 2592
rect 123864 800 123892 2858
rect 124232 2650 124260 6598
rect 124680 5228 124732 5234
rect 124680 5170 124732 5176
rect 124588 4140 124640 4146
rect 124588 4082 124640 4088
rect 124600 3398 124628 4082
rect 124588 3392 124640 3398
rect 124588 3334 124640 3340
rect 124220 2644 124272 2650
rect 124220 2586 124272 2592
rect 124220 2440 124272 2446
rect 124220 2382 124272 2388
rect 124232 2310 124260 2382
rect 124220 2304 124272 2310
rect 124220 2246 124272 2252
rect 123944 1760 123996 1766
rect 123944 1702 123996 1708
rect 123956 1426 123984 1702
rect 123944 1420 123996 1426
rect 123944 1362 123996 1368
rect 123956 882 123984 1362
rect 124128 1216 124180 1222
rect 124180 1164 124260 1170
rect 124128 1158 124260 1164
rect 124140 1142 124260 1158
rect 123944 876 123996 882
rect 123944 818 123996 824
rect 124232 800 124260 1142
rect 124600 800 124628 3334
rect 124692 2038 124720 5170
rect 124968 3738 124996 8026
rect 125612 7970 125640 8758
rect 125704 8498 125732 8774
rect 125692 8492 125744 8498
rect 125692 8434 125744 8440
rect 125704 8090 125732 8434
rect 125692 8084 125744 8090
rect 125692 8026 125744 8032
rect 125612 7942 125732 7970
rect 125416 7336 125468 7342
rect 125416 7278 125468 7284
rect 125428 6866 125456 7278
rect 125416 6860 125468 6866
rect 125416 6802 125468 6808
rect 125600 4140 125652 4146
rect 125600 4082 125652 4088
rect 124956 3732 125008 3738
rect 124956 3674 125008 3680
rect 124956 3528 125008 3534
rect 124956 3470 125008 3476
rect 124680 2032 124732 2038
rect 124680 1974 124732 1980
rect 124968 800 124996 3470
rect 125612 3398 125640 4082
rect 125704 3738 125732 7942
rect 125692 3732 125744 3738
rect 125692 3674 125744 3680
rect 125600 3392 125652 3398
rect 125600 3334 125652 3340
rect 125796 2990 125824 8978
rect 125968 8424 126020 8430
rect 125968 8366 126020 8372
rect 125876 4276 125928 4282
rect 125876 4218 125928 4224
rect 125784 2984 125836 2990
rect 125784 2926 125836 2932
rect 125888 2836 125916 4218
rect 125980 4146 126008 8366
rect 126256 7954 126284 9862
rect 126900 9654 126928 12242
rect 126978 12200 127034 13000
rect 127346 12200 127402 13000
rect 127714 12200 127770 13000
rect 128082 12200 128138 13000
rect 128450 12200 128506 13000
rect 128818 12200 128874 13000
rect 129186 12200 129242 13000
rect 129554 12200 129610 13000
rect 129922 12200 129978 13000
rect 130290 12200 130346 13000
rect 130658 12200 130714 13000
rect 131026 12200 131082 13000
rect 131394 12200 131450 13000
rect 131762 12200 131818 13000
rect 132130 12200 132186 13000
rect 132498 12200 132554 13000
rect 132866 12200 132922 13000
rect 133234 12200 133290 13000
rect 133602 12200 133658 13000
rect 133970 12200 134026 13000
rect 134338 12200 134394 13000
rect 134706 12200 134762 13000
rect 135074 12200 135130 13000
rect 135442 12200 135498 13000
rect 135810 12200 135866 13000
rect 136178 12200 136234 13000
rect 136546 12200 136602 13000
rect 136640 12504 136692 12510
rect 136640 12446 136692 12452
rect 126992 11778 127020 12200
rect 126992 11750 127112 11778
rect 126980 11688 127032 11694
rect 126980 11630 127032 11636
rect 126992 11082 127020 11630
rect 126980 11076 127032 11082
rect 126980 11018 127032 11024
rect 127084 10674 127112 11750
rect 127164 11348 127216 11354
rect 127164 11290 127216 11296
rect 127176 10810 127204 11290
rect 127164 10804 127216 10810
rect 127164 10746 127216 10752
rect 127072 10668 127124 10674
rect 127072 10610 127124 10616
rect 127360 10266 127388 12200
rect 127728 11778 127756 12200
rect 127900 12164 127952 12170
rect 127900 12106 127952 12112
rect 127544 11750 127756 11778
rect 127440 10464 127492 10470
rect 127440 10406 127492 10412
rect 127452 10266 127480 10406
rect 127348 10260 127400 10266
rect 127348 10202 127400 10208
rect 127440 10260 127492 10266
rect 127440 10202 127492 10208
rect 127360 10062 127388 10202
rect 127544 10198 127572 11750
rect 127716 11688 127768 11694
rect 127716 11630 127768 11636
rect 127728 11354 127756 11630
rect 127716 11348 127768 11354
rect 127716 11290 127768 11296
rect 127912 11082 127940 12106
rect 128096 11762 128124 12200
rect 128464 11830 128492 12200
rect 128452 11824 128504 11830
rect 128452 11766 128504 11772
rect 128084 11756 128136 11762
rect 128084 11698 128136 11704
rect 128832 11082 128860 12200
rect 127808 11076 127860 11082
rect 127808 11018 127860 11024
rect 127900 11076 127952 11082
rect 127900 11018 127952 11024
rect 128820 11076 128872 11082
rect 128820 11018 128872 11024
rect 127624 10668 127676 10674
rect 127624 10610 127676 10616
rect 127636 10470 127664 10610
rect 127624 10464 127676 10470
rect 127624 10406 127676 10412
rect 127532 10192 127584 10198
rect 127532 10134 127584 10140
rect 127348 10056 127400 10062
rect 127348 9998 127400 10004
rect 126888 9648 126940 9654
rect 126888 9590 126940 9596
rect 127072 9580 127124 9586
rect 127072 9522 127124 9528
rect 127084 9178 127112 9522
rect 127164 9512 127216 9518
rect 127164 9454 127216 9460
rect 127072 9172 127124 9178
rect 127072 9114 127124 9120
rect 126704 8900 126756 8906
rect 126704 8842 126756 8848
rect 126716 8430 126744 8842
rect 127176 8838 127204 9454
rect 127532 9376 127584 9382
rect 127532 9318 127584 9324
rect 127544 9042 127572 9318
rect 127532 9036 127584 9042
rect 127532 8978 127584 8984
rect 127164 8832 127216 8838
rect 127164 8774 127216 8780
rect 127072 8560 127124 8566
rect 127072 8502 127124 8508
rect 126704 8424 126756 8430
rect 126704 8366 126756 8372
rect 126244 7948 126296 7954
rect 126244 7890 126296 7896
rect 127084 7750 127112 8502
rect 127072 7744 127124 7750
rect 127072 7686 127124 7692
rect 126888 7404 126940 7410
rect 126888 7346 126940 7352
rect 126900 6746 126928 7346
rect 126900 6718 127020 6746
rect 126992 6662 127020 6718
rect 126980 6656 127032 6662
rect 126980 6598 127032 6604
rect 126060 5568 126112 5574
rect 126060 5510 126112 5516
rect 125968 4140 126020 4146
rect 125968 4082 126020 4088
rect 125796 2808 125916 2836
rect 125796 2666 125824 2808
rect 125704 2638 125824 2666
rect 126072 2650 126100 5510
rect 126888 4140 126940 4146
rect 126888 4082 126940 4088
rect 126428 3936 126480 3942
rect 126428 3878 126480 3884
rect 126440 3534 126468 3878
rect 126612 3596 126664 3602
rect 126612 3538 126664 3544
rect 126428 3528 126480 3534
rect 126428 3470 126480 3476
rect 126336 3392 126388 3398
rect 126388 3352 126468 3380
rect 126336 3334 126388 3340
rect 126060 2644 126112 2650
rect 125600 2440 125652 2446
rect 125600 2382 125652 2388
rect 125612 2310 125640 2382
rect 125324 2304 125376 2310
rect 125324 2246 125376 2252
rect 125600 2304 125652 2310
rect 125600 2246 125652 2252
rect 125336 800 125364 2246
rect 125612 2038 125640 2246
rect 125600 2032 125652 2038
rect 125600 1974 125652 1980
rect 125598 1048 125654 1057
rect 125598 983 125654 992
rect 125612 882 125640 983
rect 125600 876 125652 882
rect 125600 818 125652 824
rect 125704 800 125732 2638
rect 126060 2586 126112 2592
rect 126152 1896 126204 1902
rect 126152 1838 126204 1844
rect 126060 1760 126112 1766
rect 126060 1702 126112 1708
rect 125784 1352 125836 1358
rect 125784 1294 125836 1300
rect 120080 740 120132 746
rect 120080 682 120132 688
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 125796 746 125824 1294
rect 126072 800 126100 1702
rect 126164 1494 126192 1838
rect 126244 1760 126296 1766
rect 126244 1702 126296 1708
rect 126152 1488 126204 1494
rect 126152 1430 126204 1436
rect 126256 1426 126284 1702
rect 126244 1420 126296 1426
rect 126244 1362 126296 1368
rect 126150 1048 126206 1057
rect 126150 983 126206 992
rect 126164 882 126192 983
rect 126152 876 126204 882
rect 126152 818 126204 824
rect 126440 800 126468 3352
rect 126624 1902 126652 3538
rect 126900 3398 126928 4082
rect 126888 3392 126940 3398
rect 126888 3334 126940 3340
rect 126888 3052 126940 3058
rect 126888 2994 126940 3000
rect 126900 2854 126928 2994
rect 126888 2848 126940 2854
rect 126888 2790 126940 2796
rect 126900 2650 126928 2790
rect 126992 2650 127020 6598
rect 127176 4146 127204 8774
rect 127544 7954 127572 8978
rect 127532 7948 127584 7954
rect 127532 7890 127584 7896
rect 127440 7336 127492 7342
rect 127440 7278 127492 7284
rect 127452 6866 127480 7278
rect 127440 6860 127492 6866
rect 127440 6802 127492 6808
rect 127636 5370 127664 10406
rect 127820 9654 127848 11018
rect 128268 11008 128320 11014
rect 128268 10950 128320 10956
rect 128280 10810 128308 10950
rect 128268 10804 128320 10810
rect 128268 10746 128320 10752
rect 129200 10674 129228 12200
rect 129568 10690 129596 12200
rect 129740 11688 129792 11694
rect 129740 11630 129792 11636
rect 128360 10668 128412 10674
rect 128360 10610 128412 10616
rect 129188 10668 129240 10674
rect 129188 10610 129240 10616
rect 129476 10662 129596 10690
rect 128084 10464 128136 10470
rect 128084 10406 128136 10412
rect 128096 10062 128124 10406
rect 128372 10266 128400 10610
rect 129002 10296 129058 10305
rect 128360 10260 128412 10266
rect 129002 10231 129058 10240
rect 128360 10202 128412 10208
rect 129016 10130 129044 10231
rect 129004 10124 129056 10130
rect 129004 10066 129056 10072
rect 128084 10056 128136 10062
rect 128084 9998 128136 10004
rect 127808 9648 127860 9654
rect 127808 9590 127860 9596
rect 128096 8634 128124 9998
rect 129188 9716 129240 9722
rect 129188 9658 129240 9664
rect 128084 8628 128136 8634
rect 128084 8570 128136 8576
rect 127992 7744 128044 7750
rect 127992 7686 128044 7692
rect 127624 5364 127676 5370
rect 127624 5306 127676 5312
rect 127164 4140 127216 4146
rect 127164 4082 127216 4088
rect 128004 2990 128032 7686
rect 128544 6792 128596 6798
rect 128544 6734 128596 6740
rect 128360 5228 128412 5234
rect 128360 5170 128412 5176
rect 128372 4486 128400 5170
rect 128360 4480 128412 4486
rect 128360 4422 128412 4428
rect 128176 3052 128228 3058
rect 128176 2994 128228 3000
rect 127992 2984 128044 2990
rect 127992 2926 128044 2932
rect 127900 2848 127952 2854
rect 127900 2790 127952 2796
rect 126888 2644 126940 2650
rect 126888 2586 126940 2592
rect 126980 2644 127032 2650
rect 126980 2586 127032 2592
rect 127532 2440 127584 2446
rect 127532 2382 127584 2388
rect 127164 2304 127216 2310
rect 127164 2246 127216 2252
rect 126796 2032 126848 2038
rect 126796 1974 126848 1980
rect 126612 1896 126664 1902
rect 126612 1838 126664 1844
rect 126808 800 126836 1974
rect 127072 1964 127124 1970
rect 126992 1924 127072 1952
rect 126992 1222 127020 1924
rect 127072 1906 127124 1912
rect 126980 1216 127032 1222
rect 126980 1158 127032 1164
rect 125784 740 125836 746
rect 125784 682 125836 688
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 126992 678 127020 1158
rect 127176 800 127204 2246
rect 127544 800 127572 2382
rect 127912 800 127940 2790
rect 128188 2310 128216 2994
rect 128176 2304 128228 2310
rect 128176 2246 128228 2252
rect 128268 1964 128320 1970
rect 128268 1906 128320 1912
rect 128280 1222 128308 1906
rect 128556 1834 128584 6734
rect 128912 6248 128964 6254
rect 128912 6190 128964 6196
rect 128924 5914 128952 6190
rect 128912 5908 128964 5914
rect 128912 5850 128964 5856
rect 129200 4826 129228 9658
rect 129476 9586 129504 10662
rect 129556 10600 129608 10606
rect 129556 10542 129608 10548
rect 129568 10266 129596 10542
rect 129556 10260 129608 10266
rect 129556 10202 129608 10208
rect 129752 10130 129780 11630
rect 129740 10124 129792 10130
rect 129740 10066 129792 10072
rect 129936 10062 129964 12200
rect 130200 11552 130252 11558
rect 130200 11494 130252 11500
rect 130212 11150 130240 11494
rect 130304 11218 130332 12200
rect 130672 11830 130700 12200
rect 130660 11824 130712 11830
rect 130660 11766 130712 11772
rect 130476 11756 130528 11762
rect 130476 11698 130528 11704
rect 130488 11354 130516 11698
rect 130660 11620 130712 11626
rect 130660 11562 130712 11568
rect 130476 11348 130528 11354
rect 130476 11290 130528 11296
rect 130292 11212 130344 11218
rect 130292 11154 130344 11160
rect 130200 11144 130252 11150
rect 130200 11086 130252 11092
rect 130672 10674 130700 11562
rect 130660 10668 130712 10674
rect 130660 10610 130712 10616
rect 130672 10130 130700 10610
rect 130660 10124 130712 10130
rect 130660 10066 130712 10072
rect 129924 10056 129976 10062
rect 129924 9998 129976 10004
rect 130200 9920 130252 9926
rect 130200 9862 130252 9868
rect 129464 9580 129516 9586
rect 129464 9522 129516 9528
rect 129832 9512 129884 9518
rect 129832 9454 129884 9460
rect 129740 8832 129792 8838
rect 129740 8774 129792 8780
rect 129556 8424 129608 8430
rect 129556 8366 129608 8372
rect 129568 8090 129596 8366
rect 129556 8084 129608 8090
rect 129556 8026 129608 8032
rect 129752 7954 129780 8774
rect 129844 7954 129872 9454
rect 129740 7948 129792 7954
rect 129740 7890 129792 7896
rect 129832 7948 129884 7954
rect 129832 7890 129884 7896
rect 129832 7336 129884 7342
rect 129832 7278 129884 7284
rect 129844 6866 129872 7278
rect 129832 6860 129884 6866
rect 129832 6802 129884 6808
rect 130016 6384 130068 6390
rect 130016 6326 130068 6332
rect 130028 5778 130056 6326
rect 130016 5772 130068 5778
rect 130016 5714 130068 5720
rect 130212 4826 130240 9862
rect 131040 9518 131068 12200
rect 131304 11552 131356 11558
rect 131304 11494 131356 11500
rect 131120 11076 131172 11082
rect 131120 11018 131172 11024
rect 131132 9586 131160 11018
rect 131120 9580 131172 9586
rect 131120 9522 131172 9528
rect 130752 9512 130804 9518
rect 130752 9454 130804 9460
rect 131028 9512 131080 9518
rect 131028 9454 131080 9460
rect 130764 9110 130792 9454
rect 130752 9104 130804 9110
rect 130752 9046 130804 9052
rect 131118 9072 131174 9081
rect 130292 9036 130344 9042
rect 131118 9007 131120 9016
rect 130292 8978 130344 8984
rect 131172 9007 131174 9016
rect 131120 8978 131172 8984
rect 129188 4820 129240 4826
rect 129188 4762 129240 4768
rect 130200 4820 130252 4826
rect 130200 4762 130252 4768
rect 129372 4480 129424 4486
rect 129372 4422 129424 4428
rect 128636 3392 128688 3398
rect 128636 3334 128688 3340
rect 128544 1828 128596 1834
rect 128544 1770 128596 1776
rect 128268 1216 128320 1222
rect 128268 1158 128320 1164
rect 128280 800 128308 1158
rect 128648 800 128676 3334
rect 129004 2304 129056 2310
rect 129004 2246 129056 2252
rect 129016 800 129044 2246
rect 129188 1760 129240 1766
rect 129188 1702 129240 1708
rect 129200 1426 129228 1702
rect 129188 1420 129240 1426
rect 129188 1362 129240 1368
rect 129200 882 129228 1362
rect 129188 876 129240 882
rect 129188 818 129240 824
rect 129384 800 129412 4422
rect 130304 4146 130332 8978
rect 131028 8492 131080 8498
rect 131028 8434 131080 8440
rect 131040 7750 131068 8434
rect 131212 8288 131264 8294
rect 131212 8230 131264 8236
rect 131224 8022 131252 8230
rect 131212 8016 131264 8022
rect 131212 7958 131264 7964
rect 131028 7744 131080 7750
rect 131028 7686 131080 7692
rect 130936 5568 130988 5574
rect 130936 5510 130988 5516
rect 130476 4548 130528 4554
rect 130476 4490 130528 4496
rect 130200 4140 130252 4146
rect 130200 4082 130252 4088
rect 130292 4140 130344 4146
rect 130292 4082 130344 4088
rect 129832 4072 129884 4078
rect 129832 4014 129884 4020
rect 129740 3528 129792 3534
rect 129740 3470 129792 3476
rect 129752 800 129780 3470
rect 129844 1426 129872 4014
rect 130212 3602 130240 4082
rect 130200 3596 130252 3602
rect 130200 3538 130252 3544
rect 130108 2440 130160 2446
rect 130108 2382 130160 2388
rect 129832 1420 129884 1426
rect 129832 1362 129884 1368
rect 130120 800 130148 2382
rect 130488 800 130516 4490
rect 130844 4480 130896 4486
rect 130844 4422 130896 4428
rect 130660 2032 130712 2038
rect 130660 1974 130712 1980
rect 130672 1494 130700 1974
rect 130660 1488 130712 1494
rect 130660 1430 130712 1436
rect 130856 800 130884 4422
rect 130948 2106 130976 5510
rect 131040 3738 131068 7686
rect 131120 6792 131172 6798
rect 131120 6734 131172 6740
rect 131028 3732 131080 3738
rect 131028 3674 131080 3680
rect 131132 2446 131160 6734
rect 131316 4826 131344 11494
rect 131408 10826 131436 12200
rect 131776 11762 131804 12200
rect 131764 11756 131816 11762
rect 131764 11698 131816 11704
rect 131948 11280 132000 11286
rect 131948 11222 132000 11228
rect 131408 10798 131620 10826
rect 131960 10810 131988 11222
rect 131592 10742 131620 10798
rect 131948 10804 132000 10810
rect 131948 10746 132000 10752
rect 131580 10736 131632 10742
rect 131580 10678 131632 10684
rect 132144 9450 132172 12200
rect 132512 11778 132540 12200
rect 132880 12170 132908 12200
rect 132868 12164 132920 12170
rect 132868 12106 132920 12112
rect 133248 11914 133276 12200
rect 132684 11892 132736 11898
rect 133248 11886 133368 11914
rect 132684 11834 132736 11840
rect 132512 11750 132632 11778
rect 132500 11688 132552 11694
rect 132500 11630 132552 11636
rect 132512 11082 132540 11630
rect 132500 11076 132552 11082
rect 132500 11018 132552 11024
rect 132408 10464 132460 10470
rect 132408 10406 132460 10412
rect 132420 10130 132448 10406
rect 132408 10124 132460 10130
rect 132408 10066 132460 10072
rect 132420 9722 132448 10066
rect 132408 9716 132460 9722
rect 132408 9658 132460 9664
rect 132604 9586 132632 11750
rect 132696 11694 132724 11834
rect 133236 11756 133288 11762
rect 133236 11698 133288 11704
rect 132684 11688 132736 11694
rect 132684 11630 132736 11636
rect 133248 11354 133276 11698
rect 133236 11348 133288 11354
rect 133236 11290 133288 11296
rect 133144 11076 133196 11082
rect 133144 11018 133196 11024
rect 132960 10600 133012 10606
rect 132960 10542 133012 10548
rect 132972 10266 133000 10542
rect 132960 10260 133012 10266
rect 132960 10202 133012 10208
rect 133156 9654 133184 11018
rect 133340 9654 133368 11886
rect 133512 10464 133564 10470
rect 133512 10406 133564 10412
rect 133418 10160 133474 10169
rect 133418 10095 133420 10104
rect 133472 10095 133474 10104
rect 133420 10066 133472 10072
rect 133524 10062 133552 10406
rect 133512 10056 133564 10062
rect 133512 9998 133564 10004
rect 133144 9648 133196 9654
rect 133144 9590 133196 9596
rect 133328 9648 133380 9654
rect 133328 9590 133380 9596
rect 132592 9580 132644 9586
rect 132592 9522 132644 9528
rect 132132 9444 132184 9450
rect 132132 9386 132184 9392
rect 131396 8968 131448 8974
rect 131396 8910 131448 8916
rect 132406 8936 132462 8945
rect 131304 4820 131356 4826
rect 131304 4762 131356 4768
rect 131408 4146 131436 8910
rect 132406 8871 132462 8880
rect 132682 8936 132738 8945
rect 132682 8871 132738 8880
rect 132420 8616 132448 8871
rect 132696 8616 132724 8871
rect 132420 8588 132724 8616
rect 133052 8288 133104 8294
rect 133052 8230 133104 8236
rect 133064 7954 133092 8230
rect 133052 7948 133104 7954
rect 133052 7890 133104 7896
rect 133420 7880 133472 7886
rect 133420 7822 133472 7828
rect 133236 7404 133288 7410
rect 133236 7346 133288 7352
rect 132224 7336 132276 7342
rect 132224 7278 132276 7284
rect 132236 7002 132264 7278
rect 132224 6996 132276 7002
rect 132224 6938 132276 6944
rect 133248 6662 133276 7346
rect 133432 7342 133460 7822
rect 133420 7336 133472 7342
rect 133420 7278 133472 7284
rect 133236 6656 133288 6662
rect 133236 6598 133288 6604
rect 132684 4480 132736 4486
rect 132684 4422 132736 4428
rect 131304 4140 131356 4146
rect 131304 4082 131356 4088
rect 131396 4140 131448 4146
rect 131396 4082 131448 4088
rect 131316 3398 131344 4082
rect 131580 3596 131632 3602
rect 131580 3538 131632 3544
rect 131304 3392 131356 3398
rect 131304 3334 131356 3340
rect 131120 2440 131172 2446
rect 131120 2382 131172 2388
rect 131028 2372 131080 2378
rect 131028 2314 131080 2320
rect 130936 2100 130988 2106
rect 130936 2042 130988 2048
rect 131040 1902 131068 2314
rect 131212 1964 131264 1970
rect 131212 1906 131264 1912
rect 131028 1896 131080 1902
rect 131028 1838 131080 1844
rect 131040 1358 131068 1838
rect 131028 1352 131080 1358
rect 131028 1294 131080 1300
rect 131224 1222 131252 1906
rect 131212 1216 131264 1222
rect 131212 1158 131264 1164
rect 131224 800 131252 1158
rect 131592 800 131620 3538
rect 131948 3528 132000 3534
rect 131948 3470 132000 3476
rect 131762 912 131818 921
rect 131762 847 131818 856
rect 126980 672 127032 678
rect 126980 614 127032 620
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 131776 746 131804 847
rect 131960 800 131988 3470
rect 132316 3392 132368 3398
rect 132316 3334 132368 3340
rect 132040 1216 132092 1222
rect 132040 1158 132092 1164
rect 131764 740 131816 746
rect 131764 682 131816 688
rect 131946 0 132002 800
rect 132052 338 132080 1158
rect 132328 800 132356 3334
rect 132500 1760 132552 1766
rect 132500 1702 132552 1708
rect 132132 672 132184 678
rect 132132 614 132184 620
rect 132144 406 132172 614
rect 132132 400 132184 406
rect 132132 342 132184 348
rect 132040 332 132092 338
rect 132040 274 132092 280
rect 132314 0 132370 800
rect 132512 678 132540 1702
rect 132696 800 132724 4422
rect 133248 3194 133276 6598
rect 133524 3738 133552 9998
rect 133616 9382 133644 12200
rect 133604 9376 133656 9382
rect 133604 9318 133656 9324
rect 133984 9178 134012 12200
rect 134352 12170 134380 12200
rect 134340 12164 134392 12170
rect 134340 12106 134392 12112
rect 134720 11898 134748 12200
rect 134708 11892 134760 11898
rect 134708 11834 134760 11840
rect 135088 11830 135116 12200
rect 135456 12102 135484 12200
rect 135260 12096 135312 12102
rect 135260 12038 135312 12044
rect 135444 12096 135496 12102
rect 135444 12038 135496 12044
rect 135076 11824 135128 11830
rect 135076 11766 135128 11772
rect 134340 11552 134392 11558
rect 134340 11494 134392 11500
rect 134352 11150 134380 11494
rect 135272 11218 135300 12038
rect 135628 11552 135680 11558
rect 135628 11494 135680 11500
rect 135640 11286 135668 11494
rect 135628 11280 135680 11286
rect 135628 11222 135680 11228
rect 135260 11212 135312 11218
rect 135260 11154 135312 11160
rect 134340 11144 134392 11150
rect 134340 11086 134392 11092
rect 135168 11144 135220 11150
rect 135168 11086 135220 11092
rect 135076 10736 135128 10742
rect 135076 10678 135128 10684
rect 134064 10668 134116 10674
rect 134064 10610 134116 10616
rect 134076 10266 134104 10610
rect 135088 10266 135116 10678
rect 134064 10260 134116 10266
rect 134064 10202 134116 10208
rect 135076 10260 135128 10266
rect 135076 10202 135128 10208
rect 134076 9518 134104 10202
rect 134800 10056 134852 10062
rect 134800 9998 134852 10004
rect 134064 9512 134116 9518
rect 134064 9454 134116 9460
rect 134812 9450 134840 9998
rect 135180 9654 135208 11086
rect 135168 9648 135220 9654
rect 135168 9590 135220 9596
rect 134800 9444 134852 9450
rect 134800 9386 134852 9392
rect 135824 9382 135852 12200
rect 136088 11688 136140 11694
rect 136088 11630 136140 11636
rect 135996 11552 136048 11558
rect 135996 11494 136048 11500
rect 136008 11150 136036 11494
rect 136100 11354 136128 11630
rect 136088 11348 136140 11354
rect 136088 11290 136140 11296
rect 135996 11144 136048 11150
rect 135996 11086 136048 11092
rect 135812 9376 135864 9382
rect 135812 9318 135864 9324
rect 133972 9172 134024 9178
rect 133972 9114 134024 9120
rect 136192 9110 136220 12200
rect 136560 12152 136588 12200
rect 136652 12152 136680 12446
rect 136914 12200 136970 13000
rect 137008 12436 137060 12442
rect 137008 12378 137060 12384
rect 136560 12124 136680 12152
rect 136928 12152 136956 12200
rect 137020 12152 137048 12378
rect 137192 12232 137244 12238
rect 137282 12200 137338 13000
rect 137376 12300 137428 12306
rect 137376 12242 137428 12248
rect 137192 12174 137244 12180
rect 136928 12124 137048 12152
rect 137204 11762 137232 12174
rect 137296 12084 137324 12200
rect 137388 12084 137416 12242
rect 137650 12200 137706 13000
rect 137836 12232 137888 12238
rect 137296 12056 137416 12084
rect 137664 12084 137692 12200
rect 138018 12200 138074 13000
rect 138386 12200 138442 13000
rect 138754 12200 138810 13000
rect 139122 12200 139178 13000
rect 139490 12200 139546 13000
rect 139858 12200 139914 13000
rect 140226 12200 140282 13000
rect 140594 12200 140650 13000
rect 140962 12200 141018 13000
rect 141330 12200 141386 13000
rect 141698 12200 141754 13000
rect 142066 12200 142122 13000
rect 142434 12200 142490 13000
rect 142802 12200 142858 13000
rect 143170 12200 143226 13000
rect 143538 12200 143594 13000
rect 143906 12200 143962 13000
rect 144274 12200 144330 13000
rect 144642 12200 144698 13000
rect 144736 12368 144788 12374
rect 144736 12310 144788 12316
rect 137836 12174 137888 12180
rect 137848 12084 137876 12174
rect 137664 12056 137876 12084
rect 137192 11756 137244 11762
rect 137192 11698 137244 11704
rect 137204 11354 137232 11698
rect 138032 11642 138060 12200
rect 138400 11914 138428 12200
rect 138400 11886 138520 11914
rect 138388 11756 138440 11762
rect 138388 11698 138440 11704
rect 138032 11614 138244 11642
rect 137468 11552 137520 11558
rect 137468 11494 137520 11500
rect 138112 11552 138164 11558
rect 138112 11494 138164 11500
rect 137192 11348 137244 11354
rect 137192 11290 137244 11296
rect 137480 11218 137508 11494
rect 137468 11212 137520 11218
rect 137468 11154 137520 11160
rect 138124 11150 138152 11494
rect 136640 11144 136692 11150
rect 136640 11086 136692 11092
rect 138112 11144 138164 11150
rect 138112 11086 138164 11092
rect 136272 10600 136324 10606
rect 136272 10542 136324 10548
rect 136284 10130 136312 10542
rect 136272 10124 136324 10130
rect 136272 10066 136324 10072
rect 136652 9586 136680 11086
rect 137468 10668 137520 10674
rect 137468 10610 137520 10616
rect 137480 10266 137508 10610
rect 138020 10464 138072 10470
rect 138020 10406 138072 10412
rect 137468 10260 137520 10266
rect 137468 10202 137520 10208
rect 138032 10062 138060 10406
rect 138020 10056 138072 10062
rect 137834 10024 137890 10033
rect 138020 9998 138072 10004
rect 137834 9959 137836 9968
rect 137888 9959 137890 9968
rect 137836 9930 137888 9936
rect 136640 9580 136692 9586
rect 136640 9522 136692 9528
rect 136180 9104 136232 9110
rect 136180 9046 136232 9052
rect 138032 9042 138060 9998
rect 138124 9654 138152 11086
rect 138112 9648 138164 9654
rect 138112 9590 138164 9596
rect 138216 9382 138244 11614
rect 138400 9586 138428 11698
rect 138388 9580 138440 9586
rect 138388 9522 138440 9528
rect 138492 9518 138520 11886
rect 138768 9586 138796 12200
rect 139136 10826 139164 12200
rect 139504 11286 139532 12200
rect 139492 11280 139544 11286
rect 139492 11222 139544 11228
rect 139136 10798 139256 10826
rect 139124 10736 139176 10742
rect 139124 10678 139176 10684
rect 139032 10668 139084 10674
rect 139032 10610 139084 10616
rect 139044 9994 139072 10610
rect 139136 10062 139164 10678
rect 139124 10056 139176 10062
rect 139124 9998 139176 10004
rect 139032 9988 139084 9994
rect 139032 9930 139084 9936
rect 138756 9580 138808 9586
rect 138756 9522 138808 9528
rect 138480 9512 138532 9518
rect 138480 9454 138532 9460
rect 139044 9450 139072 9930
rect 139032 9444 139084 9450
rect 139032 9386 139084 9392
rect 138112 9376 138164 9382
rect 138112 9318 138164 9324
rect 138204 9376 138256 9382
rect 138204 9318 138256 9324
rect 138020 9036 138072 9042
rect 138020 8978 138072 8984
rect 138124 8566 138152 9318
rect 138112 8560 138164 8566
rect 138112 8502 138164 8508
rect 139228 8498 139256 10798
rect 139872 8906 139900 12200
rect 140240 11778 140268 12200
rect 140240 11750 140360 11778
rect 140332 11694 140360 11750
rect 140228 11688 140280 11694
rect 140228 11630 140280 11636
rect 140320 11688 140372 11694
rect 140320 11630 140372 11636
rect 140240 11082 140268 11630
rect 140228 11076 140280 11082
rect 140228 11018 140280 11024
rect 140240 9654 140268 11018
rect 140412 10464 140464 10470
rect 140412 10406 140464 10412
rect 140424 10062 140452 10406
rect 140412 10056 140464 10062
rect 140412 9998 140464 10004
rect 140228 9648 140280 9654
rect 140228 9590 140280 9596
rect 140424 9042 140452 9998
rect 140412 9036 140464 9042
rect 140412 8978 140464 8984
rect 139860 8900 139912 8906
rect 139860 8842 139912 8848
rect 139216 8492 139268 8498
rect 139216 8434 139268 8440
rect 140608 8362 140636 12200
rect 140976 11506 141004 12200
rect 141344 11642 141372 12200
rect 141344 11614 141648 11642
rect 140976 11478 141188 11506
rect 141160 11234 141188 11478
rect 141273 11452 141569 11472
rect 141329 11450 141353 11452
rect 141409 11450 141433 11452
rect 141489 11450 141513 11452
rect 141351 11398 141353 11450
rect 141415 11398 141427 11450
rect 141489 11398 141491 11450
rect 141329 11396 141353 11398
rect 141409 11396 141433 11398
rect 141489 11396 141513 11398
rect 141273 11376 141569 11396
rect 141240 11280 141292 11286
rect 141160 11228 141240 11234
rect 141160 11222 141292 11228
rect 140872 11212 140924 11218
rect 141160 11206 141280 11222
rect 140872 11154 140924 11160
rect 140688 11076 140740 11082
rect 140688 11018 140740 11024
rect 140700 8974 140728 11018
rect 140778 10568 140834 10577
rect 140778 10503 140834 10512
rect 140792 10130 140820 10503
rect 140780 10124 140832 10130
rect 140780 10066 140832 10072
rect 140884 10062 140912 11154
rect 141056 10600 141108 10606
rect 141056 10542 141108 10548
rect 140872 10056 140924 10062
rect 140872 9998 140924 10004
rect 141068 9994 141096 10542
rect 141273 10364 141569 10384
rect 141329 10362 141353 10364
rect 141409 10362 141433 10364
rect 141489 10362 141513 10364
rect 141351 10310 141353 10362
rect 141415 10310 141427 10362
rect 141489 10310 141491 10362
rect 141329 10308 141353 10310
rect 141409 10308 141433 10310
rect 141489 10308 141513 10310
rect 141273 10288 141569 10308
rect 141056 9988 141108 9994
rect 141056 9930 141108 9936
rect 141068 9722 141096 9930
rect 141056 9716 141108 9722
rect 141056 9658 141108 9664
rect 141620 9654 141648 11614
rect 141608 9648 141660 9654
rect 141608 9590 141660 9596
rect 141516 9512 141568 9518
rect 141712 9466 141740 12200
rect 142080 9738 142108 12200
rect 142344 11212 142396 11218
rect 142344 11154 142396 11160
rect 142160 10668 142212 10674
rect 142160 10610 142212 10616
rect 142172 10130 142200 10610
rect 142252 10532 142304 10538
rect 142252 10474 142304 10480
rect 142160 10124 142212 10130
rect 142160 10066 142212 10072
rect 142172 10033 142200 10066
rect 142158 10024 142214 10033
rect 142158 9959 142214 9968
rect 141988 9710 142108 9738
rect 141568 9460 141648 9466
rect 141516 9454 141648 9460
rect 141528 9438 141648 9454
rect 141712 9450 141832 9466
rect 141712 9444 141844 9450
rect 141712 9438 141792 9444
rect 141273 9276 141569 9296
rect 141329 9274 141353 9276
rect 141409 9274 141433 9276
rect 141489 9274 141513 9276
rect 141351 9222 141353 9274
rect 141415 9222 141427 9274
rect 141489 9222 141491 9274
rect 141329 9220 141353 9222
rect 141409 9220 141433 9222
rect 141489 9220 141513 9222
rect 141273 9200 141569 9220
rect 140688 8968 140740 8974
rect 140688 8910 140740 8916
rect 140872 8832 140924 8838
rect 140872 8774 140924 8780
rect 140596 8356 140648 8362
rect 140596 8298 140648 8304
rect 140884 7954 140912 8774
rect 141620 8634 141648 9438
rect 141792 9386 141844 9392
rect 141988 8838 142016 9710
rect 142068 9648 142120 9654
rect 142068 9590 142120 9596
rect 141976 8832 142028 8838
rect 141976 8774 142028 8780
rect 141608 8628 141660 8634
rect 142080 8616 142108 9590
rect 142264 9382 142292 10474
rect 142356 9586 142384 11154
rect 142448 9654 142476 12200
rect 142436 9648 142488 9654
rect 142436 9590 142488 9596
rect 142344 9580 142396 9586
rect 142344 9522 142396 9528
rect 142252 9376 142304 9382
rect 142252 9318 142304 9324
rect 142816 9042 142844 12200
rect 143184 11914 143212 12200
rect 143184 11886 143488 11914
rect 143356 11756 143408 11762
rect 143356 11698 143408 11704
rect 143368 11150 143396 11698
rect 143356 11144 143408 11150
rect 143356 11086 143408 11092
rect 143172 9580 143224 9586
rect 143172 9522 143224 9528
rect 142896 9512 142948 9518
rect 142896 9454 142948 9460
rect 142804 9036 142856 9042
rect 142804 8978 142856 8984
rect 142252 8628 142304 8634
rect 142080 8588 142252 8616
rect 141608 8570 141660 8576
rect 142252 8570 142304 8576
rect 142436 8492 142488 8498
rect 142436 8434 142488 8440
rect 141792 8424 141844 8430
rect 141792 8366 141844 8372
rect 141273 8188 141569 8208
rect 141329 8186 141353 8188
rect 141409 8186 141433 8188
rect 141489 8186 141513 8188
rect 141351 8134 141353 8186
rect 141415 8134 141427 8186
rect 141489 8134 141491 8186
rect 141329 8132 141353 8134
rect 141409 8132 141433 8134
rect 141489 8132 141513 8134
rect 141273 8112 141569 8132
rect 141804 7954 141832 8366
rect 140872 7948 140924 7954
rect 140872 7890 140924 7896
rect 141792 7948 141844 7954
rect 141792 7890 141844 7896
rect 134248 7880 134300 7886
rect 134248 7822 134300 7828
rect 133512 3732 133564 3738
rect 133512 3674 133564 3680
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 133236 3188 133288 3194
rect 133236 3130 133288 3136
rect 133052 3052 133104 3058
rect 133052 2994 133104 3000
rect 133064 2310 133092 2994
rect 133052 2304 133104 2310
rect 133052 2246 133104 2252
rect 132960 876 133012 882
rect 132960 818 133012 824
rect 132500 672 132552 678
rect 132500 614 132552 620
rect 132682 0 132738 800
rect 132972 678 133000 818
rect 133064 800 133092 2246
rect 133696 1896 133748 1902
rect 133696 1838 133748 1844
rect 133420 1760 133472 1766
rect 133420 1702 133472 1708
rect 133432 800 133460 1702
rect 133708 1018 133736 1838
rect 133696 1012 133748 1018
rect 133696 954 133748 960
rect 133708 882 133736 954
rect 133696 876 133748 882
rect 133696 818 133748 824
rect 133800 800 133828 3470
rect 134260 3194 134288 7822
rect 142448 7546 142476 8434
rect 142804 8356 142856 8362
rect 142804 8298 142856 8304
rect 142816 7954 142844 8298
rect 142804 7948 142856 7954
rect 142804 7890 142856 7896
rect 142436 7540 142488 7546
rect 142436 7482 142488 7488
rect 142804 7336 142856 7342
rect 142804 7278 142856 7284
rect 134892 7200 134944 7206
rect 134892 7142 134944 7148
rect 141792 7200 141844 7206
rect 141792 7142 141844 7148
rect 134904 6798 134932 7142
rect 141273 7100 141569 7120
rect 141329 7098 141353 7100
rect 141409 7098 141433 7100
rect 141489 7098 141513 7100
rect 141351 7046 141353 7098
rect 141415 7046 141427 7098
rect 141489 7046 141491 7098
rect 141329 7044 141353 7046
rect 141409 7044 141433 7046
rect 141489 7044 141513 7046
rect 136178 7032 136234 7041
rect 141273 7024 141569 7044
rect 136178 6967 136234 6976
rect 136192 6934 136220 6967
rect 136180 6928 136232 6934
rect 136180 6870 136232 6876
rect 141804 6866 141832 7142
rect 141792 6860 141844 6866
rect 141792 6802 141844 6808
rect 134892 6792 134944 6798
rect 134892 6734 134944 6740
rect 135996 6792 136048 6798
rect 135996 6734 136048 6740
rect 134904 6390 134932 6734
rect 134892 6384 134944 6390
rect 134892 6326 134944 6332
rect 134892 4004 134944 4010
rect 134892 3946 134944 3952
rect 134248 3188 134300 3194
rect 134248 3130 134300 3136
rect 134156 3052 134208 3058
rect 134156 2994 134208 3000
rect 134168 2310 134196 2994
rect 134524 2916 134576 2922
rect 134524 2858 134576 2864
rect 134248 2440 134300 2446
rect 134248 2382 134300 2388
rect 134156 2304 134208 2310
rect 134156 2246 134208 2252
rect 134168 1766 134196 2246
rect 134156 1760 134208 1766
rect 134156 1702 134208 1708
rect 134260 1578 134288 2382
rect 134168 1550 134288 1578
rect 133878 1048 133934 1057
rect 133878 983 133880 992
rect 133932 983 133934 992
rect 133880 954 133932 960
rect 133972 808 134024 814
rect 132960 672 133012 678
rect 132960 614 133012 620
rect 132972 338 133000 614
rect 132960 332 133012 338
rect 132960 274 133012 280
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 133972 750 134024 756
rect 134064 808 134116 814
rect 134168 800 134196 1550
rect 134340 1216 134392 1222
rect 134432 1216 134484 1222
rect 134392 1176 134432 1204
rect 134340 1158 134392 1164
rect 134432 1158 134484 1164
rect 134536 800 134564 2858
rect 134616 1420 134668 1426
rect 134616 1362 134668 1368
rect 134628 1290 134656 1362
rect 134616 1284 134668 1290
rect 134616 1226 134668 1232
rect 134904 800 134932 3946
rect 135444 2848 135496 2854
rect 135444 2790 135496 2796
rect 135352 1896 135404 1902
rect 135352 1838 135404 1844
rect 135260 1488 135312 1494
rect 135260 1430 135312 1436
rect 135272 800 135300 1430
rect 135364 1426 135392 1838
rect 135456 1426 135484 2790
rect 136008 2446 136036 6734
rect 141804 6390 141832 6802
rect 142816 6390 142844 7278
rect 142908 6934 142936 9454
rect 143184 8974 143212 9522
rect 143368 9178 143396 11086
rect 143460 9178 143488 11886
rect 143552 9382 143580 12200
rect 143920 11762 143948 12200
rect 143908 11756 143960 11762
rect 143908 11698 143960 11704
rect 144000 11552 144052 11558
rect 144000 11494 144052 11500
rect 144012 11150 144040 11494
rect 144000 11144 144052 11150
rect 144000 11086 144052 11092
rect 144184 10600 144236 10606
rect 144184 10542 144236 10548
rect 144196 9926 144224 10542
rect 144184 9920 144236 9926
rect 144184 9862 144236 9868
rect 143540 9376 143592 9382
rect 143540 9318 143592 9324
rect 143356 9172 143408 9178
rect 143356 9114 143408 9120
rect 143448 9172 143500 9178
rect 143448 9114 143500 9120
rect 144196 9042 144224 9862
rect 144288 9518 144316 12200
rect 144656 12152 144684 12200
rect 144748 12152 144776 12310
rect 145010 12200 145066 13000
rect 145104 12504 145156 12510
rect 145104 12446 145156 12452
rect 144656 12124 144776 12152
rect 144828 11756 144880 11762
rect 144828 11698 144880 11704
rect 144552 11688 144604 11694
rect 144552 11630 144604 11636
rect 144564 11354 144592 11630
rect 144840 11354 144868 11698
rect 144920 11620 144972 11626
rect 144920 11562 144972 11568
rect 144552 11348 144604 11354
rect 144552 11290 144604 11296
rect 144828 11348 144880 11354
rect 144828 11290 144880 11296
rect 144932 10674 144960 11562
rect 145024 11234 145052 12200
rect 145116 11626 145144 12446
rect 145378 12200 145434 13000
rect 145746 12200 145802 13000
rect 146114 12200 146170 13000
rect 146482 12200 146538 13000
rect 146850 12200 146906 13000
rect 147218 12200 147274 13000
rect 147586 12200 147642 13000
rect 147954 12200 148010 13000
rect 148322 12200 148378 13000
rect 148690 12200 148746 13000
rect 149058 12200 149114 13000
rect 149426 12200 149482 13000
rect 149794 12200 149850 13000
rect 150162 12200 150218 13000
rect 150530 12200 150586 13000
rect 150898 12200 150954 13000
rect 151266 12200 151322 13000
rect 151634 12200 151690 13000
rect 152002 12200 152058 13000
rect 152370 12200 152426 13000
rect 152464 12436 152516 12442
rect 152464 12378 152516 12384
rect 145104 11620 145156 11626
rect 145104 11562 145156 11568
rect 145024 11206 145236 11234
rect 145012 11144 145064 11150
rect 145012 11086 145064 11092
rect 145024 10742 145052 11086
rect 145012 10736 145064 10742
rect 145012 10678 145064 10684
rect 144920 10668 144972 10674
rect 144920 10610 144972 10616
rect 145104 10532 145156 10538
rect 145104 10474 145156 10480
rect 144552 9920 144604 9926
rect 144552 9862 144604 9868
rect 144564 9722 144592 9862
rect 144552 9716 144604 9722
rect 144552 9658 144604 9664
rect 144276 9512 144328 9518
rect 144276 9454 144328 9460
rect 145116 9450 145144 10474
rect 145104 9444 145156 9450
rect 145104 9386 145156 9392
rect 143816 9036 143868 9042
rect 143816 8978 143868 8984
rect 144184 9036 144236 9042
rect 144184 8978 144236 8984
rect 143172 8968 143224 8974
rect 143172 8910 143224 8916
rect 143264 8832 143316 8838
rect 143264 8774 143316 8780
rect 143356 8832 143408 8838
rect 143356 8774 143408 8780
rect 143276 8362 143304 8774
rect 143368 8498 143396 8774
rect 143356 8492 143408 8498
rect 143356 8434 143408 8440
rect 143264 8356 143316 8362
rect 143264 8298 143316 8304
rect 143828 7342 143856 8978
rect 145104 8628 145156 8634
rect 145104 8570 145156 8576
rect 143908 8492 143960 8498
rect 143908 8434 143960 8440
rect 143920 7818 143948 8434
rect 145012 8288 145064 8294
rect 145012 8230 145064 8236
rect 145024 7954 145052 8230
rect 145116 7954 145144 8570
rect 145208 8362 145236 11206
rect 145392 9625 145420 12200
rect 145378 9616 145434 9625
rect 145378 9551 145434 9560
rect 145656 9376 145708 9382
rect 145656 9318 145708 9324
rect 145668 9178 145696 9318
rect 145656 9172 145708 9178
rect 145656 9114 145708 9120
rect 145196 8356 145248 8362
rect 145196 8298 145248 8304
rect 145012 7948 145064 7954
rect 145012 7890 145064 7896
rect 145104 7948 145156 7954
rect 145104 7890 145156 7896
rect 143908 7812 143960 7818
rect 143908 7754 143960 7760
rect 145024 7546 145052 7890
rect 145380 7812 145432 7818
rect 145380 7754 145432 7760
rect 145012 7540 145064 7546
rect 145012 7482 145064 7488
rect 144368 7404 144420 7410
rect 144368 7346 144420 7352
rect 143816 7336 143868 7342
rect 143816 7278 143868 7284
rect 142896 6928 142948 6934
rect 142896 6870 142948 6876
rect 142896 6792 142948 6798
rect 142896 6734 142948 6740
rect 141792 6384 141844 6390
rect 141792 6326 141844 6332
rect 142804 6384 142856 6390
rect 142804 6326 142856 6332
rect 141273 6012 141569 6032
rect 141329 6010 141353 6012
rect 141409 6010 141433 6012
rect 141489 6010 141513 6012
rect 141351 5958 141353 6010
rect 141415 5958 141427 6010
rect 141489 5958 141491 6010
rect 141329 5956 141353 5958
rect 141409 5956 141433 5958
rect 141489 5956 141513 5958
rect 141273 5936 141569 5956
rect 141273 4924 141569 4944
rect 141329 4922 141353 4924
rect 141409 4922 141433 4924
rect 141489 4922 141513 4924
rect 141351 4870 141353 4922
rect 141415 4870 141427 4922
rect 141489 4870 141491 4922
rect 141329 4868 141353 4870
rect 141409 4868 141433 4870
rect 141489 4868 141513 4870
rect 141273 4848 141569 4868
rect 138664 4208 138716 4214
rect 138664 4150 138716 4156
rect 137100 3528 137152 3534
rect 137100 3470 137152 3476
rect 136640 3052 136692 3058
rect 136640 2994 136692 3000
rect 136824 3052 136876 3058
rect 136824 2994 136876 3000
rect 135996 2440 136048 2446
rect 135996 2382 136048 2388
rect 136652 2310 136680 2994
rect 136732 2848 136784 2854
rect 136732 2790 136784 2796
rect 136640 2304 136692 2310
rect 136640 2246 136692 2252
rect 136652 1850 136680 2246
rect 136376 1822 136680 1850
rect 135904 1760 135956 1766
rect 135904 1702 135956 1708
rect 135916 1562 135944 1702
rect 135904 1556 135956 1562
rect 135904 1498 135956 1504
rect 135352 1420 135404 1426
rect 135352 1362 135404 1368
rect 135444 1420 135496 1426
rect 135444 1362 135496 1368
rect 136088 1216 136140 1222
rect 136088 1158 136140 1164
rect 136100 1018 136128 1158
rect 135628 1012 135680 1018
rect 135628 954 135680 960
rect 136088 1012 136140 1018
rect 136088 954 136140 960
rect 135640 800 135668 954
rect 135994 912 136050 921
rect 135994 847 136050 856
rect 136008 800 136036 847
rect 136376 800 136404 1822
rect 136744 1714 136772 2790
rect 136652 1686 136772 1714
rect 136652 1358 136680 1686
rect 136836 1442 136864 2994
rect 136916 2848 136968 2854
rect 136916 2790 136968 2796
rect 136744 1414 136864 1442
rect 136640 1352 136692 1358
rect 136640 1294 136692 1300
rect 136744 800 136772 1414
rect 136928 882 136956 2790
rect 136916 876 136968 882
rect 136916 818 136968 824
rect 137112 800 137140 3470
rect 137284 3392 137336 3398
rect 137284 3334 137336 3340
rect 137296 1902 137324 3334
rect 138572 3188 138624 3194
rect 138572 3130 138624 3136
rect 138020 3052 138072 3058
rect 138020 2994 138072 3000
rect 137468 2440 137520 2446
rect 137468 2382 137520 2388
rect 137284 1896 137336 1902
rect 137284 1838 137336 1844
rect 137480 800 137508 2382
rect 138032 2378 138060 2994
rect 138020 2372 138072 2378
rect 138020 2314 138072 2320
rect 137652 2304 137704 2310
rect 137652 2246 137704 2252
rect 137560 1896 137612 1902
rect 137560 1838 137612 1844
rect 137572 1562 137600 1838
rect 137560 1556 137612 1562
rect 137560 1498 137612 1504
rect 137664 882 137692 2246
rect 137836 1760 137888 1766
rect 137836 1702 137888 1708
rect 137652 876 137704 882
rect 137652 818 137704 824
rect 137848 800 137876 1702
rect 138216 836 138336 864
rect 138216 800 138244 836
rect 134064 750 134116 756
rect 133984 649 134012 750
rect 133970 640 134026 649
rect 133970 575 134026 584
rect 134076 134 134104 750
rect 134064 128 134116 134
rect 134064 70 134116 76
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137744 740 137796 746
rect 137744 682 137796 688
rect 137756 474 137784 682
rect 137744 468 137796 474
rect 137744 410 137796 416
rect 137834 0 137890 800
rect 137928 740 137980 746
rect 137928 682 137980 688
rect 137940 649 137968 682
rect 137926 640 137982 649
rect 137926 575 137982 584
rect 138202 0 138258 800
rect 138308 474 138336 836
rect 138584 800 138612 3130
rect 138676 2446 138704 4150
rect 141273 3836 141569 3856
rect 141329 3834 141353 3836
rect 141409 3834 141433 3836
rect 141489 3834 141513 3836
rect 141351 3782 141353 3834
rect 141415 3782 141427 3834
rect 141489 3782 141491 3834
rect 141329 3780 141353 3782
rect 141409 3780 141433 3782
rect 141489 3780 141513 3782
rect 141273 3760 141569 3780
rect 139952 3664 140004 3670
rect 139952 3606 140004 3612
rect 138756 3392 138808 3398
rect 138756 3334 138808 3340
rect 138664 2440 138716 2446
rect 138664 2382 138716 2388
rect 138664 2100 138716 2106
rect 138664 2042 138716 2048
rect 138676 1426 138704 2042
rect 138768 1970 138796 3334
rect 139860 3052 139912 3058
rect 139860 2994 139912 3000
rect 139400 2984 139452 2990
rect 139400 2926 139452 2932
rect 139308 2440 139360 2446
rect 139308 2382 139360 2388
rect 139320 2038 139348 2382
rect 139412 2106 139440 2926
rect 139676 2916 139728 2922
rect 139676 2858 139728 2864
rect 139584 2440 139636 2446
rect 139584 2382 139636 2388
rect 139596 2106 139624 2382
rect 139400 2100 139452 2106
rect 139400 2042 139452 2048
rect 139584 2100 139636 2106
rect 139584 2042 139636 2048
rect 138940 2032 138992 2038
rect 138940 1974 138992 1980
rect 139308 2032 139360 2038
rect 139308 1974 139360 1980
rect 138756 1964 138808 1970
rect 138756 1906 138808 1912
rect 138768 1562 138796 1906
rect 138756 1556 138808 1562
rect 138756 1498 138808 1504
rect 138664 1420 138716 1426
rect 138664 1362 138716 1368
rect 138952 800 138980 1974
rect 139492 1964 139544 1970
rect 139492 1906 139544 1912
rect 139504 1766 139532 1906
rect 139492 1760 139544 1766
rect 139492 1702 139544 1708
rect 139688 1358 139716 2858
rect 139872 1494 139900 2994
rect 139860 1488 139912 1494
rect 139860 1430 139912 1436
rect 139964 1426 139992 3606
rect 141148 2984 141200 2990
rect 141148 2926 141200 2932
rect 140964 2848 141016 2854
rect 140964 2790 141016 2796
rect 140872 2372 140924 2378
rect 140872 2314 140924 2320
rect 140780 2304 140832 2310
rect 140780 2246 140832 2252
rect 139952 1420 140004 1426
rect 139952 1362 140004 1368
rect 139676 1352 139728 1358
rect 139676 1294 139728 1300
rect 140044 1284 140096 1290
rect 140044 1226 140096 1232
rect 139676 1216 139728 1222
rect 139136 1142 139348 1170
rect 139676 1158 139728 1164
rect 138296 468 138348 474
rect 138296 410 138348 416
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139136 134 139164 1142
rect 139216 1012 139268 1018
rect 139216 954 139268 960
rect 139228 814 139256 954
rect 139216 808 139268 814
rect 139320 800 139348 1142
rect 139688 800 139716 1158
rect 140056 800 140084 1226
rect 140792 1018 140820 2246
rect 140780 1012 140832 1018
rect 140780 954 140832 960
rect 140884 898 140912 2314
rect 140976 1290 141004 2790
rect 141160 2106 141188 2926
rect 142620 2916 142672 2922
rect 142620 2858 142672 2864
rect 142252 2848 142304 2854
rect 142252 2790 142304 2796
rect 141273 2748 141569 2768
rect 141329 2746 141353 2748
rect 141409 2746 141433 2748
rect 141489 2746 141513 2748
rect 141351 2694 141353 2746
rect 141415 2694 141427 2746
rect 141489 2694 141491 2746
rect 141329 2692 141353 2694
rect 141409 2692 141433 2694
rect 141489 2692 141513 2694
rect 141273 2672 141569 2692
rect 141148 2100 141200 2106
rect 141148 2042 141200 2048
rect 141056 1760 141108 1766
rect 141056 1702 141108 1708
rect 140964 1284 141016 1290
rect 140964 1226 141016 1232
rect 141068 1018 141096 1702
rect 141160 1426 141188 2042
rect 141608 1964 141660 1970
rect 141608 1906 141660 1912
rect 141273 1660 141569 1680
rect 141329 1658 141353 1660
rect 141409 1658 141433 1660
rect 141489 1658 141513 1660
rect 141351 1606 141353 1658
rect 141415 1606 141427 1658
rect 141489 1606 141491 1658
rect 141329 1604 141353 1606
rect 141409 1604 141433 1606
rect 141489 1604 141513 1606
rect 141273 1584 141569 1604
rect 141148 1420 141200 1426
rect 141148 1362 141200 1368
rect 141148 1284 141200 1290
rect 141148 1226 141200 1232
rect 141056 1012 141108 1018
rect 141056 954 141108 960
rect 140792 870 140912 898
rect 141068 882 141096 954
rect 141056 876 141108 882
rect 140332 836 140452 864
rect 139216 750 139268 756
rect 139124 128 139176 134
rect 139124 70 139176 76
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140332 406 140360 836
rect 140424 800 140452 836
rect 140792 800 140820 870
rect 141056 818 141108 824
rect 140872 808 140924 814
rect 140320 400 140372 406
rect 140320 342 140372 348
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141160 800 141188 1226
rect 141620 1204 141648 1906
rect 141528 1176 141648 1204
rect 141528 800 141556 1176
rect 141896 882 142200 898
rect 141896 876 142212 882
rect 141896 870 142160 876
rect 141896 800 141924 870
rect 142160 818 142212 824
rect 142264 800 142292 2790
rect 142632 800 142660 2858
rect 142908 2514 142936 6734
rect 144380 6662 144408 7346
rect 144368 6656 144420 6662
rect 144368 6598 144420 6604
rect 145196 6656 145248 6662
rect 145196 6598 145248 6604
rect 144092 4004 144144 4010
rect 144092 3946 144144 3952
rect 143356 3732 143408 3738
rect 143356 3674 143408 3680
rect 142988 3460 143040 3466
rect 142988 3402 143040 3408
rect 142896 2508 142948 2514
rect 142896 2450 142948 2456
rect 143000 800 143028 3402
rect 143172 2984 143224 2990
rect 143172 2926 143224 2932
rect 143184 1902 143212 2926
rect 143172 1896 143224 1902
rect 143172 1838 143224 1844
rect 143184 1562 143212 1838
rect 143172 1556 143224 1562
rect 143172 1498 143224 1504
rect 143172 1352 143224 1358
rect 143172 1294 143224 1300
rect 143184 1018 143212 1294
rect 143172 1012 143224 1018
rect 143172 954 143224 960
rect 143368 800 143396 3674
rect 143724 2984 143776 2990
rect 143724 2926 143776 2932
rect 143736 800 143764 2926
rect 144000 1216 144052 1222
rect 144000 1158 144052 1164
rect 140872 750 140924 756
rect 140884 474 140912 750
rect 140872 468 140924 474
rect 140872 410 140924 416
rect 141146 0 141202 800
rect 141514 592 141570 800
rect 141273 572 141570 592
rect 141329 570 141353 572
rect 141409 570 141433 572
rect 141489 570 141513 572
rect 141351 518 141353 570
rect 141415 518 141427 570
rect 141489 518 141491 570
rect 141329 516 141353 518
rect 141409 516 141433 518
rect 141489 516 141513 518
rect 141569 516 141570 572
rect 141273 496 141570 516
rect 141514 0 141570 496
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 144012 678 144040 1158
rect 144104 800 144132 3946
rect 144736 3596 144788 3602
rect 144736 3538 144788 3544
rect 144460 3120 144512 3126
rect 144460 3062 144512 3068
rect 144276 1964 144328 1970
rect 144276 1906 144328 1912
rect 144288 1222 144316 1906
rect 144276 1216 144328 1222
rect 144276 1158 144328 1164
rect 144472 800 144500 3062
rect 144748 1850 144776 3538
rect 144828 3392 144880 3398
rect 144828 3334 144880 3340
rect 144840 2038 144868 3334
rect 144920 3188 144972 3194
rect 144920 3130 144972 3136
rect 144828 2032 144880 2038
rect 144828 1974 144880 1980
rect 144748 1822 144868 1850
rect 144840 800 144868 1822
rect 144932 1358 144960 3130
rect 145208 2514 145236 6598
rect 145392 3194 145420 7754
rect 145760 6322 145788 12200
rect 145932 9512 145984 9518
rect 145932 9454 145984 9460
rect 145944 9178 145972 9454
rect 146128 9178 146156 12200
rect 146496 11778 146524 12200
rect 146760 12164 146812 12170
rect 146760 12106 146812 12112
rect 146496 11750 146616 11778
rect 146772 11762 146800 12106
rect 146484 11688 146536 11694
rect 146484 11630 146536 11636
rect 146496 11218 146524 11630
rect 146484 11212 146536 11218
rect 146484 11154 146536 11160
rect 145932 9172 145984 9178
rect 145932 9114 145984 9120
rect 146116 9172 146168 9178
rect 146116 9114 146168 9120
rect 146024 8968 146076 8974
rect 146024 8910 146076 8916
rect 145840 8900 145892 8906
rect 145840 8842 145892 8848
rect 145748 6316 145800 6322
rect 145748 6258 145800 6264
rect 145852 5370 145880 8842
rect 145840 5364 145892 5370
rect 145840 5306 145892 5312
rect 146036 3670 146064 8910
rect 146588 8906 146616 11750
rect 146760 11756 146812 11762
rect 146760 11698 146812 11704
rect 146864 10742 146892 12200
rect 146944 11552 146996 11558
rect 146944 11494 146996 11500
rect 146956 11150 146984 11494
rect 146944 11144 146996 11150
rect 146944 11086 146996 11092
rect 146852 10736 146904 10742
rect 146852 10678 146904 10684
rect 146944 10600 146996 10606
rect 146944 10542 146996 10548
rect 146956 9926 146984 10542
rect 147232 10198 147260 12200
rect 147496 11212 147548 11218
rect 147496 11154 147548 11160
rect 147220 10192 147272 10198
rect 147220 10134 147272 10140
rect 146668 9920 146720 9926
rect 146668 9862 146720 9868
rect 146944 9920 146996 9926
rect 146944 9862 146996 9868
rect 147128 9920 147180 9926
rect 147128 9862 147180 9868
rect 146576 8900 146628 8906
rect 146576 8842 146628 8848
rect 146300 8832 146352 8838
rect 146206 8800 146262 8809
rect 146300 8774 146352 8780
rect 146206 8735 146262 8744
rect 146220 8498 146248 8735
rect 146312 8634 146340 8774
rect 146300 8628 146352 8634
rect 146300 8570 146352 8576
rect 146208 8492 146260 8498
rect 146208 8434 146260 8440
rect 146392 8492 146444 8498
rect 146392 8434 146444 8440
rect 146404 8090 146432 8434
rect 146392 8084 146444 8090
rect 146392 8026 146444 8032
rect 146392 7880 146444 7886
rect 146392 7822 146444 7828
rect 146300 5228 146352 5234
rect 146300 5170 146352 5176
rect 146312 4554 146340 5170
rect 146300 4548 146352 4554
rect 146300 4490 146352 4496
rect 146024 3664 146076 3670
rect 146024 3606 146076 3612
rect 145380 3188 145432 3194
rect 145380 3130 145432 3136
rect 145564 3052 145616 3058
rect 145564 2994 145616 3000
rect 145196 2508 145248 2514
rect 145196 2450 145248 2456
rect 145576 2310 145604 2994
rect 145748 2848 145800 2854
rect 145748 2790 145800 2796
rect 145196 2304 145248 2310
rect 145196 2246 145248 2252
rect 145564 2304 145616 2310
rect 145564 2246 145616 2252
rect 144920 1352 144972 1358
rect 144920 1294 144972 1300
rect 145208 800 145236 2246
rect 145576 800 145604 2246
rect 145760 1358 145788 2790
rect 146300 2440 146352 2446
rect 146300 2382 146352 2388
rect 145932 2304 145984 2310
rect 145932 2246 145984 2252
rect 145748 1352 145800 1358
rect 145748 1294 145800 1300
rect 145944 800 145972 2246
rect 146024 1216 146076 1222
rect 146024 1158 146076 1164
rect 146036 882 146064 1158
rect 146024 876 146076 882
rect 146024 818 146076 824
rect 146312 800 146340 2382
rect 146404 2106 146432 7822
rect 146484 7744 146536 7750
rect 146484 7686 146536 7692
rect 146496 2514 146524 7686
rect 146680 4826 146708 9862
rect 146850 8936 146906 8945
rect 146850 8871 146906 8880
rect 146864 8566 146892 8871
rect 146852 8560 146904 8566
rect 146852 8502 146904 8508
rect 146956 6866 146984 9862
rect 147036 8084 147088 8090
rect 147036 8026 147088 8032
rect 147048 7546 147076 8026
rect 147140 7954 147168 9862
rect 147508 9654 147536 11154
rect 147600 10470 147628 12200
rect 147864 10668 147916 10674
rect 147864 10610 147916 10616
rect 147588 10464 147640 10470
rect 147588 10406 147640 10412
rect 147876 9994 147904 10610
rect 147864 9988 147916 9994
rect 147864 9930 147916 9936
rect 147496 9648 147548 9654
rect 147496 9590 147548 9596
rect 147772 9648 147824 9654
rect 147772 9590 147824 9596
rect 147784 9110 147812 9590
rect 147968 9110 147996 12200
rect 148336 10810 148364 12200
rect 148324 10804 148376 10810
rect 148324 10746 148376 10752
rect 148140 9920 148192 9926
rect 148140 9862 148192 9868
rect 148152 9586 148180 9862
rect 148232 9716 148284 9722
rect 148232 9658 148284 9664
rect 148048 9580 148100 9586
rect 148048 9522 148100 9528
rect 148140 9580 148192 9586
rect 148140 9522 148192 9528
rect 148060 9466 148088 9522
rect 148244 9466 148272 9658
rect 148704 9602 148732 12200
rect 149072 12170 149100 12200
rect 149060 12164 149112 12170
rect 149060 12106 149112 12112
rect 148784 10600 148836 10606
rect 148784 10542 148836 10548
rect 148796 9994 148824 10542
rect 148784 9988 148836 9994
rect 148784 9930 148836 9936
rect 148796 9722 148824 9930
rect 148784 9716 148836 9722
rect 148784 9658 148836 9664
rect 148612 9574 148732 9602
rect 148784 9580 148836 9586
rect 148612 9518 148640 9574
rect 148784 9522 148836 9528
rect 148060 9438 148272 9466
rect 148600 9512 148652 9518
rect 148600 9454 148652 9460
rect 147772 9104 147824 9110
rect 147772 9046 147824 9052
rect 147956 9104 148008 9110
rect 147956 9046 148008 9052
rect 147772 8492 147824 8498
rect 147772 8434 147824 8440
rect 147128 7948 147180 7954
rect 147128 7890 147180 7896
rect 147140 7546 147168 7890
rect 147036 7540 147088 7546
rect 147036 7482 147088 7488
rect 147128 7540 147180 7546
rect 147128 7482 147180 7488
rect 146944 6860 146996 6866
rect 146944 6802 146996 6808
rect 146668 4820 146720 4826
rect 146668 4762 146720 4768
rect 147404 4548 147456 4554
rect 147404 4490 147456 4496
rect 146484 2508 146536 2514
rect 146484 2450 146536 2456
rect 147036 2440 147088 2446
rect 147036 2382 147088 2388
rect 146392 2100 146444 2106
rect 146392 2042 146444 2048
rect 146668 1964 146720 1970
rect 146668 1906 146720 1912
rect 146680 1222 146708 1906
rect 146668 1216 146720 1222
rect 146668 1158 146720 1164
rect 146680 800 146708 1158
rect 147048 800 147076 2382
rect 147416 800 147444 4490
rect 147784 2514 147812 8434
rect 148048 7336 148100 7342
rect 148048 7278 148100 7284
rect 148060 6866 148088 7278
rect 148048 6860 148100 6866
rect 148048 6802 148100 6808
rect 148244 4146 148272 9438
rect 148796 9042 148824 9522
rect 149336 9512 149388 9518
rect 149336 9454 149388 9460
rect 149348 9042 149376 9454
rect 148784 9036 148836 9042
rect 148784 8978 148836 8984
rect 149336 9036 149388 9042
rect 149336 8978 149388 8984
rect 149152 8832 149204 8838
rect 149152 8774 149204 8780
rect 148322 7440 148378 7449
rect 148322 7375 148378 7384
rect 148336 7177 148364 7375
rect 148322 7168 148378 7177
rect 148322 7103 148378 7112
rect 148416 6248 148468 6254
rect 148416 6190 148468 6196
rect 148428 5914 148456 6190
rect 148876 6180 148928 6186
rect 148876 6122 148928 6128
rect 148416 5908 148468 5914
rect 148416 5850 148468 5856
rect 148888 5846 148916 6122
rect 148876 5840 148928 5846
rect 148876 5782 148928 5788
rect 148232 4140 148284 4146
rect 148232 4082 148284 4088
rect 149060 4072 149112 4078
rect 149060 4014 149112 4020
rect 148140 3528 148192 3534
rect 148140 3470 148192 3476
rect 147772 2508 147824 2514
rect 147772 2450 147824 2456
rect 147772 2372 147824 2378
rect 147772 2314 147824 2320
rect 147784 800 147812 2314
rect 147864 1896 147916 1902
rect 147864 1838 147916 1844
rect 147876 1426 147904 1838
rect 147864 1420 147916 1426
rect 147864 1362 147916 1368
rect 148152 800 148180 3470
rect 149072 3398 149100 4014
rect 149060 3392 149112 3398
rect 149060 3334 149112 3340
rect 149072 3194 149100 3334
rect 149060 3188 149112 3194
rect 149060 3130 149112 3136
rect 149060 3052 149112 3058
rect 149060 2994 149112 3000
rect 149072 2310 149100 2994
rect 149164 2854 149192 8774
rect 149244 8424 149296 8430
rect 149244 8366 149296 8372
rect 149256 7546 149284 8366
rect 149440 8022 149468 12200
rect 149808 10538 149836 12200
rect 149796 10532 149848 10538
rect 149796 10474 149848 10480
rect 149980 9920 150032 9926
rect 149980 9862 150032 9868
rect 149520 9444 149572 9450
rect 149520 9386 149572 9392
rect 149428 8016 149480 8022
rect 149428 7958 149480 7964
rect 149428 7744 149480 7750
rect 149428 7686 149480 7692
rect 149244 7540 149296 7546
rect 149244 7482 149296 7488
rect 149336 7404 149388 7410
rect 149336 7346 149388 7352
rect 149348 6662 149376 7346
rect 149336 6656 149388 6662
rect 149336 6598 149388 6604
rect 149152 2848 149204 2854
rect 149152 2790 149204 2796
rect 149244 2848 149296 2854
rect 149244 2790 149296 2796
rect 149060 2304 149112 2310
rect 149060 2246 149112 2252
rect 149152 1964 149204 1970
rect 149152 1906 149204 1912
rect 148508 1420 148560 1426
rect 148508 1362 148560 1368
rect 148520 800 148548 1362
rect 149060 1352 149112 1358
rect 148888 1300 149060 1306
rect 148888 1294 149112 1300
rect 148888 1278 149100 1294
rect 149164 1290 149192 1906
rect 149152 1284 149204 1290
rect 148888 800 148916 1278
rect 149152 1226 149204 1232
rect 149256 800 149284 2790
rect 149348 2514 149376 6598
rect 149440 2514 149468 7686
rect 149532 7342 149560 9386
rect 149520 7336 149572 7342
rect 149520 7278 149572 7284
rect 149612 4548 149664 4554
rect 149612 4490 149664 4496
rect 149336 2508 149388 2514
rect 149336 2450 149388 2456
rect 149428 2508 149480 2514
rect 149428 2450 149480 2456
rect 149624 800 149652 4490
rect 149992 3670 150020 9862
rect 150176 9738 150204 12200
rect 150440 11756 150492 11762
rect 150440 11698 150492 11704
rect 150452 11286 150480 11698
rect 150440 11280 150492 11286
rect 150440 11222 150492 11228
rect 150176 9710 150296 9738
rect 150164 9580 150216 9586
rect 150164 9522 150216 9528
rect 150072 6316 150124 6322
rect 150072 6258 150124 6264
rect 150084 5574 150112 6258
rect 150072 5568 150124 5574
rect 150072 5510 150124 5516
rect 149980 3664 150032 3670
rect 149980 3606 150032 3612
rect 149888 2304 149940 2310
rect 149888 2246 149940 2252
rect 149900 2088 149928 2246
rect 149900 2060 150020 2088
rect 149992 800 150020 2060
rect 150084 1358 150112 5510
rect 150176 4826 150204 9522
rect 150268 6186 150296 9710
rect 150544 8430 150572 12200
rect 150716 11076 150768 11082
rect 150716 11018 150768 11024
rect 150728 8809 150756 11018
rect 150912 9450 150940 12200
rect 150992 11552 151044 11558
rect 150992 11494 151044 11500
rect 151004 11218 151032 11494
rect 150992 11212 151044 11218
rect 150992 11154 151044 11160
rect 151280 10198 151308 12200
rect 151648 11778 151676 12200
rect 151452 11756 151504 11762
rect 151648 11750 151768 11778
rect 151452 11698 151504 11704
rect 151464 11082 151492 11698
rect 151636 11620 151688 11626
rect 151636 11562 151688 11568
rect 151544 11212 151596 11218
rect 151544 11154 151596 11160
rect 151452 11076 151504 11082
rect 151452 11018 151504 11024
rect 151268 10192 151320 10198
rect 151268 10134 151320 10140
rect 151084 9920 151136 9926
rect 151084 9862 151136 9868
rect 150900 9444 150952 9450
rect 150900 9386 150952 9392
rect 150714 8800 150770 8809
rect 150714 8735 150770 8744
rect 150532 8424 150584 8430
rect 150532 8366 150584 8372
rect 150900 8356 150952 8362
rect 150900 8298 150952 8304
rect 150912 7954 150940 8298
rect 150900 7948 150952 7954
rect 150900 7890 150952 7896
rect 150440 7880 150492 7886
rect 150440 7822 150492 7828
rect 150992 7880 151044 7886
rect 150992 7822 151044 7828
rect 150452 7546 150480 7822
rect 150440 7540 150492 7546
rect 150440 7482 150492 7488
rect 150808 6792 150860 6798
rect 150808 6734 150860 6740
rect 150820 6390 150848 6734
rect 150808 6384 150860 6390
rect 150808 6326 150860 6332
rect 150256 6180 150308 6186
rect 150256 6122 150308 6128
rect 150164 4820 150216 4826
rect 150164 4762 150216 4768
rect 150164 4140 150216 4146
rect 150164 4082 150216 4088
rect 150176 3670 150204 4082
rect 150164 3664 150216 3670
rect 150164 3606 150216 3612
rect 150348 3188 150400 3194
rect 150348 3130 150400 3136
rect 150256 1964 150308 1970
rect 150256 1906 150308 1912
rect 150268 1426 150296 1906
rect 150256 1420 150308 1426
rect 150256 1362 150308 1368
rect 150072 1352 150124 1358
rect 150072 1294 150124 1300
rect 150360 800 150388 3130
rect 150900 2848 150952 2854
rect 150900 2790 150952 2796
rect 150912 2446 150940 2790
rect 150900 2440 150952 2446
rect 150900 2382 150952 2388
rect 150716 2304 150768 2310
rect 150716 2246 150768 2252
rect 150728 800 150756 2246
rect 151004 2106 151032 7822
rect 151096 3942 151124 9862
rect 151556 9382 151584 11154
rect 151648 11150 151676 11562
rect 151636 11144 151688 11150
rect 151636 11086 151688 11092
rect 151636 10668 151688 10674
rect 151636 10610 151688 10616
rect 151648 9926 151676 10610
rect 151636 9920 151688 9926
rect 151636 9862 151688 9868
rect 151544 9376 151596 9382
rect 151544 9318 151596 9324
rect 151176 8492 151228 8498
rect 151176 8434 151228 8440
rect 151188 8294 151216 8434
rect 151176 8288 151228 8294
rect 151176 8230 151228 8236
rect 151084 3936 151136 3942
rect 151084 3878 151136 3884
rect 151084 3460 151136 3466
rect 151084 3402 151136 3408
rect 150992 2100 151044 2106
rect 150992 2042 151044 2048
rect 151096 800 151124 3402
rect 151188 2378 151216 8230
rect 151648 3466 151676 9862
rect 151740 9382 151768 11750
rect 151820 11076 151872 11082
rect 151820 11018 151872 11024
rect 151832 9654 151860 11018
rect 151820 9648 151872 9654
rect 151820 9590 151872 9596
rect 151728 9376 151780 9382
rect 151728 9318 151780 9324
rect 151832 9042 151860 9590
rect 152016 9110 152044 12200
rect 152096 10600 152148 10606
rect 152096 10542 152148 10548
rect 152108 10266 152136 10542
rect 152384 10538 152412 12200
rect 152476 11898 152504 12378
rect 152738 12200 152794 13000
rect 153106 12200 153162 13000
rect 153474 12200 153530 13000
rect 153842 12200 153898 13000
rect 154210 12200 154266 13000
rect 154578 12200 154634 13000
rect 154946 12200 155002 13000
rect 155314 12200 155370 13000
rect 155682 12200 155738 13000
rect 156050 12200 156106 13000
rect 156418 12200 156474 13000
rect 156786 12200 156842 13000
rect 157154 12200 157210 13000
rect 157522 12200 157578 13000
rect 157890 12200 157946 13000
rect 158258 12200 158314 13000
rect 158626 12200 158682 13000
rect 158994 12200 159050 13000
rect 159362 12200 159418 13000
rect 159730 12200 159786 13000
rect 160098 12200 160154 13000
rect 160466 12200 160522 13000
rect 160834 12200 160890 13000
rect 161202 12200 161258 13000
rect 161570 12200 161626 13000
rect 161938 12200 161994 13000
rect 162306 12200 162362 13000
rect 162674 12200 162730 13000
rect 162952 12300 163004 12306
rect 162952 12242 163004 12248
rect 152464 11892 152516 11898
rect 152464 11834 152516 11840
rect 152372 10532 152424 10538
rect 152372 10474 152424 10480
rect 152096 10260 152148 10266
rect 152096 10202 152148 10208
rect 152004 9104 152056 9110
rect 152004 9046 152056 9052
rect 151820 9036 151872 9042
rect 151820 8978 151872 8984
rect 151820 8900 151872 8906
rect 151820 8842 151872 8848
rect 151728 8832 151780 8838
rect 151728 8774 151780 8780
rect 151740 4826 151768 8774
rect 151832 6866 151860 8842
rect 152752 8634 152780 12200
rect 153014 8936 153070 8945
rect 153014 8871 153070 8880
rect 152740 8628 152792 8634
rect 152740 8570 152792 8576
rect 153028 8566 153056 8871
rect 153016 8560 153068 8566
rect 153016 8502 153068 8508
rect 152464 8492 152516 8498
rect 152464 8434 152516 8440
rect 152476 8090 152504 8434
rect 153120 8430 153148 12200
rect 153292 12164 153344 12170
rect 153292 12106 153344 12112
rect 153200 11552 153252 11558
rect 153200 11494 153252 11500
rect 153212 10674 153240 11494
rect 153304 11286 153332 12106
rect 153292 11280 153344 11286
rect 153292 11222 153344 11228
rect 153200 10668 153252 10674
rect 153200 10610 153252 10616
rect 153212 10266 153240 10610
rect 153292 10532 153344 10538
rect 153292 10474 153344 10480
rect 153200 10260 153252 10266
rect 153200 10202 153252 10208
rect 153200 9920 153252 9926
rect 153200 9862 153252 9868
rect 153212 8498 153240 9862
rect 153304 9625 153332 10474
rect 153290 9616 153346 9625
rect 153290 9551 153346 9560
rect 153200 8492 153252 8498
rect 153200 8434 153252 8440
rect 153108 8424 153160 8430
rect 153108 8366 153160 8372
rect 152464 8084 152516 8090
rect 152464 8026 152516 8032
rect 153488 7954 153516 12200
rect 153752 9376 153804 9382
rect 153752 9318 153804 9324
rect 153660 8832 153712 8838
rect 153660 8774 153712 8780
rect 153476 7948 153528 7954
rect 153476 7890 153528 7896
rect 152924 7744 152976 7750
rect 152924 7686 152976 7692
rect 152936 7478 152964 7686
rect 152924 7472 152976 7478
rect 152924 7414 152976 7420
rect 153016 7200 153068 7206
rect 153016 7142 153068 7148
rect 151820 6860 151872 6866
rect 151820 6802 151872 6808
rect 153028 6798 153056 7142
rect 152096 6792 152148 6798
rect 152096 6734 152148 6740
rect 153016 6792 153068 6798
rect 153016 6734 153068 6740
rect 152004 5568 152056 5574
rect 152004 5510 152056 5516
rect 152016 5234 152044 5510
rect 152004 5228 152056 5234
rect 152004 5170 152056 5176
rect 151728 4820 151780 4826
rect 151728 4762 151780 4768
rect 151636 3460 151688 3466
rect 151636 3402 151688 3408
rect 152004 3392 152056 3398
rect 152004 3334 152056 3340
rect 152016 2922 152044 3334
rect 151360 2916 151412 2922
rect 151360 2858 151412 2864
rect 152004 2916 152056 2922
rect 152004 2858 152056 2864
rect 151176 2372 151228 2378
rect 151176 2314 151228 2320
rect 151372 1358 151400 2858
rect 151820 2576 151872 2582
rect 151872 2524 151952 2530
rect 151820 2518 151952 2524
rect 151832 2502 151952 2518
rect 152108 2514 152136 6734
rect 153028 6390 153056 6734
rect 153016 6384 153068 6390
rect 153016 6326 153068 6332
rect 153476 6316 153528 6322
rect 153476 6258 153528 6264
rect 153384 6248 153436 6254
rect 153384 6190 153436 6196
rect 153396 5914 153424 6190
rect 153384 5908 153436 5914
rect 153384 5850 153436 5856
rect 153488 5710 153516 6258
rect 153476 5704 153528 5710
rect 153476 5646 153528 5652
rect 152924 5228 152976 5234
rect 152924 5170 152976 5176
rect 152936 4826 152964 5170
rect 152924 4820 152976 4826
rect 152924 4762 152976 4768
rect 152188 4684 152240 4690
rect 152188 4626 152240 4632
rect 151820 2440 151872 2446
rect 151820 2382 151872 2388
rect 151360 1352 151412 1358
rect 151360 1294 151412 1300
rect 151452 1352 151504 1358
rect 151452 1294 151504 1300
rect 151464 800 151492 1294
rect 151728 1216 151780 1222
rect 151728 1158 151780 1164
rect 151740 882 151768 1158
rect 151728 876 151780 882
rect 151728 818 151780 824
rect 151832 800 151860 2382
rect 151924 1494 151952 2502
rect 152096 2508 152148 2514
rect 152096 2450 152148 2456
rect 151912 1488 151964 1494
rect 151912 1430 151964 1436
rect 152200 800 152228 4626
rect 153292 4480 153344 4486
rect 153292 4422 153344 4428
rect 152556 3664 152608 3670
rect 152556 3606 152608 3612
rect 152568 800 152596 3606
rect 152648 1964 152700 1970
rect 152648 1906 152700 1912
rect 152660 1358 152688 1906
rect 152648 1352 152700 1358
rect 152648 1294 152700 1300
rect 152924 1216 152976 1222
rect 152924 1158 152976 1164
rect 152936 800 152964 1158
rect 153304 800 153332 4422
rect 153488 4282 153516 5646
rect 153672 4826 153700 8774
rect 153764 6934 153792 9318
rect 153856 9042 153884 12200
rect 154120 11076 154172 11082
rect 154120 11018 154172 11024
rect 154132 9586 154160 11018
rect 154120 9580 154172 9586
rect 154120 9522 154172 9528
rect 153844 9036 153896 9042
rect 153844 8978 153896 8984
rect 153844 8832 153896 8838
rect 153844 8774 153896 8780
rect 153752 6928 153804 6934
rect 153752 6870 153804 6876
rect 153752 6792 153804 6798
rect 153752 6734 153804 6740
rect 153660 4820 153712 4826
rect 153660 4762 153712 4768
rect 153476 4276 153528 4282
rect 153476 4218 153528 4224
rect 153568 3392 153620 3398
rect 153568 3334 153620 3340
rect 153580 1034 153608 3334
rect 153764 2106 153792 6734
rect 153856 5778 153884 8774
rect 153936 8628 153988 8634
rect 153936 8570 153988 8576
rect 153844 5772 153896 5778
rect 153844 5714 153896 5720
rect 153948 5166 153976 8570
rect 154224 8566 154252 12200
rect 154488 11756 154540 11762
rect 154488 11698 154540 11704
rect 154500 11082 154528 11698
rect 154488 11076 154540 11082
rect 154488 11018 154540 11024
rect 154212 8560 154264 8566
rect 154212 8502 154264 8508
rect 154304 8356 154356 8362
rect 154304 8298 154356 8304
rect 153936 5160 153988 5166
rect 153936 5102 153988 5108
rect 154316 3194 154344 8298
rect 154592 6474 154620 12200
rect 154960 10010 154988 12200
rect 155328 11098 155356 12200
rect 155328 11070 155448 11098
rect 155316 11008 155368 11014
rect 155316 10950 155368 10956
rect 155328 10606 155356 10950
rect 155316 10600 155368 10606
rect 155316 10542 155368 10548
rect 155328 10266 155356 10542
rect 155316 10260 155368 10266
rect 155316 10202 155368 10208
rect 154960 9982 155080 10010
rect 154856 9920 154908 9926
rect 154856 9862 154908 9868
rect 154948 9920 155000 9926
rect 154948 9862 155000 9868
rect 154868 8498 154896 9862
rect 154960 9586 154988 9862
rect 154948 9580 155000 9586
rect 154948 9522 155000 9528
rect 154960 9178 154988 9522
rect 154948 9172 155000 9178
rect 154948 9114 155000 9120
rect 154856 8492 154908 8498
rect 154856 8434 154908 8440
rect 154868 8090 154896 8434
rect 155052 8362 155080 9982
rect 155316 8560 155368 8566
rect 155316 8502 155368 8508
rect 155040 8356 155092 8362
rect 155040 8298 155092 8304
rect 154856 8084 154908 8090
rect 154856 8026 154908 8032
rect 154948 7744 155000 7750
rect 154948 7686 155000 7692
rect 154592 6446 154712 6474
rect 154580 6248 154632 6254
rect 154578 6216 154580 6225
rect 154632 6216 154634 6225
rect 154578 6151 154634 6160
rect 154684 5846 154712 6446
rect 154856 6316 154908 6322
rect 154856 6258 154908 6264
rect 154672 5840 154724 5846
rect 154672 5782 154724 5788
rect 154868 5574 154896 6258
rect 154580 5568 154632 5574
rect 154580 5510 154632 5516
rect 154856 5568 154908 5574
rect 154856 5510 154908 5516
rect 154304 3188 154356 3194
rect 154304 3130 154356 3136
rect 154396 3052 154448 3058
rect 154396 2994 154448 3000
rect 154408 2310 154436 2994
rect 154396 2304 154448 2310
rect 154396 2246 154448 2252
rect 153752 2100 153804 2106
rect 153752 2042 153804 2048
rect 153660 1964 153712 1970
rect 153660 1906 153712 1912
rect 153672 1222 153700 1906
rect 153660 1216 153712 1222
rect 153660 1158 153712 1164
rect 154028 1216 154080 1222
rect 154028 1158 154080 1164
rect 153580 1006 153700 1034
rect 153672 800 153700 1006
rect 154040 800 154068 1158
rect 154408 800 154436 2246
rect 154592 2038 154620 5510
rect 154856 5228 154908 5234
rect 154856 5170 154908 5176
rect 154868 4486 154896 5170
rect 154856 4480 154908 4486
rect 154856 4422 154908 4428
rect 154764 2304 154816 2310
rect 154764 2246 154816 2252
rect 154580 2032 154632 2038
rect 154580 1974 154632 1980
rect 154672 1964 154724 1970
rect 154672 1906 154724 1912
rect 154684 1222 154712 1906
rect 154672 1216 154724 1222
rect 154672 1158 154724 1164
rect 154776 800 154804 2246
rect 154868 2106 154896 4422
rect 154960 3194 154988 7686
rect 155328 7342 155356 8502
rect 155420 8430 155448 11070
rect 155696 9518 155724 12200
rect 155960 11552 156012 11558
rect 155960 11494 156012 11500
rect 155972 10674 156000 11494
rect 155960 10668 156012 10674
rect 155960 10610 156012 10616
rect 155972 10266 156000 10610
rect 155960 10260 156012 10266
rect 155960 10202 156012 10208
rect 155684 9512 155736 9518
rect 155684 9454 155736 9460
rect 156064 9042 156092 12200
rect 156144 11688 156196 11694
rect 156144 11630 156196 11636
rect 156156 11354 156184 11630
rect 156144 11348 156196 11354
rect 156144 11290 156196 11296
rect 156144 10600 156196 10606
rect 156144 10542 156196 10548
rect 156156 9110 156184 10542
rect 156236 9580 156288 9586
rect 156236 9522 156288 9528
rect 156248 9382 156276 9522
rect 156236 9376 156288 9382
rect 156236 9318 156288 9324
rect 156144 9104 156196 9110
rect 156144 9046 156196 9052
rect 156052 9036 156104 9042
rect 156052 8978 156104 8984
rect 155960 8968 156012 8974
rect 155960 8910 156012 8916
rect 155408 8424 155460 8430
rect 155408 8366 155460 8372
rect 155868 7404 155920 7410
rect 155868 7346 155920 7352
rect 155224 7336 155276 7342
rect 155224 7278 155276 7284
rect 155316 7336 155368 7342
rect 155316 7278 155368 7284
rect 155236 7002 155264 7278
rect 155224 6996 155276 7002
rect 155224 6938 155276 6944
rect 155880 6662 155908 7346
rect 155500 6656 155552 6662
rect 155500 6598 155552 6604
rect 155868 6656 155920 6662
rect 155868 6598 155920 6604
rect 155512 6225 155540 6598
rect 155498 6216 155554 6225
rect 155498 6151 155554 6160
rect 155776 5568 155828 5574
rect 155776 5510 155828 5516
rect 155316 5160 155368 5166
rect 155316 5102 155368 5108
rect 155328 4690 155356 5102
rect 155316 4684 155368 4690
rect 155316 4626 155368 4632
rect 155132 4548 155184 4554
rect 155132 4490 155184 4496
rect 155040 4140 155092 4146
rect 155040 4082 155092 4088
rect 155052 3466 155080 4082
rect 155040 3460 155092 3466
rect 155040 3402 155092 3408
rect 154948 3188 155000 3194
rect 154948 3130 155000 3136
rect 154856 2100 154908 2106
rect 154856 2042 154908 2048
rect 155144 800 155172 4490
rect 155224 3052 155276 3058
rect 155224 2994 155276 3000
rect 155236 2310 155264 2994
rect 155500 2440 155552 2446
rect 155500 2382 155552 2388
rect 155224 2304 155276 2310
rect 155224 2246 155276 2252
rect 155224 1284 155276 1290
rect 155224 1226 155276 1232
rect 155236 1018 155264 1226
rect 155224 1012 155276 1018
rect 155224 954 155276 960
rect 155512 800 155540 2382
rect 155788 2106 155816 5510
rect 155880 2582 155908 6598
rect 155972 4078 156000 8910
rect 156052 8492 156104 8498
rect 156052 8434 156104 8440
rect 156064 4826 156092 8434
rect 156144 7880 156196 7886
rect 156144 7822 156196 7828
rect 156156 7546 156184 7822
rect 156144 7540 156196 7546
rect 156144 7482 156196 7488
rect 156156 6866 156184 7482
rect 156144 6860 156196 6866
rect 156144 6802 156196 6808
rect 156052 4820 156104 4826
rect 156052 4762 156104 4768
rect 156248 4146 156276 9318
rect 156328 6112 156380 6118
rect 156328 6054 156380 6060
rect 156340 5710 156368 6054
rect 156432 5778 156460 12200
rect 156512 8356 156564 8362
rect 156512 8298 156564 8304
rect 156420 5772 156472 5778
rect 156420 5714 156472 5720
rect 156328 5704 156380 5710
rect 156328 5646 156380 5652
rect 156340 4690 156368 5646
rect 156524 5166 156552 8298
rect 156800 8022 156828 12200
rect 156880 11688 156932 11694
rect 156880 11630 156932 11636
rect 156892 11150 156920 11630
rect 156880 11144 156932 11150
rect 156880 11086 156932 11092
rect 157168 9654 157196 12200
rect 157432 11552 157484 11558
rect 157432 11494 157484 11500
rect 157444 11150 157472 11494
rect 157432 11144 157484 11150
rect 157432 11086 157484 11092
rect 157248 10600 157300 10606
rect 157248 10542 157300 10548
rect 157260 10470 157288 10542
rect 157248 10464 157300 10470
rect 157248 10406 157300 10412
rect 157156 9648 157208 9654
rect 157156 9590 157208 9596
rect 157156 9512 157208 9518
rect 157156 9454 157208 9460
rect 157168 9178 157196 9454
rect 157248 9376 157300 9382
rect 157248 9318 157300 9324
rect 157156 9172 157208 9178
rect 157156 9114 157208 9120
rect 157168 8634 157196 9114
rect 157260 8974 157288 9318
rect 157248 8968 157300 8974
rect 157248 8910 157300 8916
rect 157156 8628 157208 8634
rect 157156 8570 157208 8576
rect 156788 8016 156840 8022
rect 156788 7958 156840 7964
rect 157260 6390 157288 8910
rect 157536 8566 157564 12200
rect 157904 9518 157932 12200
rect 157984 10464 158036 10470
rect 157984 10406 158036 10412
rect 157996 10130 158024 10406
rect 157984 10124 158036 10130
rect 157984 10066 158036 10072
rect 157892 9512 157944 9518
rect 157892 9454 157944 9460
rect 158272 9110 158300 12200
rect 158260 9104 158312 9110
rect 158260 9046 158312 9052
rect 158640 9042 158668 12200
rect 158720 10668 158772 10674
rect 158720 10610 158772 10616
rect 158732 10266 158760 10610
rect 158720 10260 158772 10266
rect 158720 10202 158772 10208
rect 158812 9648 158864 9654
rect 158812 9590 158864 9596
rect 158628 9036 158680 9042
rect 158628 8978 158680 8984
rect 158536 8968 158588 8974
rect 158536 8910 158588 8916
rect 157524 8560 157576 8566
rect 157524 8502 157576 8508
rect 158548 8362 158576 8910
rect 158536 8356 158588 8362
rect 158536 8298 158588 8304
rect 157524 7812 157576 7818
rect 157524 7754 157576 7760
rect 157248 6384 157300 6390
rect 157248 6326 157300 6332
rect 157432 6180 157484 6186
rect 157432 6122 157484 6128
rect 157444 5914 157472 6122
rect 157536 5914 157564 7754
rect 158260 6248 158312 6254
rect 158260 6190 158312 6196
rect 157432 5908 157484 5914
rect 157432 5850 157484 5856
rect 157524 5908 157576 5914
rect 157524 5850 157576 5856
rect 157340 5704 157392 5710
rect 157340 5646 157392 5652
rect 158076 5704 158128 5710
rect 158076 5646 158128 5652
rect 156604 5228 156656 5234
rect 156604 5170 156656 5176
rect 156512 5160 156564 5166
rect 156512 5102 156564 5108
rect 156616 4826 156644 5170
rect 156604 4820 156656 4826
rect 156604 4762 156656 4768
rect 156328 4684 156380 4690
rect 156328 4626 156380 4632
rect 156420 4480 156472 4486
rect 156420 4422 156472 4428
rect 156052 4140 156104 4146
rect 156052 4082 156104 4088
rect 156236 4140 156288 4146
rect 156236 4082 156288 4088
rect 155960 4072 156012 4078
rect 155960 4014 156012 4020
rect 156064 3398 156092 4082
rect 156052 3392 156104 3398
rect 156052 3334 156104 3340
rect 156236 3052 156288 3058
rect 156236 2994 156288 3000
rect 155868 2576 155920 2582
rect 155868 2518 155920 2524
rect 156248 2446 156276 2994
rect 156236 2440 156288 2446
rect 156236 2382 156288 2388
rect 155776 2100 155828 2106
rect 155776 2042 155828 2048
rect 155868 1964 155920 1970
rect 155868 1906 155920 1912
rect 155880 1766 155908 1906
rect 155868 1760 155920 1766
rect 155868 1702 155920 1708
rect 155776 1352 155828 1358
rect 155776 1294 155828 1300
rect 155788 1018 155816 1294
rect 155776 1012 155828 1018
rect 155776 954 155828 960
rect 155880 800 155908 1702
rect 156248 800 156276 2382
rect 156432 864 156460 4422
rect 156616 3194 156644 4762
rect 157248 3460 157300 3466
rect 157248 3402 157300 3408
rect 156972 3392 157024 3398
rect 156972 3334 157024 3340
rect 156604 3188 156656 3194
rect 156604 3130 156656 3136
rect 156696 2984 156748 2990
rect 156696 2926 156748 2932
rect 156708 1970 156736 2926
rect 156696 1964 156748 1970
rect 156696 1906 156748 1912
rect 156880 1760 156932 1766
rect 156880 1702 156932 1708
rect 156786 1456 156842 1465
rect 156786 1391 156788 1400
rect 156840 1391 156842 1400
rect 156788 1362 156840 1368
rect 156892 1358 156920 1702
rect 156880 1352 156932 1358
rect 156880 1294 156932 1300
rect 156432 836 156644 864
rect 156616 800 156644 836
rect 156788 808 156840 814
rect 144000 672 144052 678
rect 144000 614 144052 620
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 151912 740 151964 746
rect 151912 682 151964 688
rect 151924 202 151952 682
rect 151912 196 151964 202
rect 151912 138 151964 144
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156984 800 157012 3334
rect 157260 2428 157288 3402
rect 157352 2582 157380 5646
rect 157340 2576 157392 2582
rect 157340 2518 157392 2524
rect 157260 2400 157380 2428
rect 157352 800 157380 2400
rect 157708 2304 157760 2310
rect 157708 2246 157760 2252
rect 157720 800 157748 2246
rect 158088 800 158116 5646
rect 158272 5234 158300 6190
rect 158260 5228 158312 5234
rect 158260 5170 158312 5176
rect 158272 4826 158300 5170
rect 158260 4820 158312 4826
rect 158260 4762 158312 4768
rect 158548 4146 158576 8298
rect 158720 7880 158772 7886
rect 158720 7822 158772 7828
rect 158732 7546 158760 7822
rect 158720 7540 158772 7546
rect 158720 7482 158772 7488
rect 158824 5166 158852 9590
rect 159008 8498 159036 12200
rect 159272 11008 159324 11014
rect 159272 10950 159324 10956
rect 159284 10674 159312 10950
rect 159272 10668 159324 10674
rect 159272 10610 159324 10616
rect 159376 10130 159404 12200
rect 159548 11620 159600 11626
rect 159548 11562 159600 11568
rect 159560 10674 159588 11562
rect 159548 10668 159600 10674
rect 159548 10610 159600 10616
rect 159560 10266 159588 10610
rect 159548 10260 159600 10266
rect 159548 10202 159600 10208
rect 159364 10124 159416 10130
rect 159364 10066 159416 10072
rect 159548 10056 159600 10062
rect 159548 9998 159600 10004
rect 159272 9580 159324 9586
rect 159272 9522 159324 9528
rect 159284 8838 159312 9522
rect 159560 9382 159588 9998
rect 159548 9376 159600 9382
rect 159548 9318 159600 9324
rect 159272 8832 159324 8838
rect 159272 8774 159324 8780
rect 158996 8492 159048 8498
rect 158996 8434 159048 8440
rect 159284 5914 159312 8774
rect 159364 8560 159416 8566
rect 159364 8502 159416 8508
rect 159376 7954 159404 8502
rect 159456 8424 159508 8430
rect 159456 8366 159508 8372
rect 159364 7948 159416 7954
rect 159364 7890 159416 7896
rect 159468 7546 159496 8366
rect 159744 8362 159772 12200
rect 160112 8566 160140 12200
rect 160376 12096 160428 12102
rect 160376 12038 160428 12044
rect 160388 11762 160416 12038
rect 160192 11756 160244 11762
rect 160192 11698 160244 11704
rect 160376 11756 160428 11762
rect 160376 11698 160428 11704
rect 160204 11354 160232 11698
rect 160192 11348 160244 11354
rect 160192 11290 160244 11296
rect 160480 10554 160508 12200
rect 160480 10526 160600 10554
rect 160468 10464 160520 10470
rect 160468 10406 160520 10412
rect 160480 10130 160508 10406
rect 160572 10130 160600 10526
rect 160468 10124 160520 10130
rect 160468 10066 160520 10072
rect 160560 10124 160612 10130
rect 160560 10066 160612 10072
rect 160480 9654 160508 10066
rect 160468 9648 160520 9654
rect 160468 9590 160520 9596
rect 160468 9512 160520 9518
rect 160468 9454 160520 9460
rect 160284 9376 160336 9382
rect 160284 9318 160336 9324
rect 160100 8560 160152 8566
rect 160100 8502 160152 8508
rect 159732 8356 159784 8362
rect 159732 8298 159784 8304
rect 159732 7880 159784 7886
rect 159732 7822 159784 7828
rect 159456 7540 159508 7546
rect 159456 7482 159508 7488
rect 159468 6458 159496 7482
rect 159456 6452 159508 6458
rect 159456 6394 159508 6400
rect 159272 5908 159324 5914
rect 159272 5850 159324 5856
rect 159180 5704 159232 5710
rect 159180 5646 159232 5652
rect 158812 5160 158864 5166
rect 158812 5102 158864 5108
rect 158536 4140 158588 4146
rect 158536 4082 158588 4088
rect 158720 4072 158772 4078
rect 158720 4014 158772 4020
rect 158168 4004 158220 4010
rect 158168 3946 158220 3952
rect 158180 1970 158208 3946
rect 158732 3466 158760 4014
rect 158720 3460 158772 3466
rect 158720 3402 158772 3408
rect 158260 2984 158312 2990
rect 158260 2926 158312 2932
rect 158168 1964 158220 1970
rect 158168 1906 158220 1912
rect 158180 1562 158208 1906
rect 158168 1556 158220 1562
rect 158168 1498 158220 1504
rect 158272 1018 158300 2926
rect 158812 2916 158864 2922
rect 158812 2858 158864 2864
rect 158444 2440 158496 2446
rect 158444 2382 158496 2388
rect 158352 1760 158404 1766
rect 158352 1702 158404 1708
rect 158364 1018 158392 1702
rect 158260 1012 158312 1018
rect 158260 954 158312 960
rect 158352 1012 158404 1018
rect 158352 954 158404 960
rect 158456 800 158484 2382
rect 158720 1760 158772 1766
rect 158720 1702 158772 1708
rect 158732 1358 158760 1702
rect 158720 1352 158772 1358
rect 158720 1294 158772 1300
rect 158824 800 158852 2858
rect 159192 800 159220 5646
rect 159548 5228 159600 5234
rect 159548 5170 159600 5176
rect 159560 4486 159588 5170
rect 159548 4480 159600 4486
rect 159548 4422 159600 4428
rect 159456 3392 159508 3398
rect 159456 3334 159508 3340
rect 159362 2544 159418 2553
rect 159362 2479 159418 2488
rect 159376 2446 159404 2479
rect 159364 2440 159416 2446
rect 159364 2382 159416 2388
rect 159468 882 159496 3334
rect 159560 2582 159588 4422
rect 159744 3194 159772 7822
rect 159916 7336 159968 7342
rect 159916 7278 159968 7284
rect 159928 6866 159956 7278
rect 159916 6860 159968 6866
rect 159916 6802 159968 6808
rect 160296 4078 160324 9318
rect 160480 9042 160508 9454
rect 160848 9382 160876 12200
rect 160836 9376 160888 9382
rect 160836 9318 160888 9324
rect 160836 9104 160888 9110
rect 160836 9046 160888 9052
rect 160468 9036 160520 9042
rect 160468 8978 160520 8984
rect 160744 8492 160796 8498
rect 160744 8434 160796 8440
rect 160756 7750 160784 8434
rect 160744 7744 160796 7750
rect 160744 7686 160796 7692
rect 160560 4140 160612 4146
rect 160560 4082 160612 4088
rect 160284 4072 160336 4078
rect 160284 4014 160336 4020
rect 159916 3460 159968 3466
rect 159916 3402 159968 3408
rect 159732 3188 159784 3194
rect 159732 3130 159784 3136
rect 159824 2848 159876 2854
rect 159824 2790 159876 2796
rect 159548 2576 159600 2582
rect 159548 2518 159600 2524
rect 159836 1970 159864 2790
rect 159824 1964 159876 1970
rect 159824 1906 159876 1912
rect 159640 1760 159692 1766
rect 159640 1702 159692 1708
rect 159652 1358 159680 1702
rect 159836 1562 159864 1906
rect 159824 1556 159876 1562
rect 159824 1498 159876 1504
rect 159640 1352 159692 1358
rect 159640 1294 159692 1300
rect 159548 1284 159600 1290
rect 159548 1226 159600 1232
rect 159456 876 159508 882
rect 159456 818 159508 824
rect 159560 800 159588 1226
rect 159928 800 159956 3402
rect 160572 3398 160600 4082
rect 160560 3392 160612 3398
rect 160560 3334 160612 3340
rect 160192 2916 160244 2922
rect 160192 2858 160244 2864
rect 160204 2582 160232 2858
rect 160192 2576 160244 2582
rect 160192 2518 160244 2524
rect 160284 2304 160336 2310
rect 160284 2246 160336 2252
rect 160296 800 160324 2246
rect 160572 2122 160600 3334
rect 160756 3194 160784 7686
rect 160848 7342 160876 9046
rect 161216 9042 161244 12200
rect 161584 10146 161612 12200
rect 161952 12084 161980 12200
rect 161952 12056 162072 12084
rect 161584 10118 161704 10146
rect 161572 10056 161624 10062
rect 161572 9998 161624 10004
rect 161204 9036 161256 9042
rect 161204 8978 161256 8984
rect 161112 8424 161164 8430
rect 161112 8366 161164 8372
rect 161124 7954 161152 8366
rect 161112 7948 161164 7954
rect 161112 7890 161164 7896
rect 160928 7404 160980 7410
rect 160928 7346 160980 7352
rect 160836 7336 160888 7342
rect 160836 7278 160888 7284
rect 160744 3188 160796 3194
rect 160744 3130 160796 3136
rect 160652 3052 160704 3058
rect 160652 2994 160704 3000
rect 160664 2310 160692 2994
rect 160652 2304 160704 2310
rect 160652 2246 160704 2252
rect 160572 2094 160692 2122
rect 160940 2106 160968 7346
rect 161480 6792 161532 6798
rect 161480 6734 161532 6740
rect 161492 6458 161520 6734
rect 161480 6452 161532 6458
rect 161480 6394 161532 6400
rect 161584 4078 161612 9998
rect 161676 8634 161704 10118
rect 162044 9110 162072 12056
rect 162216 11756 162268 11762
rect 162216 11698 162268 11704
rect 162228 11354 162256 11698
rect 162216 11348 162268 11354
rect 162216 11290 162268 11296
rect 162320 10198 162348 12200
rect 162688 10690 162716 12200
rect 162964 11762 162992 12242
rect 163042 12200 163098 13000
rect 163410 12200 163466 13000
rect 163778 12200 163834 13000
rect 163872 12368 163924 12374
rect 163872 12310 163924 12316
rect 162952 11756 163004 11762
rect 162952 11698 163004 11704
rect 163056 11642 163084 12200
rect 163056 11614 163176 11642
rect 163044 11552 163096 11558
rect 163044 11494 163096 11500
rect 163056 11150 163084 11494
rect 163044 11144 163096 11150
rect 163044 11086 163096 11092
rect 162688 10662 162808 10690
rect 162676 10600 162728 10606
rect 162676 10542 162728 10548
rect 162688 10266 162716 10542
rect 162676 10260 162728 10266
rect 162676 10202 162728 10208
rect 162308 10192 162360 10198
rect 162308 10134 162360 10140
rect 162032 9104 162084 9110
rect 162032 9046 162084 9052
rect 162308 8832 162360 8838
rect 162308 8774 162360 8780
rect 161664 8628 161716 8634
rect 161664 8570 161716 8576
rect 162124 8356 162176 8362
rect 162124 8298 162176 8304
rect 162136 7954 162164 8298
rect 162124 7948 162176 7954
rect 162124 7890 162176 7896
rect 161940 7880 161992 7886
rect 161940 7822 161992 7828
rect 161756 4140 161808 4146
rect 161756 4082 161808 4088
rect 161572 4072 161624 4078
rect 161572 4014 161624 4020
rect 161768 3398 161796 4082
rect 161756 3392 161808 3398
rect 161756 3334 161808 3340
rect 161112 3120 161164 3126
rect 161112 3062 161164 3068
rect 161020 2440 161072 2446
rect 161020 2382 161072 2388
rect 160468 808 160520 814
rect 156788 750 156840 756
rect 156800 66 156828 750
rect 156788 60 156840 66
rect 156788 2 156840 8
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160664 800 160692 2094
rect 160928 2100 160980 2106
rect 160928 2042 160980 2048
rect 160836 1964 160888 1970
rect 160836 1906 160888 1912
rect 160848 1290 160876 1906
rect 160836 1284 160888 1290
rect 160836 1226 160888 1232
rect 161032 800 161060 2382
rect 161124 1358 161152 3062
rect 161572 2644 161624 2650
rect 161572 2586 161624 2592
rect 161584 2378 161612 2586
rect 161572 2372 161624 2378
rect 161572 2314 161624 2320
rect 161112 1352 161164 1358
rect 161112 1294 161164 1300
rect 161296 1216 161348 1222
rect 161480 1216 161532 1222
rect 161296 1158 161348 1164
rect 161400 1164 161480 1170
rect 161400 1158 161532 1164
rect 161308 1018 161336 1158
rect 161400 1142 161520 1158
rect 161296 1012 161348 1018
rect 161296 954 161348 960
rect 161400 800 161428 1142
rect 161768 800 161796 3334
rect 161952 2650 161980 7822
rect 162320 4078 162348 8774
rect 162780 8566 162808 10662
rect 162860 10668 162912 10674
rect 162860 10610 162912 10616
rect 162872 10130 162900 10610
rect 162860 10124 162912 10130
rect 162860 10066 162912 10072
rect 163148 9586 163176 11614
rect 163136 9580 163188 9586
rect 163136 9522 163188 9528
rect 163228 9512 163280 9518
rect 163228 9454 163280 9460
rect 163240 8906 163268 9454
rect 163424 9450 163452 12200
rect 163412 9444 163464 9450
rect 163412 9386 163464 9392
rect 163228 8900 163280 8906
rect 163228 8842 163280 8848
rect 162400 8560 162452 8566
rect 162400 8502 162452 8508
rect 162768 8560 162820 8566
rect 162768 8502 162820 8508
rect 162412 6934 162440 8502
rect 163792 8498 163820 12200
rect 163884 11218 163912 12310
rect 164146 12200 164202 13000
rect 164514 12200 164570 13000
rect 164882 12200 164938 13000
rect 165896 12232 165948 12238
rect 163872 11212 163924 11218
rect 163872 11154 163924 11160
rect 163964 10056 164016 10062
rect 163964 9998 164016 10004
rect 163780 8492 163832 8498
rect 163780 8434 163832 8440
rect 163412 7744 163464 7750
rect 163412 7686 163464 7692
rect 163424 7546 163452 7686
rect 163412 7540 163464 7546
rect 163412 7482 163464 7488
rect 163320 7336 163372 7342
rect 163320 7278 163372 7284
rect 163332 7002 163360 7278
rect 163504 7200 163556 7206
rect 163504 7142 163556 7148
rect 163320 6996 163372 7002
rect 163320 6938 163372 6944
rect 162400 6928 162452 6934
rect 162400 6870 162452 6876
rect 163516 6866 163544 7142
rect 163504 6860 163556 6866
rect 163504 6802 163556 6808
rect 162400 6724 162452 6730
rect 162400 6666 162452 6672
rect 162308 4072 162360 4078
rect 162308 4014 162360 4020
rect 162308 3596 162360 3602
rect 162308 3538 162360 3544
rect 162032 2984 162084 2990
rect 162032 2926 162084 2932
rect 161940 2644 161992 2650
rect 161940 2586 161992 2592
rect 161940 1964 161992 1970
rect 161940 1906 161992 1912
rect 161952 1222 161980 1906
rect 161940 1216 161992 1222
rect 161940 1158 161992 1164
rect 162044 882 162072 2926
rect 162216 2440 162268 2446
rect 162136 2400 162216 2428
rect 162032 876 162084 882
rect 162032 818 162084 824
rect 162136 800 162164 2400
rect 162216 2382 162268 2388
rect 162320 1358 162348 3538
rect 162412 2106 162440 6666
rect 163516 6458 163544 6802
rect 163504 6452 163556 6458
rect 163504 6394 163556 6400
rect 163504 6248 163556 6254
rect 163504 6190 163556 6196
rect 163516 5914 163544 6190
rect 163596 6112 163648 6118
rect 163596 6054 163648 6060
rect 163504 5908 163556 5914
rect 163504 5850 163556 5856
rect 163608 5778 163636 6054
rect 163596 5772 163648 5778
rect 163596 5714 163648 5720
rect 163976 4826 164004 9998
rect 164160 8378 164188 12200
rect 164332 11620 164384 11626
rect 164332 11562 164384 11568
rect 164344 10674 164372 11562
rect 164332 10668 164384 10674
rect 164332 10610 164384 10616
rect 164344 10266 164372 10610
rect 164332 10260 164384 10266
rect 164332 10202 164384 10208
rect 164332 9580 164384 9586
rect 164332 9522 164384 9528
rect 164160 8350 164280 8378
rect 164252 7342 164280 8350
rect 164240 7336 164292 7342
rect 164240 7278 164292 7284
rect 164240 6792 164292 6798
rect 164240 6734 164292 6740
rect 163964 4820 164016 4826
rect 163964 4762 164016 4768
rect 163596 4480 163648 4486
rect 163596 4422 163648 4428
rect 162492 4140 162544 4146
rect 162492 4082 162544 4088
rect 162504 3398 162532 4082
rect 163228 3528 163280 3534
rect 163228 3470 163280 3476
rect 162492 3392 162544 3398
rect 162492 3334 162544 3340
rect 162400 2100 162452 2106
rect 162400 2042 162452 2048
rect 162308 1352 162360 1358
rect 162308 1294 162360 1300
rect 162504 800 162532 3334
rect 162860 1352 162912 1358
rect 162860 1294 162912 1300
rect 162768 1216 162820 1222
rect 162768 1158 162820 1164
rect 162780 882 162808 1158
rect 162768 876 162820 882
rect 162768 818 162820 824
rect 162872 800 162900 1294
rect 163240 800 163268 3470
rect 163608 800 163636 4422
rect 164252 3074 164280 6734
rect 164344 3194 164372 9522
rect 164424 8968 164476 8974
rect 164424 8910 164476 8916
rect 164436 3738 164464 8910
rect 164528 8378 164556 12200
rect 164896 9500 164924 12200
rect 165896 12174 165948 12180
rect 165908 11762 165936 12174
rect 165896 11756 165948 11762
rect 165896 11698 165948 11704
rect 167184 11756 167236 11762
rect 167184 11698 167236 11704
rect 165908 11354 165936 11698
rect 166080 11688 166132 11694
rect 166080 11630 166132 11636
rect 165896 11348 165948 11354
rect 165896 11290 165948 11296
rect 166092 11218 166120 11630
rect 166724 11552 166776 11558
rect 166724 11494 166776 11500
rect 166080 11212 166132 11218
rect 166080 11154 166132 11160
rect 166736 10674 166764 11494
rect 167196 11150 167224 11698
rect 167184 11144 167236 11150
rect 167184 11086 167236 11092
rect 166724 10668 166776 10674
rect 166724 10610 166776 10616
rect 165620 10600 165672 10606
rect 165620 10542 165672 10548
rect 165632 10266 165660 10542
rect 166736 10266 166764 10610
rect 165620 10260 165672 10266
rect 165620 10202 165672 10208
rect 166724 10260 166776 10266
rect 166724 10202 166776 10208
rect 165804 9580 165856 9586
rect 165804 9522 165856 9528
rect 166908 9580 166960 9586
rect 166908 9522 166960 9528
rect 164804 9472 164924 9500
rect 164804 8809 164832 9472
rect 164884 9376 164936 9382
rect 164884 9318 164936 9324
rect 164790 8800 164846 8809
rect 164790 8735 164846 8744
rect 164792 8628 164844 8634
rect 164792 8570 164844 8576
rect 164700 8492 164752 8498
rect 164700 8434 164752 8440
rect 164528 8362 164648 8378
rect 164528 8356 164660 8362
rect 164528 8350 164608 8356
rect 164608 8298 164660 8304
rect 164608 7880 164660 7886
rect 164608 7822 164660 7828
rect 164516 6656 164568 6662
rect 164516 6598 164568 6604
rect 164424 3732 164476 3738
rect 164424 3674 164476 3680
rect 164424 3392 164476 3398
rect 164424 3334 164476 3340
rect 164332 3188 164384 3194
rect 164332 3130 164384 3136
rect 164148 3052 164200 3058
rect 164252 3046 164372 3074
rect 164148 2994 164200 3000
rect 164160 2310 164188 2994
rect 164344 2650 164372 3046
rect 164332 2644 164384 2650
rect 164332 2586 164384 2592
rect 164148 2304 164200 2310
rect 164200 2252 164372 2258
rect 164148 2246 164372 2252
rect 164160 2230 164372 2246
rect 163964 1964 164016 1970
rect 163964 1906 164016 1912
rect 163976 1426 164004 1906
rect 163964 1420 164016 1426
rect 163964 1362 164016 1368
rect 163976 800 164004 1362
rect 164344 800 164372 2230
rect 164436 1222 164464 3334
rect 164528 2514 164556 6598
rect 164620 3398 164648 7822
rect 164712 5778 164740 8434
rect 164804 8022 164832 8570
rect 164792 8016 164844 8022
rect 164792 7958 164844 7964
rect 164896 6934 164924 9318
rect 165816 9178 165844 9522
rect 165804 9172 165856 9178
rect 165804 9114 165856 9120
rect 166724 9104 166776 9110
rect 166724 9046 166776 9052
rect 165160 8560 165212 8566
rect 165160 8502 165212 8508
rect 164976 7404 165028 7410
rect 164976 7346 165028 7352
rect 164884 6928 164936 6934
rect 164884 6870 164936 6876
rect 164988 6662 165016 7346
rect 164976 6656 165028 6662
rect 164976 6598 165028 6604
rect 164792 6384 164844 6390
rect 164792 6326 164844 6332
rect 164700 5772 164752 5778
rect 164700 5714 164752 5720
rect 164700 5228 164752 5234
rect 164700 5170 164752 5176
rect 164712 4486 164740 5170
rect 164700 4480 164752 4486
rect 164700 4422 164752 4428
rect 164608 3392 164660 3398
rect 164608 3334 164660 3340
rect 164608 2848 164660 2854
rect 164608 2790 164660 2796
rect 164516 2508 164568 2514
rect 164516 2450 164568 2456
rect 164620 2446 164648 2790
rect 164608 2440 164660 2446
rect 164608 2382 164660 2388
rect 164424 1216 164476 1222
rect 164424 1158 164476 1164
rect 164712 800 164740 4422
rect 164804 4026 164832 6326
rect 164976 6316 165028 6322
rect 164976 6258 165028 6264
rect 164884 6180 164936 6186
rect 164884 6122 164936 6128
rect 164896 4146 164924 6122
rect 164988 5574 165016 6258
rect 165172 6186 165200 8502
rect 165620 8492 165672 8498
rect 165620 8434 165672 8440
rect 165632 7750 165660 8434
rect 166172 8424 166224 8430
rect 166172 8366 166224 8372
rect 166184 8090 166212 8366
rect 166172 8084 166224 8090
rect 166172 8026 166224 8032
rect 166736 7954 166764 9046
rect 166920 8838 166948 9522
rect 166908 8832 166960 8838
rect 166908 8774 166960 8780
rect 166724 7948 166776 7954
rect 166724 7890 166776 7896
rect 165620 7744 165672 7750
rect 165620 7686 165672 7692
rect 165160 6180 165212 6186
rect 165160 6122 165212 6128
rect 165068 5704 165120 5710
rect 165068 5646 165120 5652
rect 164976 5568 165028 5574
rect 164976 5510 165028 5516
rect 164884 4140 164936 4146
rect 164884 4082 164936 4088
rect 164804 3998 164924 4026
rect 164896 1970 164924 3998
rect 164988 2106 165016 5510
rect 165080 3194 165108 5646
rect 165632 4146 165660 7686
rect 166920 5370 166948 8774
rect 166908 5364 166960 5370
rect 166908 5306 166960 5312
rect 165528 4140 165580 4146
rect 165528 4082 165580 4088
rect 165620 4140 165672 4146
rect 165620 4082 165672 4088
rect 165540 3738 165568 4082
rect 165528 3732 165580 3738
rect 165528 3674 165580 3680
rect 166724 3664 166776 3670
rect 166724 3606 166776 3612
rect 165068 3188 165120 3194
rect 165068 3130 165120 3136
rect 165068 3052 165120 3058
rect 165068 2994 165120 3000
rect 164976 2100 165028 2106
rect 164976 2042 165028 2048
rect 164884 1964 164936 1970
rect 164884 1906 164936 1912
rect 164896 1562 164924 1906
rect 164884 1556 164936 1562
rect 164884 1498 164936 1504
rect 165080 800 165108 2994
rect 165804 2372 165856 2378
rect 165804 2314 165856 2320
rect 165436 1420 165488 1426
rect 165436 1362 165488 1368
rect 165448 800 165476 1362
rect 165816 800 165844 2314
rect 166080 1964 166132 1970
rect 166080 1906 166132 1912
rect 166092 1562 166120 1906
rect 166172 1896 166224 1902
rect 166172 1838 166224 1844
rect 166540 1896 166592 1902
rect 166540 1838 166592 1844
rect 166080 1556 166132 1562
rect 166080 1498 166132 1504
rect 165988 808 166040 814
rect 160468 750 160520 756
rect 160480 270 160508 750
rect 160468 264 160520 270
rect 160468 206 160520 212
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 165986 776 165988 785
rect 166184 800 166212 1838
rect 166552 800 166580 1838
rect 166736 1358 166764 3606
rect 166908 1964 166960 1970
rect 166908 1906 166960 1912
rect 166724 1352 166776 1358
rect 166724 1294 166776 1300
rect 166920 1222 166948 1906
rect 166816 1216 166868 1222
rect 166816 1158 166868 1164
rect 166908 1216 166960 1222
rect 166908 1158 166960 1164
rect 166828 1018 166856 1158
rect 166816 1012 166868 1018
rect 166816 954 166868 960
rect 166040 776 166042 785
rect 165986 711 166042 720
rect 166170 0 166226 800
rect 166538 0 166594 800
<< via2 >>
rect 2870 10376 2926 10432
rect 3698 12008 3754 12064
rect 3606 10920 3662 10976
rect 3698 6024 3754 6080
rect 4066 11464 4122 11520
rect 4066 9832 4122 9888
rect 4066 8744 4122 8800
rect 4066 8200 4122 8256
rect 4066 7112 4122 7168
rect 4066 6568 4122 6624
rect 3882 5480 3938 5536
rect 3698 4936 3754 4992
rect 4710 8608 4766 8664
rect 4802 7656 4858 7712
rect 5078 9868 5080 9888
rect 5080 9868 5132 9888
rect 5132 9868 5134 9888
rect 5078 9832 5134 9868
rect 5538 9152 5594 9208
rect 5354 5636 5410 5672
rect 5354 5616 5356 5636
rect 5356 5616 5408 5636
rect 5408 5616 5410 5636
rect 5354 5228 5410 5264
rect 5354 5208 5356 5228
rect 5356 5208 5408 5228
rect 5408 5208 5410 5228
rect 5538 7112 5594 7168
rect 6090 9288 6146 9344
rect 6366 6860 6422 6896
rect 6366 6840 6368 6860
rect 6368 6840 6420 6860
rect 6420 6840 6422 6860
rect 5446 4664 5502 4720
rect 4066 4392 4122 4448
rect 938 3032 994 3088
rect 2962 2216 3018 2272
rect 4066 3848 4122 3904
rect 3790 1128 3846 1184
rect 3974 2760 4030 2816
rect 4066 1708 4068 1728
rect 4068 1708 4120 1728
rect 4120 1708 4122 1728
rect 4066 1672 4122 1708
rect 5170 1708 5172 1728
rect 5172 1708 5224 1728
rect 5224 1708 5226 1728
rect 5170 1672 5226 1708
rect 6826 7384 6882 7440
rect 6642 6160 6698 6216
rect 5906 4548 5962 4584
rect 5906 4528 5908 4548
rect 5908 4528 5960 4548
rect 5960 4528 5962 4548
rect 5906 4120 5962 4176
rect 6090 3984 6146 4040
rect 6458 3848 6514 3904
rect 6182 3304 6238 3360
rect 5630 740 5686 776
rect 5630 720 5632 740
rect 5632 720 5684 740
rect 5684 720 5686 740
rect 6642 3732 6698 3768
rect 6642 3712 6644 3732
rect 6644 3712 6696 3732
rect 6696 3712 6698 3732
rect 7654 11212 7710 11248
rect 7654 11192 7656 11212
rect 7656 11192 7708 11212
rect 7708 11192 7710 11212
rect 7378 9424 7434 9480
rect 8022 11092 8024 11112
rect 8024 11092 8076 11112
rect 8076 11092 8078 11112
rect 8022 11056 8078 11092
rect 8482 9016 8538 9072
rect 8298 8900 8354 8936
rect 8298 8880 8300 8900
rect 8300 8880 8352 8900
rect 8352 8880 8354 8900
rect 8206 7112 8262 7168
rect 8114 6432 8170 6488
rect 7746 5772 7802 5808
rect 7746 5752 7748 5772
rect 7748 5752 7800 5772
rect 7800 5752 7802 5772
rect 7194 5480 7250 5536
rect 9310 10920 9366 10976
rect 9678 10140 9680 10160
rect 9680 10140 9732 10160
rect 9732 10140 9734 10160
rect 9678 10104 9734 10140
rect 9218 6024 9274 6080
rect 7194 4256 7250 4312
rect 10874 6604 10876 6624
rect 10876 6604 10928 6624
rect 10928 6604 10930 6624
rect 10874 6568 10930 6604
rect 11794 9560 11850 9616
rect 12162 8336 12218 8392
rect 11058 5888 11114 5944
rect 10874 5072 10930 5128
rect 6274 312 6330 368
rect 8022 3732 8078 3768
rect 8022 3712 8024 3732
rect 8024 3712 8076 3732
rect 8076 3712 8078 3732
rect 9586 4392 9642 4448
rect 8114 876 8170 912
rect 8114 856 8116 876
rect 8116 856 8168 876
rect 8168 856 8170 876
rect 9034 2216 9090 2272
rect 8390 992 8446 1048
rect 9678 3304 9734 3360
rect 9770 2352 9826 2408
rect 10138 2488 10194 2544
rect 10782 2080 10838 2136
rect 10506 1264 10562 1320
rect 12898 7928 12954 7984
rect 13634 7792 13690 7848
rect 13266 7112 13322 7168
rect 12438 6976 12494 7032
rect 12438 6568 12494 6624
rect 12346 6296 12402 6352
rect 15566 9596 15568 9616
rect 15568 9596 15620 9616
rect 15620 9596 15622 9616
rect 15566 9560 15622 9596
rect 15934 8064 15990 8120
rect 16486 11736 16542 11792
rect 17314 10104 17370 10160
rect 17038 9696 17094 9752
rect 16210 8472 16266 8528
rect 17222 8336 17278 8392
rect 15658 7520 15714 7576
rect 16026 7284 16028 7304
rect 16028 7284 16080 7304
rect 16080 7284 16082 7304
rect 16026 7248 16082 7284
rect 16486 6724 16542 6760
rect 16486 6704 16488 6724
rect 16488 6704 16540 6724
rect 16540 6704 16542 6724
rect 16854 6568 16910 6624
rect 16854 6296 16910 6352
rect 17038 6296 17094 6352
rect 17038 5888 17094 5944
rect 17314 6024 17370 6080
rect 17314 5752 17370 5808
rect 12530 4392 12586 4448
rect 11518 3460 11574 3496
rect 11518 3440 11520 3460
rect 11520 3440 11572 3460
rect 11572 3440 11574 3460
rect 11242 1400 11298 1456
rect 11702 2760 11758 2816
rect 12530 4120 12586 4176
rect 12346 2896 12402 2952
rect 12714 1944 12770 2000
rect 13082 1808 13138 1864
rect 12806 1164 12808 1184
rect 12808 1164 12860 1184
rect 12860 1164 12862 1184
rect 12806 1128 12862 1164
rect 13450 1536 13506 1592
rect 19246 7656 19302 7712
rect 15842 2624 15898 2680
rect 15842 2352 15898 2408
rect 16578 3884 16580 3904
rect 16580 3884 16632 3904
rect 16632 3884 16634 3904
rect 16578 3848 16634 3884
rect 14278 40 14334 96
rect 20626 9560 20682 9616
rect 20258 9288 20314 9344
rect 21638 10668 21694 10704
rect 21638 10648 21640 10668
rect 21640 10648 21692 10668
rect 21692 10648 21694 10668
rect 22466 11464 22522 11520
rect 22834 11328 22890 11384
rect 21730 10376 21786 10432
rect 23386 10004 23388 10024
rect 23388 10004 23440 10024
rect 23440 10004 23442 10024
rect 23386 9968 23442 10004
rect 25042 12008 25098 12064
rect 24674 11872 24730 11928
rect 23938 10240 23994 10296
rect 23662 9832 23718 9888
rect 20258 2388 20260 2408
rect 20260 2388 20312 2408
rect 20312 2388 20314 2408
rect 20258 2352 20314 2388
rect 21638 9152 21694 9208
rect 22558 9288 22614 9344
rect 22190 9152 22246 9208
rect 21086 6024 21142 6080
rect 21086 3168 21142 3224
rect 21086 2388 21088 2408
rect 21088 2388 21140 2408
rect 21140 2388 21142 2408
rect 21086 2352 21142 2388
rect 21270 3848 21326 3904
rect 22190 8200 22246 8256
rect 22558 8472 22614 8528
rect 21730 3848 21786 3904
rect 21914 3596 21970 3632
rect 21914 3576 21916 3596
rect 21916 3576 21968 3596
rect 21968 3576 21970 3596
rect 21546 2760 21602 2816
rect 21546 2352 21602 2408
rect 19246 448 19302 504
rect 23846 8780 23848 8800
rect 23848 8780 23900 8800
rect 23900 8780 23902 8800
rect 23846 8744 23902 8780
rect 24674 9560 24730 9616
rect 25410 10784 25466 10840
rect 26606 12144 26662 12200
rect 26146 11600 26202 11656
rect 25778 10512 25834 10568
rect 26882 10376 26938 10432
rect 27066 10376 27122 10432
rect 26882 9696 26938 9752
rect 23294 8336 23350 8392
rect 23202 7384 23258 7440
rect 25318 9580 25374 9616
rect 25318 9560 25320 9580
rect 25320 9560 25372 9580
rect 25372 9560 25374 9580
rect 24306 6976 24362 7032
rect 24858 7656 24914 7712
rect 23938 3168 23994 3224
rect 24858 3168 24914 3224
rect 25594 6976 25650 7032
rect 25410 3168 25466 3224
rect 26422 8200 26478 8256
rect 26422 7656 26478 7712
rect 26606 7112 26662 7168
rect 27710 10376 27766 10432
rect 30654 12824 30710 12880
rect 28262 11464 28318 11520
rect 28078 11328 28134 11384
rect 27618 8336 27674 8392
rect 26974 6024 27030 6080
rect 26790 5752 26846 5808
rect 26974 5752 27030 5808
rect 26330 3168 26386 3224
rect 26238 1708 26240 1728
rect 26240 1708 26292 1728
rect 26292 1708 26294 1728
rect 26238 1672 26294 1708
rect 27802 5344 27858 5400
rect 26606 1844 26608 1864
rect 26608 1844 26660 1864
rect 26660 1844 26662 1864
rect 26606 1808 26662 1844
rect 24582 176 24638 232
rect 28430 11450 28486 11452
rect 28510 11450 28566 11452
rect 28590 11450 28646 11452
rect 28670 11450 28726 11452
rect 28430 11398 28456 11450
rect 28456 11398 28486 11450
rect 28510 11398 28520 11450
rect 28520 11398 28566 11450
rect 28590 11398 28636 11450
rect 28636 11398 28646 11450
rect 28670 11398 28700 11450
rect 28700 11398 28726 11450
rect 28430 11396 28486 11398
rect 28510 11396 28566 11398
rect 28590 11396 28646 11398
rect 28670 11396 28726 11398
rect 28430 10362 28486 10364
rect 28510 10362 28566 10364
rect 28590 10362 28646 10364
rect 28670 10362 28726 10364
rect 28430 10310 28456 10362
rect 28456 10310 28486 10362
rect 28510 10310 28520 10362
rect 28520 10310 28566 10362
rect 28590 10310 28636 10362
rect 28636 10310 28646 10362
rect 28670 10310 28700 10362
rect 28700 10310 28726 10362
rect 28430 10308 28486 10310
rect 28510 10308 28566 10310
rect 28590 10308 28646 10310
rect 28670 10308 28726 10310
rect 28262 10240 28318 10296
rect 28998 10140 29000 10160
rect 29000 10140 29052 10160
rect 29052 10140 29054 10160
rect 28998 10104 29054 10140
rect 31114 12008 31170 12064
rect 30746 10104 30802 10160
rect 31206 11872 31262 11928
rect 31482 11872 31538 11928
rect 31206 10104 31262 10160
rect 31114 9832 31170 9888
rect 31850 11328 31906 11384
rect 32126 11464 32182 11520
rect 33690 12960 33746 13016
rect 33598 12552 33654 12608
rect 31850 10104 31906 10160
rect 33414 12144 33470 12200
rect 33230 12008 33286 12064
rect 28262 9288 28318 9344
rect 28814 9288 28870 9344
rect 28430 9274 28486 9276
rect 28510 9274 28566 9276
rect 28590 9274 28646 9276
rect 28670 9274 28726 9276
rect 28430 9222 28456 9274
rect 28456 9222 28486 9274
rect 28510 9222 28520 9274
rect 28520 9222 28566 9274
rect 28590 9222 28636 9274
rect 28636 9222 28646 9274
rect 28670 9222 28700 9274
rect 28700 9222 28726 9274
rect 28430 9220 28486 9222
rect 28510 9220 28566 9222
rect 28590 9220 28646 9222
rect 28670 9220 28726 9222
rect 28262 9152 28318 9208
rect 28814 9172 28870 9208
rect 28814 9152 28816 9172
rect 28816 9152 28868 9172
rect 28868 9152 28870 9172
rect 28998 8336 29054 8392
rect 28430 8186 28486 8188
rect 28510 8186 28566 8188
rect 28590 8186 28646 8188
rect 28670 8186 28726 8188
rect 28430 8134 28456 8186
rect 28456 8134 28486 8186
rect 28510 8134 28520 8186
rect 28520 8134 28566 8186
rect 28590 8134 28636 8186
rect 28636 8134 28646 8186
rect 28670 8134 28700 8186
rect 28700 8134 28726 8186
rect 28430 8132 28486 8134
rect 28510 8132 28566 8134
rect 28590 8132 28646 8134
rect 28670 8132 28726 8134
rect 28814 7148 28816 7168
rect 28816 7148 28868 7168
rect 28868 7148 28870 7168
rect 28814 7112 28870 7148
rect 28430 7098 28486 7100
rect 28510 7098 28566 7100
rect 28590 7098 28646 7100
rect 28670 7098 28726 7100
rect 28430 7046 28456 7098
rect 28456 7046 28486 7098
rect 28510 7046 28520 7098
rect 28520 7046 28566 7098
rect 28590 7046 28636 7098
rect 28636 7046 28646 7098
rect 28670 7046 28700 7098
rect 28700 7046 28726 7098
rect 28430 7044 28486 7046
rect 28510 7044 28566 7046
rect 28590 7044 28646 7046
rect 28670 7044 28726 7046
rect 28170 6976 28226 7032
rect 28814 6996 28870 7032
rect 28814 6976 28816 6996
rect 28816 6976 28868 6996
rect 28868 6976 28870 6996
rect 31758 7112 31814 7168
rect 32034 6976 32090 7032
rect 28814 6024 28870 6080
rect 28430 6010 28486 6012
rect 28510 6010 28566 6012
rect 28590 6010 28646 6012
rect 28670 6010 28726 6012
rect 28430 5958 28456 6010
rect 28456 5958 28486 6010
rect 28510 5958 28520 6010
rect 28520 5958 28566 6010
rect 28590 5958 28636 6010
rect 28636 5958 28646 6010
rect 28670 5958 28700 6010
rect 28700 5958 28726 6010
rect 28430 5956 28486 5958
rect 28510 5956 28566 5958
rect 28590 5956 28646 5958
rect 28670 5956 28726 5958
rect 28262 5888 28318 5944
rect 28998 5752 29054 5808
rect 27250 3304 27306 3360
rect 27434 3304 27490 3360
rect 28906 5344 28962 5400
rect 29090 5344 29146 5400
rect 28998 5072 29054 5128
rect 28430 4922 28486 4924
rect 28510 4922 28566 4924
rect 28590 4922 28646 4924
rect 28670 4922 28726 4924
rect 28430 4870 28456 4922
rect 28456 4870 28486 4922
rect 28510 4870 28520 4922
rect 28520 4870 28566 4922
rect 28590 4870 28636 4922
rect 28636 4870 28646 4922
rect 28670 4870 28700 4922
rect 28700 4870 28726 4922
rect 28430 4868 28486 4870
rect 28510 4868 28566 4870
rect 28590 4868 28646 4870
rect 28670 4868 28726 4870
rect 29182 4800 29238 4856
rect 28078 3732 28134 3768
rect 28078 3712 28080 3732
rect 28080 3712 28132 3732
rect 28132 3712 28134 3732
rect 28998 3984 29054 4040
rect 28262 3848 28318 3904
rect 28814 3848 28870 3904
rect 28430 3834 28486 3836
rect 28510 3834 28566 3836
rect 28590 3834 28646 3836
rect 28670 3834 28726 3836
rect 28430 3782 28456 3834
rect 28456 3782 28486 3834
rect 28510 3782 28520 3834
rect 28520 3782 28566 3834
rect 28590 3782 28636 3834
rect 28636 3782 28646 3834
rect 28670 3782 28700 3834
rect 28700 3782 28726 3834
rect 28430 3780 28486 3782
rect 28510 3780 28566 3782
rect 28590 3780 28646 3782
rect 28670 3780 28726 3782
rect 27710 448 27766 504
rect 28262 2644 28318 2680
rect 28262 2624 28264 2644
rect 28264 2624 28316 2644
rect 28316 2624 28318 2644
rect 28906 3732 28962 3768
rect 28906 3712 28908 3732
rect 28908 3712 28960 3732
rect 28960 3712 28962 3732
rect 28814 2760 28870 2816
rect 28430 2746 28486 2748
rect 28510 2746 28566 2748
rect 28590 2746 28646 2748
rect 28670 2746 28726 2748
rect 28430 2694 28456 2746
rect 28456 2694 28486 2746
rect 28510 2694 28520 2746
rect 28520 2694 28566 2746
rect 28590 2694 28636 2746
rect 28636 2694 28646 2746
rect 28670 2694 28700 2746
rect 28700 2694 28726 2746
rect 28430 2692 28486 2694
rect 28510 2692 28566 2694
rect 28590 2692 28646 2694
rect 28670 2692 28726 2694
rect 28814 2644 28870 2680
rect 28814 2624 28816 2644
rect 28816 2624 28868 2644
rect 28868 2624 28870 2644
rect 28430 1658 28486 1660
rect 28510 1658 28566 1660
rect 28590 1658 28646 1660
rect 28670 1658 28726 1660
rect 28430 1606 28456 1658
rect 28456 1606 28486 1658
rect 28510 1606 28520 1658
rect 28520 1606 28566 1658
rect 28590 1606 28636 1658
rect 28636 1606 28646 1658
rect 28670 1606 28700 1658
rect 28700 1606 28726 1658
rect 28430 1604 28486 1606
rect 28510 1604 28566 1606
rect 28590 1604 28646 1606
rect 28670 1604 28726 1606
rect 28814 1536 28870 1592
rect 28998 1808 29054 1864
rect 28430 570 28486 572
rect 28510 570 28566 572
rect 28590 570 28646 572
rect 28670 570 28726 572
rect 28430 518 28456 570
rect 28456 518 28486 570
rect 28510 518 28520 570
rect 28520 518 28566 570
rect 28590 518 28636 570
rect 28636 518 28646 570
rect 28670 518 28700 570
rect 28700 518 28726 570
rect 28430 516 28486 518
rect 28510 516 28566 518
rect 28590 516 28646 518
rect 28670 516 28726 518
rect 31758 5208 31814 5264
rect 30838 4800 30894 4856
rect 31390 4800 31446 4856
rect 29090 448 29146 504
rect 31206 3304 31262 3360
rect 32218 4936 32274 4992
rect 31390 3032 31446 3088
rect 31942 3168 31998 3224
rect 31850 2760 31906 2816
rect 33322 8200 33378 8256
rect 33782 12280 33838 12336
rect 33966 12688 34022 12744
rect 35622 12824 35678 12880
rect 35898 12860 35900 12880
rect 35900 12860 35952 12880
rect 35952 12860 35954 12880
rect 35898 12824 35954 12860
rect 34426 12144 34482 12200
rect 35162 10260 35218 10296
rect 35162 10240 35164 10260
rect 35164 10240 35216 10260
rect 35216 10240 35218 10260
rect 32494 3848 32550 3904
rect 32770 1264 32826 1320
rect 31942 720 31998 776
rect 32862 468 32918 504
rect 32862 448 32864 468
rect 32864 448 32916 468
rect 32916 448 32918 468
rect 33138 448 33194 504
rect 36726 12416 36782 12472
rect 35990 11872 36046 11928
rect 36266 11872 36322 11928
rect 36358 11464 36414 11520
rect 36266 9016 36322 9072
rect 36634 11464 36690 11520
rect 36542 9016 36598 9072
rect 36542 8336 36598 8392
rect 37278 10104 37334 10160
rect 37462 10124 37518 10160
rect 37462 10104 37464 10124
rect 37464 10104 37516 10124
rect 37516 10104 37518 10124
rect 40406 12824 40462 12880
rect 40406 12280 40462 12336
rect 38566 9288 38622 9344
rect 36818 8336 36874 8392
rect 35162 4800 35218 4856
rect 35162 3848 35218 3904
rect 35714 3848 35770 3904
rect 35530 2388 35532 2408
rect 35532 2388 35584 2408
rect 35584 2388 35586 2408
rect 35530 2352 35586 2388
rect 35806 2896 35862 2952
rect 35990 2896 36046 2952
rect 35898 2624 35954 2680
rect 35898 2352 35954 2408
rect 34518 448 34574 504
rect 36082 2624 36138 2680
rect 36358 4800 36414 4856
rect 37002 4936 37058 4992
rect 36358 4256 36414 4312
rect 36634 3984 36690 4040
rect 39670 12008 39726 12064
rect 39854 12008 39910 12064
rect 40314 12144 40370 12200
rect 40590 12824 40646 12880
rect 40130 10104 40186 10160
rect 38750 9016 38806 9072
rect 39210 9288 39266 9344
rect 39026 9016 39082 9072
rect 39946 9424 40002 9480
rect 40774 12688 40830 12744
rect 40682 12552 40738 12608
rect 40682 12280 40738 12336
rect 41142 12960 41198 13016
rect 40958 12572 41014 12608
rect 40958 12552 40960 12572
rect 40960 12552 41012 12572
rect 41012 12552 41014 12572
rect 40682 12008 40738 12064
rect 40314 10104 40370 10160
rect 40130 9424 40186 9480
rect 36358 3848 36414 3904
rect 36542 1264 36598 1320
rect 35254 448 35310 504
rect 35806 720 35862 776
rect 35806 584 35862 640
rect 37462 2760 37518 2816
rect 38474 2760 38530 2816
rect 38750 1264 38806 1320
rect 37094 448 37150 504
rect 39210 2896 39266 2952
rect 39394 2896 39450 2952
rect 41418 12688 41474 12744
rect 41510 12572 41566 12608
rect 41510 12552 41512 12572
rect 41512 12552 41564 12572
rect 41564 12552 41566 12572
rect 41694 12588 41696 12608
rect 41696 12588 41748 12608
rect 41748 12588 41750 12608
rect 41694 12552 41750 12588
rect 41418 12144 41474 12200
rect 41602 12008 41658 12064
rect 42522 12688 42578 12744
rect 42154 12144 42210 12200
rect 42246 12008 42302 12064
rect 43166 12688 43222 12744
rect 42338 11872 42394 11928
rect 42706 9288 42762 9344
rect 42706 9016 42762 9072
rect 42890 9288 42946 9344
rect 42246 8336 42302 8392
rect 41694 6976 41750 7032
rect 41878 6976 41934 7032
rect 40222 3304 40278 3360
rect 39946 2932 39948 2952
rect 39948 2932 40000 2952
rect 40000 2932 40002 2952
rect 39946 2896 40002 2932
rect 40406 3304 40462 3360
rect 40222 2896 40278 2952
rect 45098 12280 45154 12336
rect 43718 11872 43774 11928
rect 44086 11736 44142 11792
rect 45558 11464 45614 11520
rect 45742 11736 45798 11792
rect 46294 12860 46296 12880
rect 46296 12860 46348 12880
rect 46348 12860 46350 12880
rect 46294 12824 46350 12860
rect 46478 12724 46480 12744
rect 46480 12724 46532 12744
rect 46532 12724 46534 12744
rect 46478 12688 46534 12724
rect 46478 12552 46534 12608
rect 45742 10920 45798 10976
rect 40866 4800 40922 4856
rect 41050 4800 41106 4856
rect 41510 5072 41566 5128
rect 41878 4392 41934 4448
rect 41694 4120 41750 4176
rect 41878 4120 41934 4176
rect 41786 3712 41842 3768
rect 41510 3576 41566 3632
rect 42430 4392 42486 4448
rect 40406 2760 40462 2816
rect 40774 2760 40830 2816
rect 40958 2760 41014 2816
rect 40866 1264 40922 1320
rect 41050 1264 41106 1320
rect 40498 448 40554 504
rect 41326 448 41382 504
rect 43258 4392 43314 4448
rect 43258 2896 43314 2952
rect 44086 2896 44142 2952
rect 46202 11464 46258 11520
rect 46110 10920 46166 10976
rect 46110 10512 46166 10568
rect 48502 12552 48558 12608
rect 46570 11872 46626 11928
rect 46202 9832 46258 9888
rect 46018 9560 46074 9616
rect 46202 9560 46258 9616
rect 46386 9832 46442 9888
rect 46110 8472 46166 8528
rect 43902 1128 43958 1184
rect 46570 8880 46626 8936
rect 46110 7792 46166 7848
rect 46386 7656 46442 7712
rect 46110 6568 46166 6624
rect 46386 6432 46442 6488
rect 48502 12144 48558 12200
rect 46018 6024 46074 6080
rect 46202 6024 46258 6080
rect 46202 5752 46258 5808
rect 46386 5752 46442 5808
rect 46018 4392 46074 4448
rect 46386 4528 46442 4584
rect 46386 4120 46442 4176
rect 46846 4120 46902 4176
rect 47030 4120 47086 4176
rect 45374 2760 45430 2816
rect 46846 3168 46902 3224
rect 48318 9560 48374 9616
rect 47030 2760 47086 2816
rect 47214 2760 47270 2816
rect 45190 448 45246 504
rect 46386 856 46442 912
rect 47122 1128 47178 1184
rect 47306 1128 47362 1184
rect 47030 856 47086 912
rect 46386 584 46442 640
rect 48686 9560 48742 9616
rect 49238 10648 49294 10704
rect 49790 8744 49846 8800
rect 50342 10648 50398 10704
rect 50618 12144 50674 12200
rect 50894 12980 50950 13016
rect 50894 12960 50896 12980
rect 50896 12960 50948 12980
rect 50948 12960 50950 12980
rect 50894 12416 50950 12472
rect 50710 11872 50766 11928
rect 51354 12552 51410 12608
rect 51262 12144 51318 12200
rect 51906 12008 51962 12064
rect 50618 9152 50674 9208
rect 50802 9152 50858 9208
rect 50986 8336 51042 8392
rect 48318 448 48374 504
rect 51170 7656 51226 7712
rect 50894 7520 50950 7576
rect 52458 9152 52514 9208
rect 51446 6840 51502 6896
rect 50894 5752 50950 5808
rect 51078 5752 51134 5808
rect 51354 5072 51410 5128
rect 51262 4156 51264 4176
rect 51264 4156 51316 4176
rect 51316 4156 51318 4176
rect 51262 4120 51318 4156
rect 50894 3712 50950 3768
rect 50802 3168 50858 3224
rect 51906 6568 51962 6624
rect 52458 6568 52514 6624
rect 53194 11872 53250 11928
rect 52734 10920 52790 10976
rect 52274 6024 52330 6080
rect 52458 6024 52514 6080
rect 52274 5752 52330 5808
rect 52458 5344 52514 5400
rect 53286 9560 53342 9616
rect 53102 9288 53158 9344
rect 53286 9288 53342 9344
rect 52918 8608 52974 8664
rect 53102 8608 53158 8664
rect 54022 11872 54078 11928
rect 53746 9560 53802 9616
rect 53838 9288 53894 9344
rect 54574 12144 54630 12200
rect 55678 12572 55734 12608
rect 55678 12552 55680 12572
rect 55680 12552 55732 12572
rect 55732 12552 55734 12572
rect 55770 12416 55826 12472
rect 55678 12280 55734 12336
rect 55218 12008 55274 12064
rect 54574 9832 54630 9888
rect 53746 5752 53802 5808
rect 53102 5344 53158 5400
rect 51814 5072 51870 5128
rect 52642 3576 52698 3632
rect 50802 1128 50858 1184
rect 55402 11736 55458 11792
rect 55126 10376 55182 10432
rect 54482 5072 54538 5128
rect 54850 5752 54906 5808
rect 55126 7656 55182 7712
rect 55034 5072 55090 5128
rect 56322 11872 56378 11928
rect 56322 11756 56378 11792
rect 56782 12416 56838 12472
rect 56641 11994 56697 11996
rect 56721 11994 56777 11996
rect 56801 11994 56857 11996
rect 56881 11994 56937 11996
rect 56641 11942 56667 11994
rect 56667 11942 56697 11994
rect 56721 11942 56731 11994
rect 56731 11942 56777 11994
rect 56801 11942 56847 11994
rect 56847 11942 56857 11994
rect 56881 11942 56911 11994
rect 56911 11942 56937 11994
rect 56641 11940 56697 11942
rect 56721 11940 56777 11942
rect 56801 11940 56857 11942
rect 56881 11940 56937 11942
rect 56322 11736 56324 11756
rect 56324 11736 56376 11756
rect 56376 11736 56378 11756
rect 56138 10784 56194 10840
rect 55954 9832 56010 9888
rect 55954 9696 56010 9752
rect 55494 7656 55550 7712
rect 56414 10920 56470 10976
rect 56641 10906 56697 10908
rect 56721 10906 56777 10908
rect 56801 10906 56857 10908
rect 56881 10906 56937 10908
rect 56641 10854 56667 10906
rect 56667 10854 56697 10906
rect 56721 10854 56731 10906
rect 56731 10854 56777 10906
rect 56801 10854 56847 10906
rect 56847 10854 56857 10906
rect 56881 10854 56911 10906
rect 56911 10854 56937 10906
rect 56641 10852 56697 10854
rect 56721 10852 56777 10854
rect 56801 10852 56857 10854
rect 56881 10852 56937 10854
rect 56322 9832 56378 9888
rect 57610 12144 57666 12200
rect 57150 10956 57152 10976
rect 57152 10956 57204 10976
rect 57204 10956 57206 10976
rect 57150 10920 57206 10956
rect 56641 9818 56697 9820
rect 56721 9818 56777 9820
rect 56801 9818 56857 9820
rect 56881 9818 56937 9820
rect 56641 9766 56667 9818
rect 56667 9766 56697 9818
rect 56721 9766 56731 9818
rect 56731 9766 56777 9818
rect 56801 9766 56847 9818
rect 56847 9766 56857 9818
rect 56881 9766 56911 9818
rect 56911 9766 56937 9818
rect 56641 9764 56697 9766
rect 56721 9764 56777 9766
rect 56801 9764 56857 9766
rect 56881 9764 56937 9766
rect 56414 9696 56470 9752
rect 56322 8744 56378 8800
rect 56506 8744 56562 8800
rect 55586 6432 55642 6488
rect 55494 5752 55550 5808
rect 55862 5752 55918 5808
rect 56641 8730 56697 8732
rect 56721 8730 56777 8732
rect 56801 8730 56857 8732
rect 56881 8730 56937 8732
rect 56641 8678 56667 8730
rect 56667 8678 56697 8730
rect 56721 8678 56731 8730
rect 56731 8678 56777 8730
rect 56801 8678 56847 8730
rect 56847 8678 56857 8730
rect 56881 8678 56911 8730
rect 56911 8678 56937 8730
rect 56641 8676 56697 8678
rect 56721 8676 56777 8678
rect 56801 8676 56857 8678
rect 56881 8676 56937 8678
rect 57150 9288 57206 9344
rect 57150 8744 57206 8800
rect 57426 10532 57482 10568
rect 57426 10512 57428 10532
rect 57428 10512 57480 10532
rect 57480 10512 57482 10532
rect 58070 12008 58126 12064
rect 57610 9832 57666 9888
rect 57334 8608 57390 8664
rect 56506 7692 56508 7712
rect 56508 7692 56560 7712
rect 56560 7692 56562 7712
rect 56506 7656 56562 7692
rect 56641 7642 56697 7644
rect 56721 7642 56777 7644
rect 56801 7642 56857 7644
rect 56881 7642 56937 7644
rect 56641 7590 56667 7642
rect 56667 7590 56697 7642
rect 56721 7590 56731 7642
rect 56731 7590 56777 7642
rect 56801 7590 56847 7642
rect 56847 7590 56857 7642
rect 56881 7590 56911 7642
rect 56911 7590 56937 7642
rect 56641 7588 56697 7590
rect 56721 7588 56777 7590
rect 56801 7588 56857 7590
rect 56881 7588 56937 7590
rect 56506 7520 56562 7576
rect 57058 7520 57114 7576
rect 56230 6568 56286 6624
rect 56046 6432 56102 6488
rect 55678 5208 55734 5264
rect 54942 1672 54998 1728
rect 53838 584 53894 640
rect 53654 448 53710 504
rect 55126 2352 55182 2408
rect 55126 1672 55182 1728
rect 56138 5208 56194 5264
rect 55678 4936 55734 4992
rect 56641 6554 56697 6556
rect 56721 6554 56777 6556
rect 56801 6554 56857 6556
rect 56881 6554 56937 6556
rect 56641 6502 56667 6554
rect 56667 6502 56697 6554
rect 56721 6502 56731 6554
rect 56731 6502 56777 6554
rect 56801 6502 56847 6554
rect 56847 6502 56857 6554
rect 56881 6502 56911 6554
rect 56911 6502 56937 6554
rect 56641 6500 56697 6502
rect 56721 6500 56777 6502
rect 56801 6500 56857 6502
rect 56881 6500 56937 6502
rect 56322 5480 56378 5536
rect 56641 5466 56697 5468
rect 56721 5466 56777 5468
rect 56801 5466 56857 5468
rect 56881 5466 56937 5468
rect 56641 5414 56667 5466
rect 56667 5414 56697 5466
rect 56721 5414 56731 5466
rect 56731 5414 56777 5466
rect 56801 5414 56847 5466
rect 56847 5414 56857 5466
rect 56881 5414 56911 5466
rect 56911 5414 56937 5466
rect 56641 5412 56697 5414
rect 56721 5412 56777 5414
rect 56801 5412 56857 5414
rect 56881 5412 56937 5414
rect 56506 5344 56562 5400
rect 56322 5208 56378 5264
rect 55494 4664 55550 4720
rect 55494 4528 55550 4584
rect 55494 2932 55496 2952
rect 55496 2932 55548 2952
rect 55548 2932 55550 2952
rect 55494 2896 55550 2932
rect 55402 2352 55458 2408
rect 55402 2080 55458 2136
rect 56046 3168 56102 3224
rect 56641 4378 56697 4380
rect 56721 4378 56777 4380
rect 56801 4378 56857 4380
rect 56881 4378 56937 4380
rect 56641 4326 56667 4378
rect 56667 4326 56697 4378
rect 56721 4326 56731 4378
rect 56731 4326 56777 4378
rect 56801 4326 56847 4378
rect 56847 4326 56857 4378
rect 56881 4326 56911 4378
rect 56911 4326 56937 4378
rect 56641 4324 56697 4326
rect 56721 4324 56777 4326
rect 56801 4324 56857 4326
rect 56881 4324 56937 4326
rect 55678 2216 55734 2272
rect 55678 856 55734 912
rect 55954 2080 56010 2136
rect 57242 7692 57244 7712
rect 57244 7692 57296 7712
rect 57296 7692 57298 7712
rect 57242 7656 57298 7692
rect 57610 9288 57666 9344
rect 58438 12008 58494 12064
rect 57426 6876 57428 6896
rect 57428 6876 57480 6896
rect 57480 6876 57482 6896
rect 57426 6840 57482 6876
rect 57334 6568 57390 6624
rect 57978 8064 58034 8120
rect 57426 5208 57482 5264
rect 57518 5072 57574 5128
rect 57242 4392 57298 4448
rect 56641 3290 56697 3292
rect 56721 3290 56777 3292
rect 56801 3290 56857 3292
rect 56881 3290 56937 3292
rect 56641 3238 56667 3290
rect 56667 3238 56697 3290
rect 56721 3238 56731 3290
rect 56731 3238 56777 3290
rect 56801 3238 56847 3290
rect 56847 3238 56857 3290
rect 56881 3238 56911 3290
rect 56911 3238 56937 3290
rect 56641 3236 56697 3238
rect 56721 3236 56777 3238
rect 56801 3236 56857 3238
rect 56881 3236 56937 3238
rect 57426 3032 57482 3088
rect 56641 2202 56697 2204
rect 56721 2202 56777 2204
rect 56801 2202 56857 2204
rect 56881 2202 56937 2204
rect 56641 2150 56667 2202
rect 56667 2150 56697 2202
rect 56721 2150 56731 2202
rect 56731 2150 56777 2202
rect 56801 2150 56847 2202
rect 56847 2150 56857 2202
rect 56881 2150 56911 2202
rect 56911 2150 56937 2202
rect 56641 2148 56697 2150
rect 56721 2148 56777 2150
rect 56801 2148 56857 2150
rect 56881 2148 56937 2150
rect 56230 992 56286 1048
rect 56641 1114 56697 1116
rect 56721 1114 56777 1116
rect 56801 1114 56857 1116
rect 56881 1114 56937 1116
rect 56641 1062 56667 1114
rect 56667 1062 56697 1114
rect 56721 1062 56731 1114
rect 56731 1062 56777 1114
rect 56801 1062 56847 1114
rect 56847 1062 56857 1114
rect 56881 1062 56911 1114
rect 56911 1062 56937 1114
rect 56641 1060 56697 1062
rect 56721 1060 56777 1062
rect 56801 1060 56857 1062
rect 56881 1060 56937 1062
rect 55494 584 55550 640
rect 55678 584 55734 640
rect 57242 2352 57298 2408
rect 57242 2216 57298 2272
rect 57242 1672 57298 1728
rect 57426 1672 57482 1728
rect 57334 856 57390 912
rect 58806 11872 58862 11928
rect 58346 8064 58402 8120
rect 59542 10240 59598 10296
rect 58346 2896 58402 2952
rect 59818 9288 59874 9344
rect 60554 12144 60610 12200
rect 60462 11736 60518 11792
rect 60646 11736 60702 11792
rect 60094 9832 60150 9888
rect 60278 9832 60334 9888
rect 62762 12552 62818 12608
rect 59910 3576 59966 3632
rect 60186 3576 60242 3632
rect 57334 584 57390 640
rect 61842 11872 61898 11928
rect 62302 12144 62358 12200
rect 63222 12280 63278 12336
rect 62578 9832 62634 9888
rect 63038 11464 63094 11520
rect 63038 9832 63094 9888
rect 60922 7520 60978 7576
rect 60922 7112 60978 7168
rect 60462 6976 60518 7032
rect 61474 6840 61530 6896
rect 60462 6704 60518 6760
rect 60830 6704 60886 6760
rect 60830 5888 60886 5944
rect 62118 5480 62174 5536
rect 62302 5208 62358 5264
rect 61566 2896 61622 2952
rect 60278 1128 60334 1184
rect 60646 1672 60702 1728
rect 60922 1672 60978 1728
rect 60462 620 60464 640
rect 60464 620 60516 640
rect 60516 620 60518 640
rect 60462 584 60518 620
rect 61198 1128 61254 1184
rect 61382 1128 61438 1184
rect 63590 11736 63646 11792
rect 63774 10240 63830 10296
rect 63682 9560 63738 9616
rect 64050 8472 64106 8528
rect 65522 12008 65578 12064
rect 66166 10920 66222 10976
rect 66626 8064 66682 8120
rect 69018 10376 69074 10432
rect 69294 11328 69350 11384
rect 69294 10376 69350 10432
rect 71502 9696 71558 9752
rect 72606 9016 72662 9072
rect 70766 8608 70822 8664
rect 69846 8200 69902 8256
rect 67546 7792 67602 7848
rect 64602 6432 64658 6488
rect 63866 5072 63922 5128
rect 63314 4800 63370 4856
rect 62854 4256 62910 4312
rect 62578 2896 62634 2952
rect 65522 6196 65524 6216
rect 65524 6196 65576 6216
rect 65576 6196 65578 6216
rect 65522 6160 65578 6196
rect 64694 5344 64750 5400
rect 63774 3576 63830 3632
rect 61198 584 61254 640
rect 65062 40 65118 96
rect 65522 1672 65578 1728
rect 66902 2896 66958 2952
rect 67454 3460 67510 3496
rect 67454 3440 67456 3460
rect 67456 3440 67508 3460
rect 67508 3440 67510 3460
rect 67454 3168 67510 3224
rect 72790 7948 72846 7984
rect 72790 7928 72792 7948
rect 72792 7928 72844 7948
rect 72844 7928 72846 7948
rect 69294 6704 69350 6760
rect 68006 1264 68062 1320
rect 65614 40 65670 96
rect 68374 2896 68430 2952
rect 68558 1672 68614 1728
rect 68742 1672 68798 1728
rect 70950 6296 71006 6352
rect 70030 4528 70086 4584
rect 69386 3848 69442 3904
rect 70122 3884 70124 3904
rect 70124 3884 70176 3904
rect 70176 3884 70178 3904
rect 70122 3848 70178 3884
rect 69570 3168 69626 3224
rect 70122 3188 70178 3224
rect 70122 3168 70124 3188
rect 70124 3168 70176 3188
rect 70176 3168 70178 3188
rect 70398 3188 70454 3224
rect 70398 3168 70400 3188
rect 70400 3168 70452 3188
rect 70452 3168 70454 3188
rect 70582 3712 70638 3768
rect 70582 3168 70638 3224
rect 70490 1672 70546 1728
rect 70030 1264 70086 1320
rect 70214 1128 70270 1184
rect 71042 2352 71098 2408
rect 71318 2372 71374 2408
rect 71318 2352 71320 2372
rect 71320 2352 71372 2372
rect 71372 2352 71374 2372
rect 71870 7248 71926 7304
rect 71686 1672 71742 1728
rect 74538 11192 74594 11248
rect 74538 9152 74594 9208
rect 76286 11056 76342 11112
rect 76378 10648 76434 10704
rect 77574 11636 77576 11656
rect 77576 11636 77628 11656
rect 77628 11636 77630 11656
rect 77574 11600 77630 11636
rect 77390 10784 77446 10840
rect 79414 10140 79416 10160
rect 79416 10140 79468 10160
rect 79468 10140 79470 10160
rect 79414 10104 79470 10140
rect 79874 11736 79930 11792
rect 77390 9988 77446 10024
rect 77390 9968 77392 9988
rect 77392 9968 77444 9988
rect 77444 9968 77446 9988
rect 76470 9324 76472 9344
rect 76472 9324 76524 9344
rect 76524 9324 76526 9344
rect 76470 9288 76526 9324
rect 82542 11756 82598 11792
rect 82542 11736 82544 11756
rect 82544 11736 82596 11756
rect 82596 11736 82598 11756
rect 81162 10548 81164 10568
rect 81164 10548 81216 10568
rect 81216 10548 81218 10568
rect 81162 10512 81218 10548
rect 80794 9460 80796 9480
rect 80796 9460 80848 9480
rect 80848 9460 80850 9480
rect 80794 9424 80850 9460
rect 84852 11450 84908 11452
rect 84932 11450 84988 11452
rect 85012 11450 85068 11452
rect 85092 11450 85148 11452
rect 84852 11398 84878 11450
rect 84878 11398 84908 11450
rect 84932 11398 84942 11450
rect 84942 11398 84988 11450
rect 85012 11398 85058 11450
rect 85058 11398 85068 11450
rect 85092 11398 85122 11450
rect 85122 11398 85148 11450
rect 84852 11396 84908 11398
rect 84932 11396 84988 11398
rect 85012 11396 85068 11398
rect 85092 11396 85148 11398
rect 84852 10362 84908 10364
rect 84932 10362 84988 10364
rect 85012 10362 85068 10364
rect 85092 10362 85148 10364
rect 84852 10310 84878 10362
rect 84878 10310 84908 10362
rect 84932 10310 84942 10362
rect 84942 10310 84988 10362
rect 85012 10310 85058 10362
rect 85058 10310 85068 10362
rect 85092 10310 85122 10362
rect 85122 10310 85148 10362
rect 84852 10308 84908 10310
rect 84932 10308 84988 10310
rect 85012 10308 85068 10310
rect 85092 10308 85148 10310
rect 84852 9274 84908 9276
rect 84932 9274 84988 9276
rect 85012 9274 85068 9276
rect 85092 9274 85148 9276
rect 84852 9222 84878 9274
rect 84878 9222 84908 9274
rect 84932 9222 84942 9274
rect 84942 9222 84988 9274
rect 85012 9222 85058 9274
rect 85058 9222 85068 9274
rect 85092 9222 85122 9274
rect 85122 9222 85148 9274
rect 84852 9220 84908 9222
rect 84932 9220 84988 9222
rect 85012 9220 85068 9222
rect 85092 9220 85148 9222
rect 85670 10548 85672 10568
rect 85672 10548 85724 10568
rect 85724 10548 85726 10568
rect 85670 10512 85726 10548
rect 81990 8900 82046 8936
rect 81990 8880 81992 8900
rect 81992 8880 82044 8900
rect 82044 8880 82046 8900
rect 85578 8744 85634 8800
rect 85670 8472 85726 8528
rect 74630 8336 74686 8392
rect 73526 7656 73582 7712
rect 73066 3848 73122 3904
rect 72054 2896 72110 2952
rect 72422 1264 72478 1320
rect 72974 3168 73030 3224
rect 74354 4120 74410 4176
rect 73802 3712 73858 3768
rect 73526 3304 73582 3360
rect 75918 2624 75974 2680
rect 75274 1672 75330 1728
rect 74998 992 75054 1048
rect 74998 720 75054 776
rect 77114 2352 77170 2408
rect 77574 2100 77630 2136
rect 77574 2080 77576 2100
rect 77576 2080 77628 2100
rect 77628 2080 77630 2100
rect 77298 1536 77354 1592
rect 77574 1128 77630 1184
rect 80794 7384 80850 7440
rect 80426 7112 80482 7168
rect 82266 2760 82322 2816
rect 88062 9832 88118 9888
rect 84852 8186 84908 8188
rect 84932 8186 84988 8188
rect 85012 8186 85068 8188
rect 85092 8186 85148 8188
rect 84852 8134 84878 8186
rect 84878 8134 84908 8186
rect 84932 8134 84942 8186
rect 84942 8134 84988 8186
rect 85012 8134 85058 8186
rect 85058 8134 85068 8186
rect 85092 8134 85122 8186
rect 85122 8134 85148 8186
rect 84852 8132 84908 8134
rect 84932 8132 84988 8134
rect 85012 8132 85068 8134
rect 85092 8132 85148 8134
rect 83186 6976 83242 7032
rect 83002 6568 83058 6624
rect 83462 1844 83464 1864
rect 83464 1844 83516 1864
rect 83516 1844 83518 1864
rect 83462 1808 83518 1844
rect 84198 1944 84254 2000
rect 84852 7098 84908 7100
rect 84932 7098 84988 7100
rect 85012 7098 85068 7100
rect 85092 7098 85148 7100
rect 84852 7046 84878 7098
rect 84878 7046 84908 7098
rect 84932 7046 84942 7098
rect 84942 7046 84988 7098
rect 85012 7046 85058 7098
rect 85058 7046 85068 7098
rect 85092 7046 85122 7098
rect 85122 7046 85148 7098
rect 84852 7044 84908 7046
rect 84932 7044 84988 7046
rect 85012 7044 85068 7046
rect 85092 7044 85148 7046
rect 84852 6010 84908 6012
rect 84932 6010 84988 6012
rect 85012 6010 85068 6012
rect 85092 6010 85148 6012
rect 84852 5958 84878 6010
rect 84878 5958 84908 6010
rect 84932 5958 84942 6010
rect 84942 5958 84988 6010
rect 85012 5958 85058 6010
rect 85058 5958 85068 6010
rect 85092 5958 85122 6010
rect 85122 5958 85148 6010
rect 84852 5956 84908 5958
rect 84932 5956 84988 5958
rect 85012 5956 85068 5958
rect 85092 5956 85148 5958
rect 84852 4922 84908 4924
rect 84932 4922 84988 4924
rect 85012 4922 85068 4924
rect 85092 4922 85148 4924
rect 84852 4870 84878 4922
rect 84878 4870 84908 4922
rect 84932 4870 84942 4922
rect 84942 4870 84988 4922
rect 85012 4870 85058 4922
rect 85058 4870 85068 4922
rect 85092 4870 85122 4922
rect 85122 4870 85148 4922
rect 84852 4868 84908 4870
rect 84932 4868 84988 4870
rect 85012 4868 85068 4870
rect 85092 4868 85148 4870
rect 84852 3834 84908 3836
rect 84932 3834 84988 3836
rect 85012 3834 85068 3836
rect 85092 3834 85148 3836
rect 84852 3782 84878 3834
rect 84878 3782 84908 3834
rect 84932 3782 84942 3834
rect 84942 3782 84988 3834
rect 85012 3782 85058 3834
rect 85058 3782 85068 3834
rect 85092 3782 85122 3834
rect 85122 3782 85148 3834
rect 84852 3780 84908 3782
rect 84932 3780 84988 3782
rect 85012 3780 85068 3782
rect 85092 3780 85148 3782
rect 85210 3576 85266 3632
rect 84852 2746 84908 2748
rect 84932 2746 84988 2748
rect 85012 2746 85068 2748
rect 85092 2746 85148 2748
rect 84852 2694 84878 2746
rect 84878 2694 84908 2746
rect 84932 2694 84942 2746
rect 84942 2694 84988 2746
rect 85012 2694 85058 2746
rect 85058 2694 85068 2746
rect 85092 2694 85122 2746
rect 85122 2694 85148 2746
rect 84852 2692 84908 2694
rect 84932 2692 84988 2694
rect 85012 2692 85068 2694
rect 85092 2692 85148 2694
rect 84852 1658 84908 1660
rect 84932 1658 84988 1660
rect 85012 1658 85068 1660
rect 85092 1658 85148 1660
rect 84852 1606 84878 1658
rect 84878 1606 84908 1658
rect 84932 1606 84942 1658
rect 84942 1606 84988 1658
rect 85012 1606 85058 1658
rect 85058 1606 85068 1658
rect 85092 1606 85122 1658
rect 85122 1606 85148 1658
rect 84852 1604 84908 1606
rect 84932 1604 84988 1606
rect 85012 1604 85068 1606
rect 85092 1604 85148 1606
rect 84290 312 84346 368
rect 84852 570 84908 572
rect 84932 570 84988 572
rect 85012 570 85068 572
rect 85092 570 85148 572
rect 84852 518 84878 570
rect 84878 518 84908 570
rect 84932 518 84942 570
rect 84942 518 84988 570
rect 85012 518 85058 570
rect 85058 518 85068 570
rect 85092 518 85122 570
rect 85122 518 85148 570
rect 84852 516 84908 518
rect 84932 516 84988 518
rect 85012 516 85068 518
rect 85092 516 85148 518
rect 86498 992 86554 1048
rect 86958 2896 87014 2952
rect 87326 2760 87382 2816
rect 87602 2644 87658 2680
rect 87602 2624 87604 2644
rect 87604 2624 87656 2644
rect 87656 2624 87658 2644
rect 88154 2216 88210 2272
rect 89442 3984 89498 4040
rect 89718 2624 89774 2680
rect 87602 856 87658 912
rect 90454 3032 90510 3088
rect 90822 5108 90824 5128
rect 90824 5108 90876 5128
rect 90876 5108 90878 5128
rect 90822 5072 90878 5108
rect 91374 2508 91430 2544
rect 91374 2488 91376 2508
rect 91376 2488 91428 2508
rect 91428 2488 91430 2508
rect 85486 40 85542 96
rect 86130 176 86186 232
rect 88982 740 89038 776
rect 88982 720 88984 740
rect 88984 720 89036 740
rect 89036 720 89038 740
rect 95146 8880 95202 8936
rect 95146 8472 95202 8528
rect 97538 10784 97594 10840
rect 98366 9868 98368 9888
rect 98368 9868 98420 9888
rect 98420 9868 98422 9888
rect 98366 9832 98422 9868
rect 97814 9560 97870 9616
rect 96618 6976 96674 7032
rect 99286 6432 99342 6488
rect 98274 5888 98330 5944
rect 95054 2896 95110 2952
rect 95146 2760 95202 2816
rect 99562 4120 99618 4176
rect 98826 1672 98882 1728
rect 98090 1128 98146 1184
rect 100666 5752 100722 5808
rect 100390 1672 100446 1728
rect 100942 5072 100998 5128
rect 101402 5480 101458 5536
rect 101034 4664 101090 4720
rect 102230 9832 102286 9888
rect 103242 9560 103298 9616
rect 103334 6196 103336 6216
rect 103336 6196 103388 6216
rect 103388 6196 103390 6216
rect 103334 6160 103390 6196
rect 104070 6976 104126 7032
rect 103978 6568 104034 6624
rect 103426 6024 103482 6080
rect 103426 5888 103482 5944
rect 103610 5888 103666 5944
rect 101402 992 101458 1048
rect 106186 10804 106242 10840
rect 106186 10784 106188 10804
rect 106188 10784 106240 10804
rect 106240 10784 106242 10804
rect 104714 6452 104770 6488
rect 104714 6432 104716 6452
rect 104716 6432 104768 6452
rect 104768 6432 104770 6452
rect 104714 6024 104770 6080
rect 104438 5480 104494 5536
rect 107198 10240 107254 10296
rect 106370 6432 106426 6488
rect 106370 5888 106426 5944
rect 106094 5092 106150 5128
rect 106094 5072 106096 5092
rect 106096 5072 106148 5092
rect 106148 5072 106150 5092
rect 106186 4664 106242 4720
rect 103518 1420 103574 1456
rect 103518 1400 103520 1420
rect 103520 1400 103572 1420
rect 103572 1400 103574 1420
rect 103702 584 103758 640
rect 104898 1128 104954 1184
rect 104806 992 104862 1048
rect 108210 9580 108266 9616
rect 108210 9560 108212 9580
rect 108212 9560 108264 9580
rect 108264 9560 108266 9580
rect 108118 9172 108174 9208
rect 108118 9152 108120 9172
rect 108120 9152 108172 9172
rect 108172 9152 108174 9172
rect 108854 10532 108910 10568
rect 108854 10512 108856 10532
rect 108856 10512 108908 10532
rect 108908 10512 108910 10532
rect 108670 9016 108726 9072
rect 107750 6568 107806 6624
rect 107842 6432 107898 6488
rect 106738 5888 106794 5944
rect 106646 2760 106702 2816
rect 106370 1536 106426 1592
rect 106370 856 106426 912
rect 107566 4004 107622 4040
rect 107566 3984 107568 4004
rect 107568 3984 107620 4004
rect 107620 3984 107622 4004
rect 107474 3848 107530 3904
rect 107566 3440 107622 3496
rect 108302 6196 108304 6216
rect 108304 6196 108356 6216
rect 108356 6196 108358 6216
rect 108302 6160 108358 6196
rect 108394 4120 108450 4176
rect 108026 3576 108082 3632
rect 108394 3440 108450 3496
rect 107658 2624 107714 2680
rect 108578 3032 108634 3088
rect 107290 1400 107346 1456
rect 106738 856 106794 912
rect 106370 620 106372 640
rect 106372 620 106424 640
rect 106424 620 106426 640
rect 106370 584 106426 620
rect 108946 6704 109002 6760
rect 107014 720 107070 776
rect 109314 4020 109316 4040
rect 109316 4020 109368 4040
rect 109368 4020 109370 4040
rect 109314 3984 109370 4020
rect 108946 3884 108948 3904
rect 108948 3884 109000 3904
rect 109000 3884 109002 3904
rect 108946 3848 109002 3884
rect 109038 3032 109094 3088
rect 108854 2916 108910 2952
rect 108854 2896 108856 2916
rect 108856 2896 108908 2916
rect 108908 2896 108910 2916
rect 109130 2932 109132 2952
rect 109132 2932 109184 2952
rect 109184 2932 109186 2952
rect 109130 2896 109186 2932
rect 109406 2896 109462 2952
rect 110142 10104 110198 10160
rect 110418 6976 110474 7032
rect 109038 1300 109040 1320
rect 109040 1300 109092 1320
rect 109092 1300 109094 1320
rect 109038 1264 109094 1300
rect 109038 1164 109040 1184
rect 109040 1164 109092 1184
rect 109092 1164 109094 1184
rect 109038 1128 109094 1164
rect 109038 856 109094 912
rect 109682 1164 109684 1184
rect 109684 1164 109736 1184
rect 109736 1164 109738 1184
rect 109682 1128 109738 1164
rect 108486 584 108542 640
rect 113062 11994 113118 11996
rect 113142 11994 113198 11996
rect 113222 11994 113278 11996
rect 113302 11994 113358 11996
rect 113062 11942 113088 11994
rect 113088 11942 113118 11994
rect 113142 11942 113152 11994
rect 113152 11942 113198 11994
rect 113222 11942 113268 11994
rect 113268 11942 113278 11994
rect 113302 11942 113332 11994
rect 113332 11942 113358 11994
rect 113062 11940 113118 11942
rect 113142 11940 113198 11942
rect 113222 11940 113278 11942
rect 113302 11940 113358 11942
rect 113062 10906 113118 10908
rect 113142 10906 113198 10908
rect 113222 10906 113278 10908
rect 113302 10906 113358 10908
rect 113062 10854 113088 10906
rect 113088 10854 113118 10906
rect 113142 10854 113152 10906
rect 113152 10854 113198 10906
rect 113222 10854 113268 10906
rect 113268 10854 113278 10906
rect 113302 10854 113332 10906
rect 113332 10854 113358 10906
rect 113062 10852 113118 10854
rect 113142 10852 113198 10854
rect 113222 10852 113278 10854
rect 113302 10852 113358 10854
rect 112994 10512 113050 10568
rect 111062 2896 111118 2952
rect 111062 992 111118 1048
rect 111338 992 111394 1048
rect 112166 1536 112222 1592
rect 113062 9818 113118 9820
rect 113142 9818 113198 9820
rect 113222 9818 113278 9820
rect 113302 9818 113358 9820
rect 113062 9766 113088 9818
rect 113088 9766 113118 9818
rect 113142 9766 113152 9818
rect 113152 9766 113198 9818
rect 113222 9766 113268 9818
rect 113268 9766 113278 9818
rect 113302 9766 113332 9818
rect 113332 9766 113358 9818
rect 113062 9764 113118 9766
rect 113142 9764 113198 9766
rect 113222 9764 113278 9766
rect 113302 9764 113358 9766
rect 115018 11600 115074 11656
rect 116490 11500 116492 11520
rect 116492 11500 116544 11520
rect 116544 11500 116546 11520
rect 116490 11464 116546 11500
rect 116950 11328 117006 11384
rect 117042 10648 117098 10704
rect 113546 9596 113548 9616
rect 113548 9596 113600 9616
rect 113600 9596 113602 9616
rect 113546 9560 113602 9596
rect 115662 9152 115718 9208
rect 113062 8730 113118 8732
rect 113142 8730 113198 8732
rect 113222 8730 113278 8732
rect 113302 8730 113358 8732
rect 113062 8678 113088 8730
rect 113088 8678 113118 8730
rect 113142 8678 113152 8730
rect 113152 8678 113198 8730
rect 113222 8678 113268 8730
rect 113268 8678 113278 8730
rect 113302 8678 113332 8730
rect 113332 8678 113358 8730
rect 113062 8676 113118 8678
rect 113142 8676 113198 8678
rect 113222 8676 113278 8678
rect 113302 8676 113358 8678
rect 112902 7656 112958 7712
rect 113062 7642 113118 7644
rect 113142 7642 113198 7644
rect 113222 7642 113278 7644
rect 113302 7642 113358 7644
rect 113062 7590 113088 7642
rect 113088 7590 113118 7642
rect 113142 7590 113152 7642
rect 113152 7590 113198 7642
rect 113222 7590 113268 7642
rect 113268 7590 113278 7642
rect 113302 7590 113332 7642
rect 113332 7590 113358 7642
rect 113062 7588 113118 7590
rect 113142 7588 113198 7590
rect 113222 7588 113278 7590
rect 113302 7588 113358 7590
rect 113086 7384 113142 7440
rect 114558 7520 114614 7576
rect 114374 7384 114430 7440
rect 113638 6724 113694 6760
rect 113638 6704 113640 6724
rect 113640 6704 113692 6724
rect 113692 6704 113694 6724
rect 113062 6554 113118 6556
rect 113142 6554 113198 6556
rect 113222 6554 113278 6556
rect 113302 6554 113358 6556
rect 113062 6502 113088 6554
rect 113088 6502 113118 6554
rect 113142 6502 113152 6554
rect 113152 6502 113198 6554
rect 113222 6502 113268 6554
rect 113268 6502 113278 6554
rect 113302 6502 113332 6554
rect 113332 6502 113358 6554
rect 113062 6500 113118 6502
rect 113142 6500 113198 6502
rect 113222 6500 113278 6502
rect 113302 6500 113358 6502
rect 113062 5466 113118 5468
rect 113142 5466 113198 5468
rect 113222 5466 113278 5468
rect 113302 5466 113358 5468
rect 113062 5414 113088 5466
rect 113088 5414 113118 5466
rect 113142 5414 113152 5466
rect 113152 5414 113198 5466
rect 113222 5414 113268 5466
rect 113268 5414 113278 5466
rect 113302 5414 113332 5466
rect 113332 5414 113358 5466
rect 113062 5412 113118 5414
rect 113142 5412 113198 5414
rect 113222 5412 113278 5414
rect 113302 5412 113358 5414
rect 112626 1672 112682 1728
rect 113062 4378 113118 4380
rect 113142 4378 113198 4380
rect 113222 4378 113278 4380
rect 113302 4378 113358 4380
rect 113062 4326 113088 4378
rect 113088 4326 113118 4378
rect 113142 4326 113152 4378
rect 113152 4326 113198 4378
rect 113222 4326 113268 4378
rect 113268 4326 113278 4378
rect 113302 4326 113332 4378
rect 113332 4326 113358 4378
rect 113062 4324 113118 4326
rect 113142 4324 113198 4326
rect 113222 4324 113278 4326
rect 113302 4324 113358 4326
rect 113062 3290 113118 3292
rect 113142 3290 113198 3292
rect 113222 3290 113278 3292
rect 113302 3290 113358 3292
rect 113062 3238 113088 3290
rect 113088 3238 113118 3290
rect 113142 3238 113152 3290
rect 113152 3238 113198 3290
rect 113222 3238 113268 3290
rect 113268 3238 113278 3290
rect 113302 3238 113332 3290
rect 113332 3238 113358 3290
rect 113062 3236 113118 3238
rect 113142 3236 113198 3238
rect 113222 3236 113278 3238
rect 113302 3236 113358 3238
rect 114466 2760 114522 2816
rect 113062 2202 113118 2204
rect 113142 2202 113198 2204
rect 113222 2202 113278 2204
rect 113302 2202 113358 2204
rect 113062 2150 113088 2202
rect 113088 2150 113118 2202
rect 113142 2150 113152 2202
rect 113152 2150 113198 2202
rect 113222 2150 113268 2202
rect 113268 2150 113278 2202
rect 113302 2150 113332 2202
rect 113332 2150 113358 2202
rect 113062 2148 113118 2150
rect 113142 2148 113198 2150
rect 113222 2148 113278 2150
rect 113302 2148 113358 2150
rect 113062 1114 113118 1116
rect 113142 1114 113198 1116
rect 113222 1114 113278 1116
rect 113302 1114 113358 1116
rect 113062 1062 113088 1114
rect 113088 1062 113118 1114
rect 113142 1062 113152 1114
rect 113152 1062 113198 1114
rect 113222 1062 113268 1114
rect 113268 1062 113278 1114
rect 113302 1062 113332 1114
rect 113332 1062 113358 1114
rect 113062 1060 113118 1062
rect 113142 1060 113198 1062
rect 113222 1060 113278 1062
rect 113302 1060 113358 1062
rect 113546 1264 113602 1320
rect 114466 1672 114522 1728
rect 114098 584 114154 640
rect 122562 11600 122618 11656
rect 122930 11328 122986 11384
rect 120538 10648 120594 10704
rect 121182 10512 121238 10568
rect 119250 9596 119252 9616
rect 119252 9596 119304 9616
rect 119304 9596 119306 9616
rect 119250 9560 119306 9596
rect 118146 9288 118202 9344
rect 116122 7828 116124 7848
rect 116124 7828 116176 7848
rect 116176 7828 116178 7848
rect 116122 7792 116178 7828
rect 116950 7792 117006 7848
rect 115018 3576 115074 3632
rect 115386 2624 115442 2680
rect 122470 9560 122526 9616
rect 124770 11464 124826 11520
rect 124770 9288 124826 9344
rect 118606 6740 118608 6760
rect 118608 6740 118660 6760
rect 118660 6740 118662 6760
rect 118606 6704 118662 6740
rect 118054 2524 118056 2544
rect 118056 2524 118108 2544
rect 118108 2524 118110 2544
rect 118054 2488 118110 2524
rect 118054 992 118110 1048
rect 118790 1672 118846 1728
rect 119066 992 119122 1048
rect 120722 2524 120724 2544
rect 120724 2524 120776 2544
rect 120776 2524 120778 2544
rect 120722 2488 120778 2524
rect 122746 7520 122802 7576
rect 122746 7248 122802 7304
rect 123022 6724 123078 6760
rect 123022 6704 123024 6724
rect 123024 6704 123076 6724
rect 123076 6704 123078 6724
rect 124126 6060 124128 6080
rect 124128 6060 124180 6080
rect 124180 6060 124182 6080
rect 124126 6024 124182 6060
rect 125598 992 125654 1048
rect 126150 992 126206 1048
rect 129002 10240 129058 10296
rect 131118 9036 131174 9072
rect 131118 9016 131120 9036
rect 131120 9016 131172 9036
rect 131172 9016 131174 9036
rect 133418 10124 133474 10160
rect 133418 10104 133420 10124
rect 133420 10104 133472 10124
rect 133472 10104 133474 10124
rect 132406 8880 132462 8936
rect 132682 8880 132738 8936
rect 131762 856 131818 912
rect 137834 9988 137890 10024
rect 137834 9968 137836 9988
rect 137836 9968 137888 9988
rect 137888 9968 137890 9988
rect 141273 11450 141329 11452
rect 141353 11450 141409 11452
rect 141433 11450 141489 11452
rect 141513 11450 141569 11452
rect 141273 11398 141299 11450
rect 141299 11398 141329 11450
rect 141353 11398 141363 11450
rect 141363 11398 141409 11450
rect 141433 11398 141479 11450
rect 141479 11398 141489 11450
rect 141513 11398 141543 11450
rect 141543 11398 141569 11450
rect 141273 11396 141329 11398
rect 141353 11396 141409 11398
rect 141433 11396 141489 11398
rect 141513 11396 141569 11398
rect 140778 10512 140834 10568
rect 141273 10362 141329 10364
rect 141353 10362 141409 10364
rect 141433 10362 141489 10364
rect 141513 10362 141569 10364
rect 141273 10310 141299 10362
rect 141299 10310 141329 10362
rect 141353 10310 141363 10362
rect 141363 10310 141409 10362
rect 141433 10310 141479 10362
rect 141479 10310 141489 10362
rect 141513 10310 141543 10362
rect 141543 10310 141569 10362
rect 141273 10308 141329 10310
rect 141353 10308 141409 10310
rect 141433 10308 141489 10310
rect 141513 10308 141569 10310
rect 142158 9968 142214 10024
rect 141273 9274 141329 9276
rect 141353 9274 141409 9276
rect 141433 9274 141489 9276
rect 141513 9274 141569 9276
rect 141273 9222 141299 9274
rect 141299 9222 141329 9274
rect 141353 9222 141363 9274
rect 141363 9222 141409 9274
rect 141433 9222 141479 9274
rect 141479 9222 141489 9274
rect 141513 9222 141543 9274
rect 141543 9222 141569 9274
rect 141273 9220 141329 9222
rect 141353 9220 141409 9222
rect 141433 9220 141489 9222
rect 141513 9220 141569 9222
rect 141273 8186 141329 8188
rect 141353 8186 141409 8188
rect 141433 8186 141489 8188
rect 141513 8186 141569 8188
rect 141273 8134 141299 8186
rect 141299 8134 141329 8186
rect 141353 8134 141363 8186
rect 141363 8134 141409 8186
rect 141433 8134 141479 8186
rect 141479 8134 141489 8186
rect 141513 8134 141543 8186
rect 141543 8134 141569 8186
rect 141273 8132 141329 8134
rect 141353 8132 141409 8134
rect 141433 8132 141489 8134
rect 141513 8132 141569 8134
rect 141273 7098 141329 7100
rect 141353 7098 141409 7100
rect 141433 7098 141489 7100
rect 141513 7098 141569 7100
rect 141273 7046 141299 7098
rect 141299 7046 141329 7098
rect 141353 7046 141363 7098
rect 141363 7046 141409 7098
rect 141433 7046 141479 7098
rect 141479 7046 141489 7098
rect 141513 7046 141543 7098
rect 141543 7046 141569 7098
rect 141273 7044 141329 7046
rect 141353 7044 141409 7046
rect 141433 7044 141489 7046
rect 141513 7044 141569 7046
rect 136178 6976 136234 7032
rect 133878 1012 133934 1048
rect 133878 992 133880 1012
rect 133880 992 133932 1012
rect 133932 992 133934 1012
rect 145378 9560 145434 9616
rect 141273 6010 141329 6012
rect 141353 6010 141409 6012
rect 141433 6010 141489 6012
rect 141513 6010 141569 6012
rect 141273 5958 141299 6010
rect 141299 5958 141329 6010
rect 141353 5958 141363 6010
rect 141363 5958 141409 6010
rect 141433 5958 141479 6010
rect 141479 5958 141489 6010
rect 141513 5958 141543 6010
rect 141543 5958 141569 6010
rect 141273 5956 141329 5958
rect 141353 5956 141409 5958
rect 141433 5956 141489 5958
rect 141513 5956 141569 5958
rect 141273 4922 141329 4924
rect 141353 4922 141409 4924
rect 141433 4922 141489 4924
rect 141513 4922 141569 4924
rect 141273 4870 141299 4922
rect 141299 4870 141329 4922
rect 141353 4870 141363 4922
rect 141363 4870 141409 4922
rect 141433 4870 141479 4922
rect 141479 4870 141489 4922
rect 141513 4870 141543 4922
rect 141543 4870 141569 4922
rect 141273 4868 141329 4870
rect 141353 4868 141409 4870
rect 141433 4868 141489 4870
rect 141513 4868 141569 4870
rect 135994 856 136050 912
rect 133970 584 134026 640
rect 137926 584 137982 640
rect 141273 3834 141329 3836
rect 141353 3834 141409 3836
rect 141433 3834 141489 3836
rect 141513 3834 141569 3836
rect 141273 3782 141299 3834
rect 141299 3782 141329 3834
rect 141353 3782 141363 3834
rect 141363 3782 141409 3834
rect 141433 3782 141479 3834
rect 141479 3782 141489 3834
rect 141513 3782 141543 3834
rect 141543 3782 141569 3834
rect 141273 3780 141329 3782
rect 141353 3780 141409 3782
rect 141433 3780 141489 3782
rect 141513 3780 141569 3782
rect 141273 2746 141329 2748
rect 141353 2746 141409 2748
rect 141433 2746 141489 2748
rect 141513 2746 141569 2748
rect 141273 2694 141299 2746
rect 141299 2694 141329 2746
rect 141353 2694 141363 2746
rect 141363 2694 141409 2746
rect 141433 2694 141479 2746
rect 141479 2694 141489 2746
rect 141513 2694 141543 2746
rect 141543 2694 141569 2746
rect 141273 2692 141329 2694
rect 141353 2692 141409 2694
rect 141433 2692 141489 2694
rect 141513 2692 141569 2694
rect 141273 1658 141329 1660
rect 141353 1658 141409 1660
rect 141433 1658 141489 1660
rect 141513 1658 141569 1660
rect 141273 1606 141299 1658
rect 141299 1606 141329 1658
rect 141353 1606 141363 1658
rect 141363 1606 141409 1658
rect 141433 1606 141479 1658
rect 141479 1606 141489 1658
rect 141513 1606 141543 1658
rect 141543 1606 141569 1658
rect 141273 1604 141329 1606
rect 141353 1604 141409 1606
rect 141433 1604 141489 1606
rect 141513 1604 141569 1606
rect 141273 570 141329 572
rect 141353 570 141409 572
rect 141433 570 141489 572
rect 141513 570 141569 572
rect 141273 518 141299 570
rect 141299 518 141329 570
rect 141353 518 141363 570
rect 141363 518 141409 570
rect 141433 518 141479 570
rect 141479 518 141489 570
rect 141513 518 141543 570
rect 141543 518 141569 570
rect 141273 516 141329 518
rect 141353 516 141409 518
rect 141433 516 141489 518
rect 141513 516 141569 518
rect 146206 8744 146262 8800
rect 146850 8880 146906 8936
rect 148322 7384 148378 7440
rect 148322 7112 148378 7168
rect 150714 8744 150770 8800
rect 153014 8880 153070 8936
rect 153290 9560 153346 9616
rect 154578 6196 154580 6216
rect 154580 6196 154632 6216
rect 154632 6196 154634 6216
rect 154578 6160 154634 6196
rect 155498 6160 155554 6216
rect 156786 1420 156842 1456
rect 156786 1400 156788 1420
rect 156788 1400 156840 1420
rect 156840 1400 156842 1420
rect 159362 2488 159418 2544
rect 164790 8744 164846 8800
rect 165986 756 165988 776
rect 165988 756 166040 776
rect 166040 756 166042 776
rect 165986 720 166042 756
<< metal3 >>
rect 33685 13018 33751 13021
rect 41137 13018 41203 13021
rect 33685 13016 41203 13018
rect 33685 12960 33690 13016
rect 33746 12960 41142 13016
rect 41198 12960 41203 13016
rect 33685 12958 41203 12960
rect 33685 12955 33751 12958
rect 41137 12955 41203 12958
rect 50889 13018 50955 13021
rect 60038 13018 60044 13020
rect 50889 13016 60044 13018
rect 50889 12960 50894 13016
rect 50950 12960 60044 13016
rect 50889 12958 60044 12960
rect 50889 12955 50955 12958
rect 60038 12956 60044 12958
rect 60108 12956 60114 13020
rect 30649 12882 30715 12885
rect 35617 12882 35683 12885
rect 30649 12880 35683 12882
rect 30649 12824 30654 12880
rect 30710 12824 35622 12880
rect 35678 12824 35683 12880
rect 30649 12822 35683 12824
rect 30649 12819 30715 12822
rect 35617 12819 35683 12822
rect 35893 12882 35959 12885
rect 40401 12882 40467 12885
rect 35893 12880 40467 12882
rect 35893 12824 35898 12880
rect 35954 12824 40406 12880
rect 40462 12824 40467 12880
rect 35893 12822 40467 12824
rect 35893 12819 35959 12822
rect 40401 12819 40467 12822
rect 40585 12882 40651 12885
rect 46289 12882 46355 12885
rect 40585 12880 46355 12882
rect 40585 12824 40590 12880
rect 40646 12824 46294 12880
rect 46350 12824 46355 12880
rect 40585 12822 46355 12824
rect 40585 12819 40651 12822
rect 46289 12819 46355 12822
rect 33961 12746 34027 12749
rect 40769 12746 40835 12749
rect 33961 12744 40835 12746
rect 33961 12688 33966 12744
rect 34022 12688 40774 12744
rect 40830 12688 40835 12744
rect 33961 12686 40835 12688
rect 33961 12683 34027 12686
rect 40769 12683 40835 12686
rect 41413 12746 41479 12749
rect 42517 12746 42583 12749
rect 41413 12744 42583 12746
rect 41413 12688 41418 12744
rect 41474 12688 42522 12744
rect 42578 12688 42583 12744
rect 41413 12686 42583 12688
rect 41413 12683 41479 12686
rect 42517 12683 42583 12686
rect 43161 12746 43227 12749
rect 46473 12746 46539 12749
rect 43161 12744 46539 12746
rect 43161 12688 43166 12744
rect 43222 12688 46478 12744
rect 46534 12688 46539 12744
rect 43161 12686 46539 12688
rect 43161 12683 43227 12686
rect 46473 12683 46539 12686
rect 33593 12610 33659 12613
rect 40677 12610 40743 12613
rect 33593 12608 40743 12610
rect 33593 12552 33598 12608
rect 33654 12552 40682 12608
rect 40738 12552 40743 12608
rect 33593 12550 40743 12552
rect 33593 12547 33659 12550
rect 40677 12547 40743 12550
rect 40953 12610 41019 12613
rect 41505 12610 41571 12613
rect 40953 12608 41571 12610
rect 40953 12552 40958 12608
rect 41014 12552 41510 12608
rect 41566 12552 41571 12608
rect 40953 12550 41571 12552
rect 40953 12547 41019 12550
rect 41505 12547 41571 12550
rect 41689 12610 41755 12613
rect 46473 12610 46539 12613
rect 41689 12608 46539 12610
rect 41689 12552 41694 12608
rect 41750 12552 46478 12608
rect 46534 12552 46539 12608
rect 41689 12550 46539 12552
rect 41689 12547 41755 12550
rect 46473 12547 46539 12550
rect 48497 12610 48563 12613
rect 51349 12610 51415 12613
rect 48497 12608 51415 12610
rect 48497 12552 48502 12608
rect 48558 12552 51354 12608
rect 51410 12552 51415 12608
rect 48497 12550 51415 12552
rect 48497 12547 48563 12550
rect 51349 12547 51415 12550
rect 55673 12610 55739 12613
rect 62757 12610 62823 12613
rect 55673 12608 62823 12610
rect 55673 12552 55678 12608
rect 55734 12552 62762 12608
rect 62818 12552 62823 12608
rect 55673 12550 62823 12552
rect 55673 12547 55739 12550
rect 62757 12547 62823 12550
rect 36721 12474 36787 12477
rect 50889 12474 50955 12477
rect 36721 12472 50955 12474
rect 36721 12416 36726 12472
rect 36782 12416 50894 12472
rect 50950 12416 50955 12472
rect 36721 12414 50955 12416
rect 36721 12411 36787 12414
rect 50889 12411 50955 12414
rect 55765 12474 55831 12477
rect 56777 12474 56843 12477
rect 55765 12472 56843 12474
rect 55765 12416 55770 12472
rect 55826 12416 56782 12472
rect 56838 12416 56843 12472
rect 55765 12414 56843 12416
rect 55765 12411 55831 12414
rect 56777 12411 56843 12414
rect 33777 12338 33843 12341
rect 40401 12338 40467 12341
rect 33777 12336 40467 12338
rect 33777 12280 33782 12336
rect 33838 12280 40406 12336
rect 40462 12280 40467 12336
rect 33777 12278 40467 12280
rect 33777 12275 33843 12278
rect 40401 12275 40467 12278
rect 40677 12338 40743 12341
rect 45093 12338 45159 12341
rect 40677 12336 45159 12338
rect 40677 12280 40682 12336
rect 40738 12280 45098 12336
rect 45154 12280 45159 12336
rect 40677 12278 45159 12280
rect 40677 12275 40743 12278
rect 45093 12275 45159 12278
rect 55673 12338 55739 12341
rect 63217 12338 63283 12341
rect 55673 12336 63283 12338
rect 55673 12280 55678 12336
rect 55734 12280 63222 12336
rect 63278 12280 63283 12336
rect 55673 12278 63283 12280
rect 55673 12275 55739 12278
rect 63217 12275 63283 12278
rect 26601 12202 26667 12205
rect 33409 12202 33475 12205
rect 26601 12200 33475 12202
rect 26601 12144 26606 12200
rect 26662 12144 33414 12200
rect 33470 12144 33475 12200
rect 26601 12142 33475 12144
rect 26601 12139 26667 12142
rect 33409 12139 33475 12142
rect 34421 12202 34487 12205
rect 40309 12202 40375 12205
rect 41413 12202 41479 12205
rect 34421 12200 40375 12202
rect 34421 12144 34426 12200
rect 34482 12144 40314 12200
rect 40370 12144 40375 12200
rect 34421 12142 40375 12144
rect 34421 12139 34487 12142
rect 40309 12139 40375 12142
rect 40542 12200 41479 12202
rect 40542 12144 41418 12200
rect 41474 12144 41479 12200
rect 40542 12142 41479 12144
rect 0 12066 800 12096
rect 3693 12066 3759 12069
rect 0 12064 3759 12066
rect 0 12008 3698 12064
rect 3754 12008 3759 12064
rect 0 12006 3759 12008
rect 0 11976 800 12006
rect 3693 12003 3759 12006
rect 25037 12066 25103 12069
rect 31109 12066 31175 12069
rect 25037 12064 31175 12066
rect 25037 12008 25042 12064
rect 25098 12008 31114 12064
rect 31170 12008 31175 12064
rect 25037 12006 31175 12008
rect 25037 12003 25103 12006
rect 31109 12003 31175 12006
rect 33225 12066 33291 12069
rect 39665 12066 39731 12069
rect 33225 12064 39731 12066
rect 33225 12008 33230 12064
rect 33286 12008 39670 12064
rect 39726 12008 39731 12064
rect 33225 12006 39731 12008
rect 33225 12003 33291 12006
rect 39665 12003 39731 12006
rect 39849 12066 39915 12069
rect 40542 12066 40602 12142
rect 41413 12139 41479 12142
rect 42149 12202 42215 12205
rect 48497 12202 48563 12205
rect 42149 12200 48563 12202
rect 42149 12144 42154 12200
rect 42210 12144 48502 12200
rect 48558 12144 48563 12200
rect 42149 12142 48563 12144
rect 42149 12139 42215 12142
rect 48497 12139 48563 12142
rect 50613 12202 50679 12205
rect 51257 12202 51323 12205
rect 50613 12200 51323 12202
rect 50613 12144 50618 12200
rect 50674 12144 51262 12200
rect 51318 12144 51323 12200
rect 50613 12142 51323 12144
rect 50613 12139 50679 12142
rect 51257 12139 51323 12142
rect 54569 12202 54635 12205
rect 57605 12202 57671 12205
rect 54569 12200 57671 12202
rect 54569 12144 54574 12200
rect 54630 12144 57610 12200
rect 57666 12144 57671 12200
rect 54569 12142 57671 12144
rect 54569 12139 54635 12142
rect 57605 12139 57671 12142
rect 60549 12202 60615 12205
rect 62297 12202 62363 12205
rect 60549 12200 62363 12202
rect 60549 12144 60554 12200
rect 60610 12144 62302 12200
rect 62358 12144 62363 12200
rect 60549 12142 62363 12144
rect 60549 12139 60615 12142
rect 62297 12139 62363 12142
rect 39849 12064 40602 12066
rect 39849 12008 39854 12064
rect 39910 12008 40602 12064
rect 39849 12006 40602 12008
rect 40677 12066 40743 12069
rect 41597 12066 41663 12069
rect 40677 12064 41663 12066
rect 40677 12008 40682 12064
rect 40738 12008 41602 12064
rect 41658 12008 41663 12064
rect 40677 12006 41663 12008
rect 39849 12003 39915 12006
rect 40677 12003 40743 12006
rect 41597 12003 41663 12006
rect 42241 12066 42307 12069
rect 51901 12066 51967 12069
rect 42241 12064 51967 12066
rect 42241 12008 42246 12064
rect 42302 12008 51906 12064
rect 51962 12008 51967 12064
rect 42241 12006 51967 12008
rect 42241 12003 42307 12006
rect 51901 12003 51967 12006
rect 55213 12066 55279 12069
rect 55438 12066 55444 12068
rect 55213 12064 55444 12066
rect 55213 12008 55218 12064
rect 55274 12008 55444 12064
rect 55213 12006 55444 12008
rect 55213 12003 55279 12006
rect 55438 12004 55444 12006
rect 55508 12004 55514 12068
rect 58065 12066 58131 12069
rect 58433 12066 58499 12069
rect 65517 12066 65583 12069
rect 58065 12064 65583 12066
rect 58065 12008 58070 12064
rect 58126 12008 58438 12064
rect 58494 12008 65522 12064
rect 65578 12008 65583 12064
rect 58065 12006 65583 12008
rect 58065 12003 58131 12006
rect 58433 12003 58499 12006
rect 65517 12003 65583 12006
rect 56629 12000 56949 12001
rect 56629 11936 56637 12000
rect 56701 11936 56717 12000
rect 56781 11936 56797 12000
rect 56861 11936 56877 12000
rect 56941 11936 56949 12000
rect 56629 11935 56949 11936
rect 113050 12000 113370 12001
rect 113050 11936 113058 12000
rect 113122 11936 113138 12000
rect 113202 11936 113218 12000
rect 113282 11936 113298 12000
rect 113362 11936 113370 12000
rect 113050 11935 113370 11936
rect 24669 11930 24735 11933
rect 31201 11930 31267 11933
rect 24669 11928 31267 11930
rect 24669 11872 24674 11928
rect 24730 11872 31206 11928
rect 31262 11872 31267 11928
rect 24669 11870 31267 11872
rect 24669 11867 24735 11870
rect 31201 11867 31267 11870
rect 31477 11930 31543 11933
rect 35985 11930 36051 11933
rect 31477 11928 36051 11930
rect 31477 11872 31482 11928
rect 31538 11872 35990 11928
rect 36046 11872 36051 11928
rect 31477 11870 36051 11872
rect 31477 11867 31543 11870
rect 35985 11867 36051 11870
rect 36261 11930 36327 11933
rect 42333 11930 42399 11933
rect 36261 11928 42399 11930
rect 36261 11872 36266 11928
rect 36322 11872 42338 11928
rect 42394 11872 42399 11928
rect 36261 11870 42399 11872
rect 36261 11867 36327 11870
rect 42333 11867 42399 11870
rect 43713 11930 43779 11933
rect 46565 11930 46631 11933
rect 43713 11928 46631 11930
rect 43713 11872 43718 11928
rect 43774 11872 46570 11928
rect 46626 11872 46631 11928
rect 43713 11870 46631 11872
rect 43713 11867 43779 11870
rect 46565 11867 46631 11870
rect 50705 11930 50771 11933
rect 53189 11930 53255 11933
rect 50705 11928 53255 11930
rect 50705 11872 50710 11928
rect 50766 11872 53194 11928
rect 53250 11872 53255 11928
rect 50705 11870 53255 11872
rect 50705 11867 50771 11870
rect 53189 11867 53255 11870
rect 54017 11930 54083 11933
rect 56317 11930 56383 11933
rect 54017 11928 56383 11930
rect 54017 11872 54022 11928
rect 54078 11872 56322 11928
rect 56378 11872 56383 11928
rect 54017 11870 56383 11872
rect 54017 11867 54083 11870
rect 56317 11867 56383 11870
rect 58801 11930 58867 11933
rect 61837 11930 61903 11933
rect 58801 11928 61903 11930
rect 58801 11872 58806 11928
rect 58862 11872 61842 11928
rect 61898 11872 61903 11928
rect 58801 11870 61903 11872
rect 58801 11867 58867 11870
rect 61837 11867 61903 11870
rect 16481 11794 16547 11797
rect 44081 11794 44147 11797
rect 16481 11792 44147 11794
rect 16481 11736 16486 11792
rect 16542 11736 44086 11792
rect 44142 11736 44147 11792
rect 16481 11734 44147 11736
rect 16481 11731 16547 11734
rect 44081 11731 44147 11734
rect 45737 11794 45803 11797
rect 55397 11794 55463 11797
rect 45737 11792 55463 11794
rect 45737 11736 45742 11792
rect 45798 11736 55402 11792
rect 55458 11736 55463 11792
rect 45737 11734 55463 11736
rect 45737 11731 45803 11734
rect 55397 11731 55463 11734
rect 56317 11794 56383 11797
rect 60457 11794 60523 11797
rect 56317 11792 60523 11794
rect 56317 11736 56322 11792
rect 56378 11736 60462 11792
rect 60518 11736 60523 11792
rect 56317 11734 60523 11736
rect 56317 11731 56383 11734
rect 60457 11731 60523 11734
rect 60641 11794 60707 11797
rect 63585 11794 63651 11797
rect 60641 11792 63651 11794
rect 60641 11736 60646 11792
rect 60702 11736 63590 11792
rect 63646 11736 63651 11792
rect 60641 11734 63651 11736
rect 60641 11731 60707 11734
rect 63585 11731 63651 11734
rect 79869 11794 79935 11797
rect 82537 11794 82603 11797
rect 79869 11792 82603 11794
rect 79869 11736 79874 11792
rect 79930 11736 82542 11792
rect 82598 11736 82603 11792
rect 79869 11734 82603 11736
rect 79869 11731 79935 11734
rect 82537 11731 82603 11734
rect 26141 11658 26207 11661
rect 77569 11658 77635 11661
rect 26141 11656 77635 11658
rect 26141 11600 26146 11656
rect 26202 11600 77574 11656
rect 77630 11600 77635 11656
rect 26141 11598 77635 11600
rect 26141 11595 26207 11598
rect 77569 11595 77635 11598
rect 115013 11658 115079 11661
rect 122557 11658 122623 11661
rect 115013 11656 122623 11658
rect 115013 11600 115018 11656
rect 115074 11600 122562 11656
rect 122618 11600 122623 11656
rect 115013 11598 122623 11600
rect 115013 11595 115079 11598
rect 122557 11595 122623 11598
rect 0 11522 800 11552
rect 4061 11522 4127 11525
rect 0 11520 4127 11522
rect 0 11464 4066 11520
rect 4122 11464 4127 11520
rect 0 11462 4127 11464
rect 0 11432 800 11462
rect 4061 11459 4127 11462
rect 22461 11522 22527 11525
rect 28257 11522 28323 11525
rect 22461 11520 28323 11522
rect 22461 11464 22466 11520
rect 22522 11464 28262 11520
rect 28318 11464 28323 11520
rect 22461 11462 28323 11464
rect 22461 11459 22527 11462
rect 28257 11459 28323 11462
rect 32121 11522 32187 11525
rect 36353 11522 36419 11525
rect 32121 11520 36419 11522
rect 32121 11464 32126 11520
rect 32182 11464 36358 11520
rect 36414 11464 36419 11520
rect 32121 11462 36419 11464
rect 32121 11459 32187 11462
rect 36353 11459 36419 11462
rect 36629 11522 36695 11525
rect 45553 11522 45619 11525
rect 36629 11520 45619 11522
rect 36629 11464 36634 11520
rect 36690 11464 45558 11520
rect 45614 11464 45619 11520
rect 36629 11462 45619 11464
rect 36629 11459 36695 11462
rect 45553 11459 45619 11462
rect 46197 11522 46263 11525
rect 63033 11522 63099 11525
rect 46197 11520 63099 11522
rect 46197 11464 46202 11520
rect 46258 11464 63038 11520
rect 63094 11464 63099 11520
rect 46197 11462 63099 11464
rect 46197 11459 46263 11462
rect 63033 11459 63099 11462
rect 116485 11522 116551 11525
rect 124765 11522 124831 11525
rect 116485 11520 124831 11522
rect 116485 11464 116490 11520
rect 116546 11464 124770 11520
rect 124826 11464 124831 11520
rect 116485 11462 124831 11464
rect 116485 11459 116551 11462
rect 124765 11459 124831 11462
rect 28418 11456 28738 11457
rect 28418 11392 28426 11456
rect 28490 11392 28506 11456
rect 28570 11392 28586 11456
rect 28650 11392 28666 11456
rect 28730 11392 28738 11456
rect 28418 11391 28738 11392
rect 84840 11456 85160 11457
rect 84840 11392 84848 11456
rect 84912 11392 84928 11456
rect 84992 11392 85008 11456
rect 85072 11392 85088 11456
rect 85152 11392 85160 11456
rect 84840 11391 85160 11392
rect 141261 11456 141581 11457
rect 141261 11392 141269 11456
rect 141333 11392 141349 11456
rect 141413 11392 141429 11456
rect 141493 11392 141509 11456
rect 141573 11392 141581 11456
rect 141261 11391 141581 11392
rect 22829 11386 22895 11389
rect 28073 11386 28139 11389
rect 22829 11384 28139 11386
rect 22829 11328 22834 11384
rect 22890 11328 28078 11384
rect 28134 11328 28139 11384
rect 22829 11326 28139 11328
rect 22829 11323 22895 11326
rect 28073 11323 28139 11326
rect 31845 11386 31911 11389
rect 69289 11386 69355 11389
rect 31845 11384 69355 11386
rect 31845 11328 31850 11384
rect 31906 11328 69294 11384
rect 69350 11328 69355 11384
rect 31845 11326 69355 11328
rect 31845 11323 31911 11326
rect 69289 11323 69355 11326
rect 116945 11386 117011 11389
rect 122925 11386 122991 11389
rect 116945 11384 122991 11386
rect 116945 11328 116950 11384
rect 117006 11328 122930 11384
rect 122986 11328 122991 11384
rect 116945 11326 122991 11328
rect 116945 11323 117011 11326
rect 122925 11323 122991 11326
rect 7649 11250 7715 11253
rect 74533 11250 74599 11253
rect 7649 11248 74599 11250
rect 7649 11192 7654 11248
rect 7710 11192 74538 11248
rect 74594 11192 74599 11248
rect 7649 11190 74599 11192
rect 7649 11187 7715 11190
rect 74533 11187 74599 11190
rect 8017 11114 8083 11117
rect 76281 11114 76347 11117
rect 8017 11112 76347 11114
rect 8017 11056 8022 11112
rect 8078 11056 76286 11112
rect 76342 11056 76347 11112
rect 8017 11054 76347 11056
rect 8017 11051 8083 11054
rect 76281 11051 76347 11054
rect 0 10978 800 11008
rect 3601 10978 3667 10981
rect 0 10976 3667 10978
rect 0 10920 3606 10976
rect 3662 10920 3667 10976
rect 0 10918 3667 10920
rect 0 10888 800 10918
rect 3601 10915 3667 10918
rect 9305 10978 9371 10981
rect 45737 10978 45803 10981
rect 9305 10976 45803 10978
rect 9305 10920 9310 10976
rect 9366 10920 45742 10976
rect 45798 10920 45803 10976
rect 9305 10918 45803 10920
rect 9305 10915 9371 10918
rect 45737 10915 45803 10918
rect 46105 10978 46171 10981
rect 52729 10978 52795 10981
rect 56409 10978 56475 10981
rect 46105 10976 51274 10978
rect 46105 10920 46110 10976
rect 46166 10920 51274 10976
rect 46105 10918 51274 10920
rect 46105 10915 46171 10918
rect 25405 10842 25471 10845
rect 51214 10842 51274 10918
rect 52729 10976 56475 10978
rect 52729 10920 52734 10976
rect 52790 10920 56414 10976
rect 56470 10920 56475 10976
rect 52729 10918 56475 10920
rect 52729 10915 52795 10918
rect 56409 10915 56475 10918
rect 57145 10978 57211 10981
rect 66161 10978 66227 10981
rect 57145 10976 66227 10978
rect 57145 10920 57150 10976
rect 57206 10920 66166 10976
rect 66222 10920 66227 10976
rect 57145 10918 66227 10920
rect 57145 10915 57211 10918
rect 66161 10915 66227 10918
rect 56629 10912 56949 10913
rect 56629 10848 56637 10912
rect 56701 10848 56717 10912
rect 56781 10848 56797 10912
rect 56861 10848 56877 10912
rect 56941 10848 56949 10912
rect 56629 10847 56949 10848
rect 113050 10912 113370 10913
rect 113050 10848 113058 10912
rect 113122 10848 113138 10912
rect 113202 10848 113218 10912
rect 113282 10848 113298 10912
rect 113362 10848 113370 10912
rect 113050 10847 113370 10848
rect 56133 10842 56199 10845
rect 77385 10842 77451 10845
rect 25405 10840 51090 10842
rect 25405 10784 25410 10840
rect 25466 10784 51090 10840
rect 25405 10782 51090 10784
rect 51214 10840 56199 10842
rect 51214 10784 56138 10840
rect 56194 10784 56199 10840
rect 51214 10782 56199 10784
rect 25405 10779 25471 10782
rect 21633 10706 21699 10709
rect 49233 10706 49299 10709
rect 50337 10706 50403 10709
rect 21633 10704 46306 10706
rect 21633 10648 21638 10704
rect 21694 10648 46306 10704
rect 21633 10646 46306 10648
rect 21633 10643 21699 10646
rect 25773 10570 25839 10573
rect 25773 10568 28872 10570
rect 25773 10512 25778 10568
rect 25834 10512 28872 10568
rect 25773 10510 28872 10512
rect 25773 10507 25839 10510
rect 0 10434 800 10464
rect 2865 10434 2931 10437
rect 0 10432 2931 10434
rect 0 10376 2870 10432
rect 2926 10376 2931 10432
rect 0 10374 2931 10376
rect 0 10344 800 10374
rect 2865 10371 2931 10374
rect 21725 10434 21791 10437
rect 26877 10434 26943 10437
rect 21725 10432 26943 10434
rect 21725 10376 21730 10432
rect 21786 10376 26882 10432
rect 26938 10376 26943 10432
rect 21725 10374 26943 10376
rect 21725 10371 21791 10374
rect 26877 10371 26943 10374
rect 27061 10434 27127 10437
rect 27705 10434 27771 10437
rect 27061 10432 27771 10434
rect 27061 10376 27066 10432
rect 27122 10376 27710 10432
rect 27766 10376 27771 10432
rect 27061 10374 27771 10376
rect 28812 10434 28872 10510
rect 29126 10508 29132 10572
rect 29196 10570 29202 10572
rect 46105 10570 46171 10573
rect 29196 10568 46171 10570
rect 29196 10512 46110 10568
rect 46166 10512 46171 10568
rect 29196 10510 46171 10512
rect 46246 10570 46306 10646
rect 49233 10704 50403 10706
rect 49233 10648 49238 10704
rect 49294 10648 50342 10704
rect 50398 10648 50403 10704
rect 49233 10646 50403 10648
rect 51030 10706 51090 10782
rect 56133 10779 56199 10782
rect 57102 10840 77451 10842
rect 57102 10784 77390 10840
rect 77446 10784 77451 10840
rect 57102 10782 77451 10784
rect 57102 10706 57162 10782
rect 77385 10779 77451 10782
rect 97533 10842 97599 10845
rect 106181 10842 106247 10845
rect 97533 10840 106247 10842
rect 97533 10784 97538 10840
rect 97594 10784 106186 10840
rect 106242 10784 106247 10840
rect 97533 10782 106247 10784
rect 97533 10779 97599 10782
rect 106181 10779 106247 10782
rect 76373 10706 76439 10709
rect 51030 10646 57162 10706
rect 57240 10704 76439 10706
rect 57240 10648 76378 10704
rect 76434 10648 76439 10704
rect 57240 10646 76439 10648
rect 49233 10643 49299 10646
rect 50337 10643 50403 10646
rect 57240 10570 57300 10646
rect 76373 10643 76439 10646
rect 117037 10706 117103 10709
rect 120533 10706 120599 10709
rect 117037 10704 120599 10706
rect 117037 10648 117042 10704
rect 117098 10648 120538 10704
rect 120594 10648 120599 10704
rect 117037 10646 120599 10648
rect 117037 10643 117103 10646
rect 120533 10643 120599 10646
rect 46246 10510 57300 10570
rect 57421 10570 57487 10573
rect 81157 10570 81223 10573
rect 85665 10570 85731 10573
rect 57421 10568 81223 10570
rect 57421 10512 57426 10568
rect 57482 10512 81162 10568
rect 81218 10512 81223 10568
rect 57421 10510 81223 10512
rect 29196 10508 29202 10510
rect 46105 10507 46171 10510
rect 57421 10507 57487 10510
rect 81157 10507 81223 10510
rect 81758 10568 85731 10570
rect 81758 10512 85670 10568
rect 85726 10512 85731 10568
rect 81758 10510 85731 10512
rect 55121 10434 55187 10437
rect 69013 10434 69079 10437
rect 28812 10432 55187 10434
rect 28812 10376 55126 10432
rect 55182 10376 55187 10432
rect 28812 10374 55187 10376
rect 27061 10371 27127 10374
rect 27705 10371 27771 10374
rect 55121 10371 55187 10374
rect 55262 10432 69079 10434
rect 55262 10376 69018 10432
rect 69074 10376 69079 10432
rect 55262 10374 69079 10376
rect 28418 10368 28738 10369
rect 28418 10304 28426 10368
rect 28490 10304 28506 10368
rect 28570 10304 28586 10368
rect 28650 10304 28666 10368
rect 28730 10304 28738 10368
rect 28418 10303 28738 10304
rect 23933 10298 23999 10301
rect 28257 10298 28323 10301
rect 35157 10298 35223 10301
rect 55262 10298 55322 10374
rect 69013 10371 69079 10374
rect 69289 10434 69355 10437
rect 81758 10434 81818 10510
rect 85665 10507 85731 10510
rect 108849 10570 108915 10573
rect 112989 10570 113055 10573
rect 108849 10568 113055 10570
rect 108849 10512 108854 10568
rect 108910 10512 112994 10568
rect 113050 10512 113055 10568
rect 108849 10510 113055 10512
rect 108849 10507 108915 10510
rect 112989 10507 113055 10510
rect 121177 10570 121243 10573
rect 140773 10570 140839 10573
rect 121177 10568 140839 10570
rect 121177 10512 121182 10568
rect 121238 10512 140778 10568
rect 140834 10512 140839 10568
rect 121177 10510 140839 10512
rect 121177 10507 121243 10510
rect 140773 10507 140839 10510
rect 69289 10432 81818 10434
rect 69289 10376 69294 10432
rect 69350 10376 81818 10432
rect 69289 10374 81818 10376
rect 69289 10371 69355 10374
rect 84840 10368 85160 10369
rect 84840 10304 84848 10368
rect 84912 10304 84928 10368
rect 84992 10304 85008 10368
rect 85072 10304 85088 10368
rect 85152 10304 85160 10368
rect 84840 10303 85160 10304
rect 141261 10368 141581 10369
rect 141261 10304 141269 10368
rect 141333 10304 141349 10368
rect 141413 10304 141429 10368
rect 141493 10304 141509 10368
rect 141573 10304 141581 10368
rect 141261 10303 141581 10304
rect 59537 10298 59603 10301
rect 63769 10298 63835 10301
rect 23933 10296 28323 10298
rect 23933 10240 23938 10296
rect 23994 10240 28262 10296
rect 28318 10240 28323 10296
rect 23933 10238 28323 10240
rect 23933 10235 23999 10238
rect 28257 10235 28323 10238
rect 28812 10238 35082 10298
rect 9673 10162 9739 10165
rect 17309 10162 17375 10165
rect 28812 10162 28872 10238
rect 9673 10160 17375 10162
rect 9673 10104 9678 10160
rect 9734 10104 17314 10160
rect 17370 10104 17375 10160
rect 9673 10102 17375 10104
rect 9673 10099 9739 10102
rect 17309 10099 17375 10102
rect 20302 10102 28872 10162
rect 28993 10162 29059 10165
rect 30741 10162 30807 10165
rect 28993 10160 30807 10162
rect 28993 10104 28998 10160
rect 29054 10104 30746 10160
rect 30802 10104 30807 10160
rect 28993 10102 30807 10104
rect 0 9890 800 9920
rect 4061 9890 4127 9893
rect 0 9888 4127 9890
rect 0 9832 4066 9888
rect 4122 9832 4127 9888
rect 0 9830 4127 9832
rect 0 9800 800 9830
rect 4061 9827 4127 9830
rect 5073 9890 5139 9893
rect 20302 9890 20362 10102
rect 28993 10099 29059 10102
rect 30741 10099 30807 10102
rect 31201 10162 31267 10165
rect 31845 10162 31911 10165
rect 31201 10160 31911 10162
rect 31201 10104 31206 10160
rect 31262 10104 31850 10160
rect 31906 10104 31911 10160
rect 31201 10102 31911 10104
rect 35022 10162 35082 10238
rect 35157 10296 55322 10298
rect 35157 10240 35162 10296
rect 35218 10240 55322 10296
rect 35157 10238 55322 10240
rect 55492 10238 57530 10298
rect 35157 10235 35223 10238
rect 37273 10162 37339 10165
rect 35022 10160 37339 10162
rect 35022 10104 37278 10160
rect 37334 10104 37339 10160
rect 35022 10102 37339 10104
rect 31201 10099 31267 10102
rect 31845 10099 31911 10102
rect 37273 10099 37339 10102
rect 37457 10162 37523 10165
rect 40125 10162 40191 10165
rect 37457 10160 40191 10162
rect 37457 10104 37462 10160
rect 37518 10104 40130 10160
rect 40186 10104 40191 10160
rect 37457 10102 40191 10104
rect 37457 10099 37523 10102
rect 40125 10099 40191 10102
rect 40309 10162 40375 10165
rect 55492 10162 55552 10238
rect 57470 10162 57530 10238
rect 59537 10296 63835 10298
rect 59537 10240 59542 10296
rect 59598 10240 63774 10296
rect 63830 10240 63835 10296
rect 59537 10238 63835 10240
rect 59537 10235 59603 10238
rect 63769 10235 63835 10238
rect 107193 10298 107259 10301
rect 128997 10298 129063 10301
rect 107193 10296 129063 10298
rect 107193 10240 107198 10296
rect 107254 10240 129002 10296
rect 129058 10240 129063 10296
rect 107193 10238 129063 10240
rect 107193 10235 107259 10238
rect 128997 10235 129063 10238
rect 79409 10162 79475 10165
rect 40309 10160 55552 10162
rect 40309 10104 40314 10160
rect 40370 10104 55552 10160
rect 40309 10102 55552 10104
rect 55630 10102 57300 10162
rect 57470 10160 79475 10162
rect 57470 10104 79414 10160
rect 79470 10104 79475 10160
rect 57470 10102 79475 10104
rect 40309 10099 40375 10102
rect 23381 10026 23447 10029
rect 55630 10026 55690 10102
rect 57240 10026 57300 10102
rect 79409 10099 79475 10102
rect 110137 10162 110203 10165
rect 133413 10162 133479 10165
rect 110137 10160 133479 10162
rect 110137 10104 110142 10160
rect 110198 10104 133418 10160
rect 133474 10104 133479 10160
rect 110137 10102 133479 10104
rect 110137 10099 110203 10102
rect 133413 10099 133479 10102
rect 77385 10026 77451 10029
rect 23381 10024 55690 10026
rect 23381 9968 23386 10024
rect 23442 9968 55690 10024
rect 23381 9966 55690 9968
rect 55814 9966 57162 10026
rect 57240 10024 77451 10026
rect 57240 9968 77390 10024
rect 77446 9968 77451 10024
rect 57240 9966 77451 9968
rect 23381 9963 23447 9966
rect 5073 9888 20362 9890
rect 5073 9832 5078 9888
rect 5134 9832 20362 9888
rect 5073 9830 20362 9832
rect 23657 9890 23723 9893
rect 29126 9890 29132 9892
rect 23657 9888 29132 9890
rect 23657 9832 23662 9888
rect 23718 9832 29132 9888
rect 23657 9830 29132 9832
rect 5073 9827 5139 9830
rect 23657 9827 23723 9830
rect 29126 9828 29132 9830
rect 29196 9828 29202 9892
rect 31109 9890 31175 9893
rect 46197 9890 46263 9893
rect 31109 9888 46263 9890
rect 31109 9832 31114 9888
rect 31170 9832 46202 9888
rect 46258 9832 46263 9888
rect 31109 9830 46263 9832
rect 31109 9827 31175 9830
rect 46197 9827 46263 9830
rect 46381 9890 46447 9893
rect 54569 9890 54635 9893
rect 46381 9888 54635 9890
rect 46381 9832 46386 9888
rect 46442 9832 54574 9888
rect 54630 9832 54635 9888
rect 46381 9830 54635 9832
rect 46381 9827 46447 9830
rect 54569 9827 54635 9830
rect 17033 9754 17099 9757
rect 25998 9754 26004 9756
rect 17033 9752 26004 9754
rect 17033 9696 17038 9752
rect 17094 9696 26004 9752
rect 17033 9694 26004 9696
rect 17033 9691 17099 9694
rect 25998 9692 26004 9694
rect 26068 9692 26074 9756
rect 26877 9754 26943 9757
rect 55814 9754 55874 9966
rect 55949 9890 56015 9893
rect 56317 9890 56383 9893
rect 55949 9888 56383 9890
rect 55949 9832 55954 9888
rect 56010 9832 56322 9888
rect 56378 9832 56383 9888
rect 55949 9830 56383 9832
rect 55949 9827 56015 9830
rect 56317 9827 56383 9830
rect 56629 9824 56949 9825
rect 56629 9760 56637 9824
rect 56701 9760 56717 9824
rect 56781 9760 56797 9824
rect 56861 9760 56877 9824
rect 56941 9760 56949 9824
rect 56629 9759 56949 9760
rect 26877 9752 55874 9754
rect 26877 9696 26882 9752
rect 26938 9696 55874 9752
rect 26877 9694 55874 9696
rect 55949 9754 56015 9757
rect 56409 9754 56475 9757
rect 55949 9752 56475 9754
rect 55949 9696 55954 9752
rect 56010 9696 56414 9752
rect 56470 9696 56475 9752
rect 55949 9694 56475 9696
rect 57102 9754 57162 9966
rect 77385 9963 77451 9966
rect 137829 10026 137895 10029
rect 142153 10026 142219 10029
rect 137829 10024 142219 10026
rect 137829 9968 137834 10024
rect 137890 9968 142158 10024
rect 142214 9968 142219 10024
rect 137829 9966 142219 9968
rect 137829 9963 137895 9966
rect 142153 9963 142219 9966
rect 57605 9890 57671 9893
rect 60089 9890 60155 9893
rect 57605 9888 60155 9890
rect 57605 9832 57610 9888
rect 57666 9832 60094 9888
rect 60150 9832 60155 9888
rect 57605 9830 60155 9832
rect 57605 9827 57671 9830
rect 60089 9827 60155 9830
rect 60273 9890 60339 9893
rect 62573 9890 62639 9893
rect 60273 9888 62639 9890
rect 60273 9832 60278 9888
rect 60334 9832 62578 9888
rect 62634 9832 62639 9888
rect 60273 9830 62639 9832
rect 60273 9827 60339 9830
rect 62573 9827 62639 9830
rect 63033 9890 63099 9893
rect 88057 9890 88123 9893
rect 63033 9888 88123 9890
rect 63033 9832 63038 9888
rect 63094 9832 88062 9888
rect 88118 9832 88123 9888
rect 63033 9830 88123 9832
rect 63033 9827 63099 9830
rect 88057 9827 88123 9830
rect 98361 9890 98427 9893
rect 102225 9890 102291 9893
rect 98361 9888 102291 9890
rect 98361 9832 98366 9888
rect 98422 9832 102230 9888
rect 102286 9832 102291 9888
rect 98361 9830 102291 9832
rect 98361 9827 98427 9830
rect 102225 9827 102291 9830
rect 113050 9824 113370 9825
rect 113050 9760 113058 9824
rect 113122 9760 113138 9824
rect 113202 9760 113218 9824
rect 113282 9760 113298 9824
rect 113362 9760 113370 9824
rect 113050 9759 113370 9760
rect 71497 9754 71563 9757
rect 57102 9752 71563 9754
rect 57102 9696 71502 9752
rect 71558 9696 71563 9752
rect 57102 9694 71563 9696
rect 26877 9691 26943 9694
rect 55949 9691 56015 9694
rect 56409 9691 56475 9694
rect 71497 9691 71563 9694
rect 11789 9618 11855 9621
rect 15561 9618 15627 9621
rect 11789 9616 15627 9618
rect 11789 9560 11794 9616
rect 11850 9560 15566 9616
rect 15622 9560 15627 9616
rect 11789 9558 15627 9560
rect 11789 9555 11855 9558
rect 15561 9555 15627 9558
rect 20621 9618 20687 9621
rect 24669 9618 24735 9621
rect 20621 9616 24735 9618
rect 20621 9560 20626 9616
rect 20682 9560 24674 9616
rect 24730 9560 24735 9616
rect 20621 9558 24735 9560
rect 20621 9555 20687 9558
rect 24669 9555 24735 9558
rect 25313 9618 25379 9621
rect 46013 9618 46079 9621
rect 25313 9616 46079 9618
rect 25313 9560 25318 9616
rect 25374 9560 46018 9616
rect 46074 9560 46079 9616
rect 25313 9558 46079 9560
rect 25313 9555 25379 9558
rect 46013 9555 46079 9558
rect 46197 9618 46263 9621
rect 48313 9618 48379 9621
rect 46197 9616 48379 9618
rect 46197 9560 46202 9616
rect 46258 9560 48318 9616
rect 48374 9560 48379 9616
rect 46197 9558 48379 9560
rect 46197 9555 46263 9558
rect 48313 9555 48379 9558
rect 48681 9618 48747 9621
rect 53281 9618 53347 9621
rect 48681 9616 53347 9618
rect 48681 9560 48686 9616
rect 48742 9560 53286 9616
rect 53342 9560 53347 9616
rect 48681 9558 53347 9560
rect 48681 9555 48747 9558
rect 53281 9555 53347 9558
rect 53741 9618 53807 9621
rect 63677 9618 63743 9621
rect 53741 9616 63743 9618
rect 53741 9560 53746 9616
rect 53802 9560 63682 9616
rect 63738 9560 63743 9616
rect 53741 9558 63743 9560
rect 53741 9555 53807 9558
rect 63677 9555 63743 9558
rect 97809 9618 97875 9621
rect 103237 9618 103303 9621
rect 97809 9616 103303 9618
rect 97809 9560 97814 9616
rect 97870 9560 103242 9616
rect 103298 9560 103303 9616
rect 97809 9558 103303 9560
rect 97809 9555 97875 9558
rect 103237 9555 103303 9558
rect 108205 9618 108271 9621
rect 113541 9618 113607 9621
rect 108205 9616 113607 9618
rect 108205 9560 108210 9616
rect 108266 9560 113546 9616
rect 113602 9560 113607 9616
rect 108205 9558 113607 9560
rect 108205 9555 108271 9558
rect 113541 9555 113607 9558
rect 119245 9618 119311 9621
rect 122465 9618 122531 9621
rect 119245 9616 122531 9618
rect 119245 9560 119250 9616
rect 119306 9560 122470 9616
rect 122526 9560 122531 9616
rect 119245 9558 122531 9560
rect 119245 9555 119311 9558
rect 122465 9555 122531 9558
rect 145373 9618 145439 9621
rect 153285 9618 153351 9621
rect 145373 9616 153351 9618
rect 145373 9560 145378 9616
rect 145434 9560 153290 9616
rect 153346 9560 153351 9616
rect 145373 9558 153351 9560
rect 145373 9555 145439 9558
rect 153285 9555 153351 9558
rect 7373 9482 7439 9485
rect 39941 9482 40007 9485
rect 7373 9480 40007 9482
rect 7373 9424 7378 9480
rect 7434 9424 39946 9480
rect 40002 9424 40007 9480
rect 7373 9422 40007 9424
rect 7373 9419 7439 9422
rect 39941 9419 40007 9422
rect 40125 9482 40191 9485
rect 80789 9482 80855 9485
rect 40125 9480 80855 9482
rect 40125 9424 40130 9480
rect 40186 9424 80794 9480
rect 80850 9424 80855 9480
rect 40125 9422 80855 9424
rect 40125 9419 40191 9422
rect 80789 9419 80855 9422
rect 0 9346 800 9376
rect 6085 9346 6151 9349
rect 0 9344 6151 9346
rect 0 9288 6090 9344
rect 6146 9288 6151 9344
rect 0 9286 6151 9288
rect 0 9256 800 9286
rect 6085 9283 6151 9286
rect 20253 9346 20319 9349
rect 22553 9346 22619 9349
rect 28257 9346 28323 9349
rect 20253 9344 22386 9346
rect 20253 9288 20258 9344
rect 20314 9288 22386 9344
rect 20253 9286 22386 9288
rect 20253 9283 20319 9286
rect 5533 9212 5599 9213
rect 5533 9210 5580 9212
rect 5488 9208 5580 9210
rect 5488 9152 5538 9208
rect 5488 9150 5580 9152
rect 5533 9148 5580 9150
rect 5644 9148 5650 9212
rect 21633 9210 21699 9213
rect 22185 9210 22251 9213
rect 21633 9208 22251 9210
rect 21633 9152 21638 9208
rect 21694 9152 22190 9208
rect 22246 9152 22251 9208
rect 21633 9150 22251 9152
rect 22326 9210 22386 9286
rect 22553 9344 28323 9346
rect 22553 9288 22558 9344
rect 22614 9288 28262 9344
rect 28318 9288 28323 9344
rect 22553 9286 28323 9288
rect 22553 9283 22619 9286
rect 28257 9283 28323 9286
rect 28809 9346 28875 9349
rect 38561 9346 38627 9349
rect 28809 9344 38627 9346
rect 28809 9288 28814 9344
rect 28870 9288 38566 9344
rect 38622 9288 38627 9344
rect 28809 9286 38627 9288
rect 28809 9283 28875 9286
rect 38561 9283 38627 9286
rect 39205 9346 39271 9349
rect 42701 9346 42767 9349
rect 39205 9344 42767 9346
rect 39205 9288 39210 9344
rect 39266 9288 42706 9344
rect 42762 9288 42767 9344
rect 39205 9286 42767 9288
rect 39205 9283 39271 9286
rect 42701 9283 42767 9286
rect 42885 9346 42951 9349
rect 53097 9346 53163 9349
rect 42885 9344 53163 9346
rect 42885 9288 42890 9344
rect 42946 9288 53102 9344
rect 53158 9288 53163 9344
rect 42885 9286 53163 9288
rect 42885 9283 42951 9286
rect 53097 9283 53163 9286
rect 53281 9346 53347 9349
rect 53833 9346 53899 9349
rect 57145 9346 57211 9349
rect 53281 9344 53666 9346
rect 53281 9288 53286 9344
rect 53342 9288 53666 9344
rect 53281 9286 53666 9288
rect 53281 9283 53347 9286
rect 28418 9280 28738 9281
rect 28418 9216 28426 9280
rect 28490 9216 28506 9280
rect 28570 9216 28586 9280
rect 28650 9216 28666 9280
rect 28730 9216 28738 9280
rect 28418 9215 28738 9216
rect 28257 9210 28323 9213
rect 22326 9208 28323 9210
rect 22326 9152 28262 9208
rect 28318 9152 28323 9208
rect 22326 9150 28323 9152
rect 5533 9147 5599 9148
rect 21633 9147 21699 9150
rect 22185 9147 22251 9150
rect 28257 9147 28323 9150
rect 28809 9210 28875 9213
rect 42374 9210 42380 9212
rect 28809 9208 42380 9210
rect 28809 9152 28814 9208
rect 28870 9152 42380 9208
rect 28809 9150 42380 9152
rect 28809 9147 28875 9150
rect 42374 9148 42380 9150
rect 42444 9148 42450 9212
rect 50613 9210 50679 9213
rect 42566 9208 50679 9210
rect 42566 9152 50618 9208
rect 50674 9152 50679 9208
rect 42566 9150 50679 9152
rect 8477 9074 8543 9077
rect 36261 9074 36327 9077
rect 8477 9072 36327 9074
rect 8477 9016 8482 9072
rect 8538 9016 36266 9072
rect 36322 9016 36327 9072
rect 8477 9014 36327 9016
rect 8477 9011 8543 9014
rect 36261 9011 36327 9014
rect 36537 9074 36603 9077
rect 38745 9074 38811 9077
rect 36537 9072 38811 9074
rect 36537 9016 36542 9072
rect 36598 9016 38750 9072
rect 38806 9016 38811 9072
rect 36537 9014 38811 9016
rect 36537 9011 36603 9014
rect 38745 9011 38811 9014
rect 39021 9074 39087 9077
rect 42566 9074 42626 9150
rect 50613 9147 50679 9150
rect 50797 9210 50863 9213
rect 52453 9210 52519 9213
rect 50797 9208 52519 9210
rect 50797 9152 50802 9208
rect 50858 9152 52458 9208
rect 52514 9152 52519 9208
rect 50797 9150 52519 9152
rect 53606 9210 53666 9286
rect 53833 9344 57211 9346
rect 53833 9288 53838 9344
rect 53894 9288 57150 9344
rect 57206 9288 57211 9344
rect 53833 9286 57211 9288
rect 53833 9283 53899 9286
rect 57145 9283 57211 9286
rect 57605 9346 57671 9349
rect 59813 9346 59879 9349
rect 57605 9344 59879 9346
rect 57605 9288 57610 9344
rect 57666 9288 59818 9344
rect 59874 9288 59879 9344
rect 57605 9286 59879 9288
rect 57605 9283 57671 9286
rect 59813 9283 59879 9286
rect 60038 9284 60044 9348
rect 60108 9346 60114 9348
rect 76465 9346 76531 9349
rect 60108 9344 76531 9346
rect 60108 9288 76470 9344
rect 76526 9288 76531 9344
rect 60108 9286 76531 9288
rect 60108 9284 60114 9286
rect 76465 9283 76531 9286
rect 118141 9346 118207 9349
rect 124765 9346 124831 9349
rect 118141 9344 124831 9346
rect 118141 9288 118146 9344
rect 118202 9288 124770 9344
rect 124826 9288 124831 9344
rect 118141 9286 124831 9288
rect 118141 9283 118207 9286
rect 124765 9283 124831 9286
rect 84840 9280 85160 9281
rect 84840 9216 84848 9280
rect 84912 9216 84928 9280
rect 84992 9216 85008 9280
rect 85072 9216 85088 9280
rect 85152 9216 85160 9280
rect 84840 9215 85160 9216
rect 141261 9280 141581 9281
rect 141261 9216 141269 9280
rect 141333 9216 141349 9280
rect 141413 9216 141429 9280
rect 141493 9216 141509 9280
rect 141573 9216 141581 9280
rect 141261 9215 141581 9216
rect 74533 9210 74599 9213
rect 53606 9208 74599 9210
rect 53606 9152 74538 9208
rect 74594 9152 74599 9208
rect 53606 9150 74599 9152
rect 50797 9147 50863 9150
rect 52453 9147 52519 9150
rect 74533 9147 74599 9150
rect 108113 9210 108179 9213
rect 115657 9210 115723 9213
rect 108113 9208 115723 9210
rect 108113 9152 108118 9208
rect 108174 9152 115662 9208
rect 115718 9152 115723 9208
rect 108113 9150 115723 9152
rect 108113 9147 108179 9150
rect 115657 9147 115723 9150
rect 39021 9072 42626 9074
rect 39021 9016 39026 9072
rect 39082 9016 42626 9072
rect 39021 9014 42626 9016
rect 42701 9074 42767 9077
rect 72601 9074 72667 9077
rect 42701 9072 72667 9074
rect 42701 9016 42706 9072
rect 42762 9016 72606 9072
rect 72662 9016 72667 9072
rect 42701 9014 72667 9016
rect 39021 9011 39087 9014
rect 42701 9011 42767 9014
rect 72601 9011 72667 9014
rect 108665 9074 108731 9077
rect 131113 9074 131179 9077
rect 108665 9072 131179 9074
rect 108665 9016 108670 9072
rect 108726 9016 131118 9072
rect 131174 9016 131179 9072
rect 108665 9014 131179 9016
rect 108665 9011 108731 9014
rect 131113 9011 131179 9014
rect 8293 8938 8359 8941
rect 46422 8938 46428 8940
rect 8293 8936 46428 8938
rect 8293 8880 8298 8936
rect 8354 8880 46428 8936
rect 8293 8878 46428 8880
rect 8293 8875 8359 8878
rect 46422 8876 46428 8878
rect 46492 8876 46498 8940
rect 46565 8938 46631 8941
rect 81985 8938 82051 8941
rect 46565 8936 82051 8938
rect 46565 8880 46570 8936
rect 46626 8880 81990 8936
rect 82046 8880 82051 8936
rect 46565 8878 82051 8880
rect 46565 8875 46631 8878
rect 81985 8875 82051 8878
rect 95141 8938 95207 8941
rect 132401 8938 132467 8941
rect 95141 8936 96538 8938
rect 95141 8880 95146 8936
rect 95202 8880 96538 8936
rect 95141 8878 96538 8880
rect 95141 8875 95207 8878
rect 96478 8836 96538 8878
rect 111060 8878 113604 8938
rect 0 8802 800 8832
rect 4061 8802 4127 8805
rect 0 8800 4127 8802
rect 0 8744 4066 8800
rect 4122 8744 4127 8800
rect 0 8742 4127 8744
rect 0 8712 800 8742
rect 4061 8739 4127 8742
rect 23841 8802 23907 8805
rect 49785 8802 49851 8805
rect 23841 8800 49851 8802
rect 23841 8744 23846 8800
rect 23902 8744 49790 8800
rect 49846 8744 49851 8800
rect 23841 8742 49851 8744
rect 23841 8739 23907 8742
rect 49785 8739 49851 8742
rect 50286 8740 50292 8804
rect 50356 8802 50362 8804
rect 56317 8802 56383 8805
rect 50356 8800 56383 8802
rect 50356 8744 56322 8800
rect 56378 8744 56383 8800
rect 50356 8742 56383 8744
rect 50356 8740 50362 8742
rect 56317 8739 56383 8742
rect 56501 8800 56567 8805
rect 56501 8744 56506 8800
rect 56562 8744 56567 8800
rect 56501 8739 56567 8744
rect 57145 8802 57211 8805
rect 85573 8802 85639 8805
rect 57145 8800 85639 8802
rect 57145 8744 57150 8800
rect 57206 8744 85578 8800
rect 85634 8744 85639 8800
rect 96478 8802 96722 8836
rect 111060 8802 111120 8878
rect 96478 8776 111120 8802
rect 57145 8742 85639 8744
rect 96662 8742 111120 8776
rect 113544 8802 113604 8878
rect 114694 8936 132467 8938
rect 114694 8880 132406 8936
rect 132462 8880 132467 8936
rect 114694 8878 132467 8880
rect 114694 8836 114754 8878
rect 132401 8875 132467 8878
rect 132677 8938 132743 8941
rect 146845 8938 146911 8941
rect 132677 8936 141802 8938
rect 132677 8880 132682 8936
rect 132738 8904 141802 8936
rect 142110 8936 146911 8938
rect 142110 8904 146850 8936
rect 132738 8880 146850 8904
rect 146906 8880 146911 8936
rect 132677 8878 146911 8880
rect 132677 8875 132743 8878
rect 141742 8844 142170 8878
rect 146845 8875 146911 8878
rect 153009 8938 153075 8941
rect 154438 8938 154682 8972
rect 153009 8936 157994 8938
rect 153009 8880 153014 8936
rect 153070 8912 157994 8936
rect 153070 8880 154498 8912
rect 153009 8878 154498 8880
rect 154622 8878 157994 8912
rect 153009 8875 153075 8878
rect 114510 8802 114754 8836
rect 113544 8776 114754 8802
rect 146201 8802 146267 8805
rect 150709 8802 150775 8805
rect 146201 8800 150775 8802
rect 113544 8742 114570 8776
rect 146201 8744 146206 8800
rect 146262 8744 150714 8800
rect 150770 8744 150775 8800
rect 146201 8742 150775 8744
rect 157934 8802 157994 8878
rect 164785 8802 164851 8805
rect 157934 8800 164851 8802
rect 157934 8744 164790 8800
rect 164846 8744 164851 8800
rect 157934 8742 164851 8744
rect 57145 8739 57211 8742
rect 85573 8739 85639 8742
rect 146201 8739 146267 8742
rect 150709 8739 150775 8742
rect 164785 8739 164851 8742
rect 4705 8666 4771 8669
rect 4705 8664 46306 8666
rect 4705 8608 4710 8664
rect 4766 8608 46306 8664
rect 4705 8606 46306 8608
rect 4705 8603 4771 8606
rect 16205 8530 16271 8533
rect 22553 8530 22619 8533
rect 16205 8528 22619 8530
rect 16205 8472 16210 8528
rect 16266 8472 22558 8528
rect 22614 8472 22619 8528
rect 16205 8470 22619 8472
rect 16205 8467 16271 8470
rect 22553 8467 22619 8470
rect 22694 8470 42810 8530
rect 12157 8396 12223 8397
rect 12157 8392 12204 8396
rect 12268 8394 12274 8396
rect 17217 8394 17283 8397
rect 22694 8394 22754 8470
rect 12157 8336 12162 8392
rect 12157 8332 12204 8336
rect 12268 8334 12314 8394
rect 17217 8392 22754 8394
rect 17217 8336 17222 8392
rect 17278 8336 22754 8392
rect 17217 8334 22754 8336
rect 23289 8394 23355 8397
rect 27613 8394 27679 8397
rect 28993 8394 29059 8397
rect 36537 8394 36603 8397
rect 23289 8392 27679 8394
rect 23289 8336 23294 8392
rect 23350 8336 27618 8392
rect 27674 8336 27679 8392
rect 23289 8334 27679 8336
rect 12268 8332 12274 8334
rect 12157 8331 12223 8332
rect 17217 8331 17283 8334
rect 23289 8331 23355 8334
rect 27613 8331 27679 8334
rect 28260 8334 28872 8394
rect 0 8258 800 8288
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8168 800 8198
rect 4061 8195 4127 8198
rect 22185 8258 22251 8261
rect 26417 8258 26483 8261
rect 22185 8256 26483 8258
rect 22185 8200 22190 8256
rect 22246 8200 26422 8256
rect 26478 8200 26483 8256
rect 22185 8198 26483 8200
rect 22185 8195 22251 8198
rect 26417 8195 26483 8198
rect 15929 8122 15995 8125
rect 28260 8122 28320 8334
rect 28418 8192 28738 8193
rect 28418 8128 28426 8192
rect 28490 8128 28506 8192
rect 28570 8128 28586 8192
rect 28650 8128 28666 8192
rect 28730 8128 28738 8192
rect 28418 8127 28738 8128
rect 15929 8120 28320 8122
rect 15929 8064 15934 8120
rect 15990 8064 28320 8120
rect 15929 8062 28320 8064
rect 28812 8122 28872 8334
rect 28993 8392 36603 8394
rect 28993 8336 28998 8392
rect 29054 8336 36542 8392
rect 36598 8336 36603 8392
rect 28993 8334 36603 8336
rect 28993 8331 29059 8334
rect 36537 8331 36603 8334
rect 36813 8394 36879 8397
rect 42241 8394 42307 8397
rect 36813 8392 42307 8394
rect 36813 8336 36818 8392
rect 36874 8336 42246 8392
rect 42302 8336 42307 8392
rect 36813 8334 42307 8336
rect 42750 8394 42810 8470
rect 42926 8468 42932 8532
rect 42996 8530 43002 8532
rect 46105 8530 46171 8533
rect 42996 8528 46171 8530
rect 42996 8472 46110 8528
rect 46166 8472 46171 8528
rect 42996 8470 46171 8472
rect 46246 8530 46306 8606
rect 46422 8604 46428 8668
rect 46492 8666 46498 8668
rect 52913 8666 52979 8669
rect 46492 8664 52979 8666
rect 46492 8608 52918 8664
rect 52974 8608 52979 8664
rect 46492 8606 52979 8608
rect 46492 8604 46498 8606
rect 52913 8603 52979 8606
rect 53097 8666 53163 8669
rect 56504 8666 56564 8739
rect 56629 8736 56949 8737
rect 56629 8672 56637 8736
rect 56701 8672 56717 8736
rect 56781 8672 56797 8736
rect 56861 8672 56877 8736
rect 56941 8672 56949 8736
rect 56629 8671 56949 8672
rect 113050 8736 113370 8737
rect 113050 8672 113058 8736
rect 113122 8672 113138 8736
rect 113202 8672 113218 8736
rect 113282 8672 113298 8736
rect 113362 8672 113370 8736
rect 113050 8671 113370 8672
rect 53097 8664 56564 8666
rect 53097 8608 53102 8664
rect 53158 8608 56564 8664
rect 53097 8606 56564 8608
rect 57329 8666 57395 8669
rect 70761 8666 70827 8669
rect 57329 8664 70827 8666
rect 57329 8608 57334 8664
rect 57390 8608 70766 8664
rect 70822 8608 70827 8664
rect 57329 8606 70827 8608
rect 53097 8603 53163 8606
rect 57329 8603 57395 8606
rect 70761 8603 70827 8606
rect 64045 8530 64111 8533
rect 46246 8528 64111 8530
rect 46246 8472 64050 8528
rect 64106 8472 64111 8528
rect 46246 8470 64111 8472
rect 42996 8468 43002 8470
rect 46105 8467 46171 8470
rect 64045 8467 64111 8470
rect 85665 8530 85731 8533
rect 95141 8530 95207 8533
rect 85665 8528 95207 8530
rect 85665 8472 85670 8528
rect 85726 8472 95146 8528
rect 95202 8472 95207 8528
rect 85665 8470 95207 8472
rect 85665 8467 85731 8470
rect 95141 8467 95207 8470
rect 50838 8394 50844 8396
rect 42750 8334 50844 8394
rect 36813 8331 36879 8334
rect 42241 8331 42307 8334
rect 50838 8332 50844 8334
rect 50908 8332 50914 8396
rect 50981 8394 51047 8397
rect 74625 8394 74691 8397
rect 50981 8392 74691 8394
rect 50981 8336 50986 8392
rect 51042 8336 74630 8392
rect 74686 8336 74691 8392
rect 50981 8334 74691 8336
rect 50981 8331 51047 8334
rect 74625 8331 74691 8334
rect 33317 8258 33383 8261
rect 69841 8258 69907 8261
rect 33317 8256 69907 8258
rect 33317 8200 33322 8256
rect 33378 8200 69846 8256
rect 69902 8200 69907 8256
rect 33317 8198 69907 8200
rect 33317 8195 33383 8198
rect 69841 8195 69907 8198
rect 84840 8192 85160 8193
rect 84840 8128 84848 8192
rect 84912 8128 84928 8192
rect 84992 8128 85008 8192
rect 85072 8128 85088 8192
rect 85152 8128 85160 8192
rect 84840 8127 85160 8128
rect 141261 8192 141581 8193
rect 141261 8128 141269 8192
rect 141333 8128 141349 8192
rect 141413 8128 141429 8192
rect 141493 8128 141509 8192
rect 141573 8128 141581 8192
rect 141261 8127 141581 8128
rect 57973 8122 58039 8125
rect 28812 8120 58039 8122
rect 28812 8064 57978 8120
rect 58034 8064 58039 8120
rect 28812 8062 58039 8064
rect 15929 8059 15995 8062
rect 57973 8059 58039 8062
rect 58341 8122 58407 8125
rect 66621 8122 66687 8125
rect 58341 8120 66687 8122
rect 58341 8064 58346 8120
rect 58402 8064 66626 8120
rect 66682 8064 66687 8120
rect 58341 8062 66687 8064
rect 58341 8059 58407 8062
rect 66621 8059 66687 8062
rect 12893 7986 12959 7989
rect 72785 7986 72851 7989
rect 12893 7984 72851 7986
rect 12893 7928 12898 7984
rect 12954 7928 72790 7984
rect 72846 7928 72851 7984
rect 12893 7926 72851 7928
rect 12893 7923 12959 7926
rect 72785 7923 72851 7926
rect 13629 7850 13695 7853
rect 46105 7850 46171 7853
rect 13629 7848 46171 7850
rect 13629 7792 13634 7848
rect 13690 7792 46110 7848
rect 46166 7792 46171 7848
rect 13629 7790 46171 7792
rect 13629 7787 13695 7790
rect 46105 7787 46171 7790
rect 46246 7790 56058 7850
rect 0 7714 800 7744
rect 4797 7714 4863 7717
rect 0 7712 4863 7714
rect 0 7656 4802 7712
rect 4858 7656 4863 7712
rect 0 7654 4863 7656
rect 0 7624 800 7654
rect 4797 7651 4863 7654
rect 19241 7714 19307 7717
rect 24853 7714 24919 7717
rect 19241 7712 24919 7714
rect 19241 7656 19246 7712
rect 19302 7656 24858 7712
rect 24914 7656 24919 7712
rect 19241 7654 24919 7656
rect 19241 7651 19307 7654
rect 24853 7651 24919 7654
rect 26417 7714 26483 7717
rect 46246 7714 46306 7790
rect 26417 7712 46306 7714
rect 26417 7656 26422 7712
rect 26478 7656 46306 7712
rect 26417 7654 46306 7656
rect 46381 7714 46447 7717
rect 51165 7714 51231 7717
rect 55121 7714 55187 7717
rect 55489 7716 55555 7717
rect 46381 7712 51090 7714
rect 46381 7656 46386 7712
rect 46442 7656 51090 7712
rect 46381 7654 51090 7656
rect 26417 7651 26483 7654
rect 46381 7651 46447 7654
rect 15653 7578 15719 7581
rect 50889 7578 50955 7581
rect 15653 7576 50955 7578
rect 15653 7520 15658 7576
rect 15714 7520 50894 7576
rect 50950 7520 50955 7576
rect 15653 7518 50955 7520
rect 51030 7578 51090 7654
rect 51165 7712 55187 7714
rect 51165 7656 51170 7712
rect 51226 7656 55126 7712
rect 55182 7656 55187 7712
rect 51165 7654 55187 7656
rect 51165 7651 51231 7654
rect 55121 7651 55187 7654
rect 55438 7652 55444 7716
rect 55508 7714 55555 7716
rect 55998 7714 56058 7790
rect 57278 7788 57284 7852
rect 57348 7850 57354 7852
rect 67541 7850 67607 7853
rect 57348 7848 67607 7850
rect 57348 7792 67546 7848
rect 67602 7792 67607 7848
rect 57348 7790 67607 7792
rect 57348 7788 57354 7790
rect 67541 7787 67607 7790
rect 116117 7850 116183 7853
rect 116945 7850 117011 7853
rect 116117 7848 117011 7850
rect 116117 7792 116122 7848
rect 116178 7792 116950 7848
rect 117006 7792 117011 7848
rect 116117 7790 117011 7792
rect 116117 7787 116183 7790
rect 116945 7787 117011 7790
rect 56501 7714 56567 7717
rect 55508 7712 55600 7714
rect 55550 7656 55600 7712
rect 55508 7654 55600 7656
rect 55998 7712 56567 7714
rect 55998 7656 56506 7712
rect 56562 7656 56567 7712
rect 55998 7654 56567 7656
rect 55508 7652 55555 7654
rect 55489 7651 55555 7652
rect 56501 7651 56567 7654
rect 57237 7714 57303 7717
rect 73521 7714 73587 7717
rect 57237 7712 73587 7714
rect 57237 7656 57242 7712
rect 57298 7656 73526 7712
rect 73582 7656 73587 7712
rect 57237 7654 73587 7656
rect 57237 7651 57303 7654
rect 73521 7651 73587 7654
rect 103462 7652 103468 7716
rect 103532 7714 103538 7716
rect 112897 7714 112963 7717
rect 103532 7712 112963 7714
rect 103532 7656 112902 7712
rect 112958 7656 112963 7712
rect 103532 7654 112963 7656
rect 103532 7652 103538 7654
rect 112897 7651 112963 7654
rect 56629 7648 56949 7649
rect 56629 7584 56637 7648
rect 56701 7584 56717 7648
rect 56781 7584 56797 7648
rect 56861 7584 56877 7648
rect 56941 7584 56949 7648
rect 56629 7583 56949 7584
rect 113050 7648 113370 7649
rect 113050 7584 113058 7648
rect 113122 7584 113138 7648
rect 113202 7584 113218 7648
rect 113282 7584 113298 7648
rect 113362 7584 113370 7648
rect 113050 7583 113370 7584
rect 56501 7578 56567 7581
rect 51030 7576 56567 7578
rect 51030 7520 56506 7576
rect 56562 7520 56567 7576
rect 51030 7518 56567 7520
rect 15653 7515 15719 7518
rect 50889 7515 50955 7518
rect 56501 7515 56567 7518
rect 57053 7578 57119 7581
rect 60917 7578 60983 7581
rect 57053 7576 60983 7578
rect 57053 7520 57058 7576
rect 57114 7520 60922 7576
rect 60978 7520 60983 7576
rect 57053 7518 60983 7520
rect 57053 7515 57119 7518
rect 60917 7515 60983 7518
rect 114553 7578 114619 7581
rect 122741 7578 122807 7581
rect 114553 7576 122807 7578
rect 114553 7520 114558 7576
rect 114614 7520 122746 7576
rect 122802 7520 122807 7576
rect 114553 7518 122807 7520
rect 114553 7515 114619 7518
rect 122741 7515 122807 7518
rect 6821 7442 6887 7445
rect 23197 7442 23263 7445
rect 6821 7440 23263 7442
rect 6821 7384 6826 7440
rect 6882 7384 23202 7440
rect 23258 7384 23263 7440
rect 6821 7382 23263 7384
rect 6821 7379 6887 7382
rect 23197 7379 23263 7382
rect 26136 7380 26142 7444
rect 26206 7442 26212 7444
rect 80789 7442 80855 7445
rect 26206 7440 80855 7442
rect 26206 7384 80794 7440
rect 80850 7384 80855 7440
rect 26206 7382 80855 7384
rect 26206 7380 26212 7382
rect 80789 7379 80855 7382
rect 113081 7442 113147 7445
rect 114369 7442 114435 7445
rect 113081 7440 114435 7442
rect 113081 7384 113086 7440
rect 113142 7384 114374 7440
rect 114430 7384 114435 7440
rect 113081 7382 114435 7384
rect 113081 7379 113147 7382
rect 114369 7379 114435 7382
rect 148317 7442 148383 7445
rect 153142 7442 153148 7444
rect 148317 7440 153148 7442
rect 148317 7384 148322 7440
rect 148378 7384 153148 7440
rect 148317 7382 153148 7384
rect 148317 7379 148383 7382
rect 153142 7380 153148 7382
rect 153212 7380 153218 7444
rect 16021 7306 16087 7309
rect 71865 7306 71931 7309
rect 103462 7306 103468 7308
rect 16021 7304 71931 7306
rect 16021 7248 16026 7304
rect 16082 7248 71870 7304
rect 71926 7248 71931 7304
rect 16021 7246 71931 7248
rect 16021 7243 16087 7246
rect 71865 7243 71931 7246
rect 72374 7246 91754 7306
rect 0 7170 800 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 800 7110
rect 4061 7107 4127 7110
rect 5533 7170 5599 7173
rect 8201 7170 8267 7173
rect 5533 7168 8267 7170
rect 5533 7112 5538 7168
rect 5594 7112 8206 7168
rect 8262 7112 8267 7168
rect 5533 7110 8267 7112
rect 5533 7107 5599 7110
rect 8201 7107 8267 7110
rect 13261 7170 13327 7173
rect 26601 7170 26667 7173
rect 13261 7168 26667 7170
rect 13261 7112 13266 7168
rect 13322 7112 26606 7168
rect 26662 7112 26667 7168
rect 13261 7110 26667 7112
rect 13261 7107 13327 7110
rect 26601 7107 26667 7110
rect 28809 7170 28875 7173
rect 31753 7170 31819 7173
rect 60917 7170 60983 7173
rect 72374 7170 72434 7246
rect 28809 7168 31819 7170
rect 28809 7112 28814 7168
rect 28870 7112 31758 7168
rect 31814 7112 31819 7168
rect 28809 7110 31819 7112
rect 28809 7107 28875 7110
rect 31753 7107 31819 7110
rect 31894 7110 60842 7170
rect 28418 7104 28738 7105
rect 28418 7040 28426 7104
rect 28490 7040 28506 7104
rect 28570 7040 28586 7104
rect 28650 7040 28666 7104
rect 28730 7040 28738 7104
rect 28418 7039 28738 7040
rect 12433 7034 12499 7037
rect 24301 7034 24367 7037
rect 12433 7032 24367 7034
rect 12433 6976 12438 7032
rect 12494 6976 24306 7032
rect 24362 6976 24367 7032
rect 12433 6974 24367 6976
rect 12433 6971 12499 6974
rect 24301 6971 24367 6974
rect 25589 7034 25655 7037
rect 28165 7034 28231 7037
rect 25589 7032 28231 7034
rect 25589 6976 25594 7032
rect 25650 6976 28170 7032
rect 28226 6976 28231 7032
rect 25589 6974 28231 6976
rect 25589 6971 25655 6974
rect 28165 6971 28231 6974
rect 28809 7034 28875 7037
rect 31894 7034 31954 7110
rect 28809 7032 31954 7034
rect 28809 6976 28814 7032
rect 28870 6976 31954 7032
rect 28809 6974 31954 6976
rect 32029 7034 32095 7037
rect 41689 7034 41755 7037
rect 32029 7032 41755 7034
rect 32029 6976 32034 7032
rect 32090 6976 41694 7032
rect 41750 6976 41755 7032
rect 32029 6974 41755 6976
rect 28809 6971 28875 6974
rect 32029 6971 32095 6974
rect 41689 6971 41755 6974
rect 41873 7034 41939 7037
rect 60457 7034 60523 7037
rect 41873 7032 60523 7034
rect 41873 6976 41878 7032
rect 41934 6976 60462 7032
rect 60518 6976 60523 7032
rect 41873 6974 60523 6976
rect 60782 7034 60842 7110
rect 60917 7168 72434 7170
rect 60917 7112 60922 7168
rect 60978 7112 72434 7168
rect 60917 7110 72434 7112
rect 60917 7107 60983 7110
rect 80278 7108 80284 7172
rect 80348 7170 80354 7172
rect 80421 7170 80487 7173
rect 80348 7168 80487 7170
rect 80348 7112 80426 7168
rect 80482 7112 80487 7168
rect 80348 7110 80487 7112
rect 91694 7170 91754 7246
rect 99974 7246 103468 7306
rect 99974 7170 100034 7246
rect 103462 7244 103468 7246
rect 103532 7244 103538 7308
rect 122741 7306 122807 7309
rect 125366 7306 125610 7340
rect 122741 7304 132602 7306
rect 122741 7248 122746 7304
rect 122802 7280 132602 7304
rect 122802 7248 125426 7280
rect 122741 7246 125426 7248
rect 125550 7246 132602 7280
rect 122741 7243 122807 7246
rect 91694 7110 100034 7170
rect 132542 7170 132602 7246
rect 135302 7246 144746 7306
rect 135302 7170 135362 7246
rect 132542 7110 135362 7170
rect 144686 7170 144746 7246
rect 148317 7170 148383 7173
rect 144686 7168 148383 7170
rect 144686 7112 148322 7168
rect 148378 7112 148383 7168
rect 144686 7110 148383 7112
rect 80348 7108 80354 7110
rect 80421 7107 80487 7110
rect 148317 7107 148383 7110
rect 84840 7104 85160 7105
rect 84840 7040 84848 7104
rect 84912 7040 84928 7104
rect 84992 7040 85008 7104
rect 85072 7040 85088 7104
rect 85152 7040 85160 7104
rect 84840 7039 85160 7040
rect 141261 7104 141581 7105
rect 141261 7040 141269 7104
rect 141333 7040 141349 7104
rect 141413 7040 141429 7104
rect 141493 7040 141509 7104
rect 141573 7040 141581 7104
rect 141261 7039 141581 7040
rect 83181 7034 83247 7037
rect 60782 7032 83247 7034
rect 60782 6976 83186 7032
rect 83242 6976 83247 7032
rect 60782 6974 83247 6976
rect 41873 6971 41939 6974
rect 60457 6971 60523 6974
rect 83181 6971 83247 6974
rect 96613 7034 96679 7037
rect 104065 7034 104131 7037
rect 96613 7032 104131 7034
rect 96613 6976 96618 7032
rect 96674 6976 104070 7032
rect 104126 6976 104131 7032
rect 96613 6974 104131 6976
rect 96613 6971 96679 6974
rect 104065 6971 104131 6974
rect 110413 7034 110479 7037
rect 136173 7034 136239 7037
rect 110413 7032 136239 7034
rect 110413 6976 110418 7032
rect 110474 6976 136178 7032
rect 136234 6976 136239 7032
rect 110413 6974 136239 6976
rect 110413 6971 110479 6974
rect 136173 6971 136239 6974
rect 6361 6898 6427 6901
rect 51441 6898 51507 6901
rect 6361 6896 51507 6898
rect 6361 6840 6366 6896
rect 6422 6840 51446 6896
rect 51502 6840 51507 6896
rect 6361 6838 51507 6840
rect 6361 6835 6427 6838
rect 51441 6835 51507 6838
rect 51574 6836 51580 6900
rect 51644 6898 51650 6900
rect 57421 6898 57487 6901
rect 61469 6898 61535 6901
rect 51644 6838 57300 6898
rect 51644 6836 51650 6838
rect 16481 6762 16547 6765
rect 57240 6762 57300 6838
rect 57421 6896 61535 6898
rect 57421 6840 57426 6896
rect 57482 6840 61474 6896
rect 61530 6840 61535 6896
rect 57421 6838 61535 6840
rect 57421 6835 57487 6838
rect 61469 6835 61535 6838
rect 60457 6762 60523 6765
rect 16481 6760 57162 6762
rect 16481 6704 16486 6760
rect 16542 6704 57162 6760
rect 16481 6702 57162 6704
rect 57240 6760 60523 6762
rect 57240 6704 60462 6760
rect 60518 6704 60523 6760
rect 57240 6702 60523 6704
rect 16481 6699 16547 6702
rect 0 6626 800 6656
rect 4061 6626 4127 6629
rect 0 6624 4127 6626
rect 0 6568 4066 6624
rect 4122 6568 4127 6624
rect 0 6566 4127 6568
rect 0 6536 800 6566
rect 4061 6563 4127 6566
rect 10869 6626 10935 6629
rect 12433 6626 12499 6629
rect 10869 6624 12499 6626
rect 10869 6568 10874 6624
rect 10930 6568 12438 6624
rect 12494 6568 12499 6624
rect 10869 6566 12499 6568
rect 10869 6563 10935 6566
rect 12433 6563 12499 6566
rect 16849 6626 16915 6629
rect 46105 6626 46171 6629
rect 51901 6626 51967 6629
rect 16849 6624 46171 6626
rect 16849 6568 16854 6624
rect 16910 6568 46110 6624
rect 46166 6568 46171 6624
rect 16849 6566 46171 6568
rect 16849 6563 16915 6566
rect 46105 6563 46171 6566
rect 46246 6624 51967 6626
rect 46246 6568 51906 6624
rect 51962 6568 51967 6624
rect 46246 6566 51967 6568
rect 8109 6490 8175 6493
rect 46246 6490 46306 6566
rect 51901 6563 51967 6566
rect 52453 6626 52519 6629
rect 56225 6626 56291 6629
rect 52453 6624 56291 6626
rect 52453 6568 52458 6624
rect 52514 6568 56230 6624
rect 56286 6568 56291 6624
rect 52453 6566 56291 6568
rect 52453 6563 52519 6566
rect 56225 6563 56291 6566
rect 56629 6560 56949 6561
rect 56629 6496 56637 6560
rect 56701 6496 56717 6560
rect 56781 6496 56797 6560
rect 56861 6496 56877 6560
rect 56941 6496 56949 6560
rect 56629 6495 56949 6496
rect 8109 6488 46306 6490
rect 8109 6432 8114 6488
rect 8170 6432 46306 6488
rect 8109 6430 46306 6432
rect 46381 6490 46447 6493
rect 55581 6490 55647 6493
rect 56041 6492 56107 6493
rect 55990 6490 55996 6492
rect 46381 6488 55647 6490
rect 46381 6432 46386 6488
rect 46442 6432 55586 6488
rect 55642 6432 55647 6488
rect 46381 6430 55647 6432
rect 55950 6430 55996 6490
rect 56060 6488 56107 6492
rect 56102 6432 56107 6488
rect 8109 6427 8175 6430
rect 46381 6427 46447 6430
rect 55581 6427 55647 6430
rect 55990 6428 55996 6430
rect 56060 6428 56107 6432
rect 57102 6490 57162 6702
rect 60457 6699 60523 6702
rect 60825 6762 60891 6765
rect 69289 6762 69355 6765
rect 60825 6760 69355 6762
rect 60825 6704 60830 6760
rect 60886 6704 69294 6760
rect 69350 6704 69355 6760
rect 60825 6702 69355 6704
rect 60825 6699 60891 6702
rect 69289 6699 69355 6702
rect 108941 6762 109007 6765
rect 113633 6762 113699 6765
rect 108941 6760 113699 6762
rect 108941 6704 108946 6760
rect 109002 6704 113638 6760
rect 113694 6704 113699 6760
rect 108941 6702 113699 6704
rect 108941 6699 109007 6702
rect 113633 6699 113699 6702
rect 118601 6762 118667 6765
rect 123017 6762 123083 6765
rect 118601 6760 123083 6762
rect 118601 6704 118606 6760
rect 118662 6704 123022 6760
rect 123078 6704 123083 6760
rect 118601 6702 123083 6704
rect 118601 6699 118667 6702
rect 123017 6699 123083 6702
rect 57329 6626 57395 6629
rect 82997 6626 83063 6629
rect 57329 6624 83063 6626
rect 57329 6568 57334 6624
rect 57390 6568 83002 6624
rect 83058 6568 83063 6624
rect 57329 6566 83063 6568
rect 57329 6563 57395 6566
rect 82997 6563 83063 6566
rect 103973 6626 104039 6629
rect 107745 6626 107811 6629
rect 103973 6624 107811 6626
rect 103973 6568 103978 6624
rect 104034 6568 107750 6624
rect 107806 6568 107811 6624
rect 103973 6566 107811 6568
rect 103973 6563 104039 6566
rect 107745 6563 107811 6566
rect 113050 6560 113370 6561
rect 113050 6496 113058 6560
rect 113122 6496 113138 6560
rect 113202 6496 113218 6560
rect 113282 6496 113298 6560
rect 113362 6496 113370 6560
rect 113050 6495 113370 6496
rect 64597 6490 64663 6493
rect 57102 6488 64663 6490
rect 57102 6432 64602 6488
rect 64658 6432 64663 6488
rect 57102 6430 64663 6432
rect 56041 6427 56107 6428
rect 64597 6427 64663 6430
rect 99281 6490 99347 6493
rect 104709 6490 104775 6493
rect 99281 6488 104775 6490
rect 99281 6432 99286 6488
rect 99342 6432 104714 6488
rect 104770 6432 104775 6488
rect 99281 6430 104775 6432
rect 99281 6427 99347 6430
rect 104709 6427 104775 6430
rect 106365 6490 106431 6493
rect 107837 6490 107903 6493
rect 106365 6488 107903 6490
rect 106365 6432 106370 6488
rect 106426 6432 107842 6488
rect 107898 6432 107903 6488
rect 106365 6430 107903 6432
rect 106365 6427 106431 6430
rect 107837 6427 107903 6430
rect 12341 6354 12407 6357
rect 16849 6354 16915 6357
rect 12341 6352 16915 6354
rect 12341 6296 12346 6352
rect 12402 6296 16854 6352
rect 16910 6296 16915 6352
rect 12341 6294 16915 6296
rect 12341 6291 12407 6294
rect 16849 6291 16915 6294
rect 17033 6354 17099 6357
rect 70945 6354 71011 6357
rect 17033 6352 71011 6354
rect 17033 6296 17038 6352
rect 17094 6296 70950 6352
rect 71006 6296 71011 6352
rect 17033 6294 71011 6296
rect 17033 6291 17099 6294
rect 70945 6291 71011 6294
rect 6637 6218 6703 6221
rect 65517 6218 65583 6221
rect 6637 6216 65583 6218
rect 6637 6160 6642 6216
rect 6698 6160 65522 6216
rect 65578 6160 65583 6216
rect 6637 6158 65583 6160
rect 6637 6155 6703 6158
rect 65517 6155 65583 6158
rect 103329 6218 103395 6221
rect 108297 6218 108363 6221
rect 103329 6216 108363 6218
rect 103329 6160 103334 6216
rect 103390 6160 108302 6216
rect 108358 6160 108363 6216
rect 103329 6158 108363 6160
rect 103329 6155 103395 6158
rect 108297 6155 108363 6158
rect 154573 6218 154639 6221
rect 155493 6218 155559 6221
rect 154573 6216 155559 6218
rect 154573 6160 154578 6216
rect 154634 6160 155498 6216
rect 155554 6160 155559 6216
rect 154573 6158 155559 6160
rect 154573 6155 154639 6158
rect 155493 6155 155559 6158
rect 0 6082 800 6112
rect 3693 6082 3759 6085
rect 0 6080 3759 6082
rect 0 6024 3698 6080
rect 3754 6024 3759 6080
rect 0 6022 3759 6024
rect 0 5992 800 6022
rect 3693 6019 3759 6022
rect 9213 6082 9279 6085
rect 17309 6082 17375 6085
rect 9213 6080 17375 6082
rect 9213 6024 9218 6080
rect 9274 6024 17314 6080
rect 17370 6024 17375 6080
rect 9213 6022 17375 6024
rect 9213 6019 9279 6022
rect 17309 6019 17375 6022
rect 21081 6082 21147 6085
rect 26969 6082 27035 6085
rect 21081 6080 27035 6082
rect 21081 6024 21086 6080
rect 21142 6024 26974 6080
rect 27030 6024 27035 6080
rect 21081 6022 27035 6024
rect 21081 6019 21147 6022
rect 26969 6019 27035 6022
rect 28809 6082 28875 6085
rect 46013 6082 46079 6085
rect 28809 6080 46079 6082
rect 28809 6024 28814 6080
rect 28870 6024 46018 6080
rect 46074 6024 46079 6080
rect 28809 6022 46079 6024
rect 28809 6019 28875 6022
rect 46013 6019 46079 6022
rect 46197 6082 46263 6085
rect 52269 6082 52335 6085
rect 46197 6080 52335 6082
rect 46197 6024 46202 6080
rect 46258 6024 52274 6080
rect 52330 6024 52335 6080
rect 46197 6022 52335 6024
rect 46197 6019 46263 6022
rect 52269 6019 52335 6022
rect 52453 6082 52519 6085
rect 69054 6082 69060 6084
rect 52453 6080 69060 6082
rect 52453 6024 52458 6080
rect 52514 6024 69060 6080
rect 52453 6022 69060 6024
rect 52453 6019 52519 6022
rect 69054 6020 69060 6022
rect 69124 6020 69130 6084
rect 103421 6082 103487 6085
rect 104709 6082 104775 6085
rect 124121 6082 124187 6085
rect 103421 6080 104775 6082
rect 103421 6024 103426 6080
rect 103482 6024 104714 6080
rect 104770 6024 104775 6080
rect 103421 6022 104775 6024
rect 103421 6019 103487 6022
rect 104709 6019 104775 6022
rect 104942 6080 124187 6082
rect 104942 6024 124126 6080
rect 124182 6024 124187 6080
rect 104942 6022 124187 6024
rect 28418 6016 28738 6017
rect 28418 5952 28426 6016
rect 28490 5952 28506 6016
rect 28570 5952 28586 6016
rect 28650 5952 28666 6016
rect 28730 5952 28738 6016
rect 28418 5951 28738 5952
rect 84840 6016 85160 6017
rect 84840 5952 84848 6016
rect 84912 5952 84928 6016
rect 84992 5952 85008 6016
rect 85072 5952 85088 6016
rect 85152 5952 85160 6016
rect 84840 5951 85160 5952
rect 11053 5946 11119 5949
rect 17033 5946 17099 5949
rect 28257 5946 28323 5949
rect 60825 5946 60891 5949
rect 11053 5944 17099 5946
rect 11053 5888 11058 5944
rect 11114 5888 17038 5944
rect 17094 5888 17099 5944
rect 11053 5886 17099 5888
rect 11053 5883 11119 5886
rect 17033 5883 17099 5886
rect 17174 5944 28323 5946
rect 17174 5888 28262 5944
rect 28318 5888 28323 5944
rect 17174 5886 28323 5888
rect 7741 5810 7807 5813
rect 17174 5810 17234 5886
rect 28257 5883 28323 5886
rect 28812 5944 60891 5946
rect 28812 5888 60830 5944
rect 60886 5888 60891 5944
rect 28812 5886 60891 5888
rect 7741 5808 17234 5810
rect 7741 5752 7746 5808
rect 7802 5752 17234 5808
rect 7741 5750 17234 5752
rect 17309 5810 17375 5813
rect 26785 5810 26851 5813
rect 17309 5808 26851 5810
rect 17309 5752 17314 5808
rect 17370 5752 26790 5808
rect 26846 5752 26851 5808
rect 17309 5750 26851 5752
rect 7741 5747 7807 5750
rect 17309 5747 17375 5750
rect 26785 5747 26851 5750
rect 26969 5810 27035 5813
rect 28812 5810 28872 5886
rect 60825 5883 60891 5886
rect 60958 5884 60964 5948
rect 61028 5946 61034 5948
rect 67582 5946 67588 5948
rect 61028 5886 67588 5946
rect 61028 5884 61034 5886
rect 67582 5884 67588 5886
rect 67652 5884 67658 5948
rect 98269 5946 98335 5949
rect 103421 5946 103487 5949
rect 98269 5944 103487 5946
rect 98269 5888 98274 5944
rect 98330 5888 103426 5944
rect 103482 5888 103487 5944
rect 98269 5886 103487 5888
rect 98269 5883 98335 5886
rect 103421 5883 103487 5886
rect 103605 5946 103671 5949
rect 104942 5946 105002 6022
rect 124121 6019 124187 6022
rect 141261 6016 141581 6017
rect 141261 5952 141269 6016
rect 141333 5952 141349 6016
rect 141413 5952 141429 6016
rect 141493 5952 141509 6016
rect 141573 5952 141581 6016
rect 141261 5951 141581 5952
rect 103605 5944 105002 5946
rect 103605 5888 103610 5944
rect 103666 5888 105002 5944
rect 103605 5886 105002 5888
rect 106365 5946 106431 5949
rect 106733 5946 106799 5949
rect 106365 5944 106799 5946
rect 106365 5888 106370 5944
rect 106426 5888 106738 5944
rect 106794 5888 106799 5944
rect 106365 5886 106799 5888
rect 103605 5883 103671 5886
rect 106365 5883 106431 5886
rect 106733 5883 106799 5886
rect 26969 5808 28872 5810
rect 26969 5752 26974 5808
rect 27030 5752 28872 5808
rect 26969 5750 28872 5752
rect 28993 5810 29059 5813
rect 46197 5810 46263 5813
rect 28993 5808 46263 5810
rect 28993 5752 28998 5808
rect 29054 5752 46202 5808
rect 46258 5752 46263 5808
rect 28993 5750 46263 5752
rect 26969 5747 27035 5750
rect 28993 5747 29059 5750
rect 46197 5747 46263 5750
rect 46381 5810 46447 5813
rect 50889 5810 50955 5813
rect 46381 5808 50955 5810
rect 46381 5752 46386 5808
rect 46442 5752 50894 5808
rect 50950 5752 50955 5808
rect 46381 5750 50955 5752
rect 46381 5747 46447 5750
rect 50889 5747 50955 5750
rect 51073 5810 51139 5813
rect 52269 5810 52335 5813
rect 53741 5810 53807 5813
rect 51073 5808 51642 5810
rect 51073 5752 51078 5808
rect 51134 5752 51642 5808
rect 51073 5750 51642 5752
rect 51073 5747 51139 5750
rect 5349 5674 5415 5677
rect 51390 5674 51396 5676
rect 5349 5672 51396 5674
rect 5349 5616 5354 5672
rect 5410 5616 51396 5672
rect 5349 5614 51396 5616
rect 5349 5611 5415 5614
rect 51390 5612 51396 5614
rect 51460 5612 51466 5676
rect 51582 5674 51642 5750
rect 52269 5808 53807 5810
rect 52269 5752 52274 5808
rect 52330 5752 53746 5808
rect 53802 5752 53807 5808
rect 52269 5750 53807 5752
rect 52269 5747 52335 5750
rect 53741 5747 53807 5750
rect 54845 5810 54911 5813
rect 55489 5810 55555 5813
rect 54845 5808 55555 5810
rect 54845 5752 54850 5808
rect 54906 5752 55494 5808
rect 55550 5752 55555 5808
rect 54845 5750 55555 5752
rect 54845 5747 54911 5750
rect 55489 5747 55555 5750
rect 55857 5810 55923 5813
rect 100661 5810 100727 5813
rect 55857 5808 100727 5810
rect 55857 5752 55862 5808
rect 55918 5752 100666 5808
rect 100722 5752 100727 5808
rect 55857 5750 100727 5752
rect 55857 5747 55923 5750
rect 100661 5747 100727 5750
rect 61694 5674 61700 5676
rect 51582 5614 61700 5674
rect 61694 5612 61700 5614
rect 61764 5612 61770 5676
rect 0 5538 800 5568
rect 3877 5538 3943 5541
rect 0 5536 3943 5538
rect 0 5480 3882 5536
rect 3938 5480 3943 5536
rect 0 5478 3943 5480
rect 0 5448 800 5478
rect 3877 5475 3943 5478
rect 7189 5538 7255 5541
rect 56317 5538 56383 5541
rect 62113 5538 62179 5541
rect 7189 5536 56383 5538
rect 7189 5480 7194 5536
rect 7250 5480 56322 5536
rect 56378 5480 56383 5536
rect 7189 5478 56383 5480
rect 7189 5475 7255 5478
rect 56317 5475 56383 5478
rect 57102 5536 62179 5538
rect 57102 5480 62118 5536
rect 62174 5480 62179 5536
rect 57102 5478 62179 5480
rect 56629 5472 56949 5473
rect 56629 5408 56637 5472
rect 56701 5408 56717 5472
rect 56781 5408 56797 5472
rect 56861 5408 56877 5472
rect 56941 5408 56949 5472
rect 56629 5407 56949 5408
rect 27797 5402 27863 5405
rect 28901 5402 28967 5405
rect 27797 5400 28967 5402
rect 27797 5344 27802 5400
rect 27858 5344 28906 5400
rect 28962 5344 28967 5400
rect 27797 5342 28967 5344
rect 27797 5339 27863 5342
rect 28901 5339 28967 5342
rect 29085 5402 29151 5405
rect 52453 5402 52519 5405
rect 29085 5400 52519 5402
rect 29085 5344 29090 5400
rect 29146 5344 52458 5400
rect 52514 5344 52519 5400
rect 29085 5342 52519 5344
rect 29085 5339 29151 5342
rect 52453 5339 52519 5342
rect 53097 5402 53163 5405
rect 56501 5402 56567 5405
rect 53097 5400 56567 5402
rect 53097 5344 53102 5400
rect 53158 5344 56506 5400
rect 56562 5344 56567 5400
rect 53097 5342 56567 5344
rect 53097 5339 53163 5342
rect 56501 5339 56567 5342
rect 5349 5266 5415 5269
rect 31753 5266 31819 5269
rect 55673 5266 55739 5269
rect 5349 5264 31819 5266
rect 5349 5208 5354 5264
rect 5410 5208 31758 5264
rect 31814 5208 31819 5264
rect 5349 5206 31819 5208
rect 5349 5203 5415 5206
rect 31753 5203 31819 5206
rect 31894 5264 55739 5266
rect 31894 5208 55678 5264
rect 55734 5208 55739 5264
rect 31894 5206 55739 5208
rect 10869 5130 10935 5133
rect 28993 5130 29059 5133
rect 31894 5130 31954 5206
rect 55673 5203 55739 5206
rect 55806 5204 55812 5268
rect 55876 5266 55882 5268
rect 56133 5266 56199 5269
rect 55876 5264 56199 5266
rect 55876 5208 56138 5264
rect 56194 5208 56199 5264
rect 55876 5206 56199 5208
rect 55876 5204 55882 5206
rect 56133 5203 56199 5206
rect 56317 5266 56383 5269
rect 57102 5266 57162 5478
rect 62113 5475 62179 5478
rect 101397 5538 101463 5541
rect 104433 5538 104499 5541
rect 101397 5536 104499 5538
rect 101397 5480 101402 5536
rect 101458 5480 104438 5536
rect 104494 5480 104499 5536
rect 101397 5478 104499 5480
rect 101397 5475 101463 5478
rect 104433 5475 104499 5478
rect 113050 5472 113370 5473
rect 113050 5408 113058 5472
rect 113122 5408 113138 5472
rect 113202 5408 113218 5472
rect 113282 5408 113298 5472
rect 113362 5408 113370 5472
rect 113050 5407 113370 5408
rect 64689 5402 64755 5405
rect 56317 5264 57162 5266
rect 56317 5208 56322 5264
rect 56378 5208 57162 5264
rect 56317 5206 57162 5208
rect 57240 5400 64755 5402
rect 57240 5344 64694 5400
rect 64750 5344 64755 5400
rect 57240 5342 64755 5344
rect 56317 5203 56383 5206
rect 41505 5130 41571 5133
rect 10869 5128 28872 5130
rect 10869 5072 10874 5128
rect 10930 5072 28872 5128
rect 10869 5070 28872 5072
rect 10869 5067 10935 5070
rect 0 4994 800 5024
rect 3693 4994 3759 4997
rect 0 4992 3759 4994
rect 0 4936 3698 4992
rect 3754 4936 3759 4992
rect 0 4934 3759 4936
rect 28812 4994 28872 5070
rect 28993 5128 31954 5130
rect 28993 5072 28998 5128
rect 29054 5072 31954 5128
rect 28993 5070 31954 5072
rect 32078 5128 41571 5130
rect 32078 5072 41510 5128
rect 41566 5072 41571 5128
rect 32078 5070 41571 5072
rect 28993 5067 29059 5070
rect 32078 4994 32138 5070
rect 41505 5067 41571 5070
rect 41638 5068 41644 5132
rect 41708 5130 41714 5132
rect 51349 5130 51415 5133
rect 41708 5128 51415 5130
rect 41708 5072 51354 5128
rect 51410 5072 51415 5128
rect 41708 5070 51415 5072
rect 41708 5068 41714 5070
rect 51349 5067 51415 5070
rect 51809 5130 51875 5133
rect 54477 5130 54543 5133
rect 51809 5128 54543 5130
rect 51809 5072 51814 5128
rect 51870 5072 54482 5128
rect 54538 5072 54543 5128
rect 51809 5070 54543 5072
rect 51809 5067 51875 5070
rect 54477 5067 54543 5070
rect 55029 5130 55095 5133
rect 55254 5130 55260 5132
rect 55029 5128 55260 5130
rect 55029 5072 55034 5128
rect 55090 5072 55260 5128
rect 55029 5070 55260 5072
rect 55029 5067 55095 5070
rect 55254 5068 55260 5070
rect 55324 5068 55330 5132
rect 57240 5130 57300 5342
rect 64689 5339 64755 5342
rect 57421 5266 57487 5269
rect 62297 5266 62363 5269
rect 57421 5264 62363 5266
rect 57421 5208 57426 5264
rect 57482 5208 62302 5264
rect 62358 5208 62363 5264
rect 57421 5206 62363 5208
rect 57421 5203 57487 5206
rect 62297 5203 62363 5206
rect 55492 5070 57300 5130
rect 57513 5130 57579 5133
rect 63861 5130 63927 5133
rect 90817 5130 90883 5133
rect 57513 5128 63927 5130
rect 57513 5072 57518 5128
rect 57574 5072 63866 5128
rect 63922 5072 63927 5128
rect 57513 5070 63927 5072
rect 28812 4934 32138 4994
rect 32213 4994 32279 4997
rect 36670 4994 36676 4996
rect 32213 4992 36676 4994
rect 32213 4936 32218 4992
rect 32274 4936 36676 4992
rect 32213 4934 36676 4936
rect 0 4904 800 4934
rect 3693 4931 3759 4934
rect 32213 4931 32279 4934
rect 36670 4932 36676 4934
rect 36740 4932 36746 4996
rect 36997 4994 37063 4997
rect 55492 4994 55552 5070
rect 57513 5067 57579 5070
rect 63861 5067 63927 5070
rect 72374 5128 90883 5130
rect 72374 5072 90822 5128
rect 90878 5072 90883 5128
rect 72374 5070 90883 5072
rect 36997 4992 55552 4994
rect 36997 4936 37002 4992
rect 37058 4936 55552 4992
rect 36997 4934 55552 4936
rect 55673 4994 55739 4997
rect 72374 4994 72434 5070
rect 90817 5067 90883 5070
rect 100937 5130 101003 5133
rect 106089 5130 106155 5133
rect 100937 5128 106155 5130
rect 100937 5072 100942 5128
rect 100998 5072 106094 5128
rect 106150 5072 106155 5128
rect 100937 5070 106155 5072
rect 100937 5067 101003 5070
rect 106089 5067 106155 5070
rect 55673 4992 72434 4994
rect 55673 4936 55678 4992
rect 55734 4936 72434 4992
rect 55673 4934 72434 4936
rect 36997 4931 37063 4934
rect 55673 4931 55739 4934
rect 28418 4928 28738 4929
rect 28418 4864 28426 4928
rect 28490 4864 28506 4928
rect 28570 4864 28586 4928
rect 28650 4864 28666 4928
rect 28730 4864 28738 4928
rect 28418 4863 28738 4864
rect 84840 4928 85160 4929
rect 84840 4864 84848 4928
rect 84912 4864 84928 4928
rect 84992 4864 85008 4928
rect 85072 4864 85088 4928
rect 85152 4864 85160 4928
rect 84840 4863 85160 4864
rect 141261 4928 141581 4929
rect 141261 4864 141269 4928
rect 141333 4864 141349 4928
rect 141413 4864 141429 4928
rect 141493 4864 141509 4928
rect 141573 4864 141581 4928
rect 141261 4863 141581 4864
rect 29177 4858 29243 4861
rect 30833 4858 30899 4861
rect 29177 4856 30899 4858
rect 29177 4800 29182 4856
rect 29238 4800 30838 4856
rect 30894 4800 30899 4856
rect 29177 4798 30899 4800
rect 29177 4795 29243 4798
rect 30833 4795 30899 4798
rect 31385 4858 31451 4861
rect 35157 4858 35223 4861
rect 31385 4856 35223 4858
rect 31385 4800 31390 4856
rect 31446 4800 35162 4856
rect 35218 4800 35223 4856
rect 31385 4798 35223 4800
rect 31385 4795 31451 4798
rect 35157 4795 35223 4798
rect 36353 4858 36419 4861
rect 40861 4858 40927 4861
rect 36353 4856 40927 4858
rect 36353 4800 36358 4856
rect 36414 4800 40866 4856
rect 40922 4800 40927 4856
rect 36353 4798 40927 4800
rect 36353 4795 36419 4798
rect 40861 4795 40927 4798
rect 41045 4858 41111 4861
rect 63309 4858 63375 4861
rect 41045 4856 63375 4858
rect 41045 4800 41050 4856
rect 41106 4800 63314 4856
rect 63370 4800 63375 4856
rect 41045 4798 63375 4800
rect 41045 4795 41111 4798
rect 63309 4795 63375 4798
rect 5441 4722 5507 4725
rect 55489 4722 55555 4725
rect 101029 4722 101095 4725
rect 106181 4722 106247 4725
rect 5441 4720 55555 4722
rect 5441 4664 5446 4720
rect 5502 4664 55494 4720
rect 55550 4664 55555 4720
rect 5441 4662 55555 4664
rect 5441 4659 5507 4662
rect 55489 4659 55555 4662
rect 55630 4662 57300 4722
rect 5901 4586 5967 4589
rect 46381 4586 46447 4589
rect 55489 4586 55555 4589
rect 5901 4584 46306 4586
rect 5901 4528 5906 4584
rect 5962 4528 46306 4584
rect 5901 4526 46306 4528
rect 5901 4523 5967 4526
rect 0 4450 800 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 800 4390
rect 4061 4387 4127 4390
rect 9581 4450 9647 4453
rect 12382 4450 12388 4452
rect 9581 4448 12388 4450
rect 9581 4392 9586 4448
rect 9642 4392 12388 4448
rect 9581 4390 12388 4392
rect 9581 4387 9647 4390
rect 12382 4388 12388 4390
rect 12452 4388 12458 4452
rect 12525 4450 12591 4453
rect 41638 4450 41644 4452
rect 12525 4448 41644 4450
rect 12525 4392 12530 4448
rect 12586 4392 41644 4448
rect 12525 4390 41644 4392
rect 12525 4387 12591 4390
rect 41638 4388 41644 4390
rect 41708 4388 41714 4452
rect 41873 4450 41939 4453
rect 42425 4450 42491 4453
rect 41873 4448 42491 4450
rect 41873 4392 41878 4448
rect 41934 4392 42430 4448
rect 42486 4392 42491 4448
rect 41873 4390 42491 4392
rect 41873 4387 41939 4390
rect 42425 4387 42491 4390
rect 43253 4450 43319 4453
rect 46013 4450 46079 4453
rect 43253 4448 46079 4450
rect 43253 4392 43258 4448
rect 43314 4392 46018 4448
rect 46074 4392 46079 4448
rect 43253 4390 46079 4392
rect 46246 4450 46306 4526
rect 46381 4584 55555 4586
rect 46381 4528 46386 4584
rect 46442 4528 55494 4584
rect 55550 4528 55555 4584
rect 46381 4526 55555 4528
rect 46381 4523 46447 4526
rect 55489 4523 55555 4526
rect 55630 4450 55690 4662
rect 57240 4586 57300 4662
rect 101029 4720 106247 4722
rect 101029 4664 101034 4720
rect 101090 4664 106186 4720
rect 106242 4664 106247 4720
rect 101029 4662 106247 4664
rect 101029 4659 101095 4662
rect 106181 4659 106247 4662
rect 70025 4586 70091 4589
rect 46246 4390 55690 4450
rect 55814 4526 57162 4586
rect 57240 4584 70091 4586
rect 57240 4528 70030 4584
rect 70086 4528 70091 4584
rect 57240 4526 70091 4528
rect 43253 4387 43319 4390
rect 46013 4387 46079 4390
rect 7189 4314 7255 4317
rect 36353 4314 36419 4317
rect 55814 4314 55874 4526
rect 56629 4384 56949 4385
rect 56629 4320 56637 4384
rect 56701 4320 56717 4384
rect 56781 4320 56797 4384
rect 56861 4320 56877 4384
rect 56941 4320 56949 4384
rect 56629 4319 56949 4320
rect 7189 4312 36419 4314
rect 7189 4256 7194 4312
rect 7250 4256 36358 4312
rect 36414 4256 36419 4312
rect 7189 4254 36419 4256
rect 7189 4251 7255 4254
rect 36353 4251 36419 4254
rect 36494 4254 55874 4314
rect 57102 4314 57162 4526
rect 70025 4523 70091 4526
rect 57237 4450 57303 4453
rect 89662 4450 89668 4452
rect 57237 4448 89668 4450
rect 57237 4392 57242 4448
rect 57298 4392 89668 4448
rect 57237 4390 89668 4392
rect 57237 4387 57303 4390
rect 89662 4388 89668 4390
rect 89732 4388 89738 4452
rect 113050 4384 113370 4385
rect 113050 4320 113058 4384
rect 113122 4320 113138 4384
rect 113202 4320 113218 4384
rect 113282 4320 113298 4384
rect 113362 4320 113370 4384
rect 113050 4319 113370 4320
rect 62849 4314 62915 4317
rect 57102 4312 62915 4314
rect 57102 4256 62854 4312
rect 62910 4256 62915 4312
rect 57102 4254 62915 4256
rect 5901 4178 5967 4181
rect 12525 4178 12591 4181
rect 5901 4176 12591 4178
rect 5901 4120 5906 4176
rect 5962 4120 12530 4176
rect 12586 4120 12591 4176
rect 5901 4118 12591 4120
rect 5901 4115 5967 4118
rect 12525 4115 12591 4118
rect 12750 4116 12756 4180
rect 12820 4178 12826 4180
rect 36494 4178 36554 4254
rect 62849 4251 62915 4254
rect 12820 4118 36554 4178
rect 12820 4116 12826 4118
rect 36670 4116 36676 4180
rect 36740 4178 36746 4180
rect 41689 4178 41755 4181
rect 36740 4176 41755 4178
rect 36740 4120 41694 4176
rect 41750 4120 41755 4176
rect 36740 4118 41755 4120
rect 36740 4116 36746 4118
rect 41689 4115 41755 4118
rect 41873 4178 41939 4181
rect 46381 4178 46447 4181
rect 41873 4176 46447 4178
rect 41873 4120 41878 4176
rect 41934 4120 46386 4176
rect 46442 4120 46447 4176
rect 41873 4118 46447 4120
rect 41873 4115 41939 4118
rect 46381 4115 46447 4118
rect 46606 4116 46612 4180
rect 46676 4178 46682 4180
rect 46841 4178 46907 4181
rect 46676 4176 46907 4178
rect 46676 4120 46846 4176
rect 46902 4120 46907 4176
rect 46676 4118 46907 4120
rect 46676 4116 46682 4118
rect 46841 4115 46907 4118
rect 47025 4178 47091 4181
rect 51022 4178 51028 4180
rect 47025 4176 51028 4178
rect 47025 4120 47030 4176
rect 47086 4120 51028 4176
rect 47025 4118 51028 4120
rect 47025 4115 47091 4118
rect 51022 4116 51028 4118
rect 51092 4116 51098 4180
rect 51257 4178 51323 4181
rect 74349 4178 74415 4181
rect 51257 4176 74415 4178
rect 51257 4120 51262 4176
rect 51318 4120 74354 4176
rect 74410 4120 74415 4176
rect 51257 4118 74415 4120
rect 51257 4115 51323 4118
rect 74349 4115 74415 4118
rect 99557 4178 99623 4181
rect 108389 4178 108455 4181
rect 99557 4176 108455 4178
rect 99557 4120 99562 4176
rect 99618 4120 108394 4176
rect 108450 4120 108455 4176
rect 99557 4118 108455 4120
rect 99557 4115 99623 4118
rect 108389 4115 108455 4118
rect 6085 4042 6151 4045
rect 28993 4042 29059 4045
rect 36629 4042 36695 4045
rect 89437 4042 89503 4045
rect 6085 4040 28872 4042
rect 6085 3984 6090 4040
rect 6146 3984 28872 4040
rect 6085 3982 28872 3984
rect 6085 3979 6151 3982
rect 0 3906 800 3936
rect 28812 3909 28872 3982
rect 28993 4040 36554 4042
rect 28993 3984 28998 4040
rect 29054 3984 36554 4040
rect 28993 3982 36554 3984
rect 28993 3979 29059 3982
rect 4061 3906 4127 3909
rect 0 3904 4127 3906
rect 0 3848 4066 3904
rect 4122 3848 4127 3904
rect 0 3846 4127 3848
rect 0 3816 800 3846
rect 4061 3843 4127 3846
rect 6310 3844 6316 3908
rect 6380 3906 6386 3908
rect 6453 3906 6519 3909
rect 6380 3904 6519 3906
rect 6380 3848 6458 3904
rect 6514 3848 6519 3904
rect 6380 3846 6519 3848
rect 6380 3844 6386 3846
rect 6453 3843 6519 3846
rect 16573 3906 16639 3909
rect 21265 3906 21331 3909
rect 16573 3904 21331 3906
rect 16573 3848 16578 3904
rect 16634 3848 21270 3904
rect 21326 3848 21331 3904
rect 16573 3846 21331 3848
rect 16573 3843 16639 3846
rect 21265 3843 21331 3846
rect 21725 3906 21791 3909
rect 28257 3906 28323 3909
rect 21725 3904 28323 3906
rect 21725 3848 21730 3904
rect 21786 3848 28262 3904
rect 28318 3848 28323 3904
rect 21725 3846 28323 3848
rect 21725 3843 21791 3846
rect 28257 3843 28323 3846
rect 28809 3904 28875 3909
rect 28809 3848 28814 3904
rect 28870 3848 28875 3904
rect 28809 3843 28875 3848
rect 32489 3906 32555 3909
rect 35157 3906 35223 3909
rect 32489 3904 35223 3906
rect 32489 3848 32494 3904
rect 32550 3848 35162 3904
rect 35218 3848 35223 3904
rect 32489 3846 35223 3848
rect 32489 3843 32555 3846
rect 35157 3843 35223 3846
rect 35709 3906 35775 3909
rect 36353 3906 36419 3909
rect 35709 3904 36419 3906
rect 35709 3848 35714 3904
rect 35770 3848 36358 3904
rect 36414 3848 36419 3904
rect 35709 3846 36419 3848
rect 36494 3906 36554 3982
rect 36629 4040 89503 4042
rect 36629 3984 36634 4040
rect 36690 3984 89442 4040
rect 89498 3984 89503 4040
rect 36629 3982 89503 3984
rect 36629 3979 36695 3982
rect 89437 3979 89503 3982
rect 107561 4042 107627 4045
rect 109309 4042 109375 4045
rect 107561 4040 109375 4042
rect 107561 3984 107566 4040
rect 107622 3984 109314 4040
rect 109370 3984 109375 4040
rect 107561 3982 109375 3984
rect 107561 3979 107627 3982
rect 109309 3979 109375 3982
rect 69381 3906 69447 3909
rect 36494 3904 69447 3906
rect 36494 3848 69386 3904
rect 69442 3848 69447 3904
rect 36494 3846 69447 3848
rect 35709 3843 35775 3846
rect 36353 3843 36419 3846
rect 69381 3843 69447 3846
rect 70117 3906 70183 3909
rect 73061 3906 73127 3909
rect 70117 3904 73127 3906
rect 70117 3848 70122 3904
rect 70178 3848 73066 3904
rect 73122 3848 73127 3904
rect 70117 3846 73127 3848
rect 70117 3843 70183 3846
rect 73061 3843 73127 3846
rect 107469 3906 107535 3909
rect 108941 3906 109007 3909
rect 107469 3904 109007 3906
rect 107469 3848 107474 3904
rect 107530 3848 108946 3904
rect 109002 3848 109007 3904
rect 107469 3846 109007 3848
rect 107469 3843 107535 3846
rect 108941 3843 109007 3846
rect 28418 3840 28738 3841
rect 28418 3776 28426 3840
rect 28490 3776 28506 3840
rect 28570 3776 28586 3840
rect 28650 3776 28666 3840
rect 28730 3776 28738 3840
rect 28418 3775 28738 3776
rect 84840 3840 85160 3841
rect 84840 3776 84848 3840
rect 84912 3776 84928 3840
rect 84992 3776 85008 3840
rect 85072 3776 85088 3840
rect 85152 3776 85160 3840
rect 84840 3775 85160 3776
rect 141261 3840 141581 3841
rect 141261 3776 141269 3840
rect 141333 3776 141349 3840
rect 141413 3776 141429 3840
rect 141493 3776 141509 3840
rect 141573 3776 141581 3840
rect 141261 3775 141581 3776
rect 6637 3772 6703 3773
rect 6637 3770 6684 3772
rect 6592 3768 6684 3770
rect 6592 3712 6642 3768
rect 6592 3710 6684 3712
rect 6637 3708 6684 3710
rect 6748 3708 6754 3772
rect 8017 3770 8083 3773
rect 28073 3770 28139 3773
rect 8017 3768 28139 3770
rect 8017 3712 8022 3768
rect 8078 3712 28078 3768
rect 28134 3712 28139 3768
rect 8017 3710 28139 3712
rect 6637 3707 6703 3708
rect 8017 3707 8083 3710
rect 28073 3707 28139 3710
rect 28901 3770 28967 3773
rect 41781 3770 41847 3773
rect 50889 3770 50955 3773
rect 28901 3768 41706 3770
rect 28901 3712 28906 3768
rect 28962 3712 41706 3768
rect 28901 3710 41706 3712
rect 28901 3707 28967 3710
rect 21909 3634 21975 3637
rect 41505 3634 41571 3637
rect 21909 3632 41571 3634
rect 21909 3576 21914 3632
rect 21970 3576 41510 3632
rect 41566 3576 41571 3632
rect 21909 3574 41571 3576
rect 41646 3634 41706 3710
rect 41781 3768 50955 3770
rect 41781 3712 41786 3768
rect 41842 3712 50894 3768
rect 50950 3712 50955 3768
rect 41781 3710 50955 3712
rect 41781 3707 41847 3710
rect 50889 3707 50955 3710
rect 51390 3708 51396 3772
rect 51460 3770 51466 3772
rect 70577 3770 70643 3773
rect 73797 3770 73863 3773
rect 51460 3710 70456 3770
rect 51460 3708 51466 3710
rect 51758 3634 51764 3636
rect 41646 3574 51764 3634
rect 21909 3571 21975 3574
rect 41505 3571 41571 3574
rect 51758 3572 51764 3574
rect 51828 3572 51834 3636
rect 52637 3634 52703 3637
rect 59905 3634 59971 3637
rect 52637 3632 59971 3634
rect 52637 3576 52642 3632
rect 52698 3576 59910 3632
rect 59966 3576 59971 3632
rect 52637 3574 59971 3576
rect 52637 3571 52703 3574
rect 59905 3571 59971 3574
rect 60181 3634 60247 3637
rect 63769 3634 63835 3637
rect 60181 3632 63835 3634
rect 60181 3576 60186 3632
rect 60242 3576 63774 3632
rect 63830 3576 63835 3632
rect 60181 3574 63835 3576
rect 70396 3634 70456 3710
rect 70577 3768 73863 3770
rect 70577 3712 70582 3768
rect 70638 3712 73802 3768
rect 73858 3712 73863 3768
rect 70577 3710 73863 3712
rect 70577 3707 70643 3710
rect 73797 3707 73863 3710
rect 85205 3634 85271 3637
rect 70396 3632 85271 3634
rect 70396 3576 85210 3632
rect 85266 3576 85271 3632
rect 70396 3574 85271 3576
rect 60181 3571 60247 3574
rect 63769 3571 63835 3574
rect 85205 3571 85271 3574
rect 108021 3634 108087 3637
rect 115013 3634 115079 3637
rect 108021 3632 115079 3634
rect 108021 3576 108026 3632
rect 108082 3576 115018 3632
rect 115074 3576 115079 3632
rect 108021 3574 115079 3576
rect 108021 3571 108087 3574
rect 115013 3571 115079 3574
rect 11513 3498 11579 3501
rect 67449 3498 67515 3501
rect 11513 3496 67515 3498
rect 11513 3440 11518 3496
rect 11574 3440 67454 3496
rect 67510 3440 67515 3496
rect 11513 3438 67515 3440
rect 11513 3435 11579 3438
rect 67449 3435 67515 3438
rect 107561 3498 107627 3501
rect 108389 3498 108455 3501
rect 107561 3496 108455 3498
rect 107561 3440 107566 3496
rect 107622 3440 108394 3496
rect 108450 3440 108455 3496
rect 107561 3438 108455 3440
rect 107561 3435 107627 3438
rect 108389 3435 108455 3438
rect 0 3362 800 3392
rect 6177 3362 6243 3365
rect 0 3360 6243 3362
rect 0 3304 6182 3360
rect 6238 3304 6243 3360
rect 0 3302 6243 3304
rect 0 3272 800 3302
rect 6177 3299 6243 3302
rect 9673 3362 9739 3365
rect 27245 3362 27311 3365
rect 9673 3360 27311 3362
rect 9673 3304 9678 3360
rect 9734 3304 27250 3360
rect 27306 3304 27311 3360
rect 9673 3302 27311 3304
rect 9673 3299 9739 3302
rect 27245 3299 27311 3302
rect 27429 3362 27495 3365
rect 31201 3362 31267 3365
rect 27429 3360 31267 3362
rect 27429 3304 27434 3360
rect 27490 3304 31206 3360
rect 31262 3304 31267 3360
rect 27429 3302 31267 3304
rect 27429 3299 27495 3302
rect 31201 3299 31267 3302
rect 31886 3300 31892 3364
rect 31956 3362 31962 3364
rect 40217 3362 40283 3365
rect 31956 3360 40283 3362
rect 31956 3304 40222 3360
rect 40278 3304 40283 3360
rect 31956 3302 40283 3304
rect 31956 3300 31962 3302
rect 40217 3299 40283 3302
rect 40401 3362 40467 3365
rect 73521 3362 73587 3365
rect 40401 3360 56242 3362
rect 40401 3304 40406 3360
rect 40462 3304 56242 3360
rect 40401 3302 56242 3304
rect 40401 3299 40467 3302
rect 21081 3226 21147 3229
rect 23933 3226 23999 3229
rect 21081 3224 23999 3226
rect 21081 3168 21086 3224
rect 21142 3168 23938 3224
rect 23994 3168 23999 3224
rect 21081 3166 23999 3168
rect 21081 3163 21147 3166
rect 23933 3163 23999 3166
rect 24853 3226 24919 3229
rect 25405 3226 25471 3229
rect 24853 3224 25471 3226
rect 24853 3168 24858 3224
rect 24914 3168 25410 3224
rect 25466 3168 25471 3224
rect 24853 3166 25471 3168
rect 24853 3163 24919 3166
rect 25405 3163 25471 3166
rect 26325 3226 26391 3229
rect 31937 3226 32003 3229
rect 46841 3226 46907 3229
rect 50797 3226 50863 3229
rect 26325 3224 31816 3226
rect 26325 3168 26330 3224
rect 26386 3168 31816 3224
rect 26325 3166 31816 3168
rect 26325 3163 26391 3166
rect 933 3090 999 3093
rect 31385 3090 31451 3093
rect 933 3088 31451 3090
rect 933 3032 938 3088
rect 994 3032 31390 3088
rect 31446 3032 31451 3088
rect 933 3030 31451 3032
rect 31756 3090 31816 3166
rect 31937 3224 46306 3226
rect 31937 3168 31942 3224
rect 31998 3168 46306 3224
rect 31937 3166 46306 3168
rect 31937 3163 32003 3166
rect 46246 3090 46306 3166
rect 46841 3224 50863 3226
rect 46841 3168 46846 3224
rect 46902 3168 50802 3224
rect 50858 3168 50863 3224
rect 46841 3166 50863 3168
rect 46841 3163 46907 3166
rect 50797 3163 50863 3166
rect 51022 3164 51028 3228
rect 51092 3226 51098 3228
rect 56041 3226 56107 3229
rect 51092 3224 56107 3226
rect 51092 3168 56046 3224
rect 56102 3168 56107 3224
rect 51092 3166 56107 3168
rect 51092 3164 51098 3166
rect 56041 3163 56107 3166
rect 56182 3090 56242 3302
rect 57102 3302 67650 3362
rect 56629 3296 56949 3297
rect 56629 3232 56637 3296
rect 56701 3232 56717 3296
rect 56781 3232 56797 3296
rect 56861 3232 56877 3296
rect 56941 3232 56949 3296
rect 56629 3231 56949 3232
rect 57102 3090 57162 3302
rect 67449 3226 67515 3229
rect 31756 3030 46122 3090
rect 46246 3030 55690 3090
rect 56182 3030 57162 3090
rect 57240 3224 67515 3226
rect 57240 3168 67454 3224
rect 67510 3168 67515 3224
rect 57240 3166 67515 3168
rect 67590 3226 67650 3302
rect 67958 3360 73587 3362
rect 67958 3304 73526 3360
rect 73582 3304 73587 3360
rect 67958 3302 73587 3304
rect 67958 3226 68018 3302
rect 73521 3299 73587 3302
rect 113050 3296 113370 3297
rect 113050 3232 113058 3296
rect 113122 3232 113138 3296
rect 113202 3232 113218 3296
rect 113282 3232 113298 3296
rect 113362 3232 113370 3296
rect 113050 3231 113370 3232
rect 67590 3166 68018 3226
rect 933 3027 999 3030
rect 31385 3027 31451 3030
rect 12341 2954 12407 2957
rect 35801 2954 35867 2957
rect 12341 2952 35867 2954
rect 12341 2896 12346 2952
rect 12402 2896 35806 2952
rect 35862 2896 35867 2952
rect 12341 2894 35867 2896
rect 12341 2891 12407 2894
rect 35801 2891 35867 2894
rect 35985 2954 36051 2957
rect 39205 2954 39271 2957
rect 35985 2952 39271 2954
rect 35985 2896 35990 2952
rect 36046 2896 39210 2952
rect 39266 2896 39271 2952
rect 35985 2894 39271 2896
rect 35985 2891 36051 2894
rect 39205 2891 39271 2894
rect 39389 2954 39455 2957
rect 39941 2954 40007 2957
rect 39389 2952 40007 2954
rect 39389 2896 39394 2952
rect 39450 2896 39946 2952
rect 40002 2896 40007 2952
rect 39389 2894 40007 2896
rect 39389 2891 39455 2894
rect 39941 2891 40007 2894
rect 40217 2954 40283 2957
rect 43253 2954 43319 2957
rect 40217 2952 43319 2954
rect 40217 2896 40222 2952
rect 40278 2896 43258 2952
rect 43314 2896 43319 2952
rect 40217 2894 43319 2896
rect 40217 2891 40283 2894
rect 43253 2891 43319 2894
rect 44081 2954 44147 2957
rect 46062 2954 46122 3030
rect 55489 2954 55555 2957
rect 44081 2952 45570 2954
rect 44081 2896 44086 2952
rect 44142 2896 45570 2952
rect 44081 2894 45570 2896
rect 46062 2952 55555 2954
rect 46062 2896 55494 2952
rect 55550 2896 55555 2952
rect 46062 2894 55555 2896
rect 55630 2954 55690 3030
rect 57240 2954 57300 3166
rect 67449 3163 67515 3166
rect 69054 3164 69060 3228
rect 69124 3226 69130 3228
rect 69565 3226 69631 3229
rect 69124 3224 69631 3226
rect 69124 3168 69570 3224
rect 69626 3168 69631 3224
rect 69124 3166 69631 3168
rect 69124 3164 69130 3166
rect 69565 3163 69631 3166
rect 70117 3226 70183 3229
rect 70393 3226 70459 3229
rect 70117 3224 70459 3226
rect 70117 3168 70122 3224
rect 70178 3168 70398 3224
rect 70454 3168 70459 3224
rect 70117 3166 70459 3168
rect 70117 3163 70183 3166
rect 70393 3163 70459 3166
rect 70577 3226 70643 3229
rect 72969 3226 73035 3229
rect 70577 3224 73035 3226
rect 70577 3168 70582 3224
rect 70638 3168 72974 3224
rect 73030 3168 73035 3224
rect 70577 3166 73035 3168
rect 70577 3163 70643 3166
rect 72969 3163 73035 3166
rect 57421 3090 57487 3093
rect 90449 3090 90515 3093
rect 57421 3088 90515 3090
rect 57421 3032 57426 3088
rect 57482 3032 90454 3088
rect 90510 3032 90515 3088
rect 57421 3030 90515 3032
rect 57421 3027 57487 3030
rect 90449 3027 90515 3030
rect 108573 3090 108639 3093
rect 109033 3090 109099 3093
rect 108573 3088 109099 3090
rect 108573 3032 108578 3088
rect 108634 3032 109038 3088
rect 109094 3032 109099 3088
rect 108573 3030 109099 3032
rect 108573 3027 108639 3030
rect 109033 3027 109099 3030
rect 55630 2894 57300 2954
rect 58341 2954 58407 2957
rect 61561 2954 61627 2957
rect 58341 2952 61627 2954
rect 58341 2896 58346 2952
rect 58402 2896 61566 2952
rect 61622 2896 61627 2952
rect 58341 2894 61627 2896
rect 44081 2891 44147 2894
rect 0 2818 800 2848
rect 3969 2818 4035 2821
rect 0 2816 4035 2818
rect 0 2760 3974 2816
rect 4030 2760 4035 2816
rect 0 2758 4035 2760
rect 0 2728 800 2758
rect 3969 2755 4035 2758
rect 11697 2818 11763 2821
rect 21541 2818 21607 2821
rect 11697 2816 21607 2818
rect 11697 2760 11702 2816
rect 11758 2760 21546 2816
rect 21602 2760 21607 2816
rect 11697 2758 21607 2760
rect 11697 2755 11763 2758
rect 21541 2755 21607 2758
rect 28809 2818 28875 2821
rect 31702 2818 31708 2820
rect 28809 2816 31708 2818
rect 28809 2760 28814 2816
rect 28870 2760 31708 2816
rect 28809 2758 31708 2760
rect 28809 2755 28875 2758
rect 31702 2756 31708 2758
rect 31772 2756 31778 2820
rect 31845 2818 31911 2821
rect 35934 2818 35940 2820
rect 31845 2816 35940 2818
rect 31845 2760 31850 2816
rect 31906 2760 35940 2816
rect 31845 2758 35940 2760
rect 31845 2755 31911 2758
rect 35934 2756 35940 2758
rect 36004 2756 36010 2820
rect 37457 2818 37523 2821
rect 38326 2818 38332 2820
rect 37457 2816 38332 2818
rect 37457 2760 37462 2816
rect 37518 2760 38332 2816
rect 37457 2758 38332 2760
rect 37457 2755 37523 2758
rect 38326 2756 38332 2758
rect 38396 2756 38402 2820
rect 38469 2818 38535 2821
rect 40401 2818 40467 2821
rect 38469 2816 40467 2818
rect 38469 2760 38474 2816
rect 38530 2760 40406 2816
rect 40462 2760 40467 2816
rect 38469 2758 40467 2760
rect 38469 2755 38535 2758
rect 40401 2755 40467 2758
rect 40534 2756 40540 2820
rect 40604 2818 40610 2820
rect 40769 2818 40835 2821
rect 40604 2816 40835 2818
rect 40604 2760 40774 2816
rect 40830 2760 40835 2816
rect 40604 2758 40835 2760
rect 40604 2756 40610 2758
rect 40769 2755 40835 2758
rect 40953 2818 41019 2821
rect 45369 2818 45435 2821
rect 40953 2816 45435 2818
rect 40953 2760 40958 2816
rect 41014 2760 45374 2816
rect 45430 2760 45435 2816
rect 40953 2758 45435 2760
rect 45510 2818 45570 2894
rect 55489 2891 55555 2894
rect 58341 2891 58407 2894
rect 61561 2891 61627 2894
rect 62573 2954 62639 2957
rect 66897 2954 66963 2957
rect 62573 2952 66963 2954
rect 62573 2896 62578 2952
rect 62634 2896 66902 2952
rect 66958 2896 66963 2952
rect 62573 2894 66963 2896
rect 62573 2891 62639 2894
rect 66897 2891 66963 2894
rect 68369 2954 68435 2957
rect 72049 2954 72115 2957
rect 68369 2952 72115 2954
rect 68369 2896 68374 2952
rect 68430 2896 72054 2952
rect 72110 2896 72115 2952
rect 68369 2894 72115 2896
rect 68369 2891 68435 2894
rect 72049 2891 72115 2894
rect 86953 2954 87019 2957
rect 95049 2954 95115 2957
rect 86953 2952 95115 2954
rect 86953 2896 86958 2952
rect 87014 2896 95054 2952
rect 95110 2896 95115 2952
rect 86953 2894 95115 2896
rect 86953 2891 87019 2894
rect 95049 2891 95115 2894
rect 108849 2954 108915 2957
rect 109125 2954 109191 2957
rect 108849 2952 109191 2954
rect 108849 2896 108854 2952
rect 108910 2896 109130 2952
rect 109186 2896 109191 2952
rect 108849 2894 109191 2896
rect 108849 2891 108915 2894
rect 109125 2891 109191 2894
rect 109401 2954 109467 2957
rect 111057 2954 111123 2957
rect 109401 2952 111123 2954
rect 109401 2896 109406 2952
rect 109462 2896 111062 2952
rect 111118 2896 111123 2952
rect 109401 2894 111123 2896
rect 109401 2891 109467 2894
rect 111057 2891 111123 2894
rect 47025 2818 47091 2821
rect 45510 2816 47091 2818
rect 45510 2760 47030 2816
rect 47086 2760 47091 2816
rect 45510 2758 47091 2760
rect 40953 2755 41019 2758
rect 45369 2755 45435 2758
rect 47025 2755 47091 2758
rect 47209 2818 47275 2821
rect 82261 2818 82327 2821
rect 47209 2816 82327 2818
rect 47209 2760 47214 2816
rect 47270 2760 82266 2816
rect 82322 2760 82327 2816
rect 47209 2758 82327 2760
rect 47209 2755 47275 2758
rect 82261 2755 82327 2758
rect 87321 2818 87387 2821
rect 95141 2818 95207 2821
rect 87321 2816 95207 2818
rect 87321 2760 87326 2816
rect 87382 2760 95146 2816
rect 95202 2760 95207 2816
rect 87321 2758 95207 2760
rect 87321 2755 87387 2758
rect 95141 2755 95207 2758
rect 106641 2818 106707 2821
rect 114461 2818 114527 2821
rect 106641 2816 114527 2818
rect 106641 2760 106646 2816
rect 106702 2760 114466 2816
rect 114522 2760 114527 2816
rect 106641 2758 114527 2760
rect 106641 2755 106707 2758
rect 114461 2755 114527 2758
rect 28418 2752 28738 2753
rect 28418 2688 28426 2752
rect 28490 2688 28506 2752
rect 28570 2688 28586 2752
rect 28650 2688 28666 2752
rect 28730 2688 28738 2752
rect 28418 2687 28738 2688
rect 84840 2752 85160 2753
rect 84840 2688 84848 2752
rect 84912 2688 84928 2752
rect 84992 2688 85008 2752
rect 85072 2688 85088 2752
rect 85152 2688 85160 2752
rect 84840 2687 85160 2688
rect 141261 2752 141581 2753
rect 141261 2688 141269 2752
rect 141333 2688 141349 2752
rect 141413 2688 141429 2752
rect 141493 2688 141509 2752
rect 141573 2688 141581 2752
rect 141261 2687 141581 2688
rect 15837 2682 15903 2685
rect 28257 2682 28323 2685
rect 15837 2680 28323 2682
rect 15837 2624 15842 2680
rect 15898 2624 28262 2680
rect 28318 2624 28323 2680
rect 15837 2622 28323 2624
rect 15837 2619 15903 2622
rect 28257 2619 28323 2622
rect 28809 2682 28875 2685
rect 35893 2682 35959 2685
rect 28809 2680 35959 2682
rect 28809 2624 28814 2680
rect 28870 2624 35898 2680
rect 35954 2624 35959 2680
rect 28809 2622 35959 2624
rect 28809 2619 28875 2622
rect 35893 2619 35959 2622
rect 36077 2682 36143 2685
rect 75913 2682 75979 2685
rect 36077 2680 75979 2682
rect 36077 2624 36082 2680
rect 36138 2624 75918 2680
rect 75974 2624 75979 2680
rect 36077 2622 75979 2624
rect 36077 2619 36143 2622
rect 75913 2619 75979 2622
rect 86902 2620 86908 2684
rect 86972 2682 86978 2684
rect 87597 2682 87663 2685
rect 89713 2684 89779 2685
rect 89662 2682 89668 2684
rect 86972 2680 87663 2682
rect 86972 2624 87602 2680
rect 87658 2624 87663 2680
rect 86972 2622 87663 2624
rect 89622 2622 89668 2682
rect 89732 2680 89779 2684
rect 89774 2624 89779 2680
rect 86972 2620 86978 2622
rect 87597 2619 87663 2622
rect 89662 2620 89668 2622
rect 89732 2620 89779 2624
rect 89713 2619 89779 2620
rect 107653 2682 107719 2685
rect 115381 2682 115447 2685
rect 107653 2680 115447 2682
rect 107653 2624 107658 2680
rect 107714 2624 115386 2680
rect 115442 2624 115447 2680
rect 107653 2622 115447 2624
rect 107653 2619 107719 2622
rect 115381 2619 115447 2622
rect 10133 2546 10199 2549
rect 91369 2546 91435 2549
rect 10133 2544 91435 2546
rect 10133 2488 10138 2544
rect 10194 2488 91374 2544
rect 91430 2488 91435 2544
rect 10133 2486 91435 2488
rect 10133 2483 10199 2486
rect 91369 2483 91435 2486
rect 118049 2546 118115 2549
rect 120717 2546 120783 2549
rect 118049 2544 120783 2546
rect 118049 2488 118054 2544
rect 118110 2488 120722 2544
rect 120778 2488 120783 2544
rect 118049 2486 120783 2488
rect 118049 2483 118115 2486
rect 120717 2483 120783 2486
rect 153142 2484 153148 2548
rect 153212 2546 153218 2548
rect 159357 2546 159423 2549
rect 153212 2544 159423 2546
rect 153212 2488 159362 2544
rect 159418 2488 159423 2544
rect 153212 2486 159423 2488
rect 153212 2484 153218 2486
rect 159357 2483 159423 2486
rect 9765 2410 9831 2413
rect 15837 2410 15903 2413
rect 9765 2408 15903 2410
rect 9765 2352 9770 2408
rect 9826 2352 15842 2408
rect 15898 2352 15903 2408
rect 9765 2350 15903 2352
rect 9765 2347 9831 2350
rect 15837 2347 15903 2350
rect 20253 2410 20319 2413
rect 21081 2410 21147 2413
rect 20253 2408 21147 2410
rect 20253 2352 20258 2408
rect 20314 2352 21086 2408
rect 21142 2352 21147 2408
rect 20253 2350 21147 2352
rect 20253 2347 20319 2350
rect 21081 2347 21147 2350
rect 21541 2410 21607 2413
rect 35525 2410 35591 2413
rect 21541 2408 35591 2410
rect 21541 2352 21546 2408
rect 21602 2352 35530 2408
rect 35586 2352 35591 2408
rect 21541 2350 35591 2352
rect 21541 2347 21607 2350
rect 35525 2347 35591 2350
rect 35893 2410 35959 2413
rect 35893 2408 46306 2410
rect 35893 2352 35898 2408
rect 35954 2352 46306 2408
rect 35893 2350 46306 2352
rect 35893 2347 35959 2350
rect 0 2274 800 2304
rect 2957 2274 3023 2277
rect 0 2272 3023 2274
rect 0 2216 2962 2272
rect 3018 2216 3023 2272
rect 0 2214 3023 2216
rect 0 2184 800 2214
rect 2957 2211 3023 2214
rect 9029 2274 9095 2277
rect 46054 2274 46060 2276
rect 9029 2272 46060 2274
rect 9029 2216 9034 2272
rect 9090 2216 46060 2272
rect 9029 2214 46060 2216
rect 9029 2211 9095 2214
rect 46054 2212 46060 2214
rect 46124 2212 46130 2276
rect 46246 2274 46306 2350
rect 46422 2348 46428 2412
rect 46492 2410 46498 2412
rect 55121 2410 55187 2413
rect 46492 2408 55187 2410
rect 46492 2352 55126 2408
rect 55182 2352 55187 2408
rect 46492 2350 55187 2352
rect 46492 2348 46498 2350
rect 55121 2347 55187 2350
rect 55397 2410 55463 2413
rect 57237 2410 57303 2413
rect 71037 2410 71103 2413
rect 55397 2408 57162 2410
rect 55397 2352 55402 2408
rect 55458 2352 57162 2408
rect 55397 2350 57162 2352
rect 55397 2347 55463 2350
rect 55673 2274 55739 2277
rect 46246 2272 55739 2274
rect 46246 2216 55678 2272
rect 55734 2216 55739 2272
rect 46246 2214 55739 2216
rect 55673 2211 55739 2214
rect 56629 2208 56949 2209
rect 56629 2144 56637 2208
rect 56701 2144 56717 2208
rect 56781 2144 56797 2208
rect 56861 2144 56877 2208
rect 56941 2144 56949 2208
rect 56629 2143 56949 2144
rect 10777 2138 10843 2141
rect 55397 2138 55463 2141
rect 55949 2140 56015 2141
rect 55949 2138 55996 2140
rect 10777 2136 55463 2138
rect 10777 2080 10782 2136
rect 10838 2080 55402 2136
rect 55458 2080 55463 2136
rect 10777 2078 55463 2080
rect 55904 2136 55996 2138
rect 55904 2080 55954 2136
rect 55904 2078 55996 2080
rect 10777 2075 10843 2078
rect 55397 2075 55463 2078
rect 55949 2076 55996 2078
rect 56060 2076 56066 2140
rect 57102 2138 57162 2350
rect 57237 2408 71103 2410
rect 57237 2352 57242 2408
rect 57298 2352 71042 2408
rect 71098 2352 71103 2408
rect 57237 2350 71103 2352
rect 57237 2347 57303 2350
rect 71037 2347 71103 2350
rect 71313 2410 71379 2413
rect 77109 2410 77175 2413
rect 71313 2408 77175 2410
rect 71313 2352 71318 2408
rect 71374 2352 77114 2408
rect 77170 2352 77175 2408
rect 71313 2350 77175 2352
rect 71313 2347 71379 2350
rect 77109 2347 77175 2350
rect 57237 2274 57303 2277
rect 88149 2274 88215 2277
rect 57237 2272 88215 2274
rect 57237 2216 57242 2272
rect 57298 2216 88154 2272
rect 88210 2216 88215 2272
rect 57237 2214 88215 2216
rect 57237 2211 57303 2214
rect 88149 2211 88215 2214
rect 113050 2208 113370 2209
rect 113050 2144 113058 2208
rect 113122 2144 113138 2208
rect 113202 2144 113218 2208
rect 113282 2144 113298 2208
rect 113362 2144 113370 2208
rect 113050 2143 113370 2144
rect 77569 2138 77635 2141
rect 57102 2136 77635 2138
rect 57102 2080 77574 2136
rect 77630 2080 77635 2136
rect 57102 2078 77635 2080
rect 55949 2075 56015 2076
rect 77569 2075 77635 2078
rect 12709 2002 12775 2005
rect 84193 2002 84259 2005
rect 12709 2000 84259 2002
rect 12709 1944 12714 2000
rect 12770 1944 84198 2000
rect 84254 1944 84259 2000
rect 12709 1942 84259 1944
rect 12709 1939 12775 1942
rect 84193 1939 84259 1942
rect 13077 1866 13143 1869
rect 26601 1866 26667 1869
rect 28993 1866 29059 1869
rect 83457 1866 83523 1869
rect 13077 1864 26667 1866
rect 13077 1808 13082 1864
rect 13138 1808 26606 1864
rect 26662 1808 26667 1864
rect 13077 1806 26667 1808
rect 13077 1803 13143 1806
rect 26601 1803 26667 1806
rect 28214 1806 28872 1866
rect 0 1730 800 1760
rect 4061 1730 4127 1733
rect 0 1728 4127 1730
rect 0 1672 4066 1728
rect 4122 1672 4127 1728
rect 0 1670 4127 1672
rect 0 1640 800 1670
rect 4061 1667 4127 1670
rect 5165 1730 5231 1733
rect 26233 1730 26299 1733
rect 5165 1728 26299 1730
rect 5165 1672 5170 1728
rect 5226 1672 26238 1728
rect 26294 1672 26299 1728
rect 5165 1670 26299 1672
rect 5165 1667 5231 1670
rect 26233 1667 26299 1670
rect 13445 1594 13511 1597
rect 28214 1594 28274 1806
rect 28812 1730 28872 1806
rect 28993 1864 83523 1866
rect 28993 1808 28998 1864
rect 29054 1808 83462 1864
rect 83518 1808 83523 1864
rect 28993 1806 83523 1808
rect 28993 1803 29059 1806
rect 83457 1803 83523 1806
rect 54937 1730 55003 1733
rect 28812 1728 55003 1730
rect 28812 1672 54942 1728
rect 54998 1672 55003 1728
rect 28812 1670 55003 1672
rect 54937 1667 55003 1670
rect 55121 1730 55187 1733
rect 57237 1730 57303 1733
rect 55121 1728 57303 1730
rect 55121 1672 55126 1728
rect 55182 1672 57242 1728
rect 57298 1672 57303 1728
rect 55121 1670 57303 1672
rect 55121 1667 55187 1670
rect 57237 1667 57303 1670
rect 57421 1730 57487 1733
rect 60641 1730 60707 1733
rect 57421 1728 60707 1730
rect 57421 1672 57426 1728
rect 57482 1672 60646 1728
rect 60702 1672 60707 1728
rect 57421 1670 60707 1672
rect 57421 1667 57487 1670
rect 60641 1667 60707 1670
rect 60917 1730 60983 1733
rect 65517 1730 65583 1733
rect 60917 1728 65583 1730
rect 60917 1672 60922 1728
rect 60978 1672 65522 1728
rect 65578 1672 65583 1728
rect 60917 1670 65583 1672
rect 60917 1667 60983 1670
rect 65517 1667 65583 1670
rect 67582 1668 67588 1732
rect 67652 1730 67658 1732
rect 68553 1730 68619 1733
rect 67652 1728 68619 1730
rect 67652 1672 68558 1728
rect 68614 1672 68619 1728
rect 67652 1670 68619 1672
rect 67652 1668 67658 1670
rect 68553 1667 68619 1670
rect 68737 1730 68803 1733
rect 70485 1730 70551 1733
rect 68737 1728 70551 1730
rect 68737 1672 68742 1728
rect 68798 1672 70490 1728
rect 70546 1672 70551 1728
rect 68737 1670 70551 1672
rect 68737 1667 68803 1670
rect 70485 1667 70551 1670
rect 71681 1730 71747 1733
rect 75269 1730 75335 1733
rect 71681 1728 75335 1730
rect 71681 1672 71686 1728
rect 71742 1672 75274 1728
rect 75330 1672 75335 1728
rect 71681 1670 75335 1672
rect 71681 1667 71747 1670
rect 75269 1667 75335 1670
rect 98821 1730 98887 1733
rect 100385 1730 100451 1733
rect 98821 1728 100451 1730
rect 98821 1672 98826 1728
rect 98882 1672 100390 1728
rect 100446 1672 100451 1728
rect 98821 1670 100451 1672
rect 98821 1667 98887 1670
rect 100385 1667 100451 1670
rect 111742 1668 111748 1732
rect 111812 1730 111818 1732
rect 112621 1730 112687 1733
rect 111812 1728 112687 1730
rect 111812 1672 112626 1728
rect 112682 1672 112687 1728
rect 111812 1670 112687 1672
rect 111812 1668 111818 1670
rect 112621 1667 112687 1670
rect 114461 1730 114527 1733
rect 118785 1730 118851 1733
rect 114461 1728 118851 1730
rect 114461 1672 114466 1728
rect 114522 1672 118790 1728
rect 118846 1672 118851 1728
rect 114461 1670 118851 1672
rect 114461 1667 114527 1670
rect 118785 1667 118851 1670
rect 28418 1664 28738 1665
rect 28418 1600 28426 1664
rect 28490 1600 28506 1664
rect 28570 1600 28586 1664
rect 28650 1600 28666 1664
rect 28730 1600 28738 1664
rect 28418 1599 28738 1600
rect 84840 1664 85160 1665
rect 84840 1600 84848 1664
rect 84912 1600 84928 1664
rect 84992 1600 85008 1664
rect 85072 1600 85088 1664
rect 85152 1600 85160 1664
rect 84840 1599 85160 1600
rect 141261 1664 141581 1665
rect 141261 1600 141269 1664
rect 141333 1600 141349 1664
rect 141413 1600 141429 1664
rect 141493 1600 141509 1664
rect 141573 1600 141581 1664
rect 141261 1599 141581 1600
rect 13445 1592 28274 1594
rect 13445 1536 13450 1592
rect 13506 1536 28274 1592
rect 13445 1534 28274 1536
rect 28809 1594 28875 1597
rect 77293 1594 77359 1597
rect 28809 1592 77359 1594
rect 28809 1536 28814 1592
rect 28870 1536 77298 1592
rect 77354 1536 77359 1592
rect 28809 1534 77359 1536
rect 13445 1531 13511 1534
rect 28809 1531 28875 1534
rect 77293 1531 77359 1534
rect 106365 1594 106431 1597
rect 112161 1594 112227 1597
rect 106365 1592 112227 1594
rect 106365 1536 106370 1592
rect 106426 1536 112166 1592
rect 112222 1536 112227 1592
rect 106365 1534 112227 1536
rect 106365 1531 106431 1534
rect 112161 1531 112227 1534
rect 11237 1460 11303 1461
rect 11237 1458 11284 1460
rect 11192 1456 11284 1458
rect 11192 1400 11242 1456
rect 11192 1398 11284 1400
rect 11237 1396 11284 1398
rect 11348 1396 11354 1460
rect 103513 1458 103579 1461
rect 11470 1456 103579 1458
rect 11470 1400 103518 1456
rect 103574 1400 103579 1456
rect 11470 1398 103579 1400
rect 11237 1395 11303 1396
rect 10501 1322 10567 1325
rect 11470 1322 11530 1398
rect 103513 1395 103579 1398
rect 107285 1458 107351 1461
rect 156781 1458 156847 1461
rect 107285 1456 156847 1458
rect 107285 1400 107290 1456
rect 107346 1400 156786 1456
rect 156842 1400 156847 1456
rect 107285 1398 156847 1400
rect 107285 1395 107351 1398
rect 156781 1395 156847 1398
rect 10501 1320 11530 1322
rect 10501 1264 10506 1320
rect 10562 1264 11530 1320
rect 10501 1262 11530 1264
rect 32765 1322 32831 1325
rect 36302 1322 36308 1324
rect 32765 1320 36308 1322
rect 32765 1264 32770 1320
rect 32826 1264 36308 1320
rect 32765 1262 36308 1264
rect 10501 1259 10567 1262
rect 32765 1259 32831 1262
rect 36302 1260 36308 1262
rect 36372 1260 36378 1324
rect 36537 1322 36603 1325
rect 38745 1322 38811 1325
rect 36537 1320 38811 1322
rect 36537 1264 36542 1320
rect 36598 1264 38750 1320
rect 38806 1264 38811 1320
rect 36537 1262 38811 1264
rect 36537 1259 36603 1262
rect 38745 1259 38811 1262
rect 38878 1260 38884 1324
rect 38948 1322 38954 1324
rect 40861 1322 40927 1325
rect 38948 1320 40927 1322
rect 38948 1264 40866 1320
rect 40922 1264 40927 1320
rect 38948 1262 40927 1264
rect 38948 1260 38954 1262
rect 40861 1259 40927 1262
rect 41045 1322 41111 1325
rect 68001 1322 68067 1325
rect 41045 1320 68067 1322
rect 41045 1264 41050 1320
rect 41106 1264 68006 1320
rect 68062 1264 68067 1320
rect 41045 1262 68067 1264
rect 41045 1259 41111 1262
rect 68001 1259 68067 1262
rect 70025 1322 70091 1325
rect 72417 1322 72483 1325
rect 70025 1320 72483 1322
rect 70025 1264 70030 1320
rect 70086 1264 72422 1320
rect 72478 1264 72483 1320
rect 70025 1262 72483 1264
rect 70025 1259 70091 1262
rect 72417 1259 72483 1262
rect 109033 1322 109099 1325
rect 113541 1322 113607 1325
rect 109033 1320 113607 1322
rect 109033 1264 109038 1320
rect 109094 1264 113546 1320
rect 113602 1264 113607 1320
rect 109033 1262 113607 1264
rect 109033 1259 109099 1262
rect 113541 1259 113607 1262
rect 0 1186 800 1216
rect 3785 1186 3851 1189
rect 0 1184 3851 1186
rect 0 1128 3790 1184
rect 3846 1128 3851 1184
rect 0 1126 3851 1128
rect 0 1096 800 1126
rect 3785 1123 3851 1126
rect 12801 1186 12867 1189
rect 43897 1186 43963 1189
rect 12801 1184 43963 1186
rect 12801 1128 12806 1184
rect 12862 1128 43902 1184
rect 43958 1128 43963 1184
rect 12801 1126 43963 1128
rect 12801 1123 12867 1126
rect 43897 1123 43963 1126
rect 44030 1124 44036 1188
rect 44100 1186 44106 1188
rect 47117 1186 47183 1189
rect 44100 1184 47183 1186
rect 44100 1128 47122 1184
rect 47178 1128 47183 1184
rect 44100 1126 47183 1128
rect 44100 1124 44106 1126
rect 47117 1123 47183 1126
rect 47301 1186 47367 1189
rect 50654 1186 50660 1188
rect 47301 1184 50660 1186
rect 47301 1128 47306 1184
rect 47362 1128 50660 1184
rect 47301 1126 50660 1128
rect 47301 1123 47367 1126
rect 50654 1124 50660 1126
rect 50724 1124 50730 1188
rect 50797 1186 50863 1189
rect 60273 1186 60339 1189
rect 61193 1186 61259 1189
rect 50797 1184 56288 1186
rect 50797 1128 50802 1184
rect 50858 1128 56288 1184
rect 50797 1126 56288 1128
rect 50797 1123 50863 1126
rect 56228 1053 56288 1126
rect 60273 1184 61259 1186
rect 60273 1128 60278 1184
rect 60334 1128 61198 1184
rect 61254 1128 61259 1184
rect 60273 1126 61259 1128
rect 60273 1123 60339 1126
rect 61193 1123 61259 1126
rect 61377 1186 61443 1189
rect 70209 1186 70275 1189
rect 77569 1186 77635 1189
rect 61377 1184 70275 1186
rect 61377 1128 61382 1184
rect 61438 1128 70214 1184
rect 70270 1128 70275 1184
rect 61377 1126 70275 1128
rect 61377 1123 61443 1126
rect 70209 1123 70275 1126
rect 72374 1184 77635 1186
rect 72374 1128 77574 1184
rect 77630 1128 77635 1184
rect 72374 1126 77635 1128
rect 56629 1120 56949 1121
rect 56629 1056 56637 1120
rect 56701 1056 56717 1120
rect 56781 1056 56797 1120
rect 56861 1056 56877 1120
rect 56941 1056 56949 1120
rect 56629 1055 56949 1056
rect 8385 1050 8451 1053
rect 8385 1048 55874 1050
rect 8385 992 8390 1048
rect 8446 992 55874 1048
rect 8385 990 55874 992
rect 8385 987 8451 990
rect 8109 914 8175 917
rect 46381 914 46447 917
rect 8109 912 46447 914
rect 8109 856 8114 912
rect 8170 856 46386 912
rect 46442 856 46447 912
rect 8109 854 46447 856
rect 8109 851 8175 854
rect 46381 851 46447 854
rect 47025 914 47091 917
rect 49918 914 49924 916
rect 47025 912 49924 914
rect 47025 856 47030 912
rect 47086 856 49924 912
rect 47025 854 49924 856
rect 47025 851 47091 854
rect 49918 852 49924 854
rect 49988 852 49994 916
rect 51390 852 51396 916
rect 51460 914 51466 916
rect 55673 914 55739 917
rect 51460 912 55739 914
rect 51460 856 55678 912
rect 55734 856 55739 912
rect 51460 854 55739 856
rect 55814 914 55874 990
rect 56225 1048 56291 1053
rect 72374 1050 72434 1126
rect 77569 1123 77635 1126
rect 98085 1186 98151 1189
rect 104893 1186 104959 1189
rect 98085 1184 104959 1186
rect 98085 1128 98090 1184
rect 98146 1128 104898 1184
rect 104954 1128 104959 1184
rect 98085 1126 104959 1128
rect 98085 1123 98151 1126
rect 104893 1123 104959 1126
rect 109033 1186 109099 1189
rect 109677 1186 109743 1189
rect 109033 1184 109743 1186
rect 109033 1128 109038 1184
rect 109094 1128 109682 1184
rect 109738 1128 109743 1184
rect 109033 1126 109743 1128
rect 109033 1123 109099 1126
rect 109677 1123 109743 1126
rect 113050 1120 113370 1121
rect 113050 1056 113058 1120
rect 113122 1056 113138 1120
rect 113202 1056 113218 1120
rect 113282 1056 113298 1120
rect 113362 1056 113370 1120
rect 113050 1055 113370 1056
rect 56225 992 56230 1048
rect 56286 992 56291 1048
rect 56225 987 56291 992
rect 57102 990 72434 1050
rect 74993 1050 75059 1053
rect 86493 1050 86559 1053
rect 74993 1048 86559 1050
rect 74993 992 74998 1048
rect 75054 992 86498 1048
rect 86554 992 86559 1048
rect 74993 990 86559 992
rect 57102 914 57162 990
rect 74993 987 75059 990
rect 86493 987 86559 990
rect 101397 1050 101463 1053
rect 104801 1050 104867 1053
rect 101397 1048 104867 1050
rect 101397 992 101402 1048
rect 101458 992 104806 1048
rect 104862 992 104867 1048
rect 101397 990 104867 992
rect 101397 987 101463 990
rect 104801 987 104867 990
rect 111057 1050 111123 1053
rect 111333 1050 111399 1053
rect 111057 1048 111399 1050
rect 111057 992 111062 1048
rect 111118 992 111338 1048
rect 111394 992 111399 1048
rect 111057 990 111399 992
rect 111057 987 111123 990
rect 111333 987 111399 990
rect 118049 1050 118115 1053
rect 119061 1050 119127 1053
rect 118049 1048 119127 1050
rect 118049 992 118054 1048
rect 118110 992 119066 1048
rect 119122 992 119127 1048
rect 118049 990 119127 992
rect 118049 987 118115 990
rect 119061 987 119127 990
rect 125593 1050 125659 1053
rect 126145 1050 126211 1053
rect 133873 1050 133939 1053
rect 125593 1048 133939 1050
rect 125593 992 125598 1048
rect 125654 992 126150 1048
rect 126206 992 133878 1048
rect 133934 992 133939 1048
rect 125593 990 133939 992
rect 125593 987 125659 990
rect 126145 987 126211 990
rect 133873 987 133939 990
rect 55814 854 57162 914
rect 57329 914 57395 917
rect 87597 914 87663 917
rect 57329 912 87663 914
rect 57329 856 57334 912
rect 57390 856 87602 912
rect 87658 856 87663 912
rect 57329 854 87663 856
rect 51460 852 51466 854
rect 55673 851 55739 854
rect 57329 851 57395 854
rect 87597 851 87663 854
rect 91686 852 91692 916
rect 91756 914 91762 916
rect 106365 914 106431 917
rect 91756 912 106431 914
rect 91756 856 106370 912
rect 106426 856 106431 912
rect 91756 854 106431 856
rect 91756 852 91762 854
rect 106365 851 106431 854
rect 106733 914 106799 917
rect 109033 914 109099 917
rect 106733 912 109099 914
rect 106733 856 106738 912
rect 106794 856 109038 912
rect 109094 856 109099 912
rect 106733 854 109099 856
rect 106733 851 106799 854
rect 109033 851 109099 854
rect 131757 914 131823 917
rect 135989 914 136055 917
rect 131757 912 136055 914
rect 131757 856 131762 912
rect 131818 856 135994 912
rect 136050 856 136055 912
rect 131757 854 136055 856
rect 131757 851 131823 854
rect 135989 851 136055 854
rect 5625 778 5691 781
rect 31937 778 32003 781
rect 5625 776 32003 778
rect 5625 720 5630 776
rect 5686 720 31942 776
rect 31998 720 32003 776
rect 5625 718 32003 720
rect 5625 715 5691 718
rect 31937 715 32003 718
rect 35801 778 35867 781
rect 74993 778 75059 781
rect 88977 778 89043 781
rect 35801 776 75059 778
rect 35801 720 35806 776
rect 35862 720 74998 776
rect 75054 720 75059 776
rect 35801 718 75059 720
rect 35801 715 35867 718
rect 74993 715 75059 718
rect 84518 776 89043 778
rect 84518 720 88982 776
rect 89038 720 89043 776
rect 84518 718 89043 720
rect 35801 642 35867 645
rect 46238 642 46244 644
rect 35801 640 46244 642
rect 35801 584 35806 640
rect 35862 584 46244 640
rect 35801 582 46244 584
rect 35801 579 35867 582
rect 46238 580 46244 582
rect 46308 580 46314 644
rect 46381 642 46447 645
rect 51022 642 51028 644
rect 46381 640 51028 642
rect 46381 584 46386 640
rect 46442 584 51028 640
rect 46381 582 51028 584
rect 46381 579 46447 582
rect 51022 580 51028 582
rect 51092 580 51098 644
rect 51206 580 51212 644
rect 51276 642 51282 644
rect 53833 642 53899 645
rect 51276 640 53899 642
rect 51276 584 53838 640
rect 53894 584 53899 640
rect 51276 582 53899 584
rect 51276 580 51282 582
rect 53833 579 53899 582
rect 53966 580 53972 644
rect 54036 642 54042 644
rect 55489 642 55555 645
rect 54036 640 55555 642
rect 54036 584 55494 640
rect 55550 584 55555 640
rect 54036 582 55555 584
rect 54036 580 54042 582
rect 55489 579 55555 582
rect 55673 642 55739 645
rect 57329 642 57395 645
rect 55673 640 57395 642
rect 55673 584 55678 640
rect 55734 584 57334 640
rect 57390 584 57395 640
rect 55673 582 57395 584
rect 55673 579 55739 582
rect 57329 579 57395 582
rect 60457 642 60523 645
rect 61193 642 61259 645
rect 60457 640 61259 642
rect 60457 584 60462 640
rect 60518 584 61198 640
rect 61254 584 61259 640
rect 60457 582 61259 584
rect 60457 579 60523 582
rect 61193 579 61259 582
rect 65006 580 65012 644
rect 65076 642 65082 644
rect 84518 642 84578 718
rect 88977 715 89043 718
rect 107009 778 107075 781
rect 165981 778 166047 781
rect 107009 776 166047 778
rect 107009 720 107014 776
rect 107070 720 165986 776
rect 166042 720 166047 776
rect 107009 718 166047 720
rect 107009 715 107075 718
rect 165981 715 166047 718
rect 65076 582 84578 642
rect 103697 642 103763 645
rect 106365 642 106431 645
rect 103697 640 106431 642
rect 103697 584 103702 640
rect 103758 584 106370 640
rect 106426 584 106431 640
rect 103697 582 106431 584
rect 65076 580 65082 582
rect 103697 579 103763 582
rect 106365 579 106431 582
rect 108481 642 108547 645
rect 114093 642 114159 645
rect 108481 640 114159 642
rect 108481 584 108486 640
rect 108542 584 114098 640
rect 114154 584 114159 640
rect 108481 582 114159 584
rect 108481 579 108547 582
rect 114093 579 114159 582
rect 133965 642 134031 645
rect 137921 642 137987 645
rect 133965 640 137987 642
rect 133965 584 133970 640
rect 134026 584 137926 640
rect 137982 584 137987 640
rect 133965 582 137987 584
rect 133965 579 134031 582
rect 137921 579 137987 582
rect 28418 576 28738 577
rect 28418 512 28426 576
rect 28490 512 28506 576
rect 28570 512 28586 576
rect 28650 512 28666 576
rect 28730 512 28738 576
rect 28418 511 28738 512
rect 84840 576 85160 577
rect 84840 512 84848 576
rect 84912 512 84928 576
rect 84992 512 85008 576
rect 85072 512 85088 576
rect 85152 512 85160 576
rect 84840 511 85160 512
rect 141261 576 141581 577
rect 141261 512 141269 576
rect 141333 512 141349 576
rect 141413 512 141429 576
rect 141493 512 141509 576
rect 141573 512 141581 576
rect 141261 511 141581 512
rect 19241 506 19307 509
rect 27705 506 27771 509
rect 19241 504 27771 506
rect 19241 448 19246 504
rect 19302 448 27710 504
rect 27766 448 27771 504
rect 19241 446 27771 448
rect 19241 443 19307 446
rect 27705 443 27771 446
rect 29085 506 29151 509
rect 32857 506 32923 509
rect 29085 504 32923 506
rect 29085 448 29090 504
rect 29146 448 32862 504
rect 32918 448 32923 504
rect 29085 446 32923 448
rect 29085 443 29151 446
rect 32857 443 32923 446
rect 33133 506 33199 509
rect 34513 506 34579 509
rect 33133 504 34579 506
rect 33133 448 33138 504
rect 33194 448 34518 504
rect 34574 448 34579 504
rect 33133 446 34579 448
rect 33133 443 33199 446
rect 34513 443 34579 446
rect 35249 506 35315 509
rect 36854 506 36860 508
rect 35249 504 36860 506
rect 35249 448 35254 504
rect 35310 448 36860 504
rect 35249 446 36860 448
rect 35249 443 35315 446
rect 36854 444 36860 446
rect 36924 444 36930 508
rect 37089 506 37155 509
rect 40350 506 40356 508
rect 37089 504 40356 506
rect 37089 448 37094 504
rect 37150 448 40356 504
rect 37089 446 40356 448
rect 37089 443 37155 446
rect 40350 444 40356 446
rect 40420 444 40426 508
rect 40493 506 40559 509
rect 41321 506 41387 509
rect 40493 504 41387 506
rect 40493 448 40498 504
rect 40554 448 41326 504
rect 41382 448 41387 504
rect 40493 446 41387 448
rect 40493 443 40559 446
rect 41321 443 41387 446
rect 41454 444 41460 508
rect 41524 506 41530 508
rect 45185 506 45251 509
rect 41524 504 45251 506
rect 41524 448 45190 504
rect 45246 448 45251 504
rect 41524 446 45251 448
rect 41524 444 41530 446
rect 45185 443 45251 446
rect 48313 506 48379 509
rect 53649 506 53715 509
rect 48313 504 53715 506
rect 48313 448 48318 504
rect 48374 448 53654 504
rect 53710 448 53715 504
rect 48313 446 53715 448
rect 48313 443 48379 446
rect 53649 443 53715 446
rect 58566 444 58572 508
rect 58636 506 58642 508
rect 64822 506 64828 508
rect 58636 446 64828 506
rect 58636 444 58642 446
rect 64822 444 64828 446
rect 64892 444 64898 508
rect 6269 370 6335 373
rect 84285 370 84351 373
rect 6269 368 84351 370
rect 6269 312 6274 368
rect 6330 312 84290 368
rect 84346 312 84351 368
rect 6269 310 84351 312
rect 6269 307 6335 310
rect 84285 307 84351 310
rect 24577 234 24643 237
rect 64822 234 64828 236
rect 24577 232 64828 234
rect 24577 176 24582 232
rect 24638 176 64828 232
rect 24577 174 64828 176
rect 24577 171 24643 174
rect 64822 172 64828 174
rect 64892 172 64898 236
rect 65374 172 65380 236
rect 65444 234 65450 236
rect 86125 234 86191 237
rect 65444 232 86191 234
rect 65444 176 86130 232
rect 86186 176 86191 232
rect 65444 174 86191 176
rect 65444 172 65450 174
rect 86125 171 86191 174
rect 14273 98 14339 101
rect 65057 98 65123 101
rect 14273 96 65123 98
rect 14273 40 14278 96
rect 14334 40 65062 96
rect 65118 40 65123 96
rect 14273 38 65123 40
rect 14273 35 14339 38
rect 65057 35 65123 38
rect 65609 98 65675 101
rect 85481 98 85547 101
rect 65609 96 85547 98
rect 65609 40 65614 96
rect 65670 40 85486 96
rect 85542 40 85547 96
rect 65609 38 85547 40
rect 65609 35 65675 38
rect 85481 35 85547 38
<< via3 >>
rect 60044 12956 60108 13020
rect 55444 12004 55508 12068
rect 56637 11996 56701 12000
rect 56637 11940 56641 11996
rect 56641 11940 56697 11996
rect 56697 11940 56701 11996
rect 56637 11936 56701 11940
rect 56717 11996 56781 12000
rect 56717 11940 56721 11996
rect 56721 11940 56777 11996
rect 56777 11940 56781 11996
rect 56717 11936 56781 11940
rect 56797 11996 56861 12000
rect 56797 11940 56801 11996
rect 56801 11940 56857 11996
rect 56857 11940 56861 11996
rect 56797 11936 56861 11940
rect 56877 11996 56941 12000
rect 56877 11940 56881 11996
rect 56881 11940 56937 11996
rect 56937 11940 56941 11996
rect 56877 11936 56941 11940
rect 113058 11996 113122 12000
rect 113058 11940 113062 11996
rect 113062 11940 113118 11996
rect 113118 11940 113122 11996
rect 113058 11936 113122 11940
rect 113138 11996 113202 12000
rect 113138 11940 113142 11996
rect 113142 11940 113198 11996
rect 113198 11940 113202 11996
rect 113138 11936 113202 11940
rect 113218 11996 113282 12000
rect 113218 11940 113222 11996
rect 113222 11940 113278 11996
rect 113278 11940 113282 11996
rect 113218 11936 113282 11940
rect 113298 11996 113362 12000
rect 113298 11940 113302 11996
rect 113302 11940 113358 11996
rect 113358 11940 113362 11996
rect 113298 11936 113362 11940
rect 28426 11452 28490 11456
rect 28426 11396 28430 11452
rect 28430 11396 28486 11452
rect 28486 11396 28490 11452
rect 28426 11392 28490 11396
rect 28506 11452 28570 11456
rect 28506 11396 28510 11452
rect 28510 11396 28566 11452
rect 28566 11396 28570 11452
rect 28506 11392 28570 11396
rect 28586 11452 28650 11456
rect 28586 11396 28590 11452
rect 28590 11396 28646 11452
rect 28646 11396 28650 11452
rect 28586 11392 28650 11396
rect 28666 11452 28730 11456
rect 28666 11396 28670 11452
rect 28670 11396 28726 11452
rect 28726 11396 28730 11452
rect 28666 11392 28730 11396
rect 84848 11452 84912 11456
rect 84848 11396 84852 11452
rect 84852 11396 84908 11452
rect 84908 11396 84912 11452
rect 84848 11392 84912 11396
rect 84928 11452 84992 11456
rect 84928 11396 84932 11452
rect 84932 11396 84988 11452
rect 84988 11396 84992 11452
rect 84928 11392 84992 11396
rect 85008 11452 85072 11456
rect 85008 11396 85012 11452
rect 85012 11396 85068 11452
rect 85068 11396 85072 11452
rect 85008 11392 85072 11396
rect 85088 11452 85152 11456
rect 85088 11396 85092 11452
rect 85092 11396 85148 11452
rect 85148 11396 85152 11452
rect 85088 11392 85152 11396
rect 141269 11452 141333 11456
rect 141269 11396 141273 11452
rect 141273 11396 141329 11452
rect 141329 11396 141333 11452
rect 141269 11392 141333 11396
rect 141349 11452 141413 11456
rect 141349 11396 141353 11452
rect 141353 11396 141409 11452
rect 141409 11396 141413 11452
rect 141349 11392 141413 11396
rect 141429 11452 141493 11456
rect 141429 11396 141433 11452
rect 141433 11396 141489 11452
rect 141489 11396 141493 11452
rect 141429 11392 141493 11396
rect 141509 11452 141573 11456
rect 141509 11396 141513 11452
rect 141513 11396 141569 11452
rect 141569 11396 141573 11452
rect 141509 11392 141573 11396
rect 56637 10908 56701 10912
rect 56637 10852 56641 10908
rect 56641 10852 56697 10908
rect 56697 10852 56701 10908
rect 56637 10848 56701 10852
rect 56717 10908 56781 10912
rect 56717 10852 56721 10908
rect 56721 10852 56777 10908
rect 56777 10852 56781 10908
rect 56717 10848 56781 10852
rect 56797 10908 56861 10912
rect 56797 10852 56801 10908
rect 56801 10852 56857 10908
rect 56857 10852 56861 10908
rect 56797 10848 56861 10852
rect 56877 10908 56941 10912
rect 56877 10852 56881 10908
rect 56881 10852 56937 10908
rect 56937 10852 56941 10908
rect 56877 10848 56941 10852
rect 113058 10908 113122 10912
rect 113058 10852 113062 10908
rect 113062 10852 113118 10908
rect 113118 10852 113122 10908
rect 113058 10848 113122 10852
rect 113138 10908 113202 10912
rect 113138 10852 113142 10908
rect 113142 10852 113198 10908
rect 113198 10852 113202 10908
rect 113138 10848 113202 10852
rect 113218 10908 113282 10912
rect 113218 10852 113222 10908
rect 113222 10852 113278 10908
rect 113278 10852 113282 10908
rect 113218 10848 113282 10852
rect 113298 10908 113362 10912
rect 113298 10852 113302 10908
rect 113302 10852 113358 10908
rect 113358 10852 113362 10908
rect 113298 10848 113362 10852
rect 29132 10508 29196 10572
rect 28426 10364 28490 10368
rect 28426 10308 28430 10364
rect 28430 10308 28486 10364
rect 28486 10308 28490 10364
rect 28426 10304 28490 10308
rect 28506 10364 28570 10368
rect 28506 10308 28510 10364
rect 28510 10308 28566 10364
rect 28566 10308 28570 10364
rect 28506 10304 28570 10308
rect 28586 10364 28650 10368
rect 28586 10308 28590 10364
rect 28590 10308 28646 10364
rect 28646 10308 28650 10364
rect 28586 10304 28650 10308
rect 28666 10364 28730 10368
rect 28666 10308 28670 10364
rect 28670 10308 28726 10364
rect 28726 10308 28730 10364
rect 28666 10304 28730 10308
rect 84848 10364 84912 10368
rect 84848 10308 84852 10364
rect 84852 10308 84908 10364
rect 84908 10308 84912 10364
rect 84848 10304 84912 10308
rect 84928 10364 84992 10368
rect 84928 10308 84932 10364
rect 84932 10308 84988 10364
rect 84988 10308 84992 10364
rect 84928 10304 84992 10308
rect 85008 10364 85072 10368
rect 85008 10308 85012 10364
rect 85012 10308 85068 10364
rect 85068 10308 85072 10364
rect 85008 10304 85072 10308
rect 85088 10364 85152 10368
rect 85088 10308 85092 10364
rect 85092 10308 85148 10364
rect 85148 10308 85152 10364
rect 85088 10304 85152 10308
rect 141269 10364 141333 10368
rect 141269 10308 141273 10364
rect 141273 10308 141329 10364
rect 141329 10308 141333 10364
rect 141269 10304 141333 10308
rect 141349 10364 141413 10368
rect 141349 10308 141353 10364
rect 141353 10308 141409 10364
rect 141409 10308 141413 10364
rect 141349 10304 141413 10308
rect 141429 10364 141493 10368
rect 141429 10308 141433 10364
rect 141433 10308 141489 10364
rect 141489 10308 141493 10364
rect 141429 10304 141493 10308
rect 141509 10364 141573 10368
rect 141509 10308 141513 10364
rect 141513 10308 141569 10364
rect 141569 10308 141573 10364
rect 141509 10304 141573 10308
rect 29132 9828 29196 9892
rect 26004 9692 26068 9756
rect 56637 9820 56701 9824
rect 56637 9764 56641 9820
rect 56641 9764 56697 9820
rect 56697 9764 56701 9820
rect 56637 9760 56701 9764
rect 56717 9820 56781 9824
rect 56717 9764 56721 9820
rect 56721 9764 56777 9820
rect 56777 9764 56781 9820
rect 56717 9760 56781 9764
rect 56797 9820 56861 9824
rect 56797 9764 56801 9820
rect 56801 9764 56857 9820
rect 56857 9764 56861 9820
rect 56797 9760 56861 9764
rect 56877 9820 56941 9824
rect 56877 9764 56881 9820
rect 56881 9764 56937 9820
rect 56937 9764 56941 9820
rect 56877 9760 56941 9764
rect 113058 9820 113122 9824
rect 113058 9764 113062 9820
rect 113062 9764 113118 9820
rect 113118 9764 113122 9820
rect 113058 9760 113122 9764
rect 113138 9820 113202 9824
rect 113138 9764 113142 9820
rect 113142 9764 113198 9820
rect 113198 9764 113202 9820
rect 113138 9760 113202 9764
rect 113218 9820 113282 9824
rect 113218 9764 113222 9820
rect 113222 9764 113278 9820
rect 113278 9764 113282 9820
rect 113218 9760 113282 9764
rect 113298 9820 113362 9824
rect 113298 9764 113302 9820
rect 113302 9764 113358 9820
rect 113358 9764 113362 9820
rect 113298 9760 113362 9764
rect 5580 9208 5644 9212
rect 5580 9152 5594 9208
rect 5594 9152 5644 9208
rect 5580 9148 5644 9152
rect 28426 9276 28490 9280
rect 28426 9220 28430 9276
rect 28430 9220 28486 9276
rect 28486 9220 28490 9276
rect 28426 9216 28490 9220
rect 28506 9276 28570 9280
rect 28506 9220 28510 9276
rect 28510 9220 28566 9276
rect 28566 9220 28570 9276
rect 28506 9216 28570 9220
rect 28586 9276 28650 9280
rect 28586 9220 28590 9276
rect 28590 9220 28646 9276
rect 28646 9220 28650 9276
rect 28586 9216 28650 9220
rect 28666 9276 28730 9280
rect 28666 9220 28670 9276
rect 28670 9220 28726 9276
rect 28726 9220 28730 9276
rect 28666 9216 28730 9220
rect 42380 9148 42444 9212
rect 60044 9284 60108 9348
rect 84848 9276 84912 9280
rect 84848 9220 84852 9276
rect 84852 9220 84908 9276
rect 84908 9220 84912 9276
rect 84848 9216 84912 9220
rect 84928 9276 84992 9280
rect 84928 9220 84932 9276
rect 84932 9220 84988 9276
rect 84988 9220 84992 9276
rect 84928 9216 84992 9220
rect 85008 9276 85072 9280
rect 85008 9220 85012 9276
rect 85012 9220 85068 9276
rect 85068 9220 85072 9276
rect 85008 9216 85072 9220
rect 85088 9276 85152 9280
rect 85088 9220 85092 9276
rect 85092 9220 85148 9276
rect 85148 9220 85152 9276
rect 85088 9216 85152 9220
rect 141269 9276 141333 9280
rect 141269 9220 141273 9276
rect 141273 9220 141329 9276
rect 141329 9220 141333 9276
rect 141269 9216 141333 9220
rect 141349 9276 141413 9280
rect 141349 9220 141353 9276
rect 141353 9220 141409 9276
rect 141409 9220 141413 9276
rect 141349 9216 141413 9220
rect 141429 9276 141493 9280
rect 141429 9220 141433 9276
rect 141433 9220 141489 9276
rect 141489 9220 141493 9276
rect 141429 9216 141493 9220
rect 141509 9276 141573 9280
rect 141509 9220 141513 9276
rect 141513 9220 141569 9276
rect 141569 9220 141573 9276
rect 141509 9216 141573 9220
rect 46428 8876 46492 8940
rect 50292 8740 50356 8804
rect 12204 8392 12268 8396
rect 12204 8336 12218 8392
rect 12218 8336 12268 8392
rect 12204 8332 12268 8336
rect 28426 8188 28490 8192
rect 28426 8132 28430 8188
rect 28430 8132 28486 8188
rect 28486 8132 28490 8188
rect 28426 8128 28490 8132
rect 28506 8188 28570 8192
rect 28506 8132 28510 8188
rect 28510 8132 28566 8188
rect 28566 8132 28570 8188
rect 28506 8128 28570 8132
rect 28586 8188 28650 8192
rect 28586 8132 28590 8188
rect 28590 8132 28646 8188
rect 28646 8132 28650 8188
rect 28586 8128 28650 8132
rect 28666 8188 28730 8192
rect 28666 8132 28670 8188
rect 28670 8132 28726 8188
rect 28726 8132 28730 8188
rect 28666 8128 28730 8132
rect 42932 8468 42996 8532
rect 46428 8604 46492 8668
rect 56637 8732 56701 8736
rect 56637 8676 56641 8732
rect 56641 8676 56697 8732
rect 56697 8676 56701 8732
rect 56637 8672 56701 8676
rect 56717 8732 56781 8736
rect 56717 8676 56721 8732
rect 56721 8676 56777 8732
rect 56777 8676 56781 8732
rect 56717 8672 56781 8676
rect 56797 8732 56861 8736
rect 56797 8676 56801 8732
rect 56801 8676 56857 8732
rect 56857 8676 56861 8732
rect 56797 8672 56861 8676
rect 56877 8732 56941 8736
rect 56877 8676 56881 8732
rect 56881 8676 56937 8732
rect 56937 8676 56941 8732
rect 56877 8672 56941 8676
rect 113058 8732 113122 8736
rect 113058 8676 113062 8732
rect 113062 8676 113118 8732
rect 113118 8676 113122 8732
rect 113058 8672 113122 8676
rect 113138 8732 113202 8736
rect 113138 8676 113142 8732
rect 113142 8676 113198 8732
rect 113198 8676 113202 8732
rect 113138 8672 113202 8676
rect 113218 8732 113282 8736
rect 113218 8676 113222 8732
rect 113222 8676 113278 8732
rect 113278 8676 113282 8732
rect 113218 8672 113282 8676
rect 113298 8732 113362 8736
rect 113298 8676 113302 8732
rect 113302 8676 113358 8732
rect 113358 8676 113362 8732
rect 113298 8672 113362 8676
rect 50844 8332 50908 8396
rect 84848 8188 84912 8192
rect 84848 8132 84852 8188
rect 84852 8132 84908 8188
rect 84908 8132 84912 8188
rect 84848 8128 84912 8132
rect 84928 8188 84992 8192
rect 84928 8132 84932 8188
rect 84932 8132 84988 8188
rect 84988 8132 84992 8188
rect 84928 8128 84992 8132
rect 85008 8188 85072 8192
rect 85008 8132 85012 8188
rect 85012 8132 85068 8188
rect 85068 8132 85072 8188
rect 85008 8128 85072 8132
rect 85088 8188 85152 8192
rect 85088 8132 85092 8188
rect 85092 8132 85148 8188
rect 85148 8132 85152 8188
rect 85088 8128 85152 8132
rect 141269 8188 141333 8192
rect 141269 8132 141273 8188
rect 141273 8132 141329 8188
rect 141329 8132 141333 8188
rect 141269 8128 141333 8132
rect 141349 8188 141413 8192
rect 141349 8132 141353 8188
rect 141353 8132 141409 8188
rect 141409 8132 141413 8188
rect 141349 8128 141413 8132
rect 141429 8188 141493 8192
rect 141429 8132 141433 8188
rect 141433 8132 141489 8188
rect 141489 8132 141493 8188
rect 141429 8128 141493 8132
rect 141509 8188 141573 8192
rect 141509 8132 141513 8188
rect 141513 8132 141569 8188
rect 141569 8132 141573 8188
rect 141509 8128 141573 8132
rect 55444 7712 55508 7716
rect 57284 7788 57348 7852
rect 55444 7656 55494 7712
rect 55494 7656 55508 7712
rect 55444 7652 55508 7656
rect 103468 7652 103532 7716
rect 56637 7644 56701 7648
rect 56637 7588 56641 7644
rect 56641 7588 56697 7644
rect 56697 7588 56701 7644
rect 56637 7584 56701 7588
rect 56717 7644 56781 7648
rect 56717 7588 56721 7644
rect 56721 7588 56777 7644
rect 56777 7588 56781 7644
rect 56717 7584 56781 7588
rect 56797 7644 56861 7648
rect 56797 7588 56801 7644
rect 56801 7588 56857 7644
rect 56857 7588 56861 7644
rect 56797 7584 56861 7588
rect 56877 7644 56941 7648
rect 56877 7588 56881 7644
rect 56881 7588 56937 7644
rect 56937 7588 56941 7644
rect 56877 7584 56941 7588
rect 113058 7644 113122 7648
rect 113058 7588 113062 7644
rect 113062 7588 113118 7644
rect 113118 7588 113122 7644
rect 113058 7584 113122 7588
rect 113138 7644 113202 7648
rect 113138 7588 113142 7644
rect 113142 7588 113198 7644
rect 113198 7588 113202 7644
rect 113138 7584 113202 7588
rect 113218 7644 113282 7648
rect 113218 7588 113222 7644
rect 113222 7588 113278 7644
rect 113278 7588 113282 7644
rect 113218 7584 113282 7588
rect 113298 7644 113362 7648
rect 113298 7588 113302 7644
rect 113302 7588 113358 7644
rect 113358 7588 113362 7644
rect 113298 7584 113362 7588
rect 26142 7380 26206 7444
rect 153148 7380 153212 7444
rect 28426 7100 28490 7104
rect 28426 7044 28430 7100
rect 28430 7044 28486 7100
rect 28486 7044 28490 7100
rect 28426 7040 28490 7044
rect 28506 7100 28570 7104
rect 28506 7044 28510 7100
rect 28510 7044 28566 7100
rect 28566 7044 28570 7100
rect 28506 7040 28570 7044
rect 28586 7100 28650 7104
rect 28586 7044 28590 7100
rect 28590 7044 28646 7100
rect 28646 7044 28650 7100
rect 28586 7040 28650 7044
rect 28666 7100 28730 7104
rect 28666 7044 28670 7100
rect 28670 7044 28726 7100
rect 28726 7044 28730 7100
rect 28666 7040 28730 7044
rect 80284 7108 80348 7172
rect 103468 7244 103532 7308
rect 84848 7100 84912 7104
rect 84848 7044 84852 7100
rect 84852 7044 84908 7100
rect 84908 7044 84912 7100
rect 84848 7040 84912 7044
rect 84928 7100 84992 7104
rect 84928 7044 84932 7100
rect 84932 7044 84988 7100
rect 84988 7044 84992 7100
rect 84928 7040 84992 7044
rect 85008 7100 85072 7104
rect 85008 7044 85012 7100
rect 85012 7044 85068 7100
rect 85068 7044 85072 7100
rect 85008 7040 85072 7044
rect 85088 7100 85152 7104
rect 85088 7044 85092 7100
rect 85092 7044 85148 7100
rect 85148 7044 85152 7100
rect 85088 7040 85152 7044
rect 141269 7100 141333 7104
rect 141269 7044 141273 7100
rect 141273 7044 141329 7100
rect 141329 7044 141333 7100
rect 141269 7040 141333 7044
rect 141349 7100 141413 7104
rect 141349 7044 141353 7100
rect 141353 7044 141409 7100
rect 141409 7044 141413 7100
rect 141349 7040 141413 7044
rect 141429 7100 141493 7104
rect 141429 7044 141433 7100
rect 141433 7044 141489 7100
rect 141489 7044 141493 7100
rect 141429 7040 141493 7044
rect 141509 7100 141573 7104
rect 141509 7044 141513 7100
rect 141513 7044 141569 7100
rect 141569 7044 141573 7100
rect 141509 7040 141573 7044
rect 51580 6836 51644 6900
rect 56637 6556 56701 6560
rect 56637 6500 56641 6556
rect 56641 6500 56697 6556
rect 56697 6500 56701 6556
rect 56637 6496 56701 6500
rect 56717 6556 56781 6560
rect 56717 6500 56721 6556
rect 56721 6500 56777 6556
rect 56777 6500 56781 6556
rect 56717 6496 56781 6500
rect 56797 6556 56861 6560
rect 56797 6500 56801 6556
rect 56801 6500 56857 6556
rect 56857 6500 56861 6556
rect 56797 6496 56861 6500
rect 56877 6556 56941 6560
rect 56877 6500 56881 6556
rect 56881 6500 56937 6556
rect 56937 6500 56941 6556
rect 56877 6496 56941 6500
rect 55996 6488 56060 6492
rect 55996 6432 56046 6488
rect 56046 6432 56060 6488
rect 55996 6428 56060 6432
rect 113058 6556 113122 6560
rect 113058 6500 113062 6556
rect 113062 6500 113118 6556
rect 113118 6500 113122 6556
rect 113058 6496 113122 6500
rect 113138 6556 113202 6560
rect 113138 6500 113142 6556
rect 113142 6500 113198 6556
rect 113198 6500 113202 6556
rect 113138 6496 113202 6500
rect 113218 6556 113282 6560
rect 113218 6500 113222 6556
rect 113222 6500 113278 6556
rect 113278 6500 113282 6556
rect 113218 6496 113282 6500
rect 113298 6556 113362 6560
rect 113298 6500 113302 6556
rect 113302 6500 113358 6556
rect 113358 6500 113362 6556
rect 113298 6496 113362 6500
rect 69060 6020 69124 6084
rect 28426 6012 28490 6016
rect 28426 5956 28430 6012
rect 28430 5956 28486 6012
rect 28486 5956 28490 6012
rect 28426 5952 28490 5956
rect 28506 6012 28570 6016
rect 28506 5956 28510 6012
rect 28510 5956 28566 6012
rect 28566 5956 28570 6012
rect 28506 5952 28570 5956
rect 28586 6012 28650 6016
rect 28586 5956 28590 6012
rect 28590 5956 28646 6012
rect 28646 5956 28650 6012
rect 28586 5952 28650 5956
rect 28666 6012 28730 6016
rect 28666 5956 28670 6012
rect 28670 5956 28726 6012
rect 28726 5956 28730 6012
rect 28666 5952 28730 5956
rect 84848 6012 84912 6016
rect 84848 5956 84852 6012
rect 84852 5956 84908 6012
rect 84908 5956 84912 6012
rect 84848 5952 84912 5956
rect 84928 6012 84992 6016
rect 84928 5956 84932 6012
rect 84932 5956 84988 6012
rect 84988 5956 84992 6012
rect 84928 5952 84992 5956
rect 85008 6012 85072 6016
rect 85008 5956 85012 6012
rect 85012 5956 85068 6012
rect 85068 5956 85072 6012
rect 85008 5952 85072 5956
rect 85088 6012 85152 6016
rect 85088 5956 85092 6012
rect 85092 5956 85148 6012
rect 85148 5956 85152 6012
rect 85088 5952 85152 5956
rect 60964 5884 61028 5948
rect 67588 5884 67652 5948
rect 141269 6012 141333 6016
rect 141269 5956 141273 6012
rect 141273 5956 141329 6012
rect 141329 5956 141333 6012
rect 141269 5952 141333 5956
rect 141349 6012 141413 6016
rect 141349 5956 141353 6012
rect 141353 5956 141409 6012
rect 141409 5956 141413 6012
rect 141349 5952 141413 5956
rect 141429 6012 141493 6016
rect 141429 5956 141433 6012
rect 141433 5956 141489 6012
rect 141489 5956 141493 6012
rect 141429 5952 141493 5956
rect 141509 6012 141573 6016
rect 141509 5956 141513 6012
rect 141513 5956 141569 6012
rect 141569 5956 141573 6012
rect 141509 5952 141573 5956
rect 51396 5612 51460 5676
rect 61700 5612 61764 5676
rect 56637 5468 56701 5472
rect 56637 5412 56641 5468
rect 56641 5412 56697 5468
rect 56697 5412 56701 5468
rect 56637 5408 56701 5412
rect 56717 5468 56781 5472
rect 56717 5412 56721 5468
rect 56721 5412 56777 5468
rect 56777 5412 56781 5468
rect 56717 5408 56781 5412
rect 56797 5468 56861 5472
rect 56797 5412 56801 5468
rect 56801 5412 56857 5468
rect 56857 5412 56861 5468
rect 56797 5408 56861 5412
rect 56877 5468 56941 5472
rect 56877 5412 56881 5468
rect 56881 5412 56937 5468
rect 56937 5412 56941 5468
rect 56877 5408 56941 5412
rect 55812 5204 55876 5268
rect 113058 5468 113122 5472
rect 113058 5412 113062 5468
rect 113062 5412 113118 5468
rect 113118 5412 113122 5468
rect 113058 5408 113122 5412
rect 113138 5468 113202 5472
rect 113138 5412 113142 5468
rect 113142 5412 113198 5468
rect 113198 5412 113202 5468
rect 113138 5408 113202 5412
rect 113218 5468 113282 5472
rect 113218 5412 113222 5468
rect 113222 5412 113278 5468
rect 113278 5412 113282 5468
rect 113218 5408 113282 5412
rect 113298 5468 113362 5472
rect 113298 5412 113302 5468
rect 113302 5412 113358 5468
rect 113358 5412 113362 5468
rect 113298 5408 113362 5412
rect 41644 5068 41708 5132
rect 55260 5068 55324 5132
rect 36676 4932 36740 4996
rect 28426 4924 28490 4928
rect 28426 4868 28430 4924
rect 28430 4868 28486 4924
rect 28486 4868 28490 4924
rect 28426 4864 28490 4868
rect 28506 4924 28570 4928
rect 28506 4868 28510 4924
rect 28510 4868 28566 4924
rect 28566 4868 28570 4924
rect 28506 4864 28570 4868
rect 28586 4924 28650 4928
rect 28586 4868 28590 4924
rect 28590 4868 28646 4924
rect 28646 4868 28650 4924
rect 28586 4864 28650 4868
rect 28666 4924 28730 4928
rect 28666 4868 28670 4924
rect 28670 4868 28726 4924
rect 28726 4868 28730 4924
rect 28666 4864 28730 4868
rect 84848 4924 84912 4928
rect 84848 4868 84852 4924
rect 84852 4868 84908 4924
rect 84908 4868 84912 4924
rect 84848 4864 84912 4868
rect 84928 4924 84992 4928
rect 84928 4868 84932 4924
rect 84932 4868 84988 4924
rect 84988 4868 84992 4924
rect 84928 4864 84992 4868
rect 85008 4924 85072 4928
rect 85008 4868 85012 4924
rect 85012 4868 85068 4924
rect 85068 4868 85072 4924
rect 85008 4864 85072 4868
rect 85088 4924 85152 4928
rect 85088 4868 85092 4924
rect 85092 4868 85148 4924
rect 85148 4868 85152 4924
rect 85088 4864 85152 4868
rect 141269 4924 141333 4928
rect 141269 4868 141273 4924
rect 141273 4868 141329 4924
rect 141329 4868 141333 4924
rect 141269 4864 141333 4868
rect 141349 4924 141413 4928
rect 141349 4868 141353 4924
rect 141353 4868 141409 4924
rect 141409 4868 141413 4924
rect 141349 4864 141413 4868
rect 141429 4924 141493 4928
rect 141429 4868 141433 4924
rect 141433 4868 141489 4924
rect 141489 4868 141493 4924
rect 141429 4864 141493 4868
rect 141509 4924 141573 4928
rect 141509 4868 141513 4924
rect 141513 4868 141569 4924
rect 141569 4868 141573 4924
rect 141509 4864 141573 4868
rect 12388 4388 12452 4452
rect 41644 4388 41708 4452
rect 56637 4380 56701 4384
rect 56637 4324 56641 4380
rect 56641 4324 56697 4380
rect 56697 4324 56701 4380
rect 56637 4320 56701 4324
rect 56717 4380 56781 4384
rect 56717 4324 56721 4380
rect 56721 4324 56777 4380
rect 56777 4324 56781 4380
rect 56717 4320 56781 4324
rect 56797 4380 56861 4384
rect 56797 4324 56801 4380
rect 56801 4324 56857 4380
rect 56857 4324 56861 4380
rect 56797 4320 56861 4324
rect 56877 4380 56941 4384
rect 56877 4324 56881 4380
rect 56881 4324 56937 4380
rect 56937 4324 56941 4380
rect 56877 4320 56941 4324
rect 89668 4388 89732 4452
rect 113058 4380 113122 4384
rect 113058 4324 113062 4380
rect 113062 4324 113118 4380
rect 113118 4324 113122 4380
rect 113058 4320 113122 4324
rect 113138 4380 113202 4384
rect 113138 4324 113142 4380
rect 113142 4324 113198 4380
rect 113198 4324 113202 4380
rect 113138 4320 113202 4324
rect 113218 4380 113282 4384
rect 113218 4324 113222 4380
rect 113222 4324 113278 4380
rect 113278 4324 113282 4380
rect 113218 4320 113282 4324
rect 113298 4380 113362 4384
rect 113298 4324 113302 4380
rect 113302 4324 113358 4380
rect 113358 4324 113362 4380
rect 113298 4320 113362 4324
rect 12756 4116 12820 4180
rect 36676 4116 36740 4180
rect 46612 4116 46676 4180
rect 51028 4116 51092 4180
rect 6316 3844 6380 3908
rect 28426 3836 28490 3840
rect 28426 3780 28430 3836
rect 28430 3780 28486 3836
rect 28486 3780 28490 3836
rect 28426 3776 28490 3780
rect 28506 3836 28570 3840
rect 28506 3780 28510 3836
rect 28510 3780 28566 3836
rect 28566 3780 28570 3836
rect 28506 3776 28570 3780
rect 28586 3836 28650 3840
rect 28586 3780 28590 3836
rect 28590 3780 28646 3836
rect 28646 3780 28650 3836
rect 28586 3776 28650 3780
rect 28666 3836 28730 3840
rect 28666 3780 28670 3836
rect 28670 3780 28726 3836
rect 28726 3780 28730 3836
rect 28666 3776 28730 3780
rect 84848 3836 84912 3840
rect 84848 3780 84852 3836
rect 84852 3780 84908 3836
rect 84908 3780 84912 3836
rect 84848 3776 84912 3780
rect 84928 3836 84992 3840
rect 84928 3780 84932 3836
rect 84932 3780 84988 3836
rect 84988 3780 84992 3836
rect 84928 3776 84992 3780
rect 85008 3836 85072 3840
rect 85008 3780 85012 3836
rect 85012 3780 85068 3836
rect 85068 3780 85072 3836
rect 85008 3776 85072 3780
rect 85088 3836 85152 3840
rect 85088 3780 85092 3836
rect 85092 3780 85148 3836
rect 85148 3780 85152 3836
rect 85088 3776 85152 3780
rect 141269 3836 141333 3840
rect 141269 3780 141273 3836
rect 141273 3780 141329 3836
rect 141329 3780 141333 3836
rect 141269 3776 141333 3780
rect 141349 3836 141413 3840
rect 141349 3780 141353 3836
rect 141353 3780 141409 3836
rect 141409 3780 141413 3836
rect 141349 3776 141413 3780
rect 141429 3836 141493 3840
rect 141429 3780 141433 3836
rect 141433 3780 141489 3836
rect 141489 3780 141493 3836
rect 141429 3776 141493 3780
rect 141509 3836 141573 3840
rect 141509 3780 141513 3836
rect 141513 3780 141569 3836
rect 141569 3780 141573 3836
rect 141509 3776 141573 3780
rect 6684 3768 6748 3772
rect 6684 3712 6698 3768
rect 6698 3712 6748 3768
rect 6684 3708 6748 3712
rect 51396 3708 51460 3772
rect 51764 3572 51828 3636
rect 31892 3300 31956 3364
rect 51028 3164 51092 3228
rect 56637 3292 56701 3296
rect 56637 3236 56641 3292
rect 56641 3236 56697 3292
rect 56697 3236 56701 3292
rect 56637 3232 56701 3236
rect 56717 3292 56781 3296
rect 56717 3236 56721 3292
rect 56721 3236 56777 3292
rect 56777 3236 56781 3292
rect 56717 3232 56781 3236
rect 56797 3292 56861 3296
rect 56797 3236 56801 3292
rect 56801 3236 56857 3292
rect 56857 3236 56861 3292
rect 56797 3232 56861 3236
rect 56877 3292 56941 3296
rect 56877 3236 56881 3292
rect 56881 3236 56937 3292
rect 56937 3236 56941 3292
rect 56877 3232 56941 3236
rect 113058 3292 113122 3296
rect 113058 3236 113062 3292
rect 113062 3236 113118 3292
rect 113118 3236 113122 3292
rect 113058 3232 113122 3236
rect 113138 3292 113202 3296
rect 113138 3236 113142 3292
rect 113142 3236 113198 3292
rect 113198 3236 113202 3292
rect 113138 3232 113202 3236
rect 113218 3292 113282 3296
rect 113218 3236 113222 3292
rect 113222 3236 113278 3292
rect 113278 3236 113282 3292
rect 113218 3232 113282 3236
rect 113298 3292 113362 3296
rect 113298 3236 113302 3292
rect 113302 3236 113358 3292
rect 113358 3236 113362 3292
rect 113298 3232 113362 3236
rect 69060 3164 69124 3228
rect 31708 2756 31772 2820
rect 35940 2756 36004 2820
rect 38332 2756 38396 2820
rect 40540 2756 40604 2820
rect 28426 2748 28490 2752
rect 28426 2692 28430 2748
rect 28430 2692 28486 2748
rect 28486 2692 28490 2748
rect 28426 2688 28490 2692
rect 28506 2748 28570 2752
rect 28506 2692 28510 2748
rect 28510 2692 28566 2748
rect 28566 2692 28570 2748
rect 28506 2688 28570 2692
rect 28586 2748 28650 2752
rect 28586 2692 28590 2748
rect 28590 2692 28646 2748
rect 28646 2692 28650 2748
rect 28586 2688 28650 2692
rect 28666 2748 28730 2752
rect 28666 2692 28670 2748
rect 28670 2692 28726 2748
rect 28726 2692 28730 2748
rect 28666 2688 28730 2692
rect 84848 2748 84912 2752
rect 84848 2692 84852 2748
rect 84852 2692 84908 2748
rect 84908 2692 84912 2748
rect 84848 2688 84912 2692
rect 84928 2748 84992 2752
rect 84928 2692 84932 2748
rect 84932 2692 84988 2748
rect 84988 2692 84992 2748
rect 84928 2688 84992 2692
rect 85008 2748 85072 2752
rect 85008 2692 85012 2748
rect 85012 2692 85068 2748
rect 85068 2692 85072 2748
rect 85008 2688 85072 2692
rect 85088 2748 85152 2752
rect 85088 2692 85092 2748
rect 85092 2692 85148 2748
rect 85148 2692 85152 2748
rect 85088 2688 85152 2692
rect 141269 2748 141333 2752
rect 141269 2692 141273 2748
rect 141273 2692 141329 2748
rect 141329 2692 141333 2748
rect 141269 2688 141333 2692
rect 141349 2748 141413 2752
rect 141349 2692 141353 2748
rect 141353 2692 141409 2748
rect 141409 2692 141413 2748
rect 141349 2688 141413 2692
rect 141429 2748 141493 2752
rect 141429 2692 141433 2748
rect 141433 2692 141489 2748
rect 141489 2692 141493 2748
rect 141429 2688 141493 2692
rect 141509 2748 141573 2752
rect 141509 2692 141513 2748
rect 141513 2692 141569 2748
rect 141569 2692 141573 2748
rect 141509 2688 141573 2692
rect 86908 2620 86972 2684
rect 89668 2680 89732 2684
rect 89668 2624 89718 2680
rect 89718 2624 89732 2680
rect 89668 2620 89732 2624
rect 153148 2484 153212 2548
rect 46060 2212 46124 2276
rect 46428 2348 46492 2412
rect 56637 2204 56701 2208
rect 56637 2148 56641 2204
rect 56641 2148 56697 2204
rect 56697 2148 56701 2204
rect 56637 2144 56701 2148
rect 56717 2204 56781 2208
rect 56717 2148 56721 2204
rect 56721 2148 56777 2204
rect 56777 2148 56781 2204
rect 56717 2144 56781 2148
rect 56797 2204 56861 2208
rect 56797 2148 56801 2204
rect 56801 2148 56857 2204
rect 56857 2148 56861 2204
rect 56797 2144 56861 2148
rect 56877 2204 56941 2208
rect 56877 2148 56881 2204
rect 56881 2148 56937 2204
rect 56937 2148 56941 2204
rect 56877 2144 56941 2148
rect 55996 2136 56060 2140
rect 55996 2080 56010 2136
rect 56010 2080 56060 2136
rect 55996 2076 56060 2080
rect 113058 2204 113122 2208
rect 113058 2148 113062 2204
rect 113062 2148 113118 2204
rect 113118 2148 113122 2204
rect 113058 2144 113122 2148
rect 113138 2204 113202 2208
rect 113138 2148 113142 2204
rect 113142 2148 113198 2204
rect 113198 2148 113202 2204
rect 113138 2144 113202 2148
rect 113218 2204 113282 2208
rect 113218 2148 113222 2204
rect 113222 2148 113278 2204
rect 113278 2148 113282 2204
rect 113218 2144 113282 2148
rect 113298 2204 113362 2208
rect 113298 2148 113302 2204
rect 113302 2148 113358 2204
rect 113358 2148 113362 2204
rect 113298 2144 113362 2148
rect 67588 1668 67652 1732
rect 111748 1668 111812 1732
rect 28426 1660 28490 1664
rect 28426 1604 28430 1660
rect 28430 1604 28486 1660
rect 28486 1604 28490 1660
rect 28426 1600 28490 1604
rect 28506 1660 28570 1664
rect 28506 1604 28510 1660
rect 28510 1604 28566 1660
rect 28566 1604 28570 1660
rect 28506 1600 28570 1604
rect 28586 1660 28650 1664
rect 28586 1604 28590 1660
rect 28590 1604 28646 1660
rect 28646 1604 28650 1660
rect 28586 1600 28650 1604
rect 28666 1660 28730 1664
rect 28666 1604 28670 1660
rect 28670 1604 28726 1660
rect 28726 1604 28730 1660
rect 28666 1600 28730 1604
rect 84848 1660 84912 1664
rect 84848 1604 84852 1660
rect 84852 1604 84908 1660
rect 84908 1604 84912 1660
rect 84848 1600 84912 1604
rect 84928 1660 84992 1664
rect 84928 1604 84932 1660
rect 84932 1604 84988 1660
rect 84988 1604 84992 1660
rect 84928 1600 84992 1604
rect 85008 1660 85072 1664
rect 85008 1604 85012 1660
rect 85012 1604 85068 1660
rect 85068 1604 85072 1660
rect 85008 1600 85072 1604
rect 85088 1660 85152 1664
rect 85088 1604 85092 1660
rect 85092 1604 85148 1660
rect 85148 1604 85152 1660
rect 85088 1600 85152 1604
rect 141269 1660 141333 1664
rect 141269 1604 141273 1660
rect 141273 1604 141329 1660
rect 141329 1604 141333 1660
rect 141269 1600 141333 1604
rect 141349 1660 141413 1664
rect 141349 1604 141353 1660
rect 141353 1604 141409 1660
rect 141409 1604 141413 1660
rect 141349 1600 141413 1604
rect 141429 1660 141493 1664
rect 141429 1604 141433 1660
rect 141433 1604 141489 1660
rect 141489 1604 141493 1660
rect 141429 1600 141493 1604
rect 141509 1660 141573 1664
rect 141509 1604 141513 1660
rect 141513 1604 141569 1660
rect 141569 1604 141573 1660
rect 141509 1600 141573 1604
rect 11284 1456 11348 1460
rect 11284 1400 11298 1456
rect 11298 1400 11348 1456
rect 11284 1396 11348 1400
rect 36308 1260 36372 1324
rect 38884 1260 38948 1324
rect 44036 1124 44100 1188
rect 50660 1124 50724 1188
rect 56637 1116 56701 1120
rect 56637 1060 56641 1116
rect 56641 1060 56697 1116
rect 56697 1060 56701 1116
rect 56637 1056 56701 1060
rect 56717 1116 56781 1120
rect 56717 1060 56721 1116
rect 56721 1060 56777 1116
rect 56777 1060 56781 1116
rect 56717 1056 56781 1060
rect 56797 1116 56861 1120
rect 56797 1060 56801 1116
rect 56801 1060 56857 1116
rect 56857 1060 56861 1116
rect 56797 1056 56861 1060
rect 56877 1116 56941 1120
rect 56877 1060 56881 1116
rect 56881 1060 56937 1116
rect 56937 1060 56941 1116
rect 56877 1056 56941 1060
rect 49924 852 49988 916
rect 51396 852 51460 916
rect 113058 1116 113122 1120
rect 113058 1060 113062 1116
rect 113062 1060 113118 1116
rect 113118 1060 113122 1116
rect 113058 1056 113122 1060
rect 113138 1116 113202 1120
rect 113138 1060 113142 1116
rect 113142 1060 113198 1116
rect 113198 1060 113202 1116
rect 113138 1056 113202 1060
rect 113218 1116 113282 1120
rect 113218 1060 113222 1116
rect 113222 1060 113278 1116
rect 113278 1060 113282 1116
rect 113218 1056 113282 1060
rect 113298 1116 113362 1120
rect 113298 1060 113302 1116
rect 113302 1060 113358 1116
rect 113358 1060 113362 1116
rect 113298 1056 113362 1060
rect 91692 852 91756 916
rect 46244 580 46308 644
rect 51028 580 51092 644
rect 51212 580 51276 644
rect 53972 580 54036 644
rect 65012 580 65076 644
rect 28426 572 28490 576
rect 28426 516 28430 572
rect 28430 516 28486 572
rect 28486 516 28490 572
rect 28426 512 28490 516
rect 28506 572 28570 576
rect 28506 516 28510 572
rect 28510 516 28566 572
rect 28566 516 28570 572
rect 28506 512 28570 516
rect 28586 572 28650 576
rect 28586 516 28590 572
rect 28590 516 28646 572
rect 28646 516 28650 572
rect 28586 512 28650 516
rect 28666 572 28730 576
rect 28666 516 28670 572
rect 28670 516 28726 572
rect 28726 516 28730 572
rect 28666 512 28730 516
rect 84848 572 84912 576
rect 84848 516 84852 572
rect 84852 516 84908 572
rect 84908 516 84912 572
rect 84848 512 84912 516
rect 84928 572 84992 576
rect 84928 516 84932 572
rect 84932 516 84988 572
rect 84988 516 84992 572
rect 84928 512 84992 516
rect 85008 572 85072 576
rect 85008 516 85012 572
rect 85012 516 85068 572
rect 85068 516 85072 572
rect 85008 512 85072 516
rect 85088 572 85152 576
rect 85088 516 85092 572
rect 85092 516 85148 572
rect 85148 516 85152 572
rect 85088 512 85152 516
rect 141269 572 141333 576
rect 141269 516 141273 572
rect 141273 516 141329 572
rect 141329 516 141333 572
rect 141269 512 141333 516
rect 141349 572 141413 576
rect 141349 516 141353 572
rect 141353 516 141409 572
rect 141409 516 141413 572
rect 141349 512 141413 516
rect 141429 572 141493 576
rect 141429 516 141433 572
rect 141433 516 141489 572
rect 141489 516 141493 572
rect 141429 512 141493 516
rect 141509 572 141573 576
rect 141509 516 141513 572
rect 141513 516 141569 572
rect 141569 516 141573 572
rect 141509 512 141573 516
rect 36860 444 36924 508
rect 40356 444 40420 508
rect 41460 444 41524 508
rect 58572 444 58636 508
rect 64828 444 64892 508
rect 64828 172 64892 236
rect 65380 172 65444 236
<< metal4 >>
rect 60043 13020 60109 13021
rect 60043 12956 60044 13020
rect 60108 12956 60109 13020
rect 60043 12955 60109 12956
rect 55443 12068 55509 12069
rect 28418 11456 28738 12016
rect 55443 12004 55444 12068
rect 55508 12004 55509 12068
rect 55443 12003 55509 12004
rect 28418 11392 28426 11456
rect 28490 11392 28506 11456
rect 28570 11392 28586 11456
rect 28650 11392 28666 11456
rect 28730 11392 28738 11456
rect 28418 10540 28738 11392
rect 28418 10368 28460 10540
rect 28696 10368 28738 10540
rect 29131 10572 29197 10573
rect 29131 10508 29132 10572
rect 29196 10508 29197 10572
rect 29131 10507 29197 10508
rect 28418 10304 28426 10368
rect 28730 10304 28738 10368
rect 26003 9756 26069 9757
rect 26003 9692 26004 9756
rect 26068 9692 26069 9756
rect 26003 9691 26069 9692
rect 12203 8396 12269 8397
rect 12203 8332 12204 8396
rect 12268 8332 12269 8396
rect 12203 8331 12269 8332
rect 12206 7258 12266 8331
rect 26006 7850 26066 9691
rect 28418 9280 28738 10304
rect 29134 9893 29194 10507
rect 29131 9892 29197 9893
rect 29131 9828 29132 9892
rect 29196 9828 29197 9892
rect 29131 9827 29197 9828
rect 28418 9216 28426 9280
rect 28490 9216 28506 9280
rect 28570 9216 28586 9280
rect 28650 9216 28666 9280
rect 28730 9216 28738 9280
rect 28418 8192 28738 9216
rect 42379 9212 42445 9213
rect 42379 9148 42380 9212
rect 42444 9148 42445 9212
rect 42379 9147 42445 9148
rect 42382 8530 42442 9147
rect 46427 8940 46493 8941
rect 46427 8876 46428 8940
rect 46492 8876 46493 8940
rect 46427 8875 46493 8876
rect 46430 8669 46490 8875
rect 50294 8805 50354 9062
rect 50291 8804 50357 8805
rect 50291 8740 50292 8804
rect 50356 8740 50357 8804
rect 50291 8739 50357 8740
rect 46427 8668 46493 8669
rect 46427 8604 46428 8668
rect 46492 8604 46493 8668
rect 46427 8603 46493 8604
rect 42931 8532 42997 8533
rect 42931 8530 42932 8532
rect 42382 8470 42932 8530
rect 42931 8468 42932 8470
rect 42996 8468 42997 8532
rect 42931 8467 42997 8468
rect 50843 8396 50909 8397
rect 50843 8332 50844 8396
rect 50908 8394 50909 8396
rect 51030 8394 51090 9062
rect 50908 8334 51090 8394
rect 50908 8332 50909 8334
rect 50843 8331 50909 8332
rect 28418 8128 28426 8192
rect 28490 8128 28506 8192
rect 28570 8128 28586 8192
rect 28650 8128 28666 8192
rect 28730 8128 28738 8192
rect 26006 7790 26204 7850
rect 26144 7445 26204 7790
rect 26141 7444 26207 7445
rect 26141 7380 26142 7444
rect 26206 7380 26207 7444
rect 26141 7379 26207 7380
rect 28418 7104 28738 8128
rect 55446 7717 55506 12003
rect 56629 12000 56949 12016
rect 56629 11936 56637 12000
rect 56701 11936 56717 12000
rect 56781 11936 56797 12000
rect 56861 11936 56877 12000
rect 56941 11936 56949 12000
rect 56629 10912 56949 11936
rect 56629 10848 56637 10912
rect 56701 10848 56717 10912
rect 56781 10848 56797 10912
rect 56861 10848 56877 10912
rect 56941 10848 56949 10912
rect 56629 9824 56949 10848
rect 56629 9760 56637 9824
rect 56701 9760 56717 9824
rect 56781 9760 56797 9824
rect 56861 9760 56877 9824
rect 56941 9760 56949 9824
rect 56629 8736 56949 9760
rect 60046 9349 60106 12955
rect 84840 11456 85160 12016
rect 84840 11392 84848 11456
rect 84912 11392 84928 11456
rect 84992 11392 85008 11456
rect 85072 11392 85088 11456
rect 85152 11392 85160 11456
rect 84840 10540 85160 11392
rect 84840 10368 84882 10540
rect 85118 10368 85160 10540
rect 84840 10304 84848 10368
rect 85152 10304 85160 10368
rect 60043 9348 60109 9349
rect 60043 9284 60044 9348
rect 60108 9284 60109 9348
rect 60043 9283 60109 9284
rect 84840 9280 85160 10304
rect 84840 9216 84848 9280
rect 84912 9216 84928 9280
rect 84992 9216 85008 9280
rect 85072 9216 85088 9280
rect 85152 9216 85160 9280
rect 56629 8672 56637 8736
rect 56701 8672 56717 8736
rect 56781 8672 56797 8736
rect 56861 8672 56877 8736
rect 56941 8672 56949 8736
rect 56629 8555 56949 8672
rect 56629 8319 56671 8555
rect 56907 8319 56949 8555
rect 55443 7716 55509 7717
rect 55443 7652 55444 7716
rect 55508 7652 55509 7716
rect 55443 7651 55509 7652
rect 28418 7040 28426 7104
rect 28490 7040 28506 7104
rect 28570 7040 28586 7104
rect 28650 7040 28666 7104
rect 28730 7040 28738 7104
rect 28418 6570 28738 7040
rect 56629 7648 56949 8319
rect 57286 7853 57346 9062
rect 84840 8192 85160 9216
rect 84840 8128 84848 8192
rect 84912 8128 84928 8192
rect 84992 8128 85008 8192
rect 85072 8128 85088 8192
rect 85152 8128 85160 8192
rect 57283 7852 57349 7853
rect 57283 7788 57284 7852
rect 57348 7788 57349 7852
rect 57283 7787 57349 7788
rect 56629 7584 56637 7648
rect 56701 7584 56717 7648
rect 56781 7584 56797 7648
rect 56861 7584 56877 7648
rect 56941 7584 56949 7648
rect 51579 6900 51645 6901
rect 51579 6836 51580 6900
rect 51644 6836 51645 6900
rect 51579 6835 51645 6836
rect 28418 6334 28460 6570
rect 28696 6334 28738 6570
rect 28418 6016 28738 6334
rect 28418 5952 28426 6016
rect 28490 5952 28506 6016
rect 28570 5952 28586 6016
rect 28650 5952 28666 6016
rect 28730 5952 28738 6016
rect 6318 3909 6378 5662
rect 28418 4928 28738 5952
rect 51582 5810 51642 6835
rect 56629 6560 56949 7584
rect 84840 7104 85160 8128
rect 113050 12000 113370 12016
rect 113050 11936 113058 12000
rect 113122 11936 113138 12000
rect 113202 11936 113218 12000
rect 113282 11936 113298 12000
rect 113362 11936 113370 12000
rect 113050 10912 113370 11936
rect 113050 10848 113058 10912
rect 113122 10848 113138 10912
rect 113202 10848 113218 10912
rect 113282 10848 113298 10912
rect 113362 10848 113370 10912
rect 113050 9824 113370 10848
rect 113050 9760 113058 9824
rect 113122 9760 113138 9824
rect 113202 9760 113218 9824
rect 113282 9760 113298 9824
rect 113362 9760 113370 9824
rect 113050 8736 113370 9760
rect 113050 8672 113058 8736
rect 113122 8672 113138 8736
rect 113202 8672 113218 8736
rect 113282 8672 113298 8736
rect 113362 8672 113370 8736
rect 113050 8555 113370 8672
rect 113050 8319 113092 8555
rect 113328 8319 113370 8555
rect 103467 7716 103533 7717
rect 103467 7652 103468 7716
rect 103532 7652 103533 7716
rect 103467 7651 103533 7652
rect 103470 7309 103530 7651
rect 113050 7648 113370 8319
rect 113050 7584 113058 7648
rect 113122 7584 113138 7648
rect 113202 7584 113218 7648
rect 113282 7584 113298 7648
rect 113362 7584 113370 7648
rect 103467 7308 103533 7309
rect 103467 7244 103468 7308
rect 103532 7244 103533 7308
rect 103467 7243 103533 7244
rect 84840 7040 84848 7104
rect 84912 7040 84928 7104
rect 84992 7040 85008 7104
rect 85072 7040 85088 7104
rect 85152 7040 85160 7104
rect 56629 6496 56637 6560
rect 56701 6496 56717 6560
rect 56781 6496 56797 6560
rect 56861 6496 56877 6560
rect 56941 6496 56949 6560
rect 55995 6492 56061 6493
rect 55995 6428 55996 6492
rect 56060 6428 56061 6492
rect 55995 6427 56061 6428
rect 51398 5750 51642 5810
rect 51398 5677 51458 5750
rect 51395 5676 51461 5677
rect 51395 5612 51396 5676
rect 51460 5612 51461 5676
rect 51395 5611 51461 5612
rect 55811 5268 55877 5269
rect 55811 5204 55812 5268
rect 55876 5204 55877 5268
rect 55811 5203 55877 5204
rect 41643 5132 41709 5133
rect 41643 5068 41644 5132
rect 41708 5068 41709 5132
rect 41643 5067 41709 5068
rect 55259 5132 55325 5133
rect 55259 5068 55260 5132
rect 55324 5130 55325 5132
rect 55814 5130 55874 5203
rect 55324 5070 55874 5130
rect 55324 5068 55325 5070
rect 55259 5067 55325 5068
rect 36675 4996 36741 4997
rect 36675 4932 36676 4996
rect 36740 4932 36741 4996
rect 36675 4931 36741 4932
rect 28418 4864 28426 4928
rect 28490 4864 28506 4928
rect 28570 4864 28586 4928
rect 28650 4864 28666 4928
rect 28730 4864 28738 4928
rect 12387 4452 12453 4453
rect 12387 4388 12388 4452
rect 12452 4450 12453 4452
rect 12452 4390 12818 4450
rect 12452 4388 12453 4390
rect 12387 4387 12453 4388
rect 12758 4181 12818 4390
rect 12755 4180 12821 4181
rect 12755 4116 12756 4180
rect 12820 4116 12821 4180
rect 12755 4115 12821 4116
rect 6315 3908 6381 3909
rect 6315 3844 6316 3908
rect 6380 3844 6381 3908
rect 6315 3843 6381 3844
rect 28418 3840 28738 4864
rect 36678 4181 36738 4931
rect 41646 4453 41706 5067
rect 41643 4452 41709 4453
rect 41643 4388 41644 4452
rect 41708 4388 41709 4452
rect 41643 4387 41709 4388
rect 36675 4180 36741 4181
rect 36675 4116 36676 4180
rect 36740 4116 36741 4180
rect 36675 4115 36741 4116
rect 46611 4180 46677 4181
rect 46611 4116 46612 4180
rect 46676 4116 46677 4180
rect 46611 4115 46677 4116
rect 51027 4180 51093 4181
rect 51027 4116 51028 4180
rect 51092 4178 51093 4180
rect 51092 4118 51458 4178
rect 51092 4116 51093 4118
rect 51027 4115 51093 4116
rect 28418 3776 28426 3840
rect 28490 3776 28506 3840
rect 28570 3776 28586 3840
rect 28650 3776 28666 3840
rect 28730 3776 28738 3840
rect 28418 2752 28738 3776
rect 31891 3364 31957 3365
rect 31891 3300 31892 3364
rect 31956 3300 31957 3364
rect 31891 3299 31957 3300
rect 31707 2820 31773 2821
rect 31707 2756 31708 2820
rect 31772 2818 31773 2820
rect 31894 2818 31954 3299
rect 31772 2758 31954 2818
rect 35939 2820 36005 2821
rect 31772 2756 31773 2758
rect 31707 2755 31773 2756
rect 35939 2756 35940 2820
rect 36004 2756 36005 2820
rect 35939 2755 36005 2756
rect 38331 2820 38397 2821
rect 38331 2756 38332 2820
rect 38396 2818 38397 2820
rect 40539 2820 40605 2821
rect 40539 2818 40540 2820
rect 38396 2758 40540 2818
rect 38396 2756 38397 2758
rect 38331 2755 38397 2756
rect 40539 2756 40540 2758
rect 40604 2756 40605 2820
rect 40539 2755 40605 2756
rect 28418 2688 28426 2752
rect 28490 2688 28506 2752
rect 28570 2688 28586 2752
rect 28650 2688 28666 2752
rect 28730 2688 28738 2752
rect 28418 2599 28738 2688
rect 28418 2363 28460 2599
rect 28696 2363 28738 2599
rect 28418 1664 28738 2363
rect 28418 1600 28426 1664
rect 28490 1600 28506 1664
rect 28570 1600 28586 1664
rect 28650 1600 28666 1664
rect 28730 1600 28738 1664
rect 11286 1461 11346 1582
rect 11283 1460 11349 1461
rect 11283 1396 11284 1460
rect 11348 1396 11349 1460
rect 11283 1395 11349 1396
rect 28418 576 28738 1600
rect 35942 1138 36002 2755
rect 46427 2412 46493 2413
rect 46427 2410 46428 2412
rect 46062 2350 46428 2410
rect 46062 2277 46122 2350
rect 46427 2348 46428 2350
rect 46492 2348 46493 2412
rect 46427 2347 46493 2348
rect 46059 2276 46125 2277
rect 46059 2212 46060 2276
rect 46124 2212 46125 2276
rect 46059 2211 46125 2212
rect 36307 1324 36373 1325
rect 36307 1260 36308 1324
rect 36372 1322 36373 1324
rect 38883 1324 38949 1325
rect 38883 1322 38884 1324
rect 36372 1262 38884 1322
rect 36372 1260 36373 1262
rect 36307 1259 36373 1260
rect 38883 1260 38884 1262
rect 38948 1260 38949 1324
rect 38883 1259 38949 1260
rect 44035 1188 44101 1189
rect 44035 1124 44036 1188
rect 44100 1124 44101 1188
rect 46614 1138 46674 4115
rect 51398 3773 51458 4118
rect 51395 3772 51461 3773
rect 51395 3708 51396 3772
rect 51460 3708 51461 3772
rect 51395 3707 51461 3708
rect 51030 3229 51090 3622
rect 51763 3572 51764 3622
rect 51828 3572 51829 3622
rect 51763 3571 51829 3572
rect 51027 3228 51093 3229
rect 51027 3164 51028 3228
rect 51092 3164 51093 3228
rect 51027 3163 51093 3164
rect 55998 2141 56058 6427
rect 56629 5472 56949 6496
rect 84840 6570 85160 7040
rect 84840 6334 84882 6570
rect 85118 6334 85160 6570
rect 69059 6084 69125 6085
rect 69059 6020 69060 6084
rect 69124 6020 69125 6084
rect 69059 6019 69125 6020
rect 60963 5948 61029 5949
rect 60963 5898 60964 5948
rect 61028 5898 61029 5948
rect 67587 5948 67653 5949
rect 67587 5884 67588 5948
rect 67652 5884 67653 5948
rect 67587 5883 67653 5884
rect 61699 5612 61700 5662
rect 61764 5612 61765 5662
rect 61699 5611 61765 5612
rect 56629 5408 56637 5472
rect 56701 5408 56717 5472
rect 56781 5408 56797 5472
rect 56861 5408 56877 5472
rect 56941 5408 56949 5472
rect 56629 4584 56949 5408
rect 56629 4384 56671 4584
rect 56907 4384 56949 4584
rect 56629 4320 56637 4384
rect 56701 4320 56717 4348
rect 56781 4320 56797 4348
rect 56861 4320 56877 4348
rect 56941 4320 56949 4384
rect 56629 3296 56949 4320
rect 56629 3232 56637 3296
rect 56701 3232 56717 3296
rect 56781 3232 56797 3296
rect 56861 3232 56877 3296
rect 56941 3232 56949 3296
rect 56629 2208 56949 3232
rect 56629 2144 56637 2208
rect 56701 2144 56717 2208
rect 56781 2144 56797 2208
rect 56861 2144 56877 2208
rect 56941 2144 56949 2208
rect 55995 2140 56061 2141
rect 55995 2076 55996 2140
rect 56060 2076 56061 2140
rect 55995 2075 56061 2076
rect 50659 1188 50725 1189
rect 50659 1138 50660 1188
rect 50724 1138 50725 1188
rect 44035 1123 44101 1124
rect 36862 990 38762 1050
rect 28418 512 28426 576
rect 28490 512 28506 576
rect 28570 512 28586 576
rect 28650 512 28666 576
rect 28730 512 28738 576
rect 28418 496 28738 512
rect 36862 509 36922 990
rect 36859 508 36925 509
rect 36859 444 36860 508
rect 36924 444 36925 508
rect 38702 458 38762 990
rect 40355 508 40421 509
rect 36859 443 36925 444
rect 40355 444 40356 508
rect 40420 506 40421 508
rect 41459 508 41525 509
rect 41459 506 41460 508
rect 40420 446 41460 506
rect 40420 444 40421 446
rect 40355 443 40421 444
rect 41459 444 41460 446
rect 41524 444 41525 508
rect 44038 458 44098 1123
rect 49923 916 49989 917
rect 49923 852 49924 916
rect 49988 852 49989 916
rect 51030 990 51458 1050
rect 49923 851 49989 852
rect 46243 644 46309 645
rect 46243 580 46244 644
rect 46308 580 46309 644
rect 46243 579 46309 580
rect 46246 458 46306 579
rect 41459 443 41525 444
rect 49926 370 49986 851
rect 51030 645 51090 990
rect 51398 917 51458 990
rect 51395 916 51461 917
rect 51395 852 51396 916
rect 51460 852 51461 916
rect 56629 1120 56949 2144
rect 67590 1733 67650 5883
rect 69062 3229 69122 6019
rect 84840 6016 85160 6334
rect 84840 5952 84848 6016
rect 84912 5952 84928 6016
rect 84992 5952 85008 6016
rect 85072 5952 85088 6016
rect 85152 5952 85160 6016
rect 84840 4928 85160 5952
rect 113050 6560 113370 7584
rect 113050 6496 113058 6560
rect 113122 6496 113138 6560
rect 113202 6496 113218 6560
rect 113282 6496 113298 6560
rect 113362 6496 113370 6560
rect 84840 4864 84848 4928
rect 84912 4864 84928 4928
rect 84992 4864 85008 4928
rect 85072 4864 85088 4928
rect 85152 4864 85160 4928
rect 84840 3840 85160 4864
rect 89667 4452 89733 4453
rect 89667 4388 89668 4452
rect 89732 4388 89733 4452
rect 89667 4387 89733 4388
rect 84840 3776 84848 3840
rect 84912 3776 84928 3840
rect 84992 3776 85008 3840
rect 85072 3776 85088 3840
rect 85152 3776 85160 3840
rect 69059 3228 69125 3229
rect 69059 3164 69060 3228
rect 69124 3164 69125 3228
rect 69059 3163 69125 3164
rect 84840 2752 85160 3776
rect 84840 2688 84848 2752
rect 84912 2688 84928 2752
rect 84992 2688 85008 2752
rect 85072 2688 85088 2752
rect 85152 2688 85160 2752
rect 84840 2599 85160 2688
rect 86910 2685 86970 3622
rect 89670 2685 89730 4387
rect 86907 2684 86973 2685
rect 86907 2620 86908 2684
rect 86972 2620 86973 2684
rect 86907 2619 86973 2620
rect 89667 2684 89733 2685
rect 89667 2620 89668 2684
rect 89732 2620 89733 2684
rect 89667 2619 89733 2620
rect 84840 2363 84882 2599
rect 85118 2363 85160 2599
rect 67587 1732 67653 1733
rect 67587 1668 67588 1732
rect 67652 1668 67653 1732
rect 67587 1667 67653 1668
rect 56629 1056 56637 1120
rect 56701 1056 56717 1120
rect 56781 1056 56797 1120
rect 56861 1056 56877 1120
rect 56941 1056 56949 1120
rect 51395 851 51461 852
rect 53974 645 54034 902
rect 51027 644 51093 645
rect 51027 580 51028 644
rect 51092 580 51093 644
rect 51027 579 51093 580
rect 51211 644 51277 645
rect 51211 580 51212 644
rect 51276 580 51277 644
rect 51211 579 51277 580
rect 53971 644 54037 645
rect 53971 580 53972 644
rect 54036 580 54037 644
rect 53971 579 54037 580
rect 51214 370 51274 579
rect 56629 496 56949 1056
rect 84840 1664 85160 2363
rect 84840 1600 84848 1664
rect 84912 1600 84928 1664
rect 84992 1600 85008 1664
rect 85072 1600 85088 1664
rect 85152 1600 85160 1664
rect 64830 990 65074 1050
rect 64830 509 64890 990
rect 65014 645 65074 990
rect 65011 644 65077 645
rect 65011 580 65012 644
rect 65076 580 65077 644
rect 65011 579 65077 580
rect 84840 576 85160 1600
rect 91694 917 91754 5662
rect 113050 5472 113370 6496
rect 113050 5408 113058 5472
rect 113122 5408 113138 5472
rect 113202 5408 113218 5472
rect 113282 5408 113298 5472
rect 113362 5408 113370 5472
rect 113050 4584 113370 5408
rect 113050 4384 113092 4584
rect 113328 4384 113370 4584
rect 113050 4320 113058 4384
rect 113122 4320 113138 4348
rect 113202 4320 113218 4348
rect 113282 4320 113298 4348
rect 113362 4320 113370 4384
rect 113050 3296 113370 4320
rect 113050 3232 113058 3296
rect 113122 3232 113138 3296
rect 113202 3232 113218 3296
rect 113282 3232 113298 3296
rect 113362 3232 113370 3296
rect 113050 2208 113370 3232
rect 113050 2144 113058 2208
rect 113122 2144 113138 2208
rect 113202 2144 113218 2208
rect 113282 2144 113298 2208
rect 113362 2144 113370 2208
rect 113050 1120 113370 2144
rect 113050 1056 113058 1120
rect 113122 1056 113138 1120
rect 113202 1056 113218 1120
rect 113282 1056 113298 1120
rect 113362 1056 113370 1120
rect 91691 916 91757 917
rect 91691 852 91692 916
rect 91756 852 91757 916
rect 91691 851 91757 852
rect 84840 512 84848 576
rect 84912 512 84928 576
rect 84992 512 85008 576
rect 85072 512 85088 576
rect 85152 512 85160 576
rect 58571 508 58637 509
rect 58571 458 58572 508
rect 58636 458 58637 508
rect 64827 508 64893 509
rect 49926 310 51274 370
rect 64827 444 64828 508
rect 64892 444 64893 508
rect 84840 496 85160 512
rect 113050 496 113370 1056
rect 141261 11456 141581 12016
rect 141261 11392 141269 11456
rect 141333 11392 141349 11456
rect 141413 11392 141429 11456
rect 141493 11392 141509 11456
rect 141573 11392 141581 11456
rect 141261 10540 141581 11392
rect 141261 10368 141303 10540
rect 141539 10368 141581 10540
rect 141261 10304 141269 10368
rect 141573 10304 141581 10368
rect 141261 9280 141581 10304
rect 141261 9216 141269 9280
rect 141333 9216 141349 9280
rect 141413 9216 141429 9280
rect 141493 9216 141509 9280
rect 141573 9216 141581 9280
rect 141261 8192 141581 9216
rect 141261 8128 141269 8192
rect 141333 8128 141349 8192
rect 141413 8128 141429 8192
rect 141493 8128 141509 8192
rect 141573 8128 141581 8192
rect 141261 7104 141581 8128
rect 153147 7444 153213 7445
rect 153147 7380 153148 7444
rect 153212 7380 153213 7444
rect 153147 7379 153213 7380
rect 141261 7040 141269 7104
rect 141333 7040 141349 7104
rect 141413 7040 141429 7104
rect 141493 7040 141509 7104
rect 141573 7040 141581 7104
rect 141261 6570 141581 7040
rect 141261 6334 141303 6570
rect 141539 6334 141581 6570
rect 141261 6016 141581 6334
rect 141261 5952 141269 6016
rect 141333 5952 141349 6016
rect 141413 5952 141429 6016
rect 141493 5952 141509 6016
rect 141573 5952 141581 6016
rect 141261 4928 141581 5952
rect 141261 4864 141269 4928
rect 141333 4864 141349 4928
rect 141413 4864 141429 4928
rect 141493 4864 141509 4928
rect 141573 4864 141581 4928
rect 141261 3840 141581 4864
rect 141261 3776 141269 3840
rect 141333 3776 141349 3840
rect 141413 3776 141429 3840
rect 141493 3776 141509 3840
rect 141573 3776 141581 3840
rect 141261 2752 141581 3776
rect 141261 2688 141269 2752
rect 141333 2688 141349 2752
rect 141413 2688 141429 2752
rect 141493 2688 141509 2752
rect 141573 2688 141581 2752
rect 141261 2599 141581 2688
rect 141261 2363 141303 2599
rect 141539 2363 141581 2599
rect 153150 2549 153210 7379
rect 153147 2548 153213 2549
rect 153147 2484 153148 2548
rect 153212 2484 153213 2548
rect 153147 2483 153213 2484
rect 141261 1664 141581 2363
rect 141261 1600 141269 1664
rect 141333 1600 141349 1664
rect 141413 1600 141429 1664
rect 141493 1600 141509 1664
rect 141573 1600 141581 1664
rect 141261 576 141581 1600
rect 141261 512 141269 576
rect 141333 512 141349 576
rect 141413 512 141429 576
rect 141493 512 141509 576
rect 141573 512 141581 576
rect 141261 496 141581 512
rect 64827 443 64893 444
rect 64830 310 65442 370
rect 64830 237 64890 310
rect 65382 237 65442 310
rect 64827 236 64893 237
rect 64827 172 64828 236
rect 64892 172 64893 236
rect 64827 171 64893 172
rect 65379 236 65445 237
rect 65379 172 65380 236
rect 65444 172 65445 236
rect 65379 171 65445 172
<< via4 >>
rect 28460 10368 28696 10540
rect 28460 10304 28490 10368
rect 28490 10304 28506 10368
rect 28506 10304 28570 10368
rect 28570 10304 28586 10368
rect 28586 10304 28650 10368
rect 28650 10304 28666 10368
rect 28666 10304 28696 10368
rect 5494 9212 5730 9298
rect 5494 9148 5580 9212
rect 5580 9148 5644 9212
rect 5644 9148 5730 9212
rect 5494 9062 5730 9148
rect 50206 9062 50442 9298
rect 50942 9062 51178 9298
rect 12118 7022 12354 7258
rect 84882 10368 85118 10540
rect 84882 10304 84912 10368
rect 84912 10304 84928 10368
rect 84928 10304 84992 10368
rect 84992 10304 85008 10368
rect 85008 10304 85072 10368
rect 85072 10304 85088 10368
rect 85088 10304 85118 10368
rect 57198 9062 57434 9298
rect 56671 8319 56907 8555
rect 28460 6334 28696 6570
rect 6230 5662 6466 5898
rect 80198 7172 80434 7258
rect 80198 7108 80284 7172
rect 80284 7108 80348 7172
rect 80348 7108 80434 7172
rect 80198 7022 80434 7108
rect 113092 8319 113328 8555
rect 6598 3772 6834 3858
rect 6598 3708 6684 3772
rect 6684 3708 6748 3772
rect 6748 3708 6834 3772
rect 6598 3622 6834 3708
rect 28460 2363 28696 2599
rect 11198 1582 11434 1818
rect 35854 902 36090 1138
rect 50942 3622 51178 3858
rect 51678 3636 51914 3858
rect 51678 3622 51764 3636
rect 51764 3622 51828 3636
rect 51828 3622 51914 3636
rect 84882 6334 85118 6570
rect 60878 5884 60964 5898
rect 60964 5884 61028 5898
rect 61028 5884 61114 5898
rect 60878 5662 61114 5884
rect 61614 5676 61850 5898
rect 61614 5662 61700 5676
rect 61700 5662 61764 5676
rect 61764 5662 61850 5676
rect 56671 4384 56907 4584
rect 56671 4348 56701 4384
rect 56701 4348 56717 4384
rect 56717 4348 56781 4384
rect 56781 4348 56797 4384
rect 56797 4348 56861 4384
rect 56861 4348 56877 4384
rect 56877 4348 56907 4384
rect 38614 222 38850 458
rect 46526 902 46762 1138
rect 50574 1124 50660 1138
rect 50660 1124 50724 1138
rect 50724 1124 50810 1138
rect 50574 902 50810 1124
rect 43950 222 44186 458
rect 46158 222 46394 458
rect 53886 902 54122 1138
rect 91606 5662 91842 5898
rect 86822 3622 87058 3858
rect 84882 2363 85118 2599
rect 113092 4384 113328 4584
rect 113092 4348 113122 4384
rect 113122 4348 113138 4384
rect 113138 4348 113202 4384
rect 113202 4348 113218 4384
rect 113218 4348 113282 4384
rect 113282 4348 113298 4384
rect 113298 4348 113328 4384
rect 111662 1732 111898 1818
rect 111662 1668 111748 1732
rect 111748 1668 111812 1732
rect 111812 1668 111898 1732
rect 111662 1582 111898 1668
rect 58486 444 58572 458
rect 58572 444 58636 458
rect 58636 444 58722 458
rect 58486 222 58722 444
rect 141303 10368 141539 10540
rect 141303 10304 141333 10368
rect 141333 10304 141349 10368
rect 141349 10304 141413 10368
rect 141413 10304 141429 10368
rect 141429 10304 141493 10368
rect 141493 10304 141509 10368
rect 141509 10304 141539 10368
rect 141303 6334 141539 6570
rect 141303 2363 141539 2599
<< metal5 >>
rect 368 10540 169556 10582
rect 368 10304 28460 10540
rect 28696 10304 84882 10540
rect 85118 10304 141303 10540
rect 141539 10304 169556 10540
rect 368 10262 169556 10304
rect 5452 9298 50484 9340
rect 5452 9062 5494 9298
rect 5730 9062 50206 9298
rect 50442 9062 50484 9298
rect 5452 9020 50484 9062
rect 50900 9298 57476 9340
rect 50900 9062 50942 9298
rect 51178 9062 57198 9298
rect 57434 9062 57476 9298
rect 50900 9020 57476 9062
rect 368 8555 169556 8597
rect 368 8319 56671 8555
rect 56907 8319 113092 8555
rect 113328 8319 169556 8555
rect 368 8277 169556 8319
rect 12076 7258 80476 7300
rect 12076 7022 12118 7258
rect 12354 7022 80198 7258
rect 80434 7022 80476 7258
rect 12076 6980 80476 7022
rect 368 6570 169556 6612
rect 368 6334 28460 6570
rect 28696 6334 84882 6570
rect 85118 6334 141303 6570
rect 141539 6334 169556 6570
rect 368 6292 169556 6334
rect 6188 5898 61156 5940
rect 6188 5662 6230 5898
rect 6466 5662 60878 5898
rect 61114 5662 61156 5898
rect 6188 5620 61156 5662
rect 61572 5898 91884 5940
rect 61572 5662 61614 5898
rect 61850 5662 91606 5898
rect 91842 5662 91884 5898
rect 61572 5620 91884 5662
rect 368 4584 169556 4626
rect 368 4348 56671 4584
rect 56907 4348 113092 4584
rect 113328 4348 169556 4584
rect 368 4306 169556 4348
rect 6556 3858 51220 3900
rect 6556 3622 6598 3858
rect 6834 3622 50942 3858
rect 51178 3622 51220 3858
rect 6556 3580 51220 3622
rect 51636 3858 87100 3900
rect 51636 3622 51678 3858
rect 51914 3622 86822 3858
rect 87058 3622 87100 3858
rect 51636 3580 87100 3622
rect 368 2599 169556 2641
rect 368 2363 28460 2599
rect 28696 2363 84882 2599
rect 85118 2363 141303 2599
rect 141539 2363 169556 2599
rect 368 2321 169556 2363
rect 11156 1818 111940 1860
rect 11156 1582 11198 1818
rect 11434 1582 111662 1818
rect 111898 1582 111940 1818
rect 11156 1540 111940 1582
rect 35812 1138 46804 1180
rect 35812 902 35854 1138
rect 36090 902 46526 1138
rect 46762 902 46804 1138
rect 35812 860 46804 902
rect 50532 1138 54164 1180
rect 50532 902 50574 1138
rect 50810 902 53886 1138
rect 54122 902 54164 1138
rect 50532 860 54164 902
rect 38572 458 44228 500
rect 38572 222 38614 458
rect 38850 222 43950 458
rect 44186 222 44228 458
rect 38572 180 44228 222
rect 46116 458 58764 500
rect 46116 222 46158 458
rect 46394 222 58486 458
rect 58722 222 58764 458
rect 46116 180 58764 222
use sky130_fd_sc_hd__decap_3  FILLER_20_1826
timestamp 1606716760
transform 1 0 168360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606716760
transform -1 0 169556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606716760
transform -1 0 169556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1606716760
transform 1 0 168636 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1835
timestamp 1606716760
transform 1 0 169188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1830
timestamp 1606716760
transform 1 0 168728 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1818
timestamp 1606716760
transform 1 0 167624 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1606716760
transform 1 0 165876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1606716760
transform 1 0 165784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[8\]_TE
timestamp 1606716760
transform 1 0 166336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1802
timestamp 1606716760
transform 1 0 166152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1806
timestamp 1606716760
transform 1 0 166520 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1790
timestamp 1606716760
transform 1 0 165048 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[18\]
timestamp 1606716760
transform 1 0 164772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1775
timestamp 1606716760
transform 1 0 163668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1606716760
transform 1 0 163484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1771
timestamp 1606716760
transform 1 0 163300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[8\]_A
timestamp 1606716760
transform 1 0 167900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1819
timestamp 1606716760
transform 1 0 167716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1823
timestamp 1606716760
transform 1 0 168084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[8\]
timestamp 1606716760
transform 1 0 166060 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1606716760
transform 1 0 165968 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1606716760
transform 1 0 165784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1796
timestamp 1606716760
transform 1 0 165600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[26\]_A
timestamp 1606716760
transform 1 0 164680 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1784
timestamp 1606716760
transform 1 0 164496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1788
timestamp 1606716760
transform 1 0 164864 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1606716760
transform 1 0 163024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1606716760
transform 1 0 162932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1606716760
transform 1 0 161920 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1759
timestamp 1606716760
transform 1 0 162196 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1752
timestamp 1606716760
transform 1 0 161552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1606716760
transform 1 0 160172 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1606716760
transform 1 0 160080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1740
timestamp 1606716760
transform 1 0 160448 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1732
timestamp 1606716760
transform 1 0 159712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[34\]
timestamp 1606716760
transform 1 0 158332 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1720
timestamp 1606716760
transform 1 0 158608 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[26\]
timestamp 1606716760
transform 1 0 162840 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1606716760
transform 1 0 162288 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[26\]_TE
timestamp 1606716760
transform 1 0 162656 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1762
timestamp 1606716760
transform 1 0 162472 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[36\]
timestamp 1606716760
transform 1 0 161828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1758
timestamp 1606716760
transform 1 0 162104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1752
timestamp 1606716760
transform 1 0 161552 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1606716760
transform 1 0 160356 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1606716760
transform 1 0 160172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1736
timestamp 1606716760
transform 1 0 160080 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1740
timestamp 1606716760
transform 1 0 160448 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[41\]
timestamp 1606716760
transform 1 0 159252 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1723
timestamp 1606716760
transform 1 0 158884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1730
timestamp 1606716760
transform 1 0 159528 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[24\]_A
timestamp 1606716760
transform 1 0 158700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1719
timestamp 1606716760
transform 1 0 158516 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1606716760
transform 1 0 157780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1709
timestamp 1606716760
transform 1 0 157596 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1713
timestamp 1606716760
transform 1 0 157964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1606716760
transform 1 0 157320 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1606716760
transform 1 0 157228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[24\]_TE
timestamp 1606716760
transform 1 0 156860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1703
timestamp 1606716760
transform 1 0 157044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1606716760
transform 1 0 156216 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1690
timestamp 1606716760
transform 1 0 155848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1697
timestamp 1606716760
transform 1 0 156492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1606716760
transform 1 0 154468 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1606716760
transform 1 0 154376 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1671
timestamp 1606716760
transform 1 0 154100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1678
timestamp 1606716760
transform 1 0 154744 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1663
timestamp 1606716760
transform 1 0 153364 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[24\]
timestamp 1606716760
transform 1 0 156860 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1700
timestamp 1606716760
transform 1 0 156768 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A
timestamp 1606716760
transform 1 0 156216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1693
timestamp 1606716760
transform 1 0 156124 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1696
timestamp 1606716760
transform 1 0 156400 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[12\]
timestamp 1606716760
transform 1 0 155112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1685
timestamp 1606716760
transform 1 0 155388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1606716760
transform 1 0 154744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1606716760
transform 1 0 154468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1673
timestamp 1606716760
transform 1 0 154284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1677
timestamp 1606716760
transform 1 0 154652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1679
timestamp 1606716760
transform 1 0 154836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[22\]_A
timestamp 1606716760
transform 1 0 152076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1647
timestamp 1606716760
transform 1 0 151892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1651
timestamp 1606716760
transform 1 0 152260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1606716760
transform 1 0 151616 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1606716760
transform 1 0 151524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[22\]_TE
timestamp 1606716760
transform 1 0 150972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1639
timestamp 1606716760
transform 1 0 151156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1606716760
transform 1 0 150512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1628
timestamp 1606716760
transform 1 0 150144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1635
timestamp 1606716760
transform 1 0 150788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[30\]
timestamp 1606716760
transform 1 0 148764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1606716760
transform 1 0 148672 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1611
timestamp 1606716760
transform 1 0 148580 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1616
timestamp 1606716760
transform 1 0 149040 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[61\]
timestamp 1606716760
transform 1 0 152904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1661
timestamp 1606716760
transform 1 0 153180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1606716760
transform 1 0 152352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1650
timestamp 1606716760
transform 1 0 152168 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1654
timestamp 1606716760
transform 1 0 152536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[22\]
timestamp 1606716760
transform 1 0 150512 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1606716760
transform 1 0 150328 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[32\]
timestamp 1606716760
transform 1 0 149500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1618
timestamp 1606716760
transform 1 0 149224 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1624
timestamp 1606716760
transform 1 0 149776 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1606716760
transform 1 0 149132 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1610
timestamp 1606716760
transform 1 0 148488 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1616
timestamp 1606716760
transform 1 0 149040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1606716760
transform 1 0 147292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1595
timestamp 1606716760
transform 1 0 147108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1599
timestamp 1606716760
transform 1 0 147476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1606716760
transform 1 0 146832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[20\]_TE
timestamp 1606716760
transform 1 0 146464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1590
timestamp 1606716760
transform 1 0 146648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1606716760
transform 1 0 145820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1578
timestamp 1606716760
transform 1 0 145544 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1582
timestamp 1606716760
transform 1 0 145912 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[21\]
timestamp 1606716760
transform 1 0 144532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1570
timestamp 1606716760
transform 1 0 144808 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1606716760
transform 1 0 143520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[17\]_TE
timestamp 1606716760
transform 1 0 143980 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1555
timestamp 1606716760
transform 1 0 143428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1559
timestamp 1606716760
transform 1 0 143796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1563
timestamp 1606716760
transform 1 0 144164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[20\]_A
timestamp 1606716760
transform 1 0 148304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1606
timestamp 1606716760
transform 1 0 148120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[20\]
timestamp 1606716760
transform 1 0 146464 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1587
timestamp 1606716760
transform 1 0 146372 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[17\]_A
timestamp 1606716760
transform 1 0 145452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1575
timestamp 1606716760
transform 1 0 145268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1579
timestamp 1606716760
transform 1 0 145636 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[17\]
timestamp 1606716760
transform 1 0 143612 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1606716760
transform 1 0 143520 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1606716760
transform 1 0 142968 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[15\]_A
timestamp 1606716760
transform 1 0 142048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1542
timestamp 1606716760
transform 1 0 142232 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1551
timestamp 1606716760
transform 1 0 143060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1538
timestamp 1606716760
transform 1 0 141864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[15\]
timestamp 1606716760
transform 1 0 140208 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1606716760
transform 1 0 140116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1606716760
transform 1 0 138828 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1503
timestamp 1606716760
transform 1 0 138644 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1507
timestamp 1606716760
transform 1 0 139012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1606716760
transform 1 0 143336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1552
timestamp 1606716760
transform 1 0 143152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[11\]_A
timestamp 1606716760
transform 1 0 142968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1548
timestamp 1606716760
transform 1 0 142784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[11\]
timestamp 1606716760
transform 1 0 141128 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[11\]_TE
timestamp 1606716760
transform 1 0 140944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1522
timestamp 1606716760
transform 1 0 140392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[13\]_A
timestamp 1606716760
transform 1 0 139840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[15\]_TE
timestamp 1606716760
transform 1 0 140208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1514
timestamp 1606716760
transform 1 0 139656 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1518
timestamp 1606716760
transform 1 0 140024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1606716760
transform 1 0 138368 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1606716760
transform 1 0 137356 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1606716760
transform 1 0 137264 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[13\]_TE
timestamp 1606716760
transform 1 0 138000 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1492
timestamp 1606716760
transform 1 0 137632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1498
timestamp 1606716760
transform 1 0 138184 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1606716760
transform 1 0 135516 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[93\]_A
timestamp 1606716760
transform 1 0 135976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1472
timestamp 1606716760
transform 1 0 135792 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1476
timestamp 1606716760
transform 1 0 136160 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1606716760
transform 1 0 134964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1465
timestamp 1606716760
transform 1 0 135148 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1606716760
transform 1 0 134504 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1606716760
transform 1 0 134412 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[93\]_TE
timestamp 1606716760
transform 1 0 134228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1453
timestamp 1606716760
transform 1 0 134044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1461
timestamp 1606716760
transform 1 0 134780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[13\]
timestamp 1606716760
transform 1 0 138000 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1606716760
transform 1 0 137908 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1606716760
transform 1 0 137080 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1606716760
transform 1 0 137448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1488
timestamp 1606716760
transform 1 0 137264 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1492
timestamp 1606716760
transform 1 0 137632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1606716760
transform 1 0 136620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1484
timestamp 1606716760
transform 1 0 136896 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1606716760
transform 1 0 136068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1473
timestamp 1606716760
transform 1 0 135884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1477
timestamp 1606716760
transform 1 0 136252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[93\]
timestamp 1606716760
transform 1 0 134228 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1454
timestamp 1606716760
transform 1 0 134136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1445
timestamp 1606716760
transform 1 0 133308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[91\]
timestamp 1606716760
transform 1 0 131652 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1606716760
transform 1 0 131560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1414
timestamp 1606716760
transform 1 0 130456 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[43\]_A
timestamp 1606716760
transform 1 0 130272 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1410
timestamp 1606716760
transform 1 0 130088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1606716760
transform 1 0 128800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1606716760
transform 1 0 129812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1606716760
transform 1 0 128708 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1606716760
transform 1 0 129260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1399
timestamp 1606716760
transform 1 0 129076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1403
timestamp 1606716760
transform 1 0 129444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1606716760
transform 1 0 132388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1606716760
transform 1 0 132296 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1606716760
transform 1 0 132848 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[91\]_A
timestamp 1606716760
transform 1 0 133216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1438
timestamp 1606716760
transform 1 0 132664 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1442
timestamp 1606716760
transform 1 0 133032 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1446
timestamp 1606716760
transform 1 0 133400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[91\]_TE
timestamp 1606716760
transform 1 0 131836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1431
timestamp 1606716760
transform 1 0 132020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1606716760
transform 1 0 131008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1606716760
transform 1 0 130456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1606716760
transform 1 0 131468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1416
timestamp 1606716760
transform 1 0 130640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1423
timestamp 1606716760
transform 1 0 131284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1427
timestamp 1606716760
transform 1 0 131652 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1412
timestamp 1606716760
transform 1 0 130272 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1387
timestamp 1606716760
transform 1 0 127972 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[8\]
timestamp 1606716760
transform 1 0 126316 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1606716760
transform 1 0 125856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1365
timestamp 1606716760
transform 1 0 125948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1606716760
transform 1 0 124108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[80\]_TE
timestamp 1606716760
transform 1 0 124568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1348
timestamp 1606716760
transform 1 0 124384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1352
timestamp 1606716760
transform 1 0 124752 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[43\]
timestamp 1606716760
transform 1 0 128616 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1606716760
transform 1 0 127236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[8\]_A
timestamp 1606716760
transform 1 0 127604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[43\]_TE
timestamp 1606716760
transform 1 0 128432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1381
timestamp 1606716760
transform 1 0 127420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1385
timestamp 1606716760
transform 1 0 127788 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1391
timestamp 1606716760
transform 1 0 128340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1377
timestamp 1606716760
transform 1 0 127052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1606716760
transform 1 0 126776 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1606716760
transform 1 0 126684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[80\]_A
timestamp 1606716760
transform 1 0 126132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[8\]_TE
timestamp 1606716760
transform 1 0 126500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1365
timestamp 1606716760
transform 1 0 125948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1369
timestamp 1606716760
transform 1 0 126316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[80\]
timestamp 1606716760
transform 1 0 124292 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1606716760
transform 1 0 124108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1343
timestamp 1606716760
transform 1 0 123924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1606716760
transform 1 0 123740 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1606716760
transform 1 0 123096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1606716760
transform 1 0 123004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1337
timestamp 1606716760
transform 1 0 123372 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1321
timestamp 1606716760
transform 1 0 121900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[88\]
timestamp 1606716760
transform 1 0 120244 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1606716760
transform 1 0 120152 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1300
timestamp 1606716760
transform 1 0 119968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1288
timestamp 1606716760
transform 1 0 118864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1606716760
transform 1 0 123280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1606716760
transform 1 0 123096 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1327
timestamp 1606716760
transform 1 0 122452 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1333
timestamp 1606716760
transform 1 0 123004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1339
timestamp 1606716760
transform 1 0 123556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[238\]
timestamp 1606716760
transform 1 0 122176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1606716760
transform 1 0 121164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1606716760
transform 1 0 121072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1606716760
transform 1 0 121624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[88\]_A
timestamp 1606716760
transform 1 0 121992 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1311
timestamp 1606716760
transform 1 0 120980 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1316
timestamp 1606716760
transform 1 0 121440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1320
timestamp 1606716760
transform 1 0 121808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1305
timestamp 1606716760
transform 1 0 120428 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[86\]_A
timestamp 1606716760
transform 1 0 119784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[88\]_TE
timestamp 1606716760
transform 1 0 120244 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1296
timestamp 1606716760
transform 1 0 119600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1300
timestamp 1606716760
transform 1 0 119968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _659_
timestamp 1606716760
transform 1 0 118220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__A
timestamp 1606716760
transform 1 0 118680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[86\]_TE
timestamp 1606716760
transform 1 0 117944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1272
timestamp 1606716760
transform 1 0 117392 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1280
timestamp 1606716760
transform 1 0 118128 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1284
timestamp 1606716760
transform 1 0 118496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1606716760
transform 1 0 117300 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[75\]_A
timestamp 1606716760
transform 1 0 116380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1259
timestamp 1606716760
transform 1 0 116196 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1263
timestamp 1606716760
transform 1 0 116564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[75\]
timestamp 1606716760
transform 1 0 114540 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1606716760
transform 1 0 114448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[86\]
timestamp 1606716760
transform 1 0 117944 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[6\]_A
timestamp 1606716760
transform 1 0 117392 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1274
timestamp 1606716760
transform 1 0 117576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1270
timestamp 1606716760
transform 1 0 117208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1606716760
transform 1 0 114448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[6\]
timestamp 1606716760
transform 1 0 115552 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1606716760
transform 1 0 115460 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__652__A
timestamp 1606716760
transform 1 0 114908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[6\]_TE
timestamp 1606716760
transform 1 0 115276 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[75\]_TE
timestamp 1606716760
transform 1 0 114264 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1243
timestamp 1606716760
transform 1 0 114724 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1247
timestamp 1606716760
transform 1 0 115092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1237
timestamp 1606716760
transform 1 0 114172 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1228
timestamp 1606716760
transform 1 0 113344 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[71\]
timestamp 1606716760
transform 1 0 111688 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1606716760
transform 1 0 111596 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[66\]_TE
timestamp 1606716760
transform 1 0 111228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1204
timestamp 1606716760
transform 1 0 111136 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1207
timestamp 1606716760
transform 1 0 111412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1198
timestamp 1606716760
transform 1 0 110584 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[64\]
timestamp 1606716760
transform 1 0 108928 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[66\]_A
timestamp 1606716760
transform 1 0 113068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[71\]_A
timestamp 1606716760
transform 1 0 113436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1223
timestamp 1606716760
transform 1 0 112884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1227
timestamp 1606716760
transform 1 0 113252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1231
timestamp 1606716760
transform 1 0 113620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[66\]
timestamp 1606716760
transform 1 0 111228 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1202
timestamp 1606716760
transform 1 0 110952 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[64\]_A
timestamp 1606716760
transform 1 0 110768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _658_
timestamp 1606716760
transform 1 0 109940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1606716760
transform 1 0 109848 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__658__A
timestamp 1606716760
transform 1 0 110400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1194
timestamp 1606716760
transform 1 0 110216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1198
timestamp 1606716760
transform 1 0 110584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[64\]_TE
timestamp 1606716760
transform 1 0 108928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1182
timestamp 1606716760
transform 1 0 109112 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _656_
timestamp 1606716760
transform 1 0 107732 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1606716760
transform 1 0 108744 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[62\]_A
timestamp 1606716760
transform 1 0 108192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1170
timestamp 1606716760
transform 1 0 108008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1174
timestamp 1606716760
transform 1 0 108376 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1179
timestamp 1606716760
transform 1 0 108836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1166
timestamp 1606716760
transform 1 0 107640 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _654_
timestamp 1606716760
transform 1 0 106628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[62\]_TE
timestamp 1606716760
transform 1 0 107088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1154
timestamp 1606716760
transform 1 0 106536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1158
timestamp 1606716760
transform 1 0 106904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1162
timestamp 1606716760
transform 1 0 107272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1606716760
transform 1 0 105892 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1148
timestamp 1606716760
transform 1 0 105984 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1135
timestamp 1606716760
transform 1 0 104788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__656__A
timestamp 1606716760
transform 1 0 108468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1173
timestamp 1606716760
transform 1 0 108284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1177
timestamp 1606716760
transform 1 0 108652 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[62\]
timestamp 1606716760
transform 1 0 106628 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__654__A
timestamp 1606716760
transform 1 0 106444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1147
timestamp 1606716760
transform 1 0 105892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[264\]
timestamp 1606716760
transform 1 0 105616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__650__A
timestamp 1606716760
transform 1 0 104788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[55\]_A
timestamp 1606716760
transform 1 0 105156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1137
timestamp 1606716760
transform 1 0 104972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1141
timestamp 1606716760
transform 1 0 105340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _650_
timestamp 1606716760
transform 1 0 104328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1606716760
transform 1 0 104236 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[55\]_TE
timestamp 1606716760
transform 1 0 104052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1133
timestamp 1606716760
transform 1 0 104604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[55\]
timestamp 1606716760
transform 1 0 103132 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1606716760
transform 1 0 103040 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[253\]
timestamp 1606716760
transform 1 0 102028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[51\]_TE
timestamp 1606716760
transform 1 0 101844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1097
timestamp 1606716760
transform 1 0 101292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1108
timestamp 1606716760
transform 1 0 102304 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[257\]
timestamp 1606716760
transform 1 0 101016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1606716760
transform 1 0 100188 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1086
timestamp 1606716760
transform 1 0 100280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[262\]
timestamp 1606716760
transform 1 0 99176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[60\]_TE
timestamp 1606716760
transform 1 0 99636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1077
timestamp 1606716760
transform 1 0 99452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1081
timestamp 1606716760
transform 1 0 99820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[51\]_A
timestamp 1606716760
transform 1 0 103684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1121
timestamp 1606716760
transform 1 0 103500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1125
timestamp 1606716760
transform 1 0 103868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[51\]
timestamp 1606716760
transform 1 0 101844 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[60\]_A
timestamp 1606716760
transform 1 0 101292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1099
timestamp 1606716760
transform 1 0 101476 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1095
timestamp 1606716760
transform 1 0 101108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[60\]
timestamp 1606716760
transform 1 0 99452 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _603_
timestamp 1606716760
transform 1 0 98164 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1066
timestamp 1606716760
transform 1 0 98440 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1606716760
transform 1 0 97336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__647__A
timestamp 1606716760
transform 1 0 96784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1046
timestamp 1606716760
transform 1 0 96600 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1050
timestamp 1606716760
transform 1 0 96968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1055
timestamp 1606716760
transform 1 0 97428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _647_
timestamp 1606716760
transform 1 0 96324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1042
timestamp 1606716760
transform 1 0 96232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[48\]_TE
timestamp 1606716760
transform 1 0 95496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1033
timestamp 1606716760
transform 1 0 95404 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1036
timestamp 1606716760
transform 1 0 95680 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[322\]
timestamp 1606716760
transform 1 0 94576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1606716760
transform 1 0 94484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1027
timestamp 1606716760
transform 1 0 94852 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1606716760
transform 1 0 98624 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__A
timestamp 1606716760
transform 1 0 98164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_1065
timestamp 1606716760
transform 1 0 98348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1069
timestamp 1606716760
transform 1 0 98716 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1062
timestamp 1606716760
transform 1 0 98072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[48\]_A
timestamp 1606716760
transform 1 0 97336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1052
timestamp 1606716760
transform 1 0 97152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1056
timestamp 1606716760
transform 1 0 97520 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[48\]
timestamp 1606716760
transform 1 0 95496 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1030
timestamp 1606716760
transform 1 0 95128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[120\]_A
timestamp 1606716760
transform 1 0 94944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1026
timestamp 1606716760
transform 1 0 94760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[120\]_TE
timestamp 1606716760
transform 1 0 93564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1011
timestamp 1606716760
transform 1 0 93380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1015
timestamp 1606716760
transform 1 0 93748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[11\]
timestamp 1606716760
transform 1 0 91724 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1606716760
transform 1 0 91632 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_984
timestamp 1606716760
transform 1 0 90896 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[321\]
timestamp 1606716760
transform 1 0 90620 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_980
timestamp 1606716760
transform 1 0 90528 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_974
timestamp 1606716760
transform 1 0 89976 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[120\]
timestamp 1606716760
transform 1 0 93104 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1606716760
transform 1 0 93012 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[11\]_A
timestamp 1606716760
transform 1 0 92828 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[318\]
timestamp 1606716760
transform 1 0 92000 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[11\]_TE
timestamp 1606716760
transform 1 0 91724 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_995
timestamp 1606716760
transform 1 0 91908 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_999
timestamp 1606716760
transform 1 0 92276 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[320\]
timestamp 1606716760
transform 1 0 90344 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_981
timestamp 1606716760
transform 1 0 90620 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_974
timestamp 1606716760
transform 1 0 89976 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1606716760
transform 1 0 88780 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_962
timestamp 1606716760
transform 1 0 88872 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_958
timestamp 1606716760
transform 1 0 88504 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_962
timestamp 1606716760
transform 1 0 88872 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _479_
timestamp 1606716760
transform 1 0 87124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[305\]
timestamp 1606716760
transform 1 0 87492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1606716760
transform 1 0 87400 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__A
timestamp 1606716760
transform 1 0 87124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_941
timestamp 1606716760
transform 1 0 86940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_945
timestamp 1606716760
transform 1 0 87308 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_950
timestamp 1606716760
transform 1 0 87768 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_942
timestamp 1606716760
transform 1 0 87032 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_946
timestamp 1606716760
transform 1 0 87400 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[82\]
timestamp 1606716760
transform 1 0 86020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1606716760
transform 1 0 85928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_926
timestamp 1606716760
transform 1 0 85560 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_934
timestamp 1606716760
transform 1 0 86296 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[202\]
timestamp 1606716760
transform 1 0 85928 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_926
timestamp 1606716760
transform 1 0 85560 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_933
timestamp 1606716760
transform 1 0 86204 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_914
timestamp 1606716760
transform 1 0 84456 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _559_
timestamp 1606716760
transform 1 0 84916 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A
timestamp 1606716760
transform 1 0 84364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A
timestamp 1606716760
transform 1 0 84732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__A
timestamp 1606716760
transform 1 0 85376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_915
timestamp 1606716760
transform 1 0 84548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_922
timestamp 1606716760
transform 1 0 85192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _546_
timestamp 1606716760
transform 1 0 83168 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _557_
timestamp 1606716760
transform 1 0 84180 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_903
timestamp 1606716760
transform 1 0 83444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1606716760
transform 1 0 83076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_897
timestamp 1606716760
transform 1 0 82892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_889
timestamp 1606716760
transform 1 0 82156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[86\]
timestamp 1606716760
transform 1 0 80500 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1606716760
transform 1 0 80224 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[84\]_TE
timestamp 1606716760
transform 1 0 79396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[86\]_TE
timestamp 1606716760
transform 1 0 80040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_861
timestamp 1606716760
transform 1 0 79580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_865
timestamp 1606716760
transform 1 0 79948 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_869
timestamp 1606716760
transform 1 0 80316 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _555_
timestamp 1606716760
transform 1 0 83904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1606716760
transform 1 0 83352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1606716760
transform 1 0 83720 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_900
timestamp 1606716760
transform 1 0 83168 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_904
timestamp 1606716760
transform 1 0 83536 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_911
timestamp 1606716760
transform 1 0 84180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _548_
timestamp 1606716760
transform 1 0 82892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__A
timestamp 1606716760
transform 1 0 82340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_889
timestamp 1606716760
transform 1 0 82156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_893
timestamp 1606716760
transform 1 0 82524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _542_
timestamp 1606716760
transform 1 0 81880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1606716760
transform 1 0 81788 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[84\]_A
timestamp 1606716760
transform 1 0 81236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[86\]_A
timestamp 1606716760
transform 1 0 81604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_877
timestamp 1606716760
transform 1 0 81052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_881
timestamp 1606716760
transform 1 0 81420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[84\]
timestamp 1606716760
transform 1 0 79396 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_20_857
timestamp 1606716760
transform 1 0 79212 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _477_
timestamp 1606716760
transform 1 0 78936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_853
timestamp 1606716760
transform 1 0 78844 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _526_
timestamp 1606716760
transform 1 0 77464 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1606716760
transform 1 0 77372 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_835
timestamp 1606716760
transform 1 0 77188 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_841
timestamp 1606716760
transform 1 0 77740 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[97\]_B
timestamp 1606716760
transform 1 0 77004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_831
timestamp 1606716760
transform 1 0 76820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _524_
timestamp 1606716760
transform 1 0 76176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1606716760
transform 1 0 76636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_827
timestamp 1606716760
transform 1 0 76452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[93\]
timestamp 1606716760
transform 1 0 74612 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1606716760
transform 1 0 74520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_816
timestamp 1606716760
transform 1 0 75440 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_856
timestamp 1606716760
transform 1 0 79120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__A
timestamp 1606716760
transform 1 0 78936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__A
timestamp 1606716760
transform 1 0 78292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_845
timestamp 1606716760
transform 1 0 78108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_849
timestamp 1606716760
transform 1 0 78476 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_853
timestamp 1606716760
transform 1 0 78844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _528_
timestamp 1606716760
transform 1 0 77832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[97\]_A
timestamp 1606716760
transform 1 0 77280 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A
timestamp 1606716760
transform 1 0 77648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_838
timestamp 1606716760
transform 1 0 77464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_834
timestamp 1606716760
transform 1 0 77096 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[97\]
timestamp 1606716760
transform 1 0 76268 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1606716760
transform 1 0 76176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_821
timestamp 1606716760
transform 1 0 75900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__A
timestamp 1606716760
transform 1 0 75716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1606716760
transform 1 0 74888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[93\]_A
timestamp 1606716760
transform 1 0 75348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[93\]_B
timestamp 1606716760
transform 1 0 74704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_806
timestamp 1606716760
transform 1 0 74520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_813
timestamp 1606716760
transform 1 0 75164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_817
timestamp 1606716760
transform 1 0 75532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _519_
timestamp 1606716760
transform 1 0 73324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__A
timestamp 1606716760
transform 1 0 73784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_789
timestamp 1606716760
transform 1 0 72956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_796
timestamp 1606716760
transform 1 0 73600 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_800
timestamp 1606716760
transform 1 0 73968 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[71\]_TE
timestamp 1606716760
transform 1 0 72772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_785
timestamp 1606716760
transform 1 0 72588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[88\]
timestamp 1606716760
transform 1 0 71760 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1606716760
transform 1 0 71668 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[147\]
timestamp 1606716760
transform 1 0 70472 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[84\]_B
timestamp 1606716760
transform 1 0 70932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_765
timestamp 1606716760
transform 1 0 70748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_769
timestamp 1606716760
transform 1 0 71116 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[80\]_B
timestamp 1606716760
transform 1 0 69920 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_754
timestamp 1606716760
transform 1 0 69736 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_758
timestamp 1606716760
transform 1 0 70104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[71\]_A
timestamp 1606716760
transform 1 0 74336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_802
timestamp 1606716760
transform 1 0 74152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[71\]
timestamp 1606716760
transform 1 0 72496 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[88\]_A
timestamp 1606716760
transform 1 0 72312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_781
timestamp 1606716760
transform 1 0 72220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[84\]_A
timestamp 1606716760
transform 1 0 71668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_773
timestamp 1606716760
transform 1 0 71484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_777
timestamp 1606716760
transform 1 0 71852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[84\]
timestamp 1606716760
transform 1 0 70656 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1606716760
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[79\]_A
timestamp 1606716760
transform 1 0 69644 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[80\]_A
timestamp 1606716760
transform 1 0 70012 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_751
timestamp 1606716760
transform 1 0 69460 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_755
timestamp 1606716760
transform 1 0 69828 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_759
timestamp 1606716760
transform 1 0 70196 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[79\]
timestamp 1606716760
transform 1 0 68632 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[80\]
timestamp 1606716760
transform 1 0 68908 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1606716760
transform 1 0 68816 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[79\]_B
timestamp 1606716760
transform 1 0 68448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_736
timestamp 1606716760
transform 1 0 68080 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[410\]
timestamp 1606716760
transform 1 0 67620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[412\]
timestamp 1606716760
transform 1 0 67804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_734
timestamp 1606716760
transform 1 0 67896 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_732
timestamp 1606716760
transform 1 0 67712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_729
timestamp 1606716760
transform 1 0 67436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_726
timestamp 1606716760
transform 1 0 67160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_717
timestamp 1606716760
transform 1 0 66332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[407\]
timestamp 1606716760
transform 1 0 66056 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1606716760
transform 1 0 65964 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_710
timestamp 1606716760
transform 1 0 65688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_714
timestamp 1606716760
transform 1 0 66056 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[77\]_A
timestamp 1606716760
transform 1 0 65504 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_706
timestamp 1606716760
transform 1 0 65320 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_705
timestamp 1606716760
transform 1 0 65228 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[167\]
timestamp 1606716760
transform 1 0 65044 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1606716760
transform 1 0 64952 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[77\]_B
timestamp 1606716760
transform 1 0 64584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_700
timestamp 1606716760
transform 1 0 64768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[77\]
timestamp 1606716760
transform 1 0 64400 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_694
timestamp 1606716760
transform 1 0 64216 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[394\]
timestamp 1606716760
transform 1 0 63572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[401\]
timestamp 1606716760
transform 1 0 63204 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1606716760
transform 1 0 63112 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_690
timestamp 1606716760
transform 1 0 63848 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_686
timestamp 1606716760
transform 1 0 63480 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_679
timestamp 1606716760
transform 1 0 62836 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[387\]
timestamp 1606716760
transform 1 0 62560 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[73\]_A
timestamp 1606716760
transform 1 0 62008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[75\]_A
timestamp 1606716760
transform 1 0 62376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_672
timestamp 1606716760
transform 1 0 62192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_670
timestamp 1606716760
transform 1 0 62008 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_668
timestamp 1606716760
transform 1 0 61824 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[73\]
timestamp 1606716760
transform 1 0 60996 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[75\]
timestamp 1606716760
transform 1 0 61180 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[73\]_B
timestamp 1606716760
transform 1 0 60812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_660
timestamp 1606716760
transform 1 0 61088 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[59\]_A
timestamp 1606716760
transform 1 0 60444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_655
timestamp 1606716760
transform 1 0 60628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_652
timestamp 1606716760
transform 1 0 60352 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1606716760
transform 1 0 60260 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[59\]_B
timestamp 1606716760
transform 1 0 59616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_651
timestamp 1606716760
transform 1 0 60260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_646
timestamp 1606716760
transform 1 0 59800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_650
timestamp 1606716760
transform 1 0 60168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[59\]
timestamp 1606716760
transform 1 0 59432 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1606716760
transform 1 0 59340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_640
timestamp 1606716760
transform 1 0 59248 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_641
timestamp 1606716760
transform 1 0 59340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[366\]
timestamp 1606716760
transform 1 0 59064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[57\]_A
timestamp 1606716760
transform 1 0 58512 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_630
timestamp 1606716760
transform 1 0 58328 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_634
timestamp 1606716760
transform 1 0 58696 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_630
timestamp 1606716760
transform 1 0 58328 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[363\]
timestamp 1606716760
transform 1 0 58052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[57\]_B
timestamp 1606716760
transform 1 0 57868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[57\]
timestamp 1606716760
transform 1 0 57500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1606716760
transform 1 0 57408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[36\]_A
timestamp 1606716760
transform 1 0 57500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_623
timestamp 1606716760
transform 1 0 57684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[36\]_B
timestamp 1606716760
transform 1 0 56856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_619
timestamp 1606716760
transform 1 0 57316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_616
timestamp 1606716760
transform 1 0 57040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[36\]
timestamp 1606716760
transform 1 0 56488 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_612
timestamp 1606716760
transform 1 0 56672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[60\]_A
timestamp 1606716760
transform 1 0 56304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[62\]_A
timestamp 1606716760
transform 1 0 55936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_606
timestamp 1606716760
transform 1 0 56120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[60\]
timestamp 1606716760
transform 1 0 55844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_602
timestamp 1606716760
transform 1 0 55752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[62\]_B
timestamp 1606716760
transform 1 0 55292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_595
timestamp 1606716760
transform 1 0 55108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_599
timestamp 1606716760
transform 1 0 55476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[362\]
timestamp 1606716760
transform 1 0 54832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[62\]
timestamp 1606716760
transform 1 0 54924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_590
timestamp 1606716760
transform 1 0 54648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1606716760
transform 1 0 54556 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[66\]_A
timestamp 1606716760
transform 1 0 54372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_589
timestamp 1606716760
transform 1 0 54556 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_585
timestamp 1606716760
transform 1 0 54188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[336\]
timestamp 1606716760
transform 1 0 53912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1606716760
transform 1 0 53728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[66\]_B
timestamp 1606716760
transform 1 0 53544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_576
timestamp 1606716760
transform 1 0 53360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_581
timestamp 1606716760
transform 1 0 53820 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_581
timestamp 1606716760
transform 1 0 53820 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[66\]
timestamp 1606716760
transform 1 0 52992 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_567
timestamp 1606716760
transform 1 0 52532 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_571
timestamp 1606716760
transform 1 0 52900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[68\]_A
timestamp 1606716760
transform 1 0 53176 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_572
timestamp 1606716760
transform 1 0 52992 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[68\]_B
timestamp 1606716760
transform 1 0 52348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_562
timestamp 1606716760
transform 1 0 52072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[358\]
timestamp 1606716760
transform 1 0 51796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1606716760
transform 1 0 51704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_556
timestamp 1606716760
transform 1 0 51520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[68\]
timestamp 1606716760
transform 1 0 52164 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_562
timestamp 1606716760
transform 1 0 52072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[95\]_A
timestamp 1606716760
transform 1 0 51520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_558
timestamp 1606716760
transform 1 0 51704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_548
timestamp 1606716760
transform 1 0 50784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_554
timestamp 1606716760
transform 1 0 51336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[169\]
timestamp 1606716760
transform 1 0 50508 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_541
timestamp 1606716760
transform 1 0 50140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[95\]_TE
timestamp 1606716760
transform 1 0 49956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_537
timestamp 1606716760
transform 1 0 49772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[55\]
timestamp 1606716760
transform 1 0 48944 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1606716760
transform 1 0 48852 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1606716760
transform 1 0 48668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[385\]
timestamp 1606716760
transform 1 0 47656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_517
timestamp 1606716760
transform 1 0 47932 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_506
timestamp 1606716760
transform 1 0 46920 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[99\]
timestamp 1606716760
transform 1 0 46092 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1606716760
transform 1 0 46000 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[51\]_B
timestamp 1606716760
transform 1 0 45816 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_490
timestamp 1606716760
transform 1 0 45448 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[95\]
timestamp 1606716760
transform 1 0 49680 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[55\]_A
timestamp 1606716760
transform 1 0 49496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[55\]_B
timestamp 1606716760
transform 1 0 49128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_523
timestamp 1606716760
transform 1 0 48484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_529
timestamp 1606716760
transform 1 0 49036 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_532
timestamp 1606716760
transform 1 0 49312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[140\]
timestamp 1606716760
transform 1 0 48208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1606716760
transform 1 0 48116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_509
timestamp 1606716760
transform 1 0 47196 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_517
timestamp 1606716760
transform 1 0 47932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[51\]_A
timestamp 1606716760
transform 1 0 46644 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[99\]_A
timestamp 1606716760
transform 1 0 47012 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_505
timestamp 1606716760
transform 1 0 46828 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_501
timestamp 1606716760
transform 1 0 46460 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[51\]
timestamp 1606716760
transform 1 0 45632 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_484
timestamp 1606716760
transform 1 0 44896 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[383\]
timestamp 1606716760
transform 1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[97\]_A
timestamp 1606716760
transform 1 0 43608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_472
timestamp 1606716760
transform 1 0 43792 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_480
timestamp 1606716760
transform 1 0 44528 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_478
timestamp 1606716760
transform 1 0 44344 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_468
timestamp 1606716760
transform 1 0 43424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[97\]
timestamp 1606716760
transform 1 0 42596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1606716760
transform 1 0 42504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1606716760
transform 1 0 43148 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_463
timestamp 1606716760
transform 1 0 42964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_466
timestamp 1606716760
transform 1 0 43240 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_455
timestamp 1606716760
transform 1 0 42228 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[149\]
timestamp 1606716760
transform 1 0 41952 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[91\]_A
timestamp 1606716760
transform 1 0 41952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_450
timestamp 1606716760
transform 1 0 41768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_454
timestamp 1606716760
transform 1 0 42136 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_444
timestamp 1606716760
transform 1 0 41216 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[88\]
timestamp 1606716760
transform 1 0 40388 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[91\]
timestamp 1606716760
transform 1 0 40940 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1606716760
transform 1 0 40296 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[86\]_A
timestamp 1606716760
transform 1 0 40388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[88\]_A
timestamp 1606716760
transform 1 0 40756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_433
timestamp 1606716760
transform 1 0 40204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_437
timestamp 1606716760
transform 1 0 40572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_433
timestamp 1606716760
transform 1 0 40204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_429
timestamp 1606716760
transform 1 0 39836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[82\]_A
timestamp 1606716760
transform 1 0 38548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_417
timestamp 1606716760
transform 1 0 38732 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[82\]
timestamp 1606716760
transform 1 0 37536 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1606716760
transform 1 0 37444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_413
timestamp 1606716760
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[80\]_TE
timestamp 1606716760
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_397
timestamp 1606716760
transform 1 0 36892 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_400
timestamp 1606716760
transform 1 0 37168 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[154\]
timestamp 1606716760
transform 1 0 36248 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_386
timestamp 1606716760
transform 1 0 35880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_393
timestamp 1606716760
transform 1 0 36524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[79\]_A
timestamp 1606716760
transform 1 0 35696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_382
timestamp 1606716760
transform 1 0 35512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[86\]
timestamp 1606716760
transform 1 0 39376 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[80\]_A
timestamp 1606716760
transform 1 0 38824 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_420
timestamp 1606716760
transform 1 0 39008 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_416
timestamp 1606716760
transform 1 0 38640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[80\]
timestamp 1606716760
transform 1 0 36984 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1606716760
transform 1 0 36892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[99\]_A
timestamp 1606716760
transform 1 0 36340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_389
timestamp 1606716760
transform 1 0 36156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1606716760
transform 1 0 36524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[79\]
timestamp 1606716760
transform 1 0 34684 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1606716760
transform 1 0 34592 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_371
timestamp 1606716760
transform 1 0 34500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_363
timestamp 1606716760
transform 1 0 33764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[71\]
timestamp 1606716760
transform 1 0 31832 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1606716760
transform 1 0 31740 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_351
timestamp 1606716760
transform 1 0 32660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_340
timestamp 1606716760
transform 1 0 31648 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_332
timestamp 1606716760
transform 1 0 30912 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[99\]
timestamp 1606716760
transform 1 0 34500 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[99\]_TE
timestamp 1606716760
transform 1 0 34316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_367
timestamp 1606716760
transform 1 0 34132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[77\]_A
timestamp 1606716760
transform 1 0 33948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_363
timestamp 1606716760
transform 1 0 33764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[77\]
timestamp 1606716760
transform 1 0 32936 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[71\]_A
timestamp 1606716760
transform 1 0 32384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_346
timestamp 1606716760
transform 1 0 32200 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_350
timestamp 1606716760
transform 1 0 32568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[73\]
timestamp 1606716760
transform 1 0 31372 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1606716760
transform 1 0 31280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[68\]_A
timestamp 1606716760
transform 1 0 30636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[73\]_A
timestamp 1606716760
transform 1 0 31096 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_327
timestamp 1606716760
transform 1 0 30452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_331
timestamp 1606716760
transform 1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_320
timestamp 1606716760
transform 1 0 29808 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[66\]
timestamp 1606716760
transform 1 0 28980 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1606716760
transform 1 0 28888 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_308
timestamp 1606716760
transform 1 0 28704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1606716760
transform 1 0 27968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[448\]
timestamp 1606716760
transform 1 0 27692 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[77\]_TE
timestamp 1606716760
transform 1 0 27232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_289
timestamp 1606716760
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_294
timestamp 1606716760
transform 1 0 27416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[57\]
timestamp 1606716760
transform 1 0 26128 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1606716760
transform 1 0 26036 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_271
timestamp 1606716760
transform 1 0 25300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[68\]
timestamp 1606716760
transform 1 0 29624 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[66\]_A
timestamp 1606716760
transform 1 0 29440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_314
timestamp 1606716760
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[77\]_A
timestamp 1606716760
transform 1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_310
timestamp 1606716760
transform 1 0 28888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[77\]
timestamp 1606716760
transform 1 0 27232 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[57\]_A
timestamp 1606716760
transform 1 0 26496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_283
timestamp 1606716760
transform 1 0 26404 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_286
timestamp 1606716760
transform 1 0 26680 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[341\]
timestamp 1606716760
transform 1 0 25760 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1606716760
transform 1 0 25668 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_279
timestamp 1606716760
transform 1 0 26036 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1606716760
transform 1 0 24196 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[53\]
timestamp 1606716760
transform 1 0 23368 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1606716760
transform 1 0 23184 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_249
timestamp 1606716760
transform 1 0 23276 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_240
timestamp 1606716760
transform 1 0 22448 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[68\]
timestamp 1606716760
transform 1 0 20792 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1606716760
transform 1 0 20332 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[60\]_TE
timestamp 1606716760
transform 1 0 20148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1606716760
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[446\]
timestamp 1606716760
transform 1 0 24656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[53\]_A
timestamp 1606716760
transform 1 0 24472 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_267
timestamp 1606716760
transform 1 0 24932 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[51\]_A
timestamp 1606716760
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_256
timestamp 1606716760
transform 1 0 23920 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_260
timestamp 1606716760
transform 1 0 24288 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[51\]
timestamp 1606716760
transform 1 0 23092 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[60\]_A
timestamp 1606716760
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[68\]_A
timestamp 1606716760
transform 1 0 22356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_237
timestamp 1606716760
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_241
timestamp 1606716760
transform 1 0 22540 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_233
timestamp 1606716760
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[60\]
timestamp 1606716760
transform 1 0 20148 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_20_214
timestamp 1606716760
transform 1 0 20056 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1606716760
transform 1 0 20056 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[68\]_TE
timestamp 1606716760
transform 1 0 19872 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[133\]
timestamp 1606716760
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[136\]
timestamp 1606716760
transform 1 0 19228 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_204
timestamp 1606716760
transform 1 0 19136 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1606716760
transform 1 0 19504 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_200
timestamp 1606716760
transform 1 0 18768 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_188
timestamp 1606716760
transform 1 0 17664 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_199
timestamp 1606716760
transform 1 0 18676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1606716760
transform 1 0 17480 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_187
timestamp 1606716760
transform 1 0 17572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[64\]_A
timestamp 1606716760
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_176
timestamp 1606716760
transform 1 0 16560 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_180
timestamp 1606716760
transform 1 0 16928 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1606716760
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1606716760
transform 1 0 15824 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1606716760
transform 1 0 14628 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_149
timestamp 1606716760
transform 1 0 14076 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1606716760
transform 1 0 14720 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_137
timestamp 1606716760
transform 1 0 12972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1606716760
transform 1 0 11776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_125
timestamp 1606716760
transform 1 0 11868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_113
timestamp 1606716760
transform 1 0 10764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_121
timestamp 1606716760
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[64\]
timestamp 1606716760
transform 1 0 14536 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1606716760
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[64\]_TE
timestamp 1606716760
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_145
timestamp 1606716760
transform 1 0 13708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[138\]
timestamp 1606716760
transform 1 0 13432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_129
timestamp 1606716760
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_141
timestamp 1606716760
transform 1 0 13340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[129\]
timestamp 1606716760
transform 1 0 11960 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_125
timestamp 1606716760
transform 1 0 11868 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[4\]_A
timestamp 1606716760
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1606716760
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 1606716760
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1606716760
transform 1 0 8924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[4\]_TE
timestamp 1606716760
transform 1 0 9476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1606716760
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_98
timestamp 1606716760
transform 1 0 9384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_101
timestamp 1606716760
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_81
timestamp 1606716760
transform 1 0 7820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[53\]
timestamp 1606716760
transform 1 0 6164 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1606716760
transform 1 0 6072 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[51\]_TE
timestamp 1606716760
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1606716760
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[4\]
timestamp 1606716760
transform 1 0 9476 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1606716760
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_93
timestamp 1606716760
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[51\]_A
timestamp 1606716760
transform 1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[53\]_A
timestamp 1606716760
transform 1 0 7912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_76
timestamp 1606716760
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1606716760
transform 1 0 7728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_84
timestamp 1606716760
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[51\]
timestamp 1606716760
transform 1 0 5704 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_20_52
timestamp 1606716760
transform 1 0 5152 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[48\]
timestamp 1606716760
transform 1 0 4324 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[48\]_A
timestamp 1606716760
transform 1 0 4784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[4\]_A
timestamp 1606716760
transform 1 0 4140 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_46
timestamp 1606716760
transform 1 0 4600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_50
timestamp 1606716760
transform 1 0 4968 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[127\]
timestamp 1606716760
transform 1 0 3312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[4\]
timestamp 1606716760
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1606716760
transform 1 0 3220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1606716760
transform 1 0 3220 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_32
timestamp 1606716760
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_36
timestamp 1606716760
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606716760
transform 1 0 2852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_35
timestamp 1606716760
transform 1 0 3588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[378\]
timestamp 1606716760
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1606716760
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_19
timestamp 1606716760
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_23
timestamp 1606716760
transform 1 0 2484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606716760
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606716760
transform 1 0 368 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606716760
transform 1 0 368 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606716760
transform 1 0 644 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606716760
transform 1 0 644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606716760
transform -1 0 169556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606716760
transform -1 0 169556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1606716760
transform 1 0 168728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1831
timestamp 1606716760
transform 1 0 168820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1835
timestamp 1606716760
transform 1 0 169188 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1826
timestamp 1606716760
transform 1 0 168360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1824
timestamp 1606716760
transform 1 0 168176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606716760
transform -1 0 169556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606716760
transform -1 0 169556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1606716760
transform 1 0 168728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1831
timestamp 1606716760
transform 1 0 168820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1835
timestamp 1606716760
transform 1 0 169188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1826
timestamp 1606716760
transform 1 0 168360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1824
timestamp 1606716760
transform 1 0 168176 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606716760
transform -1 0 169556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1606716760
transform -1 0 169556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1606716760
transform 1 0 168728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1831
timestamp 1606716760
transform 1 0 168820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1835
timestamp 1606716760
transform 1 0 169188 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1835
timestamp 1606716760
transform 1 0 169188 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1826
timestamp 1606716760
transform 1 0 168360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1606716760
transform -1 0 169556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1830
timestamp 1606716760
transform 1 0 168728 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606716760
transform -1 0 169556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606716760
transform -1 0 169556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1830
timestamp 1606716760
transform 1 0 168728 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1832
timestamp 1606716760
transform 1 0 168912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1814
timestamp 1606716760
transform 1 0 167256 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[6\]
timestamp 1606716760
transform 1 0 165600 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1788
timestamp 1606716760
transform 1 0 164864 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[4\]
timestamp 1606716760
transform 1 0 163208 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1812
timestamp 1606716760
transform 1 0 167072 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[6\]_A
timestamp 1606716760
transform 1 0 166888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[16\]
timestamp 1606716760
transform 1 0 166060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1606716760
transform 1 0 165968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[6\]_TE
timestamp 1606716760
transform 1 0 165600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1798
timestamp 1606716760
transform 1 0 165784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1804
timestamp 1606716760
transform 1 0 166336 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[4\]_A
timestamp 1606716760
transform 1 0 165048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1792
timestamp 1606716760
transform 1 0 165232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_sel_buf\[1\]_A
timestamp 1606716760
transform 1 0 164680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1784
timestamp 1606716760
transform 1 0 164496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1788
timestamp 1606716760
transform 1 0 164864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1814
timestamp 1606716760
transform 1 0 167256 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_stb_buf
timestamp 1606716760
transform 1 0 165600 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_sel_buf\[3\]_A
timestamp 1606716760
transform 1 0 165048 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1792
timestamp 1606716760
transform 1 0 165232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1788
timestamp 1606716760
transform 1 0 164864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_sel_buf\[3\]
timestamp 1606716760
transform 1 0 163208 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1814
timestamp 1606716760
transform 1 0 167256 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1812
timestamp 1606716760
transform 1 0 167072 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_stb_buf_A
timestamp 1606716760
transform 1 0 166888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[9\]
timestamp 1606716760
transform 1 0 166060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1606716760
transform 1 0 165968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_sel_buf\[0\]_A
timestamp 1606716760
transform 1 0 165416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_stb_buf_TE
timestamp 1606716760
transform 1 0 165784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1802
timestamp 1606716760
transform 1 0 166152 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1796
timestamp 1606716760
transform 1 0 165600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1804
timestamp 1606716760
transform 1 0 166336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1792
timestamp 1606716760
transform 1 0 165232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_clk2_buf
timestamp 1606716760
transform 1 0 164496 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1776
timestamp 1606716760
transform 1 0 163760 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_sel_buf\[0\]
timestamp 1606716760
transform 1 0 163576 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1770
timestamp 1606716760
transform 1 0 163208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1770
timestamp 1606716760
transform 1 0 163208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_sel_buf\[0\]_TE
timestamp 1606716760
transform 1 0 163392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[2\]
timestamp 1606716760
transform 1 0 163484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1823
timestamp 1606716760
transform 1 0 168084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[6\]
timestamp 1606716760
transform 1 0 166704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1811
timestamp 1606716760
transform 1 0 166980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1606716760
transform 1 0 166612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_clk2_buf_A
timestamp 1606716760
transform 1 0 165784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_clk2_buf_TE
timestamp 1606716760
transform 1 0 166152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1795
timestamp 1606716760
transform 1 0 165508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1800
timestamp 1606716760
transform 1 0 165968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1804
timestamp 1606716760
transform 1 0 166336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[9\]_A
timestamp 1606716760
transform 1 0 165324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1791
timestamp 1606716760
transform 1 0 165140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[9\]
timestamp 1606716760
transform 1 0 163484 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[9\]_TE
timestamp 1606716760
transform 1 0 163300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1818
timestamp 1606716760
transform 1 0 167624 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[51\]
timestamp 1606716760
transform 1 0 166244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1795
timestamp 1606716760
transform 1 0 165508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1806
timestamp 1606716760
transform 1 0 166520 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_clk_buf
timestamp 1606716760
transform 1 0 163852 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1606716760
transform 1 0 163760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1775
timestamp 1606716760
transform 1 0 163668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[7\]_TE
timestamp 1606716760
transform 1 0 163484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1772
timestamp 1606716760
transform 1 0 163392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1820
timestamp 1606716760
transform 1 0 167808 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1808
timestamp 1606716760
transform 1 0 166704 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1606716760
transform 1 0 166612 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[7\]_A
timestamp 1606716760
transform 1 0 165692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1795
timestamp 1606716760
transform 1 0 165508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1799
timestamp 1606716760
transform 1 0 165876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_clk_buf_A
timestamp 1606716760
transform 1 0 165324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1791
timestamp 1606716760
transform 1 0 165140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[7\]
timestamp 1606716760
transform 1 0 163484 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_clk_buf_TE
timestamp 1606716760
transform 1 0 163300 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1818
timestamp 1606716760
transform 1 0 167624 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[8\]
timestamp 1606716760
transform 1 0 166244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1795
timestamp 1606716760
transform 1 0 165508 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1806
timestamp 1606716760
transform 1 0 166520 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_sel_buf\[2\]
timestamp 1606716760
transform 1 0 163852 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1606716760
transform 1 0 163760 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_we_buf_TE
timestamp 1606716760
transform 1 0 163576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1773
timestamp 1606716760
transform 1 0 163484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1606716760
transform 1 0 163116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_sel_buf\[1\]_TE
timestamp 1606716760
transform 1 0 162840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1761
timestamp 1606716760
transform 1 0 162380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1765
timestamp 1606716760
transform 1 0 162748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1768
timestamp 1606716760
transform 1 0 163024 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[14\]
timestamp 1606716760
transform 1 0 162104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[7\]
timestamp 1606716760
transform 1 0 161092 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1742
timestamp 1606716760
transform 1 0 160632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1746
timestamp 1606716760
transform 1 0 161000 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1750
timestamp 1606716760
transform 1 0 161368 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[6\]_TE
timestamp 1606716760
transform 1 0 160448 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1736
timestamp 1606716760
transform 1 0 160080 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[31\]
timestamp 1606716760
transform 1 0 158424 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  mprj_sel_buf\[1\]
timestamp 1606716760
transform 1 0 162840 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[6\]_A
timestamp 1606716760
transform 1 0 162288 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[4\]_TE
timestamp 1606716760
transform 1 0 162656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1762
timestamp 1606716760
transform 1 0 162472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1758
timestamp 1606716760
transform 1 0 162104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[6\]
timestamp 1606716760
transform 1 0 160448 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1606716760
transform 1 0 160356 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1735
timestamp 1606716760
transform 1 0 159988 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[31\]_A
timestamp 1606716760
transform 1 0 159804 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1731
timestamp 1606716760
transform 1 0 159620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1606716760
transform 1 0 163116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1761
timestamp 1606716760
transform 1 0 162380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[4\]
timestamp 1606716760
transform 1 0 162104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1757
timestamp 1606716760
transform 1 0 162012 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[50\]
timestamp 1606716760
transform 1 0 161000 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1742
timestamp 1606716760
transform 1 0 160632 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1749
timestamp 1606716760
transform 1 0 161276 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[48\]
timestamp 1606716760
transform 1 0 159988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[8\]_TE
timestamp 1606716760
transform 1 0 160448 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1738
timestamp 1606716760
transform 1 0 160264 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[3\]_A
timestamp 1606716760
transform 1 0 159436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1727
timestamp 1606716760
transform 1 0 159252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1731
timestamp 1606716760
transform 1 0 159620 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1762
timestamp 1606716760
transform 1 0 162472 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1766
timestamp 1606716760
transform 1 0 162840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_sel_buf\[3\]_TE
timestamp 1606716760
transform 1 0 163024 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[8\]_A
timestamp 1606716760
transform 1 0 162288 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1606716760
transform 1 0 163116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[46\]
timestamp 1606716760
transform 1 0 161828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1758
timestamp 1606716760
transform 1 0 162104 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1758
timestamp 1606716760
transform 1 0 162104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[4\]_TE
timestamp 1606716760
transform 1 0 161276 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1747
timestamp 1606716760
transform 1 0 161092 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1751
timestamp 1606716760
transform 1 0 161460 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[8\]
timestamp 1606716760
transform 1 0 160448 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1606716760
transform 1 0 160356 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[31\]
timestamp 1606716760
transform 1 0 159436 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[29\]_A
timestamp 1606716760
transform 1 0 159068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1723
timestamp 1606716760
transform 1 0 158884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1727
timestamp 1606716760
transform 1 0 159252 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[30\]_A
timestamp 1606716760
transform 1 0 158516 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1718
timestamp 1606716760
transform 1 0 158424 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1721
timestamp 1606716760
transform 1 0 158700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[4\]_A
timestamp 1606716760
transform 1 0 162932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1765
timestamp 1606716760
transform 1 0 162748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1769
timestamp 1606716760
transform 1 0 163116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[4\]
timestamp 1606716760
transform 1 0 161092 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1606716760
transform 1 0 161000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[31\]_A
timestamp 1606716760
transform 1 0 160724 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1745
timestamp 1606716760
transform 1 0 160908 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[28\]_A
timestamp 1606716760
transform 1 0 160172 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1735
timestamp 1606716760
transform 1 0 159988 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1739
timestamp 1606716760
transform 1 0 160356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[28\]
timestamp 1606716760
transform 1 0 158332 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[1\]
timestamp 1606716760
transform 1 0 162748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1764
timestamp 1606716760
transform 1 0 162656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1768
timestamp 1606716760
transform 1 0 163024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[2\]_A
timestamp 1606716760
transform 1 0 161736 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1756
timestamp 1606716760
transform 1 0 161920 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1752
timestamp 1606716760
transform 1 0 161552 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[2\]
timestamp 1606716760
transform 1 0 159896 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[31\]_TE
timestamp 1606716760
transform 1 0 159436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1724
timestamp 1606716760
transform 1 0 158976 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1728
timestamp 1606716760
transform 1 0 159344 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1731
timestamp 1606716760
transform 1 0 159620 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[70\]
timestamp 1606716760
transform 1 0 158700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1716
timestamp 1606716760
transform 1 0 158240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1720
timestamp 1606716760
transform 1 0 158608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[5\]_A
timestamp 1606716760
transform 1 0 162932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1765
timestamp 1606716760
transform 1 0 162748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1769
timestamp 1606716760
transform 1 0 163116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[5\]
timestamp 1606716760
transform 1 0 161092 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1606716760
transform 1 0 161000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[5\]_TE
timestamp 1606716760
transform 1 0 160816 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1742
timestamp 1606716760
transform 1 0 160632 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[44\]
timestamp 1606716760
transform 1 0 159988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[2\]_TE
timestamp 1606716760
transform 1 0 160448 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1738
timestamp 1606716760
transform 1 0 160264 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1724
timestamp 1606716760
transform 1 0 158976 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1732
timestamp 1606716760
transform 1 0 159712 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[49\]
timestamp 1606716760
transform 1 0 162472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1765
timestamp 1606716760
transform 1 0 162748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1754
timestamp 1606716760
transform 1 0 161736 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[47\]
timestamp 1606716760
transform 1 0 161460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1747
timestamp 1606716760
transform 1 0 161092 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1735
timestamp 1606716760
transform 1 0 159988 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[73\]
timestamp 1606716760
transform 1 0 159712 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1731
timestamp 1606716760
transform 1 0 159620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[69\]
timestamp 1606716760
transform 1 0 158240 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1719
timestamp 1606716760
transform 1 0 158516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1606716760
transform 1 0 157504 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[3\]_TE
timestamp 1606716760
transform 1 0 157964 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1709
timestamp 1606716760
transform 1 0 157596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1715
timestamp 1606716760
transform 1 0 158148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1696
timestamp 1606716760
transform 1 0 156400 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[2\]
timestamp 1606716760
transform 1 0 154744 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1666
timestamp 1606716760
transform 1 0 153640 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[3\]
timestamp 1606716760
transform 1 0 157964 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[31\]_TE
timestamp 1606716760
transform 1 0 157780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[45\]
timestamp 1606716760
transform 1 0 156952 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1701
timestamp 1606716760
transform 1 0 156860 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1705
timestamp 1606716760
transform 1 0 157228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[65\]
timestamp 1606716760
transform 1 0 155848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[2\]_A
timestamp 1606716760
transform 1 0 156308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1693
timestamp 1606716760
transform 1 0 156124 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1697
timestamp 1606716760
transform 1 0 156492 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[2\]_TE
timestamp 1606716760
transform 1 0 155296 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1682
timestamp 1606716760
transform 1 0 155112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1686
timestamp 1606716760
transform 1 0 155480 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[64\]
timestamp 1606716760
transform 1 0 154836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1606716760
transform 1 0 154744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1677
timestamp 1606716760
transform 1 0 154652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[59\]
timestamp 1606716760
transform 1 0 153640 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1664
timestamp 1606716760
transform 1 0 153456 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1669
timestamp 1606716760
transform 1 0 153916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[29\]
timestamp 1606716760
transform 1 0 157596 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1606716760
transform 1 0 157504 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[30\]_TE
timestamp 1606716760
transform 1 0 157228 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1703
timestamp 1606716760
transform 1 0 157044 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1707
timestamp 1606716760
transform 1 0 157412 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[23\]_A
timestamp 1606716760
transform 1 0 156124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1691
timestamp 1606716760
transform 1 0 155940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1695
timestamp 1606716760
transform 1 0 156308 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[23\]
timestamp 1606716760
transform 1 0 154284 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_16_1670
timestamp 1606716760
transform 1 0 154008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[71\]
timestamp 1606716760
transform 1 0 157596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1606716760
transform 1 0 157504 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1712
timestamp 1606716760
transform 1 0 157872 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[30\]
timestamp 1606716760
transform 1 0 157228 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[29\]_TE
timestamp 1606716760
transform 1 0 157044 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1700
timestamp 1606716760
transform 1 0 156768 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1701
timestamp 1606716760
transform 1 0 156860 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[22\]_A
timestamp 1606716760
transform 1 0 156584 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[24\]_A
timestamp 1606716760
transform 1 0 156676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1696
timestamp 1606716760
transform 1 0 156400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1697
timestamp 1606716760
transform 1 0 156492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[24\]
timestamp 1606716760
transform 1 0 154836 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[22\]
timestamp 1606716760
transform 1 0 154744 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1675
timestamp 1606716760
transform 1 0 154468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1674
timestamp 1606716760
transform 1 0 154376 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[23\]_TE
timestamp 1606716760
transform 1 0 154284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[17\]_A
timestamp 1606716760
transform 1 0 154192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1606716760
transform 1 0 154744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1667
timestamp 1606716760
transform 1 0 153732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1663
timestamp 1606716760
transform 1 0 153364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[24\]_TE
timestamp 1606716760
transform 1 0 153916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[19\]_A
timestamp 1606716760
transform 1 0 153548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1671
timestamp 1606716760
transform 1 0 154100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1670
timestamp 1606716760
transform 1 0 154008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[28\]_TE
timestamp 1606716760
transform 1 0 158148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1708
timestamp 1606716760
transform 1 0 157504 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1714
timestamp 1606716760
transform 1 0 158056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[26\]_A
timestamp 1606716760
transform 1 0 157320 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1704
timestamp 1606716760
transform 1 0 157136 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[26\]
timestamp 1606716760
transform 1 0 155480 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1606716760
transform 1 0 155388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[22\]_TE
timestamp 1606716760
transform 1 0 155204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[18\]_A
timestamp 1606716760
transform 1 0 154836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1677
timestamp 1606716760
transform 1 0 154652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1681
timestamp 1606716760
transform 1 0 155020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1606716760
transform 1 0 158148 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1714
timestamp 1606716760
transform 1 0 158056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1702
timestamp 1606716760
transform 1 0 156952 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[60\]
timestamp 1606716760
transform 1 0 156676 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[26\]_TE
timestamp 1606716760
transform 1 0 156124 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1691
timestamp 1606716760
transform 1 0 155940 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1695
timestamp 1606716760
transform 1 0 156308 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[1\]
timestamp 1606716760
transform 1 0 154284 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1665
timestamp 1606716760
transform 1 0 153548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1712
timestamp 1606716760
transform 1 0 157872 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1700
timestamp 1606716760
transform 1 0 156768 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[68\]
timestamp 1606716760
transform 1 0 156492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[1\]_A
timestamp 1606716760
transform 1 0 155940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1689
timestamp 1606716760
transform 1 0 155756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1693
timestamp 1606716760
transform 1 0 156124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[42\]
timestamp 1606716760
transform 1 0 155480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1606716760
transform 1 0 155388 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[1\]_TE
timestamp 1606716760
transform 1 0 155204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[13\]_A
timestamp 1606716760
transform 1 0 154836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1677
timestamp 1606716760
transform 1 0 154652 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1681
timestamp 1606716760
transform 1 0 155020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1606716760
transform 1 0 158148 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[72\]
timestamp 1606716760
transform 1 0 156768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1703
timestamp 1606716760
transform 1 0 157044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[55\]
timestamp 1606716760
transform 1 0 155756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[25\]_TE
timestamp 1606716760
transform 1 0 156216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1692
timestamp 1606716760
transform 1 0 156032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1696
timestamp 1606716760
transform 1 0 156400 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1681
timestamp 1606716760
transform 1 0 155020 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[0\]
timestamp 1606716760
transform 1 0 153364 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[28\]
timestamp 1606716760
transform 1 0 151984 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1606716760
transform 1 0 151892 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1637
timestamp 1606716760
transform 1 0 150972 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1645
timestamp 1606716760
transform 1 0 151708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[15\]
timestamp 1606716760
transform 1 0 149316 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1617
timestamp 1606716760
transform 1 0 149132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[28\]_A
timestamp 1606716760
transform 1 0 153272 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1658
timestamp 1606716760
transform 1 0 152904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[54\]
timestamp 1606716760
transform 1 0 152628 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[28\]_TE
timestamp 1606716760
transform 1 0 152076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1647
timestamp 1606716760
transform 1 0 151892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1651
timestamp 1606716760
transform 1 0 152260 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[38\]
timestamp 1606716760
transform 1 0 151616 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[12\]_A
timestamp 1606716760
transform 1 0 151064 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[15\]_A
timestamp 1606716760
transform 1 0 151432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1640
timestamp 1606716760
transform 1 0 151248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1636
timestamp 1606716760
transform 1 0 150880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[12\]
timestamp 1606716760
transform 1 0 149224 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1606716760
transform 1 0 149132 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[12\]_TE
timestamp 1606716760
transform 1 0 148948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[15\]_TE
timestamp 1606716760
transform 1 0 148580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1609
timestamp 1606716760
transform 1 0 148396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1613
timestamp 1606716760
transform 1 0 148764 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[57\]
timestamp 1606716760
transform 1 0 152996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1662
timestamp 1606716760
transform 1 0 153272 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[56\]
timestamp 1606716760
transform 1 0 151984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1606716760
transform 1 0 151892 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1651
timestamp 1606716760
transform 1 0 152260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[19\]_TE
timestamp 1606716760
transform 1 0 151708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1643
timestamp 1606716760
transform 1 0 151524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[11\]_A
timestamp 1606716760
transform 1 0 150604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1631
timestamp 1606716760
transform 1 0 150420 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1635
timestamp 1606716760
transform 1 0 150788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[11\]
timestamp 1606716760
transform 1 0 148764 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[14\]_TE
timestamp 1606716760
transform 1 0 148580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1609
timestamp 1606716760
transform 1 0 148396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[17\]
timestamp 1606716760
transform 1 0 152352 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1648
timestamp 1606716760
transform 1 0 151984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1606716760
transform 1 0 151892 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[19\]
timestamp 1606716760
transform 1 0 151708 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1646
timestamp 1606716760
transform 1 0 151800 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1641
timestamp 1606716760
transform 1 0 151340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1637
timestamp 1606716760
transform 1 0 150972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1640
timestamp 1606716760
transform 1 0 151248 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[14\]_A
timestamp 1606716760
transform 1 0 151156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[10\]_A
timestamp 1606716760
transform 1 0 151064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1636
timestamp 1606716760
transform 1 0 150880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[10\]
timestamp 1606716760
transform 1 0 149224 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[14\]
timestamp 1606716760
transform 1 0 149316 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1618
timestamp 1606716760
transform 1 0 149224 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1615
timestamp 1606716760
transform 1 0 148948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1617
timestamp 1606716760
transform 1 0 149132 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[11\]_TE
timestamp 1606716760
transform 1 0 148764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1606716760
transform 1 0 149132 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1610
timestamp 1606716760
transform 1 0 148488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1609
timestamp 1606716760
transform 1 0 148396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[18\]
timestamp 1606716760
transform 1 0 152996 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[18\]_TE
timestamp 1606716760
transform 1 0 152812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[17\]_TE
timestamp 1606716760
transform 1 0 152352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1647
timestamp 1606716760
transform 1 0 151892 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1651
timestamp 1606716760
transform 1 0 152260 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1654
timestamp 1606716760
transform 1 0 152536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[27\]_A
timestamp 1606716760
transform 1 0 151708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1643
timestamp 1606716760
transform 1 0 151524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[27\]
timestamp 1606716760
transform 1 0 149868 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1606716760
transform 1 0 149776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[9\]_A
timestamp 1606716760
transform 1 0 149224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[27\]_TE
timestamp 1606716760
transform 1 0 149592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1620
timestamp 1606716760
transform 1 0 149408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1616
timestamp 1606716760
transform 1 0 149040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[43\]
timestamp 1606716760
transform 1 0 153272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[13\]_TE
timestamp 1606716760
transform 1 0 152996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1661
timestamp 1606716760
transform 1 0 153180 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1606716760
transform 1 0 152536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1653
timestamp 1606716760
transform 1 0 152444 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1655
timestamp 1606716760
transform 1 0 152628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[52\]
timestamp 1606716760
transform 1 0 151432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1645
timestamp 1606716760
transform 1 0 151708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[37\]
timestamp 1606716760
transform 1 0 150420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1634
timestamp 1606716760
transform 1 0 150696 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[10\]_TE
timestamp 1606716760
transform 1 0 149868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1623
timestamp 1606716760
transform 1 0 149684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1627
timestamp 1606716760
transform 1 0 150052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[13\]
timestamp 1606716760
transform 1 0 152996 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[30\]_A
timestamp 1606716760
transform 1 0 152444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1651
timestamp 1606716760
transform 1 0 152260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1655
timestamp 1606716760
transform 1 0 152628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[30\]
timestamp 1606716760
transform 1 0 150604 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[30\]_TE
timestamp 1606716760
transform 1 0 150420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1606716760
transform 1 0 149776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[23\]_A
timestamp 1606716760
transform 1 0 149316 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1621
timestamp 1606716760
transform 1 0 149500 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1625
timestamp 1606716760
transform 1 0 149868 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[23\]_TE
timestamp 1606716760
transform 1 0 148580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1609
timestamp 1606716760
transform 1 0 148396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1613
timestamp 1606716760
transform 1 0 148764 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[20\]_TE
timestamp 1606716760
transform 1 0 152996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1661
timestamp 1606716760
transform 1 0 153180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1606716760
transform 1 0 152536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1650
timestamp 1606716760
transform 1 0 152168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1655
timestamp 1606716760
transform 1 0 152628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1638
timestamp 1606716760
transform 1 0 151064 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[40\]
timestamp 1606716760
transform 1 0 150788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1627
timestamp 1606716760
transform 1 0 150052 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[29\]
timestamp 1606716760
transform 1 0 148396 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1605
timestamp 1606716760
transform 1 0 148028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_cyc_buf
timestamp 1606716760
transform 1 0 146372 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1606716760
transform 1 0 146280 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1585
timestamp 1606716760
transform 1 0 146188 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[19\]_A
timestamp 1606716760
transform 1 0 145636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1577
timestamp 1606716760
transform 1 0 145452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1581
timestamp 1606716760
transform 1 0 145820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[19\]
timestamp 1606716760
transform 1 0 143796 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1558
timestamp 1606716760
transform 1 0 143704 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[53\]
timestamp 1606716760
transform 1 0 148120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[19\]
timestamp 1606716760
transform 1 0 147108 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_cyc_buf_A
timestamp 1606716760
transform 1 0 147660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_cyc_buf_TE
timestamp 1606716760
transform 1 0 146924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1598
timestamp 1606716760
transform 1 0 147384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1603
timestamp 1606716760
transform 1 0 147844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[3\]_A
timestamp 1606716760
transform 1 0 146556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1587
timestamp 1606716760
transform 1 0 146372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1591
timestamp 1606716760
transform 1 0 146740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[3\]
timestamp 1606716760
transform 1 0 144716 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[3\]_TE
timestamp 1606716760
transform 1 0 144532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[10\]
timestamp 1606716760
transform 1 0 143612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1606716760
transform 1 0 143520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[19\]_TE
timestamp 1606716760
transform 1 0 144072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1560
timestamp 1606716760
transform 1 0 143888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1564
timestamp 1606716760
transform 1 0 144256 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[7\]_A
timestamp 1606716760
transform 1 0 148212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1605
timestamp 1606716760
transform 1 0 148028 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[7\]
timestamp 1606716760
transform 1 0 146372 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1606716760
transform 1 0 146280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1575
timestamp 1606716760
transform 1 0 145268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_1583
timestamp 1606716760
transform 1 0 146004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[17\]
timestamp 1606716760
transform 1 0 144992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[13\]
timestamp 1606716760
transform 1 0 143980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1564
timestamp 1606716760
transform 1 0 144256 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1606
timestamp 1606716760
transform 1 0 148120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1605
timestamp 1606716760
transform 1 0 148028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[5\]_A
timestamp 1606716760
transform 1 0 148304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[1\]_A
timestamp 1606716760
transform 1 0 148212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[5\]
timestamp 1606716760
transform 1 0 146464 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[1\]
timestamp 1606716760
transform 1 0 146372 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1584
timestamp 1606716760
transform 1 0 146096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[5\]_TE
timestamp 1606716760
transform 1 0 146280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1606716760
transform 1 0 146280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1574
timestamp 1606716760
transform 1 0 145176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[15\]
timestamp 1606716760
transform 1 0 145268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[7\]_TE
timestamp 1606716760
transform 1 0 145912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1578
timestamp 1606716760
transform 1 0 145544 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1579
timestamp 1606716760
transform 1 0 145636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1571
timestamp 1606716760
transform 1 0 144900 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1569
timestamp 1606716760
transform 1 0 144716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[18\]_TE
timestamp 1606716760
transform 1 0 144992 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[29\]
timestamp 1606716760
transform 1 0 144624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[22\]
timestamp 1606716760
transform 1 0 143612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1606716760
transform 1 0 143520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1561
timestamp 1606716760
transform 1 0 143980 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1555
timestamp 1606716760
transform 1 0 143428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1560
timestamp 1606716760
transform 1 0 143888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[9\]
timestamp 1606716760
transform 1 0 147384 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[1\]_TE
timestamp 1606716760
transform 1 0 147200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1594
timestamp 1606716760
transform 1 0 147016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[18\]_A
timestamp 1606716760
transform 1 0 146832 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1590
timestamp 1606716760
transform 1 0 146648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[18\]
timestamp 1606716760
transform 1 0 144992 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1606716760
transform 1 0 144164 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[12\]_A
timestamp 1606716760
transform 1 0 143612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[16\]_A
timestamp 1606716760
transform 1 0 143980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1555
timestamp 1606716760
transform 1 0 143428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1559
timestamp 1606716760
transform 1 0 143796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1564
timestamp 1606716760
transform 1 0 144256 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[23\]
timestamp 1606716760
transform 1 0 148028 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[11\]
timestamp 1606716760
transform 1 0 147016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1606716760
transform 1 0 146924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[9\]_TE
timestamp 1606716760
transform 1 0 147476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1597
timestamp 1606716760
transform 1 0 147292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1601
timestamp 1606716760
transform 1 0 147660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1589
timestamp 1606716760
transform 1 0 146556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[28\]
timestamp 1606716760
transform 1 0 145176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1577
timestamp 1606716760
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1566
timestamp 1606716760
transform 1 0 144440 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[33\]
timestamp 1606716760
transform 1 0 148120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1598
timestamp 1606716760
transform 1 0 147384 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1586
timestamp 1606716760
transform 1 0 146280 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[3\]
timestamp 1606716760
transform 1 0 146004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1580
timestamp 1606716760
transform 1 0 145728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[14\]_A
timestamp 1606716760
transform 1 0 144440 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1568
timestamp 1606716760
transform 1 0 144624 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1606716760
transform 1 0 144164 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[10\]_A
timestamp 1606716760
transform 1 0 143612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1555
timestamp 1606716760
transform 1 0 143428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1559
timestamp 1606716760
transform 1 0 143796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1564
timestamp 1606716760
transform 1 0 144256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1606
timestamp 1606716760
transform 1 0 148120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1606716760
transform 1 0 146924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1594
timestamp 1606716760
transform 1 0 147016 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1591
timestamp 1606716760
transform 1 0 146740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1579
timestamp 1606716760
transform 1 0 145636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1567
timestamp 1606716760
transform 1 0 144532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1555
timestamp 1606716760
transform 1 0 143428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1546
timestamp 1606716760
transform 1 0 142600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[0\]
timestamp 1606716760
transform 1 0 140944 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1606716760
transform 1 0 140668 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[99\]_TE
timestamp 1606716760
transform 1 0 140392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1524
timestamp 1606716760
transform 1 0 140576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1526
timestamp 1606716760
transform 1 0 140760 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1514
timestamp 1606716760
transform 1 0 139656 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1606716760
transform 1 0 139012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[97\]_A
timestamp 1606716760
transform 1 0 139472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1506
timestamp 1606716760
transform 1 0 138920 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1510
timestamp 1606716760
transform 1 0 139288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[0\]_A
timestamp 1606716760
transform 1 0 142232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[99\]_A
timestamp 1606716760
transform 1 0 142600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1540
timestamp 1606716760
transform 1 0 142048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1544
timestamp 1606716760
transform 1 0 142416 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1548
timestamp 1606716760
transform 1 0 142784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[99\]
timestamp 1606716760
transform 1 0 140392 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1606716760
transform 1 0 139840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1514
timestamp 1606716760
transform 1 0 139656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1518
timestamp 1606716760
transform 1 0 140024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1553
timestamp 1606716760
transform 1 0 143244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[25\]
timestamp 1606716760
transform 1 0 141588 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1534
timestamp 1606716760
transform 1 0 141496 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1606716760
transform 1 0 140668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[0\]_TE
timestamp 1606716760
transform 1 0 140944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1524
timestamp 1606716760
transform 1 0 140576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1526
timestamp 1606716760
transform 1 0 140760 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1530
timestamp 1606716760
transform 1 0 141128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[25\]
timestamp 1606716760
transform 1 0 139196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1508
timestamp 1606716760
transform 1 0 139104 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1512
timestamp 1606716760
transform 1 0 139472 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[25\]_A
timestamp 1606716760
transform 1 0 143244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[12\]
timestamp 1606716760
transform 1 0 142324 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[21\]_A
timestamp 1606716760
transform 1 0 142876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[25\]_TE
timestamp 1606716760
transform 1 0 142140 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1547
timestamp 1606716760
transform 1 0 142692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1551
timestamp 1606716760
transform 1 0 143060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[16\]_TE
timestamp 1606716760
transform 1 0 141772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1535
timestamp 1606716760
transform 1 0 141588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1539
timestamp 1606716760
transform 1 0 141956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[21\]
timestamp 1606716760
transform 1 0 141036 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[26\]
timestamp 1606716760
transform 1 0 141312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1606716760
transform 1 0 140668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[21\]_TE
timestamp 1606716760
transform 1 0 140852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1526
timestamp 1606716760
transform 1 0 140760 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1521
timestamp 1606716760
transform 1 0 140300 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[27\]
timestamp 1606716760
transform 1 0 140024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[35\]
timestamp 1606716760
transform 1 0 139656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1517
timestamp 1606716760
transform 1 0 139932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[301\]
timestamp 1606716760
transform 1 0 139012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1513
timestamp 1606716760
transform 1 0 139564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1510
timestamp 1606716760
transform 1 0 139288 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[16\]
timestamp 1606716760
transform 1 0 141772 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1536
timestamp 1606716760
transform 1 0 141680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[31\]
timestamp 1606716760
transform 1 0 140668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1523
timestamp 1606716760
transform 1 0 140484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1528
timestamp 1606716760
transform 1 0 140944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1515
timestamp 1606716760
transform 1 0 139748 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1606716760
transform 1 0 138552 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1503
timestamp 1606716760
transform 1 0 138644 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[14\]
timestamp 1606716760
transform 1 0 142784 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[12\]_TE
timestamp 1606716760
transform 1 0 142324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1545
timestamp 1606716760
transform 1 0 142508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[10\]_TE
timestamp 1606716760
transform 1 0 141772 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1533
timestamp 1606716760
transform 1 0 141404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1539
timestamp 1606716760
transform 1 0 141956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1606716760
transform 1 0 141312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1520
timestamp 1606716760
transform 1 0 140208 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1508
timestamp 1606716760
transform 1 0 139104 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[10\]
timestamp 1606716760
transform 1 0 141772 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1535
timestamp 1606716760
transform 1 0 141588 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1527
timestamp 1606716760
transform 1 0 140852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1515
timestamp 1606716760
transform 1 0 139748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1606716760
transform 1 0 138552 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1503
timestamp 1606716760
transform 1 0 138644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[24\]
timestamp 1606716760
transform 1 0 143152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[20\]
timestamp 1606716760
transform 1 0 142140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[14\]_TE
timestamp 1606716760
transform 1 0 142784 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1544
timestamp 1606716760
transform 1 0 142416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1550
timestamp 1606716760
transform 1 0 142968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1533
timestamp 1606716760
transform 1 0 141404 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1606716760
transform 1 0 141312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1523
timestamp 1606716760
transform 1 0 140484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1531
timestamp 1606716760
transform 1 0 141220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1511
timestamp 1606716760
transform 1 0 139380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[97\]_TE
timestamp 1606716760
transform 1 0 138000 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1494
timestamp 1606716760
transform 1 0 137816 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1498
timestamp 1606716760
transform 1 0 138184 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[95\]
timestamp 1606716760
transform 1 0 136160 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1468
timestamp 1606716760
transform 1 0 135424 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1606716760
transform 1 0 135148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1606716760
transform 1 0 135056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1606716760
transform 1 0 134044 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[46\]_A
timestamp 1606716760
transform 1 0 133676 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1448
timestamp 1606716760
transform 1 0 133584 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1451
timestamp 1606716760
transform 1 0 133860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1456
timestamp 1606716760
transform 1 0 134320 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[97\]
timestamp 1606716760
transform 1 0 138000 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1606716760
transform 1 0 137908 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[95\]_A
timestamp 1606716760
transform 1 0 137448 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1492
timestamp 1606716760
transform 1 0 137632 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[95\]_TE
timestamp 1606716760
transform 1 0 136712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1484
timestamp 1606716760
transform 1 0 136896 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[297\]
timestamp 1606716760
transform 1 0 136252 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1606716760
transform 1 0 135608 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1468
timestamp 1606716760
transform 1 0 135424 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1472
timestamp 1606716760
transform 1 0 135792 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1476
timestamp 1606716760
transform 1 0 136160 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1480
timestamp 1606716760
transform 1 0 136528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1606716760
transform 1 0 135240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1464
timestamp 1606716760
transform 1 0 135056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1606716760
transform 1 0 134780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1606716760
transform 1 0 134228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1453
timestamp 1606716760
transform 1 0 134044 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1457
timestamp 1606716760
transform 1 0 134412 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[23\]
timestamp 1606716760
transform 1 0 137724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1492
timestamp 1606716760
transform 1 0 137632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1496
timestamp 1606716760
transform 1 0 138000 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1468
timestamp 1606716760
transform 1 0 135424 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1480
timestamp 1606716760
transform 1 0 136528 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[295\]
timestamp 1606716760
transform 1 0 135148 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1606716760
transform 1 0 135056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1458
timestamp 1606716760
transform 1 0 134504 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1501
timestamp 1606716760
transform 1 0 138460 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1499
timestamp 1606716760
transform 1 0 138276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[299\]
timestamp 1606716760
transform 1 0 138000 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1606716760
transform 1 0 137908 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1489
timestamp 1606716760
transform 1 0 137356 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1483
timestamp 1606716760
transform 1 0 136804 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1477
timestamp 1606716760
transform 1 0 136252 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1471
timestamp 1606716760
transform 1 0 135700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1606716760
transform 1 0 135056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1463
timestamp 1606716760
transform 1 0 134964 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1465
timestamp 1606716760
transform 1 0 135148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1457
timestamp 1606716760
transform 1 0 134412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1459
timestamp 1606716760
transform 1 0 134596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1500
timestamp 1606716760
transform 1 0 138368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1488
timestamp 1606716760
transform 1 0 137264 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1476
timestamp 1606716760
transform 1 0 136160 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[45\]_A
timestamp 1606716760
transform 1 0 134872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1464
timestamp 1606716760
transform 1 0 135056 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1460
timestamp 1606716760
transform 1 0 134688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1496
timestamp 1606716760
transform 1 0 138000 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1484
timestamp 1606716760
transform 1 0 136896 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1606716760
transform 1 0 135700 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1470
timestamp 1606716760
transform 1 0 135608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1472
timestamp 1606716760
transform 1 0 135792 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[47\]_TE
timestamp 1606716760
transform 1 0 134872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1464
timestamp 1606716760
transform 1 0 135056 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1451
timestamp 1606716760
transform 1 0 133860 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1459
timestamp 1606716760
transform 1 0 134596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1496
timestamp 1606716760
transform 1 0 138000 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[47\]_A
timestamp 1606716760
transform 1 0 136712 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1484
timestamp 1606716760
transform 1 0 136896 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1480
timestamp 1606716760
transform 1 0 136528 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[47\]
timestamp 1606716760
transform 1 0 134872 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1449
timestamp 1606716760
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1461
timestamp 1606716760
transform 1 0 134780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1499
timestamp 1606716760
transform 1 0 138276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1487
timestamp 1606716760
transform 1 0 137172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[249\]
timestamp 1606716760
transform 1 0 135792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1606716760
transform 1 0 135700 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1475
timestamp 1606716760
transform 1 0 136068 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1459
timestamp 1606716760
transform 1 0 134596 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[284\]
timestamp 1606716760
transform 1 0 132940 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[46\]_TE
timestamp 1606716760
transform 1 0 132388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1433
timestamp 1606716760
transform 1 0 132204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1437
timestamp 1606716760
transform 1 0 132572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1444
timestamp 1606716760
transform 1 0 133216 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[245\]
timestamp 1606716760
transform 1 0 131928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1422
timestamp 1606716760
transform 1 0 131192 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[82\]
timestamp 1606716760
transform 1 0 129536 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1606716760
transform 1 0 129444 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1395
timestamp 1606716760
transform 1 0 128708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[46\]
timestamp 1606716760
transform 1 0 132388 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1606716760
transform 1 0 132296 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1432
timestamp 1606716760
transform 1 0 132112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _607_
timestamp 1606716760
transform 1 0 130364 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__A
timestamp 1606716760
transform 1 0 130824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[82\]_A
timestamp 1606716760
transform 1 0 131192 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1416
timestamp 1606716760
transform 1 0 130640 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1420
timestamp 1606716760
transform 1 0 131008 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1424
timestamp 1606716760
transform 1 0 131376 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[82\]_TE
timestamp 1606716760
transform 1 0 130180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1409
timestamp 1606716760
transform 1 0 129996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[39\]_A
timestamp 1606716760
transform 1 0 129812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1405
timestamp 1606716760
transform 1 0 129628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[248\]
timestamp 1606716760
transform 1 0 132112 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[293\]
timestamp 1606716760
transform 1 0 133124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1435
timestamp 1606716760
transform 1 0 132388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1446
timestamp 1606716760
transform 1 0 133400 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1428
timestamp 1606716760
transform 1 0 131744 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[84\]_A
timestamp 1606716760
transform 1 0 131560 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1424
timestamp 1606716760
transform 1 0 131376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[84\]
timestamp 1606716760
transform 1 0 129720 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1606716760
transform 1 0 129444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[84\]_TE
timestamp 1606716760
transform 1 0 129260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1400
timestamp 1606716760
transform 1 0 129168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1404
timestamp 1606716760
transform 1 0 129536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1447
timestamp 1606716760
transform 1 0 133492 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[247\]
timestamp 1606716760
transform 1 0 132664 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1606716760
transform 1 0 132296 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[45\]_TE
timestamp 1606716760
transform 1 0 133124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1434
timestamp 1606716760
transform 1 0 132296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1441
timestamp 1606716760
transform 1 0 132940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1445
timestamp 1606716760
transform 1 0 133308 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1435
timestamp 1606716760
transform 1 0 132388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[42\]_A
timestamp 1606716760
transform 1 0 131744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1430
timestamp 1606716760
transform 1 0 131928 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1422
timestamp 1606716760
transform 1 0 131192 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1426
timestamp 1606716760
transform 1 0 131560 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[41\]
timestamp 1606716760
transform 1 0 129536 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[42\]
timestamp 1606716760
transform 1 0 129904 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1606716760
transform 1 0 129444 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[40\]_A
timestamp 1606716760
transform 1 0 129352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[42\]_TE
timestamp 1606716760
transform 1 0 129720 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1400
timestamp 1606716760
transform 1 0 129168 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1404
timestamp 1606716760
transform 1 0 129536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[45\]
timestamp 1606716760
transform 1 0 133032 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1606716760
transform 1 0 132940 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1436
timestamp 1606716760
transform 1 0 132480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1440
timestamp 1606716760
transform 1 0 132848 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[286\]
timestamp 1606716760
transform 1 0 130732 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[41\]_A
timestamp 1606716760
transform 1 0 131192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1420
timestamp 1606716760
transform 1 0 131008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1424
timestamp 1606716760
transform 1 0 131376 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1409
timestamp 1606716760
transform 1 0 129996 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[243\]
timestamp 1606716760
transform 1 0 128708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[244\]
timestamp 1606716760
transform 1 0 129720 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[41\]_TE
timestamp 1606716760
transform 1 0 129536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1398
timestamp 1606716760
transform 1 0 128984 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[44\]
timestamp 1606716760
transform 1 0 132204 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1432
timestamp 1606716760
transform 1 0 132112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1414
timestamp 1606716760
transform 1 0 130456 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1426
timestamp 1606716760
transform 1 0 131560 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[239\]
timestamp 1606716760
transform 1 0 130180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1606716760
transform 1 0 130088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1409
timestamp 1606716760
transform 1 0 129996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[37\]_TE
timestamp 1606716760
transform 1 0 129812 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1400
timestamp 1606716760
transform 1 0 129168 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1406
timestamp 1606716760
transform 1 0 129720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[44\]_A
timestamp 1606716760
transform 1 0 133492 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[246\]
timestamp 1606716760
transform 1 0 133032 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1606716760
transform 1 0 132940 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[44\]_TE
timestamp 1606716760
transform 1 0 132204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1435
timestamp 1606716760
transform 1 0 132388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1445
timestamp 1606716760
transform 1 0 133308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1429
timestamp 1606716760
transform 1 0 131836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[37\]_A
timestamp 1606716760
transform 1 0 131652 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1425
timestamp 1606716760
transform 1 0 131468 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[37\]
timestamp 1606716760
transform 1 0 129812 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[32\]_A
timestamp 1606716760
transform 1 0 129260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1399
timestamp 1606716760
transform 1 0 129076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1403
timestamp 1606716760
transform 1 0 129444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1447
timestamp 1606716760
transform 1 0 133492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1435
timestamp 1606716760
transform 1 0 132388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1423
timestamp 1606716760
transform 1 0 131284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1606716760
transform 1 0 130088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1411
timestamp 1606716760
transform 1 0 130180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[205\]
timestamp 1606716760
transform 1 0 129076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1398
timestamp 1606716760
transform 1 0 128984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1402
timestamp 1606716760
transform 1 0 129352 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1606716760
transform 1 0 128064 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[35\]_A
timestamp 1606716760
transform 1 0 127512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[39\]_TE
timestamp 1606716760
transform 1 0 128524 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1380
timestamp 1606716760
transform 1 0 127328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1384
timestamp 1606716760
transform 1 0 127696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1391
timestamp 1606716760
transform 1 0 128340 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[35\]
timestamp 1606716760
transform 1 0 125672 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1606716760
transform 1 0 124660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1343
timestamp 1606716760
transform 1 0 123924 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1354
timestamp 1606716760
transform 1 0 124936 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1606716760
transform 1 0 123832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[39\]
timestamp 1606716760
transform 1 0 127972 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A
timestamp 1606716760
transform 1 0 127236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1606716760
transform 1 0 127788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1381
timestamp 1606716760
transform 1 0 127420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1377
timestamp 1606716760
transform 1 0 127052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1606716760
transform 1 0 126776 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1606716760
transform 1 0 126684 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1606716760
transform 1 0 125856 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[35\]_TE
timestamp 1606716760
transform 1 0 126224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1362
timestamp 1606716760
transform 1 0 125672 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1366
timestamp 1606716760
transform 1 0 126040 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1370
timestamp 1606716760
transform 1 0 126408 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1606716760
transform 1 0 125396 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1606716760
transform 1 0 125212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1606716760
transform 1 0 124384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1606716760
transform 1 0 124844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1347
timestamp 1606716760
transform 1 0 124292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1351
timestamp 1606716760
transform 1 0 124660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1355
timestamp 1606716760
transform 1 0 125028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[210\]
timestamp 1606716760
transform 1 0 127788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[40\]_TE
timestamp 1606716760
transform 1 0 127512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1381
timestamp 1606716760
transform 1 0 127420 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1384
timestamp 1606716760
transform 1 0 127696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1388
timestamp 1606716760
transform 1 0 128064 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1377
timestamp 1606716760
transform 1 0 127052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1606716760
transform 1 0 126776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1366
timestamp 1606716760
transform 1 0 126040 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[33\]
timestamp 1606716760
transform 1 0 124384 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1343
timestamp 1606716760
transform 1 0 123924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1347
timestamp 1606716760
transform 1 0 124292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1606716760
transform 1 0 123832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[241\]
timestamp 1606716760
transform 1 0 128064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[40\]
timestamp 1606716760
transform 1 0 127512 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1380
timestamp 1606716760
transform 1 0 127328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1391
timestamp 1606716760
transform 1 0 128340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1606716760
transform 1 0 126960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1378
timestamp 1606716760
transform 1 0 127144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[34\]
timestamp 1606716760
transform 1 0 125672 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1606716760
transform 1 0 126684 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[33\]_A
timestamp 1606716760
transform 1 0 125856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1362
timestamp 1606716760
transform 1 0 125672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1366
timestamp 1606716760
transform 1 0 126040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1372
timestamp 1606716760
transform 1 0 126592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1374
timestamp 1606716760
transform 1 0 126776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[236\]
timestamp 1606716760
transform 1 0 125396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1352
timestamp 1606716760
transform 1 0 124752 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1354
timestamp 1606716760
transform 1 0 124936 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[33\]_TE
timestamp 1606716760
transform 1 0 124568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[282\]
timestamp 1606716760
transform 1 0 124660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1358
timestamp 1606716760
transform 1 0 125304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1606716760
transform 1 0 123832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1348
timestamp 1606716760
transform 1 0 124384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1344
timestamp 1606716760
transform 1 0 124016 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1343
timestamp 1606716760
transform 1 0 123924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[235\]
timestamp 1606716760
transform 1 0 124108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[242\]
timestamp 1606716760
transform 1 0 127420 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1606716760
transform 1 0 127328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1384
timestamp 1606716760
transform 1 0 127696 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1392
timestamp 1606716760
transform 1 0 128432 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[34\]_A
timestamp 1606716760
transform 1 0 126960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1378
timestamp 1606716760
transform 1 0 127144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[237\]
timestamp 1606716760
transform 1 0 125488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[34\]_TE
timestamp 1606716760
transform 1 0 125948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1363
timestamp 1606716760
transform 1 0 125764 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1367
timestamp 1606716760
transform 1 0 126132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1375
timestamp 1606716760
transform 1 0 126868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1359
timestamp 1606716760
transform 1 0 125396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1347
timestamp 1606716760
transform 1 0 124292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[234\]
timestamp 1606716760
transform 1 0 127788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[32\]_TE
timestamp 1606716760
transform 1 0 127420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1383
timestamp 1606716760
transform 1 0 127604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1388
timestamp 1606716760
transform 1 0 128064 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1377
timestamp 1606716760
transform 1 0 127052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[30\]
timestamp 1606716760
transform 1 0 125396 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1358
timestamp 1606716760
transform 1 0 125304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1606716760
transform 1 0 124476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1350
timestamp 1606716760
transform 1 0 124568 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[32\]
timestamp 1606716760
transform 1 0 127420 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1606716760
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1379
timestamp 1606716760
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[30\]_A
timestamp 1606716760
transform 1 0 126684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[30\]_TE
timestamp 1606716760
transform 1 0 125856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1362
timestamp 1606716760
transform 1 0 125672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1366
timestamp 1606716760
transform 1 0 126040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1372
timestamp 1606716760
transform 1 0 126592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1375
timestamp 1606716760
transform 1 0 126868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[232\]
timestamp 1606716760
transform 1 0 125396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1358
timestamp 1606716760
transform 1 0 125304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1354
timestamp 1606716760
transform 1 0 124936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1342
timestamp 1606716760
transform 1 0 123832 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1386
timestamp 1606716760
transform 1 0 127880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1362
timestamp 1606716760
transform 1 0 125672 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1374
timestamp 1606716760
transform 1 0 126776 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1606716760
transform 1 0 124476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1347
timestamp 1606716760
transform 1 0 124292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1350
timestamp 1606716760
transform 1 0 124568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _605_
timestamp 1606716760
transform 1 0 122820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[38\]_A
timestamp 1606716760
transform 1 0 122452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1325
timestamp 1606716760
transform 1 0 122268 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1329
timestamp 1606716760
transform 1 0 122636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1334
timestamp 1606716760
transform 1 0 123096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[38\]_TE
timestamp 1606716760
transform 1 0 121348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1313
timestamp 1606716760
transform 1 0 121164 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1317
timestamp 1606716760
transform 1 0 121532 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[79\]
timestamp 1606716760
transform 1 0 119508 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1287
timestamp 1606716760
transform 1 0 118772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__A
timestamp 1606716760
transform 1 0 123004 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1331
timestamp 1606716760
transform 1 0 122820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1335
timestamp 1606716760
transform 1 0 123188 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[38\]
timestamp 1606716760
transform 1 0 121164 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1606716760
transform 1 0 121072 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[79\]_A
timestamp 1606716760
transform 1 0 120796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1308
timestamp 1606716760
transform 1 0 120704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1311
timestamp 1606716760
transform 1 0 120980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[240\]
timestamp 1606716760
transform 1 0 120060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[79\]_TE
timestamp 1606716760
transform 1 0 119508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1293
timestamp 1606716760
transform 1 0 119324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1297
timestamp 1606716760
transform 1 0 119692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1304
timestamp 1606716760
transform 1 0 120336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[281\]
timestamp 1606716760
transform 1 0 119048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1289
timestamp 1606716760
transform 1 0 118956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1334
timestamp 1606716760
transform 1 0 123096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[36\]
timestamp 1606716760
transform 1 0 121440 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[31\]_TE
timestamp 1606716760
transform 1 0 121256 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1306
timestamp 1606716760
transform 1 0 120520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[28\]
timestamp 1606716760
transform 1 0 118864 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[233\]
timestamp 1606716760
transform 1 0 122268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[31\]_A
timestamp 1606716760
transform 1 0 123096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[36\]_A
timestamp 1606716760
transform 1 0 123464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1328
timestamp 1606716760
transform 1 0 122544 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1340
timestamp 1606716760
transform 1 0 123648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1332
timestamp 1606716760
transform 1 0 122912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1336
timestamp 1606716760
transform 1 0 123280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1340
timestamp 1606716760
transform 1 0 123648 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[31\]
timestamp 1606716760
transform 1 0 121256 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1606716760
transform 1 0 121072 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[36\]_TE
timestamp 1606716760
transform 1 0 120888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1317
timestamp 1606716760
transform 1 0 121532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1313
timestamp 1606716760
transform 1 0 121164 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[21\]
timestamp 1606716760
transform 1 0 119876 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[28\]_A
timestamp 1606716760
transform 1 0 120152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[28\]_TE
timestamp 1606716760
transform 1 0 119232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1294
timestamp 1606716760
transform 1 0 119416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1298
timestamp 1606716760
transform 1 0 119784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1294
timestamp 1606716760
transform 1 0 119416 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1304
timestamp 1606716760
transform 1 0 120336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[230\]
timestamp 1606716760
transform 1 0 118772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1290
timestamp 1606716760
transform 1 0 119048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1335
timestamp 1606716760
transform 1 0 123188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[227\]
timestamp 1606716760
transform 1 0 121808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1606716760
transform 1 0 121716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[21\]_A
timestamp 1606716760
transform 1 0 121164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1307
timestamp 1606716760
transform 1 0 120612 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1315
timestamp 1606716760
transform 1 0 121348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1323
timestamp 1606716760
transform 1 0 122084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[21\]_TE
timestamp 1606716760
transform 1 0 120428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[223\]
timestamp 1606716760
transform 1 0 119968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1292
timestamp 1606716760
transform 1 0 119232 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1303
timestamp 1606716760
transform 1 0 120244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[220\]
timestamp 1606716760
transform 1 0 118956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1288
timestamp 1606716760
transform 1 0 118864 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[22\]_A
timestamp 1606716760
transform 1 0 123188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1333
timestamp 1606716760
transform 1 0 123004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1337
timestamp 1606716760
transform 1 0 123372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[22\]
timestamp 1606716760
transform 1 0 121348 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1307
timestamp 1606716760
transform 1 0 120612 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[18\]
timestamp 1606716760
transform 1 0 118956 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1606716760
transform 1 0 118864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[29\]_A
timestamp 1606716760
transform 1 0 123648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1338
timestamp 1606716760
transform 1 0 123464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[29\]
timestamp 1606716760
transform 1 0 121808 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1606716760
transform 1 0 121716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[18\]_A
timestamp 1606716760
transform 1 0 120520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[22\]_TE
timestamp 1606716760
transform 1 0 121348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[29\]_TE
timestamp 1606716760
transform 1 0 120980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1308
timestamp 1606716760
transform 1 0 120704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1313
timestamp 1606716760
transform 1 0 121164 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1317
timestamp 1606716760
transform 1 0 121532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[224\]
timestamp 1606716760
transform 1 0 120060 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1291
timestamp 1606716760
transform 1 0 119140 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1299
timestamp 1606716760
transform 1 0 119876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1304
timestamp 1606716760
transform 1 0 120336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[18\]_TE
timestamp 1606716760
transform 1 0 118956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1288
timestamp 1606716760
transform 1 0 118864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[204\]
timestamp 1606716760
transform 1 0 123280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[2\]_TE
timestamp 1606716760
transform 1 0 122820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1328
timestamp 1606716760
transform 1 0 122544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1333
timestamp 1606716760
transform 1 0 123004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1339
timestamp 1606716760
transform 1 0 123556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[25\]
timestamp 1606716760
transform 1 0 120888 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1309
timestamp 1606716760
transform 1 0 120796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1301
timestamp 1606716760
transform 1 0 120060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1606716760
transform 1 0 118864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1287
timestamp 1606716760
transform 1 0 118772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1289
timestamp 1606716760
transform 1 0 118956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[290\]
timestamp 1606716760
transform 1 0 118496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1606716760
transform 1 0 118220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1279
timestamp 1606716760
transform 1 0 118036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1282
timestamp 1606716760
transform 1 0 118312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1271
timestamp 1606716760
transform 1 0 117300 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[77\]
timestamp 1606716760
transform 1 0 115644 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1245
timestamp 1606716760
transform 1 0 114908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[288\]
timestamp 1606716760
transform 1 0 117576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1277
timestamp 1606716760
transform 1 0 117852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[277\]
timestamp 1606716760
transform 1 0 116564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[77\]_A
timestamp 1606716760
transform 1 0 117024 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[77\]_TE
timestamp 1606716760
transform 1 0 116012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1255
timestamp 1606716760
transform 1 0 115828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1259
timestamp 1606716760
transform 1 0 116196 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1266
timestamp 1606716760
transform 1 0 116840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1270
timestamp 1606716760
transform 1 0 117208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[208\]
timestamp 1606716760
transform 1 0 115552 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1606716760
transform 1 0 115460 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[68\]_A
timestamp 1606716760
transform 1 0 114724 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[73\]_A
timestamp 1606716760
transform 1 0 115092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1241
timestamp 1606716760
transform 1 0 114540 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1245
timestamp 1606716760
transform 1 0 114908 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1249
timestamp 1606716760
transform 1 0 115276 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1606716760
transform 1 0 118220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1276
timestamp 1606716760
transform 1 0 117760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1280
timestamp 1606716760
transform 1 0 118128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1282
timestamp 1606716760
transform 1 0 118312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[222\]
timestamp 1606716760
transform 1 0 116380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[20\]_TE
timestamp 1606716760
transform 1 0 115828 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1253
timestamp 1606716760
transform 1 0 115644 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1257
timestamp 1606716760
transform 1 0 116012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1264
timestamp 1606716760
transform 1 0 116656 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[26\]
timestamp 1606716760
transform 1 0 113988 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1606716760
transform 1 0 118220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[20\]_A
timestamp 1606716760
transform 1 0 117392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1275
timestamp 1606716760
transform 1 0 117668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1282
timestamp 1606716760
transform 1 0 118312 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1274
timestamp 1606716760
transform 1 0 117576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1286
timestamp 1606716760
transform 1 0 118680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[216\]
timestamp 1606716760
transform 1 0 115920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[14\]_TE
timestamp 1606716760
transform 1 0 116380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1254
timestamp 1606716760
transform 1 0 115736 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1259
timestamp 1606716760
transform 1 0 116196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1263
timestamp 1606716760
transform 1 0 116564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1270
timestamp 1606716760
transform 1 0 117208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[279\]
timestamp 1606716760
transform 1 0 114356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[20\]
timestamp 1606716760
transform 1 0 115552 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1606716760
transform 1 0 115460 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[26\]_A
timestamp 1606716760
transform 1 0 115276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[26\]_TE
timestamp 1606716760
transform 1 0 114356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1242
timestamp 1606716760
transform 1 0 114632 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1241
timestamp 1606716760
transform 1 0 114540 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[228\]
timestamp 1606716760
transform 1 0 113896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1237
timestamp 1606716760
transform 1 0 114172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[14\]_A
timestamp 1606716760
transform 1 0 118128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1278
timestamp 1606716760
transform 1 0 117944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1282
timestamp 1606716760
transform 1 0 118312 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[14\]
timestamp 1606716760
transform 1 0 116288 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1606716760
transform 1 0 116104 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1259
timestamp 1606716760
transform 1 0 116196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1238
timestamp 1606716760
transform 1 0 114264 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1250
timestamp 1606716760
transform 1 0 115368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[17\]_A
timestamp 1606716760
transform 1 0 114080 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1234
timestamp 1606716760
transform 1 0 113896 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1272
timestamp 1606716760
transform 1 0 117392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1284
timestamp 1606716760
transform 1 0 118496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[27\]
timestamp 1606716760
transform 1 0 115736 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[13\]_A
timestamp 1606716760
transform 1 0 115184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1246
timestamp 1606716760
transform 1 0 115000 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1250
timestamp 1606716760
transform 1 0 115368 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1282
timestamp 1606716760
transform 1 0 118312 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1606716760
transform 1 0 116104 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[27\]_A
timestamp 1606716760
transform 1 0 117024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[27\]_TE
timestamp 1606716760
transform 1 0 115736 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1256
timestamp 1606716760
transform 1 0 115920 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1259
timestamp 1606716760
transform 1 0 116196 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1267
timestamp 1606716760
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1270
timestamp 1606716760
transform 1 0 117208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[125\]_A
timestamp 1606716760
transform 1 0 115276 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1247
timestamp 1606716760
transform 1 0 115092 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1251
timestamp 1606716760
transform 1 0 115460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1275
timestamp 1606716760
transform 1 0 117668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1263
timestamp 1606716760
transform 1 0 116564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[229\]
timestamp 1606716760
transform 1 0 115184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1243
timestamp 1606716760
transform 1 0 114724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1247
timestamp 1606716760
transform 1 0 115092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1251
timestamp 1606716760
transform 1 0 115460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[68\]
timestamp 1606716760
transform 1 0 113252 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1606716760
transform 1 0 112608 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[73\]_TE
timestamp 1606716760
transform 1 0 112884 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1221
timestamp 1606716760
transform 1 0 112700 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1225
timestamp 1606716760
transform 1 0 113068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[71\]_TE
timestamp 1606716760
transform 1 0 111872 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1210
timestamp 1606716760
transform 1 0 111688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1214
timestamp 1606716760
transform 1 0 112056 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[59\]
timestamp 1606716760
transform 1 0 110032 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1184
timestamp 1606716760
transform 1 0 109296 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[73\]
timestamp 1606716760
transform 1 0 112884 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1221
timestamp 1606716760
transform 1 0 112700 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[268\]
timestamp 1606716760
transform 1 0 110952 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[59\]_A
timestamp 1606716760
transform 1 0 111412 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1205
timestamp 1606716760
transform 1 0 111228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1209
timestamp 1606716760
transform 1 0 111596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[266\]
timestamp 1606716760
transform 1 0 109940 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1606716760
transform 1 0 109848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[59\]_TE
timestamp 1606716760
transform 1 0 110400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1194
timestamp 1606716760
transform 1 0 110216 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1198
timestamp 1606716760
transform 1 0 110584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[57\]_A
timestamp 1606716760
transform 1 0 108928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1182
timestamp 1606716760
transform 1 0 109112 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[270\]
timestamp 1606716760
transform 1 0 112792 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1606716760
transform 1 0 112608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[68\]_TE
timestamp 1606716760
transform 1 0 113252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1221
timestamp 1606716760
transform 1 0 112700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1225
timestamp 1606716760
transform 1 0 113068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1229
timestamp 1606716760
transform 1 0 113436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1219
timestamp 1606716760
transform 1 0 112516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[273\]
timestamp 1606716760
transform 1 0 111136 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_1201
timestamp 1606716760
transform 1 0 110860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1207
timestamp 1606716760
transform 1 0 111412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1189
timestamp 1606716760
transform 1 0 109756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[215\]
timestamp 1606716760
transform 1 0 113344 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1606716760
transform 1 0 112608 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1221
timestamp 1606716760
transform 1 0 112700 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1227
timestamp 1606716760
transform 1 0 113252 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1231
timestamp 1606716760
transform 1 0 113620 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1231
timestamp 1606716760
transform 1 0 113620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1218
timestamp 1606716760
transform 1 0 112424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1219
timestamp 1606716760
transform 1 0 112516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[275\]
timestamp 1606716760
transform 1 0 112240 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[17\]_TE
timestamp 1606716760
transform 1 0 112240 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1202
timestamp 1606716760
transform 1 0 110952 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1214
timestamp 1606716760
transform 1 0 112056 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1203
timestamp 1606716760
transform 1 0 111044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1215
timestamp 1606716760
transform 1 0 112148 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1606716760
transform 1 0 109848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1190
timestamp 1606716760
transform 1 0 109848 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1187
timestamp 1606716760
transform 1 0 109572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1191
timestamp 1606716760
transform 1 0 109940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[23\]_A
timestamp 1606716760
transform 1 0 109388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1183
timestamp 1606716760
transform 1 0 109204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[17\]
timestamp 1606716760
transform 1 0 112240 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1210
timestamp 1606716760
transform 1 0 111688 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1606716760
transform 1 0 110492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1188
timestamp 1606716760
transform 1 0 109664 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1196
timestamp 1606716760
transform 1 0 110400 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1198
timestamp 1606716760
transform 1 0 110584 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[13\]
timestamp 1606716760
transform 1 0 113344 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1606716760
transform 1 0 113252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1203
timestamp 1606716760
transform 1 0 111044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1215
timestamp 1606716760
transform 1 0 112148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1191
timestamp 1606716760
transform 1 0 109940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[125\]
timestamp 1606716760
transform 1 0 113436 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[13\]_TE
timestamp 1606716760
transform 1 0 113252 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[125\]_TE
timestamp 1606716760
transform 1 0 112884 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1222
timestamp 1606716760
transform 1 0 112792 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1225
timestamp 1606716760
transform 1 0 113068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1218
timestamp 1606716760
transform 1 0 112424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[219\]
timestamp 1606716760
transform 1 0 112148 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1210
timestamp 1606716760
transform 1 0 111688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1214
timestamp 1606716760
transform 1 0 112056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1606716760
transform 1 0 110492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1198
timestamp 1606716760
transform 1 0 110584 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1185
timestamp 1606716760
transform 1 0 109388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[327\]
timestamp 1606716760
transform 1 0 113344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1606716760
transform 1 0 113252 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1231
timestamp 1606716760
transform 1 0 113620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1203
timestamp 1606716760
transform 1 0 111044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1215
timestamp 1606716760
transform 1 0 112148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1191
timestamp 1606716760
transform 1 0 109940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[57\]
timestamp 1606716760
transform 1 0 107640 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1606716760
transform 1 0 106996 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1151
timestamp 1606716760
transform 1 0 106260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1160
timestamp 1606716760
transform 1 0 107088 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[53\]
timestamp 1606716760
transform 1 0 104604 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[261\]
timestamp 1606716760
transform 1 0 108100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1168
timestamp 1606716760
transform 1 0 107824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1174
timestamp 1606716760
transform 1 0 108376 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[57\]_TE
timestamp 1606716760
transform 1 0 107640 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[259\]
timestamp 1606716760
transform 1 0 106996 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1149
timestamp 1606716760
transform 1 0 106076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1157
timestamp 1606716760
transform 1 0 106812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1162
timestamp 1606716760
transform 1 0 107272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[53\]_A
timestamp 1606716760
transform 1 0 105892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1135
timestamp 1606716760
transform 1 0 104788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1606716760
transform 1 0 104236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[53\]_TE
timestamp 1606716760
transform 1 0 104604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_1130
timestamp 1606716760
transform 1 0 104328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[23\]
timestamp 1606716760
transform 1 0 108100 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_16_1168
timestamp 1606716760
transform 1 0 107824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1606716760
transform 1 0 106996 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1160
timestamp 1606716760
transform 1 0 107088 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1147
timestamp 1606716760
transform 1 0 105892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1135
timestamp 1606716760
transform 1 0 104788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[225\]
timestamp 1606716760
transform 1 0 107824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[23\]_TE
timestamp 1606716760
transform 1 0 108284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1178
timestamp 1606716760
transform 1 0 108744 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1171
timestamp 1606716760
transform 1 0 108100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1175
timestamp 1606716760
transform 1 0 108468 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[226\]
timestamp 1606716760
transform 1 0 106444 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[24\]
timestamp 1606716760
transform 1 0 107088 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1606716760
transform 1 0 106996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1158
timestamp 1606716760
transform 1 0 106904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1149
timestamp 1606716760
transform 1 0 106076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1156
timestamp 1606716760
transform 1 0 106720 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1146
timestamp 1606716760
transform 1 0 105800 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[19\]_A
timestamp 1606716760
transform 1 0 104788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1134
timestamp 1606716760
transform 1 0 104696 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1137
timestamp 1606716760
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[328\]
timestamp 1606716760
transform 1 0 104328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1606716760
transform 1 0 104236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1133
timestamp 1606716760
transform 1 0 104604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[24\]_A
timestamp 1606716760
transform 1 0 108376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1176
timestamp 1606716760
transform 1 0 108560 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[24\]_TE
timestamp 1606716760
transform 1 0 107088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1149
timestamp 1606716760
transform 1 0 106076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1157
timestamp 1606716760
transform 1 0 106812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1162
timestamp 1606716760
transform 1 0 107272 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1606716760
transform 1 0 104880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1137
timestamp 1606716760
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[1\]_A
timestamp 1606716760
transform 1 0 104328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1132
timestamp 1606716760
transform 1 0 104512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1167
timestamp 1606716760
transform 1 0 107732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1179
timestamp 1606716760
transform 1 0 108836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1606716760
transform 1 0 107640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1165
timestamp 1606716760
transform 1 0 107548 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1153
timestamp 1606716760
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1141
timestamp 1606716760
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1129
timestamp 1606716760
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1173
timestamp 1606716760
transform 1 0 108284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1149
timestamp 1606716760
transform 1 0 106076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1161
timestamp 1606716760
transform 1 0 107180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1606716760
transform 1 0 104880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1135
timestamp 1606716760
transform 1 0 104788 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1137
timestamp 1606716760
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1127
timestamp 1606716760
transform 1 0 104052 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1167
timestamp 1606716760
transform 1 0 107732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1179
timestamp 1606716760
transform 1 0 108836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1606716760
transform 1 0 107640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1164
timestamp 1606716760
transform 1 0 107456 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1156
timestamp 1606716760
transform 1 0 106720 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1144
timestamp 1606716760
transform 1 0 105616 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1132
timestamp 1606716760
transform 1 0 104512 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1125
timestamp 1606716760
transform 1 0 103868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[16\]
timestamp 1606716760
transform 1 0 102212 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1606716760
transform 1 0 101384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1099
timestamp 1606716760
transform 1 0 101476 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1095
timestamp 1606716760
transform 1 0 101108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1083
timestamp 1606716760
transform 1 0 100004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[217\]
timestamp 1606716760
transform 1 0 99728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[221\]
timestamp 1606716760
transform 1 0 103224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[16\]_A
timestamp 1606716760
transform 1 0 103684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1121
timestamp 1606716760
transform 1 0 103500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1125
timestamp 1606716760
transform 1 0 103868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[16\]_TE
timestamp 1606716760
transform 1 0 102672 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1114
timestamp 1606716760
transform 1 0 102856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[218\]
timestamp 1606716760
transform 1 0 102212 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[15\]_A
timestamp 1606716760
transform 1 0 101476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1097
timestamp 1606716760
transform 1 0 101292 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1101
timestamp 1606716760
transform 1 0 101660 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1110
timestamp 1606716760
transform 1 0 102488 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[15\]
timestamp 1606716760
transform 1 0 99636 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[15\]_TE
timestamp 1606716760
transform 1 0 99452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1073
timestamp 1606716760
transform 1 0 99084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[19\]
timestamp 1606716760
transform 1 0 103132 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1115
timestamp 1606716760
transform 1 0 102948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[255\]
timestamp 1606716760
transform 1 0 101568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1606716760
transform 1 0 101384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1096
timestamp 1606716760
transform 1 0 101200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1099
timestamp 1606716760
transform 1 0 101476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1103
timestamp 1606716760
transform 1 0 101844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1088
timestamp 1606716760
transform 1 0 100464 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[1\]
timestamp 1606716760
transform 1 0 103040 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[19\]_TE
timestamp 1606716760
transform 1 0 103316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1117
timestamp 1606716760
transform 1 0 103132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1121
timestamp 1606716760
transform 1 0 103500 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[203\]
timestamp 1606716760
transform 1 0 102856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1114
timestamp 1606716760
transform 1 0 102856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[324\]
timestamp 1606716760
transform 1 0 101476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1606716760
transform 1 0 101384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1096
timestamp 1606716760
transform 1 0 101200 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1102
timestamp 1606716760
transform 1 0 101752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1098
timestamp 1606716760
transform 1 0 101384 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1110
timestamp 1606716760
transform 1 0 102488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[323\]
timestamp 1606716760
transform 1 0 101108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[126\]_A
timestamp 1606716760
transform 1 0 100924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[121\]_A
timestamp 1606716760
transform 1 0 100556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[124\]_A
timestamp 1606716760
transform 1 0 100280 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1084
timestamp 1606716760
transform 1 0 100096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1088
timestamp 1606716760
transform 1 0 100464 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1087
timestamp 1606716760
transform 1 0 100372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1091
timestamp 1606716760
transform 1 0 100740 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[326\]
timestamp 1606716760
transform 1 0 103316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[1\]_TE
timestamp 1606716760
transform 1 0 103040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1115
timestamp 1606716760
transform 1 0 102948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1118
timestamp 1606716760
transform 1 0 103224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1122
timestamp 1606716760
transform 1 0 103592 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1111
timestamp 1606716760
transform 1 0 102580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[214\]
timestamp 1606716760
transform 1 0 102304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1606716760
transform 1 0 102028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[12\]
timestamp 1606716760
transform 1 0 102580 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1606716760
transform 1 0 102028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1108
timestamp 1606716760
transform 1 0 102304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[12\]_A
timestamp 1606716760
transform 1 0 103868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1115
timestamp 1606716760
transform 1 0 102948 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1123
timestamp 1606716760
transform 1 0 103684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[12\]_TE
timestamp 1606716760
transform 1 0 102764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1111
timestamp 1606716760
transform 1 0 102580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[329\]
timestamp 1606716760
transform 1 0 102304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606716760
transform 1 0 102028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1120
timestamp 1606716760
transform 1 0 103408 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606716760
transform 1 0 102028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1108
timestamp 1606716760
transform 1 0 102304 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1072
timestamp 1606716760
transform 1 0 98992 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[127\]
timestamp 1606716760
transform 1 0 97336 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1053
timestamp 1606716760
transform 1 0 97244 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[206\]
timestamp 1606716760
transform 1 0 95864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1041
timestamp 1606716760
transform 1 0 96140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1606716760
transform 1 0 95772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1035
timestamp 1606716760
transform 1 0 95588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[250\]
timestamp 1606716760
transform 1 0 94576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1020
timestamp 1606716760
transform 1 0 94208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1027
timestamp 1606716760
transform 1 0 94852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1606716760
transform 1 0 98624 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[127\]_A
timestamp 1606716760
transform 1 0 98900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[127\]_TE
timestamp 1606716760
transform 1 0 98256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1066
timestamp 1606716760
transform 1 0 98440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1069
timestamp 1606716760
transform 1 0 98716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[4\]_A
timestamp 1606716760
transform 1 0 97888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1058
timestamp 1606716760
transform 1 0 97704 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1062
timestamp 1606716760
transform 1 0 98072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[4\]
timestamp 1606716760
transform 1 0 96048 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[4\]_TE
timestamp 1606716760
transform 1 0 95864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1030
timestamp 1606716760
transform 1 0 95128 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[119\]_A
timestamp 1606716760
transform 1 0 94944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1026
timestamp 1606716760
transform 1 0 94760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[126\]
timestamp 1606716760
transform 1 0 98808 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1062
timestamp 1606716760
transform 1 0 98072 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[122\]
timestamp 1606716760
transform 1 0 96416 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1038
timestamp 1606716760
transform 1 0 95864 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1606716760
transform 1 0 95772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1035
timestamp 1606716760
transform 1 0 95588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[111\]_TE
timestamp 1606716760
transform 1 0 94300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1019
timestamp 1606716760
transform 1 0 94116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1023
timestamp 1606716760
transform 1 0 94484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[124\]
timestamp 1606716760
transform 1 0 98440 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[121\]
timestamp 1606716760
transform 1 0 98716 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[121\]_TE
timestamp 1606716760
transform 1 0 98440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1606716760
transform 1 0 98624 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[122\]_A
timestamp 1606716760
transform 1 0 97704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1058
timestamp 1606716760
transform 1 0 97704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[123\]_A
timestamp 1606716760
transform 1 0 97888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[126\]_TE
timestamp 1606716760
transform 1 0 98072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1062
timestamp 1606716760
transform 1 0 98072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1060
timestamp 1606716760
transform 1 0 97888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1064
timestamp 1606716760
transform 1 0 98256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[124\]_TE
timestamp 1606716760
transform 1 0 98256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[123\]
timestamp 1606716760
transform 1 0 96048 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__A
timestamp 1606716760
transform 1 0 97152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1050
timestamp 1606716760
transform 1 0 96968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1054
timestamp 1606716760
transform 1 0 97336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1043
timestamp 1606716760
transform 1 0 96324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1039
timestamp 1606716760
transform 1 0 95956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1038
timestamp 1606716760
transform 1 0 95864 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[111\]_A
timestamp 1606716760
transform 1 0 96140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _610_
timestamp 1606716760
transform 1 0 96692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[122\]_TE
timestamp 1606716760
transform 1 0 96508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1606716760
transform 1 0 95772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[123\]_TE
timestamp 1606716760
transform 1 0 95588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[111\]
timestamp 1606716760
transform 1 0 94300 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[117\]_A
timestamp 1606716760
transform 1 0 94668 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1023
timestamp 1606716760
transform 1 0 94484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1027
timestamp 1606716760
transform 1 0 94852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1019
timestamp 1606716760
transform 1 0 94116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[114\]_A
timestamp 1606716760
transform 1 0 94024 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1016
timestamp 1606716760
transform 1 0 93840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[114\]
timestamp 1606716760
transform 1 0 92184 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_18_996
timestamp 1606716760
transform 1 0 92000 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[213\]
timestamp 1606716760
transform 1 0 90988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_988
timestamp 1606716760
transform 1 0 91264 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[118\]_TE
timestamp 1606716760
transform 1 0 90436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_977
timestamp 1606716760
transform 1 0 90252 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_981
timestamp 1606716760
transform 1 0 90620 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1606716760
transform 1 0 90160 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[119\]
timestamp 1606716760
transform 1 0 93104 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1606716760
transform 1 0 93012 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[114\]_TE
timestamp 1606716760
transform 1 0 92644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1005
timestamp 1606716760
transform 1 0 92828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[118\]_A
timestamp 1606716760
transform 1 0 92276 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_997
timestamp 1606716760
transform 1 0 92092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1001
timestamp 1606716760
transform 1 0 92460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[118\]
timestamp 1606716760
transform 1 0 90436 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_17_977
timestamp 1606716760
transform 1 0 90252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[105\]_A
timestamp 1606716760
transform 1 0 89332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_969
timestamp 1606716760
transform 1 0 89516 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[319\]
timestamp 1606716760
transform 1 0 93840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1012
timestamp 1606716760
transform 1 0 93472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[119\]_TE
timestamp 1606716760
transform 1 0 93288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1008
timestamp 1606716760
transform 1 0 93104 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[116\]
timestamp 1606716760
transform 1 0 91448 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_16_988
timestamp 1606716760
transform 1 0 91264 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[309\]
timestamp 1606716760
transform 1 0 90252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_980
timestamp 1606716760
transform 1 0 90528 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1606716760
transform 1 0 90160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[102\]_TE
timestamp 1606716760
transform 1 0 89884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_966
timestamp 1606716760
transform 1 0 89240 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_972
timestamp 1606716760
transform 1 0 89792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_975
timestamp 1606716760
transform 1 0 90068 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1011
timestamp 1606716760
transform 1 0 93380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[117\]
timestamp 1606716760
transform 1 0 92828 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1006
timestamp 1606716760
transform 1 0 92920 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1003
timestamp 1606716760
transform 1 0 92644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1003
timestamp 1606716760
transform 1 0 92644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[116\]_A
timestamp 1606716760
transform 1 0 92736 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1606716760
transform 1 0 93012 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[316\]
timestamp 1606716760
transform 1 0 93104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_999
timestamp 1606716760
transform 1 0 92276 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_995
timestamp 1606716760
transform 1 0 91908 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_995
timestamp 1606716760
transform 1 0 91908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[116\]_TE
timestamp 1606716760
transform 1 0 92092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[102\]_A
timestamp 1606716760
transform 1 0 91724 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_991
timestamp 1606716760
transform 1 0 91540 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[106\]
timestamp 1606716760
transform 1 0 90252 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[102\]
timestamp 1606716760
transform 1 0 89884 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1606716760
transform 1 0 90160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[100\]_A
timestamp 1606716760
transform 1 0 89332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[107\]_TE
timestamp 1606716760
transform 1 0 89884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_967
timestamp 1606716760
transform 1 0 89332 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_975
timestamp 1606716760
transform 1 0 90068 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_969
timestamp 1606716760
transform 1 0 89516 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606716760
transform -1 0 93012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[106\]_A
timestamp 1606716760
transform 1 0 91724 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[117\]_TE
timestamp 1606716760
transform 1 0 92552 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_995
timestamp 1606716760
transform 1 0 91908 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1001
timestamp 1606716760
transform 1 0 92460 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_991
timestamp 1606716760
transform 1 0 91540 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[107\]
timestamp 1606716760
transform 1 0 89884 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[101\]_A
timestamp 1606716760
transform 1 0 89332 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[104\]_A
timestamp 1606716760
transform 1 0 89700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_969
timestamp 1606716760
transform 1 0 89516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606716760
transform -1 0 93012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[313\]
timestamp 1606716760
transform 1 0 91724 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_996
timestamp 1606716760
transform 1 0 92000 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[107\]_A
timestamp 1606716760
transform 1 0 91172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_989
timestamp 1606716760
transform 1 0 91356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[106\]_TE
timestamp 1606716760
transform 1 0 90436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_977
timestamp 1606716760
transform 1 0 90252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_981
timestamp 1606716760
transform 1 0 90620 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1606716760
transform 1 0 90160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[10\]_A
timestamp 1606716760
transform 1 0 89608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_968
timestamp 1606716760
transform 1 0 89424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_972
timestamp 1606716760
transform 1 0 89792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606716760
transform -1 0 93012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[325\]
timestamp 1606716760
transform 1 0 91724 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_996
timestamp 1606716760
transform 1 0 92000 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_990
timestamp 1606716760
transform 1 0 91448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_978
timestamp 1606716760
transform 1 0 90344 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[108\]_A
timestamp 1606716760
transform 1 0 90160 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_974
timestamp 1606716760
transform 1 0 89976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606716760
transform -1 0 93012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1003
timestamp 1606716760
transform 1 0 92644 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_995
timestamp 1606716760
transform 1 0 91908 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[112\]
timestamp 1606716760
transform 1 0 90252 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1606716760
transform 1 0 90160 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_966
timestamp 1606716760
transform 1 0 89240 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_974
timestamp 1606716760
transform 1 0 89976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[8\]_A
timestamp 1606716760
transform 1 0 88872 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_960
timestamp 1606716760
transform 1 0 88688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_964
timestamp 1606716760
transform 1 0 89056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[8\]
timestamp 1606716760
transform 1 0 87032 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[8\]_TE
timestamp 1606716760
transform 1 0 86848 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[88\]_A
timestamp 1606716760
transform 1 0 86480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_934
timestamp 1606716760
transform 1 0 86296 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_938
timestamp 1606716760
transform 1 0 86664 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[88\]
timestamp 1606716760
transform 1 0 84640 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1606716760
transform 1 0 84548 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_965
timestamp 1606716760
transform 1 0 89148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[105\]
timestamp 1606716760
transform 1 0 87492 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1606716760
transform 1 0 87400 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[0\]_A
timestamp 1606716760
transform 1 0 86848 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[105\]_TE
timestamp 1606716760
transform 1 0 87216 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_942
timestamp 1606716760
transform 1 0 87032 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_938
timestamp 1606716760
transform 1 0 86664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[0\]
timestamp 1606716760
transform 1 0 85008 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[88\]_TE
timestamp 1606716760
transform 1 0 84640 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_915
timestamp 1606716760
transform 1 0 84548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_918
timestamp 1606716760
transform 1 0 84824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[304\]
timestamp 1606716760
transform 1 0 88964 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_959
timestamp 1606716760
transform 1 0 88596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[103\]_A
timestamp 1606716760
transform 1 0 88412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_955
timestamp 1606716760
transform 1 0 88228 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[103\]
timestamp 1606716760
transform 1 0 86572 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_16_934
timestamp 1606716760
transform 1 0 86296 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1606716760
transform 1 0 84548 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[0\]_TE
timestamp 1606716760
transform 1 0 85008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_912
timestamp 1606716760
transform 1 0 84272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_916
timestamp 1606716760
transform 1 0 84640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_922
timestamp 1606716760
transform 1 0 85192 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_965
timestamp 1606716760
transform 1 0 89148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[104\]
timestamp 1606716760
transform 1 0 87676 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[100\]
timestamp 1606716760
transform 1 0 87492 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_15_942
timestamp 1606716760
transform 1 0 87032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_941
timestamp 1606716760
transform 1 0 86940 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[103\]_TE
timestamp 1606716760
transform 1 0 86848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[101\]_TE
timestamp 1606716760
transform 1 0 87492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[100\]_TE
timestamp 1606716760
transform 1 0 87216 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1606716760
transform 1 0 87400 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_938
timestamp 1606716760
transform 1 0 86664 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[306\]
timestamp 1606716760
transform 1 0 86664 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[302\]
timestamp 1606716760
transform 1 0 86388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[308\]
timestamp 1606716760
transform 1 0 85652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_930
timestamp 1606716760
transform 1 0 85928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_927
timestamp 1606716760
transform 1 0 85652 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[307\]
timestamp 1606716760
transform 1 0 85376 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1606716760
transform 1 0 84548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_916
timestamp 1606716760
transform 1 0 84640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_924
timestamp 1606716760
transform 1 0 85376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_913
timestamp 1606716760
transform 1 0 84364 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_921
timestamp 1606716760
transform 1 0 85100 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_965
timestamp 1606716760
transform 1 0 89148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[101\]
timestamp 1606716760
transform 1 0 87492 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1606716760
transform 1 0 87400 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[104\]_TE
timestamp 1606716760
transform 1 0 87216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[303\]
timestamp 1606716760
transform 1 0 86388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_933
timestamp 1606716760
transform 1 0 86204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_938
timestamp 1606716760
transform 1 0 86664 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_925
timestamp 1606716760
transform 1 0 85468 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[16\]_A
timestamp 1606716760
transform 1 0 85284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_921
timestamp 1606716760
transform 1 0 85100 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[10\]
timestamp 1606716760
transform 1 0 87768 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_942
timestamp 1606716760
transform 1 0 87032 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[310\]
timestamp 1606716760
transform 1 0 86756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_936
timestamp 1606716760
transform 1 0 86480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_928
timestamp 1606716760
transform 1 0 85744 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1606716760
transform 1 0 84548 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_913
timestamp 1606716760
transform 1 0 84364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_916
timestamp 1606716760
transform 1 0 84640 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[108\]
timestamp 1606716760
transform 1 0 88320 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[10\]_TE
timestamp 1606716760
transform 1 0 87768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[108\]_TE
timestamp 1606716760
transform 1 0 88136 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_952
timestamp 1606716760
transform 1 0 87952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1606716760
transform 1 0 87400 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_944
timestamp 1606716760
transform 1 0 87216 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_947
timestamp 1606716760
transform 1 0 87492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_932
timestamp 1606716760
transform 1 0 86112 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_920
timestamp 1606716760
transform 1 0 85008 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[314\]
timestamp 1606716760
transform 1 0 88964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[212\]
timestamp 1606716760
transform 1 0 87952 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_955
timestamp 1606716760
transform 1 0 88228 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[109\]_TE
timestamp 1606716760
transform 1 0 87492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_949
timestamp 1606716760
transform 1 0 87676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[311\]
timestamp 1606716760
transform 1 0 86480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_939
timestamp 1606716760
transform 1 0 86756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_928
timestamp 1606716760
transform 1 0 85744 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1606716760
transform 1 0 84548 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_916
timestamp 1606716760
transform 1 0 84640 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_907
timestamp 1606716760
transform 1 0 83812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _562_
timestamp 1606716760
transform 1 0 83536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1606716760
transform 1 0 82984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_896
timestamp 1606716760
transform 1 0 82800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_900
timestamp 1606716760
transform 1 0 83168 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _553_
timestamp 1606716760
transform 1 0 82524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_885
timestamp 1606716760
transform 1 0 81788 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[82\]
timestamp 1606716760
transform 1 0 80132 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_858
timestamp 1606716760
transform 1 0 79304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_866
timestamp 1606716760
transform 1 0 80040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[162\]
timestamp 1606716760
transform 1 0 83904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_906
timestamp 1606716760
transform 1 0 83720 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_911
timestamp 1606716760
transform 1 0 84180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _566_
timestamp 1606716760
transform 1 0 82892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A
timestamp 1606716760
transform 1 0 83536 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_900
timestamp 1606716760
transform 1 0 83168 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__A
timestamp 1606716760
transform 1 0 82340 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__553__A
timestamp 1606716760
transform 1 0 82708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_889
timestamp 1606716760
transform 1 0 82156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_893
timestamp 1606716760
transform 1 0 82524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _551_
timestamp 1606716760
transform 1 0 81880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1606716760
transform 1 0 81788 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[82\]_A
timestamp 1606716760
transform 1 0 81420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_880
timestamp 1606716760
transform 1 0 81328 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_883
timestamp 1606716760
transform 1 0 81604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1606716760
transform 1 0 80776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_876
timestamp 1606716760
transform 1 0 80960 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_872
timestamp 1606716760
transform 1 0 80592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[82\]_TE
timestamp 1606716760
transform 1 0 80132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _544_
timestamp 1606716760
transform 1 0 80316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_865
timestamp 1606716760
transform 1 0 79948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A
timestamp 1606716760
transform 1 0 79764 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_861
timestamp 1606716760
transform 1 0 79580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _539_
timestamp 1606716760
transform 1 0 79304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _570_
timestamp 1606716760
transform 1 0 82892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_900
timestamp 1606716760
transform 1 0 83168 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_889
timestamp 1606716760
transform 1 0 82156 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _564_
timestamp 1606716760
transform 1 0 81880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_884
timestamp 1606716760
transform 1 0 81696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _550_
timestamp 1606716760
transform 1 0 80684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_876
timestamp 1606716760
transform 1 0 80960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[156\]
timestamp 1606716760
transform 1 0 79672 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_861
timestamp 1606716760
transform 1 0 79580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_865
timestamp 1606716760
transform 1 0 79948 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[16\]_TE
timestamp 1606716760
transform 1 0 83812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_909
timestamp 1606716760
transform 1 0 83996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__A
timestamp 1606716760
transform 1 0 83076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_905
timestamp 1606716760
transform 1 0 83628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_897
timestamp 1606716760
transform 1 0 82892 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_901
timestamp 1606716760
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[40\]
timestamp 1606716760
transform 1 0 81972 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_15_893
timestamp 1606716760
transform 1 0 82524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_889
timestamp 1606716760
transform 1 0 82156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A
timestamp 1606716760
transform 1 0 82708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1606716760
transform 1 0 82340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_883
timestamp 1606716760
transform 1 0 81604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_886
timestamp 1606716760
transform 1 0 81880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_882
timestamp 1606716760
transform 1 0 81512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1606716760
transform 1 0 81788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _568_
timestamp 1606716760
transform 1 0 81880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_870
timestamp 1606716760
transform 1 0 80408 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_869
timestamp 1606716760
transform 1 0 80316 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_875
timestamp 1606716760
transform 1 0 80868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__A
timestamp 1606716760
transform 1 0 80684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[30\]_TE
timestamp 1606716760
transform 1 0 79488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_858
timestamp 1606716760
transform 1 0 79304 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_862
timestamp 1606716760
transform 1 0 79672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[158\]
timestamp 1606716760
transform 1 0 80040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[160\]
timestamp 1606716760
transform 1 0 80132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_866
timestamp 1606716760
transform 1 0 80040 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_864
timestamp 1606716760
transform 1 0 79856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[16\]
timestamp 1606716760
transform 1 0 83444 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[40\]_A
timestamp 1606716760
transform 1 0 83260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[40\]_TE
timestamp 1606716760
transform 1 0 82340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_889
timestamp 1606716760
transform 1 0 82156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_893
timestamp 1606716760
transform 1 0 82524 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[114\]
timestamp 1606716760
transform 1 0 81880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1606716760
transform 1 0 81788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[30\]_A
timestamp 1606716760
transform 1 0 81236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_877
timestamp 1606716760
transform 1 0 81052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_881
timestamp 1606716760
transform 1 0 81420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[30\]
timestamp 1606716760
transform 1 0 79396 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[90\]
timestamp 1606716760
transform 1 0 83352 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_900
timestamp 1606716760
transform 1 0 83168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_905
timestamp 1606716760
transform 1 0 83628 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_888
timestamp 1606716760
transform 1 0 82064 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[33\]_TE
timestamp 1606716760
transform 1 0 81880 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_881
timestamp 1606716760
transform 1 0 81420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_885
timestamp 1606716760
transform 1 0 81788 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  la_buf\[31\]
timestamp 1606716760
transform 1 0 79764 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[33\]_A
timestamp 1606716760
transform 1 0 83720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_908
timestamp 1606716760
transform 1 0 83904 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_904
timestamp 1606716760
transform 1 0 83536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[33\]
timestamp 1606716760
transform 1 0 81880 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1606716760
transform 1 0 81788 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[31\]_A
timestamp 1606716760
transform 1 0 81052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_879
timestamp 1606716760
transform 1 0 81236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_876
timestamp 1606716760
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[105\]
timestamp 1606716760
transform 1 0 79580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[31\]_TE
timestamp 1606716760
transform 1 0 80040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_864
timestamp 1606716760
transform 1 0 79856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_868
timestamp 1606716760
transform 1 0 80224 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_907
timestamp 1606716760
transform 1 0 83812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_895
timestamp 1606716760
transform 1 0 82708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[107\]
timestamp 1606716760
transform 1 0 81328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_879
timestamp 1606716760
transform 1 0 81236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_883
timestamp 1606716760
transform 1 0 81604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_867
timestamp 1606716760
transform 1 0 80132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _535_
timestamp 1606716760
transform 1 0 79028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1606716760
transform 1 0 78936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__A
timestamp 1606716760
transform 1 0 78292 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_842
timestamp 1606716760
transform 1 0 77832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_846
timestamp 1606716760
transform 1 0 78200 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_849
timestamp 1606716760
transform 1 0 78476 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_853
timestamp 1606716760
transform 1 0 78844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  la_buf\[91\]
timestamp 1606716760
transform 1 0 76176 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_18_822
timestamp 1606716760
transform 1 0 75992 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _522_
timestamp 1606716760
transform 1 0 74980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[95\]_B
timestamp 1606716760
transform 1 0 74428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_807
timestamp 1606716760
transform 1 0 74612 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_814
timestamp 1606716760
transform 1 0 75256 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_857
timestamp 1606716760
transform 1 0 79212 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_854
timestamp 1606716760
transform 1 0 78936 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__A
timestamp 1606716760
transform 1 0 79028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _537_
timestamp 1606716760
transform 1 0 78292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[91\]_A
timestamp 1606716760
transform 1 0 78108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_843
timestamp 1606716760
transform 1 0 77924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_850
timestamp 1606716760
transform 1 0 78568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _533_
timestamp 1606716760
transform 1 0 77280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__A
timestamp 1606716760
transform 1 0 77740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_839
timestamp 1606716760
transform 1 0 77556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _530_
timestamp 1606716760
transform 1 0 76268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1606716760
transform 1 0 76176 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__A
timestamp 1606716760
transform 1 0 76728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_828
timestamp 1606716760
transform 1 0 76544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_832
timestamp 1606716760
transform 1 0 76912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[91\]_TE
timestamp 1606716760
transform 1 0 75992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[91\]_A
timestamp 1606716760
transform 1 0 74796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[95\]_A
timestamp 1606716760
transform 1 0 75164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A
timestamp 1606716760
transform 1 0 75532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_807
timestamp 1606716760
transform 1 0 74612 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_811
timestamp 1606716760
transform 1 0 74980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_815
timestamp 1606716760
transform 1 0 75348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_819
timestamp 1606716760
transform 1 0 75716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1606716760
transform 1 0 78936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_855
timestamp 1606716760
transform 1 0 79028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_853
timestamp 1606716760
transform 1 0 78844 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_841
timestamp 1606716760
transform 1 0 77740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _531_
timestamp 1606716760
transform 1 0 76360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_829
timestamp 1606716760
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_823
timestamp 1606716760
transform 1 0 76084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_811
timestamp 1606716760
transform 1 0 74980 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_856
timestamp 1606716760
transform 1 0 79120 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1606716760
transform 1 0 78936 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[104\]
timestamp 1606716760
transform 1 0 79028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_844
timestamp 1606716760
transform 1 0 78016 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_852
timestamp 1606716760
transform 1 0 78752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_844
timestamp 1606716760
transform 1 0 78016 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[165\]
timestamp 1606716760
transform 1 0 76268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1606716760
transform 1 0 76176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__531__A
timestamp 1606716760
transform 1 0 76728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_832
timestamp 1606716760
transform 1 0 76912 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_828
timestamp 1606716760
transform 1 0 76544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_832
timestamp 1606716760
transform 1 0 76912 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_823
timestamp 1606716760
transform 1 0 76084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_820
timestamp 1606716760
transform 1 0 75808 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_808
timestamp 1606716760
transform 1 0 74704 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_817
timestamp 1606716760
transform 1 0 75532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_813
timestamp 1606716760
transform 1 0 75164 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[99\]_A
timestamp 1606716760
transform 1 0 75348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_806
timestamp 1606716760
transform 1 0 74520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[429\]
timestamp 1606716760
transform 1 0 74428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[427\]
timestamp 1606716760
transform 1 0 74888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_857
timestamp 1606716760
transform 1 0 79212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_849
timestamp 1606716760
transform 1 0 78476 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_837
timestamp 1606716760
transform 1 0 77372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1606716760
transform 1 0 76176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_825
timestamp 1606716760
transform 1 0 76268 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_822
timestamp 1606716760
transform 1 0 75992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_810
timestamp 1606716760
transform 1 0 74888 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1606716760
transform 1 0 78936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_855
timestamp 1606716760
transform 1 0 79028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_842
timestamp 1606716760
transform 1 0 77832 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_830
timestamp 1606716760
transform 1 0 76728 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_806
timestamp 1606716760
transform 1 0 74520 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_818
timestamp 1606716760
transform 1 0 75624 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_849
timestamp 1606716760
transform 1 0 78476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_837
timestamp 1606716760
transform 1 0 77372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1606716760
transform 1 0 76176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_825
timestamp 1606716760
transform 1 0 76268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_812
timestamp 1606716760
transform 1 0 75072 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1606716760
transform 1 0 78936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_855
timestamp 1606716760
transform 1 0 79028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_842
timestamp 1606716760
transform 1 0 77832 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_830
timestamp 1606716760
transform 1 0 76728 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_806
timestamp 1606716760
transform 1 0 74520 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_818
timestamp 1606716760
transform 1 0 75624 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_803
timestamp 1606716760
transform 1 0 74244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[91\]
timestamp 1606716760
transform 1 0 73416 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1606716760
transform 1 0 73324 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[8\]_B
timestamp 1606716760
transform 1 0 72404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_785
timestamp 1606716760
transform 1 0 72588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[88\]_B
timestamp 1606716760
transform 1 0 72036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_777
timestamp 1606716760
transform 1 0 71852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_781
timestamp 1606716760
transform 1 0 72220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[73\]
timestamp 1606716760
transform 1 0 70196 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_751
timestamp 1606716760
transform 1 0 69460 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[95\]
timestamp 1606716760
transform 1 0 73784 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[8\]_A
timestamp 1606716760
transform 1 0 73232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[91\]_B
timestamp 1606716760
transform 1 0 73600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_790
timestamp 1606716760
transform 1 0 73048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_794
timestamp 1606716760
transform 1 0 73416 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[8\]
timestamp 1606716760
transform 1 0 72220 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[86\]_A
timestamp 1606716760
transform 1 0 71668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[73\]_A
timestamp 1606716760
transform 1 0 72036 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_773
timestamp 1606716760
transform 1 0 71484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_777
timestamp 1606716760
transform 1 0 71852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[86\]
timestamp 1606716760
transform 1 0 70656 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1606716760
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[73\]_TE
timestamp 1606716760
transform 1 0 70196 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_752
timestamp 1606716760
transform 1 0 69552 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_758
timestamp 1606716760
transform 1 0 70104 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_761
timestamp 1606716760
transform 1 0 70380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[99\]
timestamp 1606716760
transform 1 0 74152 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1606716760
transform 1 0 73324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_794
timestamp 1606716760
transform 1 0 73416 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_785
timestamp 1606716760
transform 1 0 72588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[145\]
timestamp 1606716760
transform 1 0 72312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[418\]
timestamp 1606716760
transform 1 0 71208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_773
timestamp 1606716760
transform 1 0 71484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_781
timestamp 1606716760
transform 1 0 72220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[416\]
timestamp 1606716760
transform 1 0 70196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[86\]_B
timestamp 1606716760
transform 1 0 70840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_751
timestamp 1606716760
transform 1 0 69460 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_762
timestamp 1606716760
transform 1 0 70472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_768
timestamp 1606716760
transform 1 0 71024 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_802
timestamp 1606716760
transform 1 0 74152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[99\]_B
timestamp 1606716760
transform 1 0 74336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[423\]
timestamp 1606716760
transform 1 0 73876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[425\]
timestamp 1606716760
transform 1 0 73416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1606716760
transform 1 0 73324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_791
timestamp 1606716760
transform 1 0 73140 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_797
timestamp 1606716760
transform 1 0 73692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_791
timestamp 1606716760
transform 1 0 73140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[421\]
timestamp 1606716760
transform 1 0 72864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[106\]
timestamp 1606716760
transform 1 0 71760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[338\]
timestamp 1606716760
transform 1 0 71852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_775
timestamp 1606716760
transform 1 0 71668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_779
timestamp 1606716760
transform 1 0 72036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_776
timestamp 1606716760
transform 1 0 71760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_780
timestamp 1606716760
transform 1 0 72128 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_769
timestamp 1606716760
transform 1 0 71116 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1606716760
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_757
timestamp 1606716760
transform 1 0 70012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_751
timestamp 1606716760
transform 1 0 69460 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_764
timestamp 1606716760
transform 1 0 70656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[32\]_A
timestamp 1606716760
transform 1 0 73600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_794
timestamp 1606716760
transform 1 0 73416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_798
timestamp 1606716760
transform 1 0 73784 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[32\]
timestamp 1606716760
transform 1 0 71760 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[32\]_TE
timestamp 1606716760
transform 1 0 71576 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_772
timestamp 1606716760
transform 1 0 71392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1606716760
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_759
timestamp 1606716760
transform 1 0 70196 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_764
timestamp 1606716760
transform 1 0 70656 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1606716760
transform 1 0 73324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_792
timestamp 1606716760
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_794
timestamp 1606716760
transform 1 0 73416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_786
timestamp 1606716760
transform 1 0 72680 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_774
timestamp 1606716760
transform 1 0 71576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_762
timestamp 1606716760
transform 1 0 70472 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_800
timestamp 1606716760
transform 1 0 73968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_788
timestamp 1606716760
transform 1 0 72864 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_776
timestamp 1606716760
transform 1 0 71760 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[101\]
timestamp 1606716760
transform 1 0 69552 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1606716760
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[2\]_A
timestamp 1606716760
transform 1 0 70104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_755
timestamp 1606716760
transform 1 0 69828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_760
timestamp 1606716760
transform 1 0 70288 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_764
timestamp 1606716760
transform 1 0 70656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1606716760
transform 1 0 73324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_792
timestamp 1606716760
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_794
timestamp 1606716760
transform 1 0 73416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_786
timestamp 1606716760
transform 1 0 72680 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_774
timestamp 1606716760
transform 1 0 71576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[27\]
timestamp 1606716760
transform 1 0 69920 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_10_753
timestamp 1606716760
transform 1 0 69644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[82\]
timestamp 1606716760
transform 1 0 68632 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_741
timestamp 1606716760
transform 1 0 68540 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1606716760
transform 1 0 67712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_731
timestamp 1606716760
transform 1 0 67620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_733
timestamp 1606716760
transform 1 0 67804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_719
timestamp 1606716760
transform 1 0 66516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[93\]
timestamp 1606716760
transform 1 0 64860 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_18_698
timestamp 1606716760
transform 1 0 64584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[82\]_A
timestamp 1606716760
transform 1 0 69368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[409\]
timestamp 1606716760
transform 1 0 68908 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[82\]_B
timestamp 1606716760
transform 1 0 68724 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_741
timestamp 1606716760
transform 1 0 68540 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_748
timestamp 1606716760
transform 1 0 69184 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_717
timestamp 1606716760
transform 1 0 66332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_729
timestamp 1606716760
transform 1 0 67436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1606716760
transform 1 0 64952 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[93\]_A
timestamp 1606716760
transform 1 0 66148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[93\]_TE
timestamp 1606716760
transform 1 0 65228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_703
timestamp 1606716760
transform 1 0 65044 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_707
timestamp 1606716760
transform 1 0 65412 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[414\]
timestamp 1606716760
transform 1 0 69184 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_745
timestamp 1606716760
transform 1 0 68908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1606716760
transform 1 0 67712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_733
timestamp 1606716760
transform 1 0 67804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_721
timestamp 1606716760
transform 1 0 66700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_729
timestamp 1606716760
transform 1 0 67436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_709
timestamp 1606716760
transform 1 0 65596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_745
timestamp 1606716760
transform 1 0 68908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_739
timestamp 1606716760
transform 1 0 68356 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1606716760
transform 1 0 67712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_733
timestamp 1606716760
transform 1 0 67804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_720
timestamp 1606716760
transform 1 0 66608 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_727
timestamp 1606716760
transform 1 0 67252 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[377\]
timestamp 1606716760
transform 1 0 65228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1606716760
transform 1 0 64952 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_708
timestamp 1606716760
transform 1 0 65504 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_701
timestamp 1606716760
transform 1 0 64860 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_703
timestamp 1606716760
transform 1 0 65044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_715
timestamp 1606716760
transform 1 0 66148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[76\]
timestamp 1606716760
transform 1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_739
timestamp 1606716760
transform 1 0 68356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_743
timestamp 1606716760
transform 1 0 68724 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_747
timestamp 1606716760
transform 1 0 69092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_727
timestamp 1606716760
transform 1 0 67252 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1606716760
transform 1 0 64952 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_701
timestamp 1606716760
transform 1 0 64860 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_703
timestamp 1606716760
transform 1 0 65044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_715
timestamp 1606716760
transform 1 0 66148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[2\]
timestamp 1606716760
transform 1 0 68816 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_12_741
timestamp 1606716760
transform 1 0 68540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1606716760
transform 1 0 67712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_733
timestamp 1606716760
transform 1 0 67804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_720
timestamp 1606716760
transform 1 0 66608 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_708
timestamp 1606716760
transform 1 0 65504 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[2\]_TE
timestamp 1606716760
transform 1 0 68816 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_742
timestamp 1606716760
transform 1 0 68632 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_746
timestamp 1606716760
transform 1 0 69000 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_718
timestamp 1606716760
transform 1 0 66424 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_730
timestamp 1606716760
transform 1 0 67528 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[198\]
timestamp 1606716760
transform 1 0 65044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1606716760
transform 1 0 64952 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_701
timestamp 1606716760
transform 1 0 64860 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_706
timestamp 1606716760
transform 1 0 65320 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_745
timestamp 1606716760
transform 1 0 68908 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1606716760
transform 1 0 67712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_731
timestamp 1606716760
transform 1 0 67620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_733
timestamp 1606716760
transform 1 0 67804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_727
timestamp 1606716760
transform 1 0 67252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_715
timestamp 1606716760
transform 1 0 66148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[390\]
timestamp 1606716760
transform 1 0 63204 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_686
timestamp 1606716760
transform 1 0 63480 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[389\]
timestamp 1606716760
transform 1 0 62192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1606716760
transform 1 0 62100 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[75\]_B
timestamp 1606716760
transform 1 0 61548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_667
timestamp 1606716760
transform 1 0 61732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_675
timestamp 1606716760
transform 1 0 62468 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_663
timestamp 1606716760
transform 1 0 61364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[375\]
timestamp 1606716760
transform 1 0 61088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[64\]_B
timestamp 1606716760
transform 1 0 60536 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_652
timestamp 1606716760
transform 1 0 60352 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_656
timestamp 1606716760
transform 1 0 60720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_684
timestamp 1606716760
transform 1 0 63296 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_696
timestamp 1606716760
transform 1 0 64400 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[403\]
timestamp 1606716760
transform 1 0 63020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[376\]
timestamp 1606716760
transform 1 0 62008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_673
timestamp 1606716760
transform 1 0 62284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[374\]
timestamp 1606716760
transform 1 0 60996 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[46\]_A
timestamp 1606716760
transform 1 0 60444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[64\]_A
timestamp 1606716760
transform 1 0 60812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_651
timestamp 1606716760
transform 1 0 60260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_655
timestamp 1606716760
transform 1 0 60628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_662
timestamp 1606716760
transform 1 0 61272 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[405\]
timestamp 1606716760
transform 1 0 63204 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[80\]
timestamp 1606716760
transform 1 0 64216 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_686
timestamp 1606716760
transform 1 0 63480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_697
timestamp 1606716760
transform 1 0 64492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[392\]
timestamp 1606716760
transform 1 0 62192 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1606716760
transform 1 0 62100 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_670
timestamp 1606716760
transform 1 0 62008 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_675
timestamp 1606716760
transform 1 0 62468 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[373\]
timestamp 1606716760
transform 1 0 60628 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_647
timestamp 1606716760
transform 1 0 59892 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_658
timestamp 1606716760
transform 1 0 60904 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[47\]
timestamp 1606716760
transform 1 0 63112 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[47\]_A
timestamp 1606716760
transform 1 0 64124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_697
timestamp 1606716760
transform 1 0 64492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_691
timestamp 1606716760
transform 1 0 63940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_695
timestamp 1606716760
transform 1 0 64308 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  la_buf\[46\]
timestamp 1606716760
transform 1 0 62836 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[47\]_B
timestamp 1606716760
transform 1 0 62928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_679
timestamp 1606716760
transform 1 0 62836 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[372\]
timestamp 1606716760
transform 1 0 61456 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1606716760
transform 1 0 62100 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_669
timestamp 1606716760
transform 1 0 61916 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_672
timestamp 1606716760
transform 1 0 62192 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_678
timestamp 1606716760
transform 1 0 62744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_667
timestamp 1606716760
transform 1 0 61732 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[369\]
timestamp 1606716760
transform 1 0 60444 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[39\]
timestamp 1606716760
transform 1 0 59892 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[44\]_A
timestamp 1606716760
transform 1 0 59892 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[126\]_TE
timestamp 1606716760
transform 1 0 60996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_656
timestamp 1606716760
transform 1 0 60720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_661
timestamp 1606716760
transform 1 0 61180 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_649
timestamp 1606716760
transform 1 0 60076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_656
timestamp 1606716760
transform 1 0 60720 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_645
timestamp 1606716760
transform 1 0 59708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[120\]
timestamp 1606716760
transform 1 0 63388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[46\]_A
timestamp 1606716760
transform 1 0 64124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[46\]_TE
timestamp 1606716760
transform 1 0 63204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_688
timestamp 1606716760
transform 1 0 63664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_692
timestamp 1606716760
transform 1 0 64032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_695
timestamp 1606716760
transform 1 0 64308 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[126\]_A
timestamp 1606716760
transform 1 0 62836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_681
timestamp 1606716760
transform 1 0 63020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_677
timestamp 1606716760
transform 1 0 62652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[126\]
timestamp 1606716760
transform 1 0 60996 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[39\]_A
timestamp 1606716760
transform 1 0 60536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[39\]_B
timestamp 1606716760
transform 1 0 60076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_651
timestamp 1606716760
transform 1 0 60260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_656
timestamp 1606716760
transform 1 0 60720 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_645
timestamp 1606716760
transform 1 0 59708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_684
timestamp 1606716760
transform 1 0 63296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_696
timestamp 1606716760
transform 1 0 64400 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1606716760
transform 1 0 62100 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_669
timestamp 1606716760
transform 1 0 61916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_672
timestamp 1606716760
transform 1 0 62192 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[200\]
timestamp 1606716760
transform 1 0 60904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[29\]_TE
timestamp 1606716760
transform 1 0 60260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_649
timestamp 1606716760
transform 1 0 60076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_653
timestamp 1606716760
transform 1 0 60444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_657
timestamp 1606716760
transform 1 0 60812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_661
timestamp 1606716760
transform 1 0 61180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_693
timestamp 1606716760
transform 1 0 64124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_681
timestamp 1606716760
transform 1 0 63020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[29\]_A
timestamp 1606716760
transform 1 0 61732 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_665
timestamp 1606716760
transform 1 0 61548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_669
timestamp 1606716760
transform 1 0 61916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[29\]
timestamp 1606716760
transform 1 0 59892 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[34\]_A
timestamp 1606716760
transform 1 0 59708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[124\]
timestamp 1606716760
transform 1 0 64492 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_10_684
timestamp 1606716760
transform 1 0 63296 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_696
timestamp 1606716760
transform 1 0 64400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1606716760
transform 1 0 62100 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_664
timestamp 1606716760
transform 1 0 61456 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_670
timestamp 1606716760
transform 1 0 62008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_672
timestamp 1606716760
transform 1 0 62192 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[103\]
timestamp 1606716760
transform 1 0 60076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_652
timestamp 1606716760
transform 1 0 60352 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[64\]
timestamp 1606716760
transform 1 0 59524 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_635
timestamp 1606716760
transform 1 0 58788 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[6\]
timestamp 1606716760
transform 1 0 57132 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1606716760
transform 1 0 56488 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_611
timestamp 1606716760
transform 1 0 56580 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[32\]
timestamp 1606716760
transform 1 0 54924 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[33\]_B
timestamp 1606716760
transform 1 0 55936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[60\]_B
timestamp 1606716760
transform 1 0 56304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_602
timestamp 1606716760
transform 1 0 55752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_606
timestamp 1606716760
transform 1 0 56120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_592
timestamp 1606716760
transform 1 0 54832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[46\]
timestamp 1606716760
transform 1 0 59432 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1606716760
transform 1 0 59340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[6\]_A
timestamp 1606716760
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[46\]_B
timestamp 1606716760
transform 1 0 59156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[6\]_TE
timestamp 1606716760
transform 1 0 58788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_633
timestamp 1606716760
transform 1 0 58604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_637
timestamp 1606716760
transform 1 0 58972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_627
timestamp 1606716760
transform 1 0 58052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[45\]
timestamp 1606716760
transform 1 0 56856 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[33\]_A
timestamp 1606716760
transform 1 0 56672 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[45\]_A
timestamp 1606716760
transform 1 0 57868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_623
timestamp 1606716760
transform 1 0 57684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_610
timestamp 1606716760
transform 1 0 56488 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[33\]
timestamp 1606716760
transform 1 0 55292 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[32\]_A
timestamp 1606716760
transform 1 0 56304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[32\]_B
timestamp 1606716760
transform 1 0 55108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_606
timestamp 1606716760
transform 1 0 56120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[44\]
timestamp 1606716760
transform 1 0 59064 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[43\]_A
timestamp 1606716760
transform 1 0 58512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_630
timestamp 1606716760
transform 1 0 58328 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_634
timestamp 1606716760
transform 1 0 58696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[43\]
timestamp 1606716760
transform 1 0 57500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[40\]_B
timestamp 1606716760
transform 1 0 56764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[45\]_B
timestamp 1606716760
transform 1 0 57132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_615
timestamp 1606716760
transform 1 0 56948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_619
timestamp 1606716760
transform 1 0 57316 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1606716760
transform 1 0 56488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_609
timestamp 1606716760
transform 1 0 56396 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_611
timestamp 1606716760
transform 1 0 56580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_601
timestamp 1606716760
transform 1 0 55660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[31\]
timestamp 1606716760
transform 1 0 54832 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[6\]_B
timestamp 1606716760
transform 1 0 54648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[37\]
timestamp 1606716760
transform 1 0 58328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[367\]
timestamp 1606716760
transform 1 0 59432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1606716760
transform 1 0 59340 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[37\]_B
timestamp 1606716760
transform 1 0 59340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[44\]_B
timestamp 1606716760
transform 1 0 59156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_639
timestamp 1606716760
transform 1 0 59156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_643
timestamp 1606716760
transform 1 0 59524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_637
timestamp 1606716760
transform 1 0 58972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[42\]_A
timestamp 1606716760
transform 1 0 58788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_628
timestamp 1606716760
transform 1 0 58144 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_633
timestamp 1606716760
transform 1 0 58604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[38\]
timestamp 1606716760
transform 1 0 56580 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[42\]
timestamp 1606716760
transform 1 0 57776 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_620
timestamp 1606716760
transform 1 0 57408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_624
timestamp 1606716760
transform 1 0 57776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_620
timestamp 1606716760
transform 1 0 57408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[43\]_B
timestamp 1606716760
transform 1 0 57960 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[42\]_B
timestamp 1606716760
transform 1 0 57592 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[38\]_A
timestamp 1606716760
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1606716760
transform 1 0 56488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_609
timestamp 1606716760
transform 1 0 56396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_616
timestamp 1606716760
transform 1 0 57040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[40\]_A
timestamp 1606716760
transform 1 0 57224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[3\]
timestamp 1606716760
transform 1 0 54832 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[40\]
timestamp 1606716760
transform 1 0 56212 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_601
timestamp 1606716760
transform 1 0 55660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_601
timestamp 1606716760
transform 1 0 55660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[3\]_B
timestamp 1606716760
transform 1 0 55844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[31\]_B
timestamp 1606716760
transform 1 0 55844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_605
timestamp 1606716760
transform 1 0 56028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_605
timestamp 1606716760
transform 1 0 56028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_592
timestamp 1606716760
transform 1 0 54832 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[31\]_A
timestamp 1606716760
transform 1 0 55476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[6\]_A
timestamp 1606716760
transform 1 0 55016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_596
timestamp 1606716760
transform 1 0 55200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[108\]
timestamp 1606716760
transform 1 0 59432 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1606716760
transform 1 0 59340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[37\]_A
timestamp 1606716760
transform 1 0 58972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_633
timestamp 1606716760
transform 1 0 58604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_639
timestamp 1606716760
transform 1 0 59156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[44\]
timestamp 1606716760
transform 1 0 56948 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[44\]_TE
timestamp 1606716760
transform 1 0 56764 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[38\]_B
timestamp 1606716760
transform 1 0 56396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_611
timestamp 1606716760
transform 1 0 56580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[118\]
timestamp 1606716760
transform 1 0 55936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[35\]_A
timestamp 1606716760
transform 1 0 55200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[3\]_A
timestamp 1606716760
transform 1 0 55568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_594
timestamp 1606716760
transform 1 0 55016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_598
timestamp 1606716760
transform 1 0 55384 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_602
timestamp 1606716760
transform 1 0 55752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_607
timestamp 1606716760
transform 1 0 56212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[34\]
timestamp 1606716760
transform 1 0 58420 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[44\]_A
timestamp 1606716760
transform 1 0 58236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_628
timestamp 1606716760
transform 1 0 58144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[34\]_B
timestamp 1606716760
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_620
timestamp 1606716760
transform 1 0 57408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_624
timestamp 1606716760
transform 1 0 57776 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[41\]
timestamp 1606716760
transform 1 0 56580 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1606716760
transform 1 0 56488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_595
timestamp 1606716760
transform 1 0 55108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_607
timestamp 1606716760
transform 1 0 56212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[333\]
timestamp 1606716760
transform 1 0 54832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1606716760
transform 1 0 59340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[34\]_A
timestamp 1606716760
transform 1 0 58420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[34\]_TE
timestamp 1606716760
transform 1 0 58788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_629
timestamp 1606716760
transform 1 0 58236 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_633
timestamp 1606716760
transform 1 0 58604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_637
timestamp 1606716760
transform 1 0 58972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_642
timestamp 1606716760
transform 1 0 59432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[34\]
timestamp 1606716760
transform 1 0 57408 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[41\]_A
timestamp 1606716760
transform 1 0 57224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[41\]_B
timestamp 1606716760
transform 1 0 56856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_612
timestamp 1606716760
transform 1 0 56672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_616
timestamp 1606716760
transform 1 0 57040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[196\]
timestamp 1606716760
transform 1 0 56396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[368\]
timestamp 1606716760
transform 1 0 55384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_601
timestamp 1606716760
transform 1 0 55660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_590
timestamp 1606716760
transform 1 0 54648 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_641
timestamp 1606716760
transform 1 0 59340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[122\]
timestamp 1606716760
transform 1 0 57684 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[364\]
timestamp 1606716760
transform 1 0 56672 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_615
timestamp 1606716760
transform 1 0 56948 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1606716760
transform 1 0 56488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_611
timestamp 1606716760
transform 1 0 56580 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[370\]
timestamp 1606716760
transform 1 0 55476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_597
timestamp 1606716760
transform 1 0 55292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_602
timestamp 1606716760
transform 1 0 55752 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_576
timestamp 1606716760
transform 1 0 53360 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_588
timestamp 1606716760
transform 1 0 54464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[28\]
timestamp 1606716760
transform 1 0 52532 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[25\]_B
timestamp 1606716760
transform 1 0 51980 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_563
timestamp 1606716760
transform 1 0 52164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_559
timestamp 1606716760
transform 1 0 51796 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[22\]
timestamp 1606716760
transform 1 0 50968 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1606716760
transform 1 0 50876 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_541
timestamp 1606716760
transform 1 0 50140 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[21\]_B
timestamp 1606716760
transform 1 0 49956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[361\]
timestamp 1606716760
transform 1 0 54280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1606716760
transform 1 0 53728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[28\]_B
timestamp 1606716760
transform 1 0 53544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_576
timestamp 1606716760
transform 1 0 53360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_581
timestamp 1606716760
transform 1 0 53820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_585
timestamp 1606716760
transform 1 0 54188 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_589
timestamp 1606716760
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[28\]_A
timestamp 1606716760
transform 1 0 53176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[22\]_A
timestamp 1606716760
transform 1 0 52348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[25\]_A
timestamp 1606716760
transform 1 0 52716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_563
timestamp 1606716760
transform 1 0 52164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_567
timestamp 1606716760
transform 1 0 52532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_571
timestamp 1606716760
transform 1 0 52900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[25\]
timestamp 1606716760
transform 1 0 51336 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[21\]_A
timestamp 1606716760
transform 1 0 50784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[22\]_B
timestamp 1606716760
transform 1 0 51152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_546
timestamp 1606716760
transform 1 0 50600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_550
timestamp 1606716760
transform 1 0 50968 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[21\]
timestamp 1606716760
transform 1 0 49772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[71\]
timestamp 1606716760
transform 1 0 53268 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[71\]_A
timestamp 1606716760
transform 1 0 54280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_584
timestamp 1606716760
transform 1 0 54096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_588
timestamp 1606716760
transform 1 0 54464 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_571
timestamp 1606716760
transform 1 0 52900 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_559
timestamp 1606716760
transform 1 0 51796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[24\]
timestamp 1606716760
transform 1 0 50968 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1606716760
transform 1 0 50876 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_548
timestamp 1606716760
transform 1 0 50784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[351\]
timestamp 1606716760
transform 1 0 49772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_540
timestamp 1606716760
transform 1 0 50048 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[6\]
timestamp 1606716760
transform 1 0 54004 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_589
timestamp 1606716760
transform 1 0 54556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[35\]_B
timestamp 1606716760
transform 1 0 54372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_581
timestamp 1606716760
transform 1 0 53820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_579
timestamp 1606716760
transform 1 0 53636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1606716760
transform 1 0 53820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[71\]_B
timestamp 1606716760
transform 1 0 53452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1606716760
transform 1 0 53728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[356\]
timestamp 1606716760
transform 1 0 53544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[26\]
timestamp 1606716760
transform 1 0 51980 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_571
timestamp 1606716760
transform 1 0 52900 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_570
timestamp 1606716760
transform 1 0 52808 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[24\]_A
timestamp 1606716760
transform 1 0 52440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[353\]
timestamp 1606716760
transform 1 0 52624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[27\]_B
timestamp 1606716760
transform 1 0 51520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_558
timestamp 1606716760
transform 1 0 51704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_564
timestamp 1606716760
transform 1 0 52256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_560
timestamp 1606716760
transform 1 0 51888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[23\]_A
timestamp 1606716760
transform 1 0 52072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_537
timestamp 1606716760
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[23\]
timestamp 1606716760
transform 1 0 51060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[355\]
timestamp 1606716760
transform 1 0 50968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1606716760
transform 1 0 50876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[23\]_B
timestamp 1606716760
transform 1 0 50876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_547
timestamp 1606716760
transform 1 0 50692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_553
timestamp 1606716760
transform 1 0 51244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_537
timestamp 1606716760
transform 1 0 49772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[352\]
timestamp 1606716760
transform 1 0 50048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[24\]_B
timestamp 1606716760
transform 1 0 50508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_543
timestamp 1606716760
transform 1 0 50324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[35\]
timestamp 1606716760
transform 1 0 54188 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1606716760
transform 1 0 53728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_581
timestamp 1606716760
transform 1 0 53820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_574
timestamp 1606716760
transform 1 0 53176 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[26\]_A
timestamp 1606716760
transform 1 0 52624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[26\]_B
timestamp 1606716760
transform 1 0 52992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_563
timestamp 1606716760
transform 1 0 52164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_567
timestamp 1606716760
transform 1 0 52532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_570
timestamp 1606716760
transform 1 0 52808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[27\]
timestamp 1606716760
transform 1 0 51336 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_543
timestamp 1606716760
transform 1 0 50324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_551
timestamp 1606716760
transform 1 0 51060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[354\]
timestamp 1606716760
transform 1 0 50048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[20\]_A
timestamp 1606716760
transform 1 0 49864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[365\]
timestamp 1606716760
transform 1 0 53820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_584
timestamp 1606716760
transform 1 0 54096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[396\]
timestamp 1606716760
transform 1 0 52808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[27\]_A
timestamp 1606716760
transform 1 0 51980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_563
timestamp 1606716760
transform 1 0 52164 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_569
timestamp 1606716760
transform 1 0 52716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_573
timestamp 1606716760
transform 1 0 53084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_557
timestamp 1606716760
transform 1 0 51612 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[357\]
timestamp 1606716760
transform 1 0 50968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1606716760
transform 1 0 50876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[30\]_B
timestamp 1606716760
transform 1 0 51428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_546
timestamp 1606716760
transform 1 0 50600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_553
timestamp 1606716760
transform 1 0 51244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[371\]
timestamp 1606716760
transform 1 0 54372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1606716760
transform 1 0 53728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_575
timestamp 1606716760
transform 1 0 53268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_579
timestamp 1606716760
transform 1 0 53636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_581
timestamp 1606716760
transform 1 0 53820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[30\]_A
timestamp 1606716760
transform 1 0 51980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_563
timestamp 1606716760
transform 1 0 52164 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_559
timestamp 1606716760
transform 1 0 51796 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[30\]
timestamp 1606716760
transform 1 0 50968 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_542
timestamp 1606716760
transform 1 0 50232 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[360\]
timestamp 1606716760
transform 1 0 49956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[398\]
timestamp 1606716760
transform 1 0 53912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_579
timestamp 1606716760
transform 1 0 53636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_585
timestamp 1606716760
transform 1 0 54188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_571
timestamp 1606716760
transform 1 0 52900 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[15\]
timestamp 1606716760
transform 1 0 51244 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1606716760
transform 1 0 50876 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_546
timestamp 1606716760
transform 1 0 50600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_550
timestamp 1606716760
transform 1 0 50968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_535
timestamp 1606716760
transform 1 0 49588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[66\]
timestamp 1606716760
transform 1 0 47932 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[53\]_B
timestamp 1606716760
transform 1 0 47380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_509
timestamp 1606716760
transform 1 0 47196 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_513
timestamp 1606716760
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[381\]
timestamp 1606716760
transform 1 0 45356 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[53\]
timestamp 1606716760
transform 1 0 46368 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[126\]_B
timestamp 1606716760
transform 1 0 46000 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_492
timestamp 1606716760
transform 1 0 45632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_498
timestamp 1606716760
transform 1 0 46184 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1606716760
transform 1 0 45264 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[16\]_A
timestamp 1606716760
transform 1 0 49220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[66\]_A
timestamp 1606716760
transform 1 0 49588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_529
timestamp 1606716760
transform 1 0 49036 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_533
timestamp 1606716760
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[16\]
timestamp 1606716760
transform 1 0 48208 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1606716760
transform 1 0 48116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[53\]_A
timestamp 1606716760
transform 1 0 47196 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[66\]_TE
timestamp 1606716760
transform 1 0 47932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_511
timestamp 1606716760
transform 1 0 47380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[126\]_A
timestamp 1606716760
transform 1 0 46828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_503
timestamp 1606716760
transform 1 0 46644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_507
timestamp 1606716760
transform 1 0 47012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[126\]
timestamp 1606716760
transform 1 0 45816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_490
timestamp 1606716760
transform 1 0 45448 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[16\]_B
timestamp 1606716760
transform 1 0 48484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_525
timestamp 1606716760
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_521
timestamp 1606716760
transform 1 0 48300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[346\]
timestamp 1606716760
transform 1 0 48024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_510
timestamp 1606716760
transform 1 0 47288 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[17\]
timestamp 1606716760
transform 1 0 46460 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1606716760
transform 1 0 45356 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1606716760
transform 1 0 45264 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_487
timestamp 1606716760
transform 1 0 45172 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[350\]
timestamp 1606716760
transform 1 0 48392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[20\]
timestamp 1606716760
transform 1 0 48576 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[20\]_B
timestamp 1606716760
transform 1 0 49588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_533
timestamp 1606716760
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_525
timestamp 1606716760
transform 1 0 48668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_506
timestamp 1606716760
transform 1 0 46920 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_520
timestamp 1606716760
transform 1 0 48208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_518
timestamp 1606716760
transform 1 0 48024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_514
timestamp 1606716760
transform 1 0 47656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_518
timestamp 1606716760
transform 1 0 48024 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[17\]_B
timestamp 1606716760
transform 1 0 47472 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1606716760
transform 1 0 48116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_507
timestamp 1606716760
transform 1 0 47012 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_503
timestamp 1606716760
transform 1 0 46644 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[201\]
timestamp 1606716760
transform 1 0 46644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_510
timestamp 1606716760
transform 1 0 47288 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[17\]_A
timestamp 1606716760
transform 1 0 47104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[347\]
timestamp 1606716760
transform 1 0 46368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[35\]_TE
timestamp 1606716760
transform 1 0 45724 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_489
timestamp 1606716760
transform 1 0 45356 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_495
timestamp 1606716760
transform 1 0 45908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_496
timestamp 1606716760
transform 1 0 46000 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1606716760
transform 1 0 45264 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_485
timestamp 1606716760
transform 1 0 44988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_484
timestamp 1606716760
transform 1 0 44896 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[14\]
timestamp 1606716760
transform 1 0 48484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[14\]_A
timestamp 1606716760
transform 1 0 49496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_532
timestamp 1606716760
transform 1 0 49312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_536
timestamp 1606716760
transform 1 0 49680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1606716760
transform 1 0 48116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[35\]_A
timestamp 1606716760
transform 1 0 47564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_511
timestamp 1606716760
transform 1 0 47380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_515
timestamp 1606716760
transform 1 0 47748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_520
timestamp 1606716760
transform 1 0 48208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[35\]
timestamp 1606716760
transform 1 0 45724 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_13_492
timestamp 1606716760
transform 1 0 45632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_486
timestamp 1606716760
transform 1 0 45080 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[344\]
timestamp 1606716760
transform 1 0 49220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[14\]_B
timestamp 1606716760
transform 1 0 48668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_523
timestamp 1606716760
transform 1 0 48484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_527
timestamp 1606716760
transform 1 0 48852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_534
timestamp 1606716760
transform 1 0 49496 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[127\]
timestamp 1606716760
transform 1 0 46828 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[109\]
timestamp 1606716760
transform 1 0 45816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_489
timestamp 1606716760
transform 1 0 45356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_493
timestamp 1606716760
transform 1 0 45724 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_497
timestamp 1606716760
transform 1 0 46092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1606716760
transform 1 0 45264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[2\]_B
timestamp 1606716760
transform 1 0 44896 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_486
timestamp 1606716760
transform 1 0 45080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[127\]_A
timestamp 1606716760
transform 1 0 48392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_524
timestamp 1606716760
transform 1 0 48576 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_536
timestamp 1606716760
transform 1 0 49680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1606716760
transform 1 0 48116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_520
timestamp 1606716760
transform 1 0 48208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[127\]_TE
timestamp 1606716760
transform 1 0 46828 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_502
timestamp 1606716760
transform 1 0 46552 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_507
timestamp 1606716760
transform 1 0 47012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[191\]
timestamp 1606716760
transform 1 0 46276 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[2\]_A
timestamp 1606716760
transform 1 0 45724 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_491
timestamp 1606716760
transform 1 0 45540 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_495
timestamp 1606716760
transform 1 0 45908 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_522
timestamp 1606716760
transform 1 0 48392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_534
timestamp 1606716760
transform 1 0 49496 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_510
timestamp 1606716760
transform 1 0 47288 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[117\]
timestamp 1606716760
transform 1 0 45632 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_10_489
timestamp 1606716760
transform 1 0 45356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1606716760
transform 1 0 45264 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_487
timestamp 1606716760
transform 1 0 45172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[456\]
timestamp 1606716760
transform 1 0 44252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_473
timestamp 1606716760
transform 1 0 43884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_480
timestamp 1606716760
transform 1 0 44528 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_461
timestamp 1606716760
transform 1 0 42780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[75\]
timestamp 1606716760
transform 1 0 41124 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_18_440
timestamp 1606716760
transform 1 0 40848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_478
timestamp 1606716760
transform 1 0 44344 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[349\]
timestamp 1606716760
transform 1 0 42596 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1606716760
transform 1 0 42504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[75\]_A
timestamp 1606716760
transform 1 0 43056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_456
timestamp 1606716760
transform 1 0 42320 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_462
timestamp 1606716760
transform 1 0 42872 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_466
timestamp 1606716760
transform 1 0 43240 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_448
timestamp 1606716760
transform 1 0 41584 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[95\]_A
timestamp 1606716760
transform 1 0 41032 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[75\]_TE
timestamp 1606716760
transform 1 0 41400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_440
timestamp 1606716760
transform 1 0 40848 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_444
timestamp 1606716760
transform 1 0 41216 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[95\]
timestamp 1606716760
transform 1 0 40020 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_475
timestamp 1606716760
transform 1 0 44068 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[1\]_B
timestamp 1606716760
transform 1 0 42780 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_458
timestamp 1606716760
transform 1 0 42504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_463
timestamp 1606716760
transform 1 0 42964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[13\]
timestamp 1606716760
transform 1 0 41676 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[19\]_B
timestamp 1606716760
transform 1 0 41124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_441
timestamp 1606716760
transform 1 0 40940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_445
timestamp 1606716760
transform 1 0 41308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[19\]
timestamp 1606716760
transform 1 0 40112 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[1\]_A
timestamp 1606716760
transform 1 0 43608 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_473
timestamp 1606716760
transform 1 0 43884 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_472
timestamp 1606716760
transform 1 0 43792 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_468
timestamp 1606716760
transform 1 0 43424 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[331\]
timestamp 1606716760
transform 1 0 42504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[1\]
timestamp 1606716760
transform 1 0 42596 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1606716760
transform 1 0 42504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[13\]_A
timestamp 1606716760
transform 1 0 42320 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_461
timestamp 1606716760
transform 1 0 42780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_453
timestamp 1606716760
transform 1 0 42044 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_448
timestamp 1606716760
transform 1 0 41584 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_450
timestamp 1606716760
transform 1 0 41768 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[13\]_B
timestamp 1606716760
transform 1 0 41860 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[19\]_A
timestamp 1606716760
transform 1 0 41400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[343\]
timestamp 1606716760
transform 1 0 41492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_444
timestamp 1606716760
transform 1 0 41216 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_440
timestamp 1606716760
transform 1 0 40848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_445
timestamp 1606716760
transform 1 0 41308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_437
timestamp 1606716760
transform 1 0 40572 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[18\]_A
timestamp 1606716760
transform 1 0 41032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[18\]
timestamp 1606716760
transform 1 0 40020 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[18\]_B
timestamp 1606716760
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_474
timestamp 1606716760
transform 1 0 43976 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[348\]
timestamp 1606716760
transform 1 0 42596 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1606716760
transform 1 0 42504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_457
timestamp 1606716760
transform 1 0 42412 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_462
timestamp 1606716760
transform 1 0 42872 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_449
timestamp 1606716760
transform 1 0 41676 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[342\]
timestamp 1606716760
transform 1 0 41400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[12\]_A
timestamp 1606716760
transform 1 0 40848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[15\]_A
timestamp 1606716760
transform 1 0 41216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_438
timestamp 1606716760
transform 1 0 40664 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_442
timestamp 1606716760
transform 1 0 41032 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[12\]
timestamp 1606716760
transform 1 0 39836 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[332\]
timestamp 1606716760
transform 1 0 44252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_476
timestamp 1606716760
transform 1 0 44160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_480
timestamp 1606716760
transform 1 0 44528 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[359\]
timestamp 1606716760
transform 1 0 42412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[29\]_B
timestamp 1606716760
transform 1 0 42872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_456
timestamp 1606716760
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_460
timestamp 1606716760
transform 1 0 42688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_464
timestamp 1606716760
transform 1 0 43056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[42\]_A
timestamp 1606716760
transform 1 0 41584 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_450
timestamp 1606716760
transform 1 0 41768 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_446
timestamp 1606716760
transform 1 0 41400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[2\]
timestamp 1606716760
transform 1 0 44712 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[29\]_A
timestamp 1606716760
transform 1 0 43608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_472
timestamp 1606716760
transform 1 0 43792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_480
timestamp 1606716760
transform 1 0 44528 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_468
timestamp 1606716760
transform 1 0 43424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[29\]
timestamp 1606716760
transform 1 0 42596 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1606716760
transform 1 0 42504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_457
timestamp 1606716760
transform 1 0 42412 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[10\]_A
timestamp 1606716760
transform 1 0 41676 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_451
timestamp 1606716760
transform 1 0 41860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_447
timestamp 1606716760
transform 1 0 41492 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[42\]
timestamp 1606716760
transform 1 0 39836 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_10_479
timestamp 1606716760
transform 1 0 44436 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_467
timestamp 1606716760
transform 1 0 43332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[25\]
timestamp 1606716760
transform 1 0 41676 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_10_443
timestamp 1606716760
transform 1 0 41124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_431
timestamp 1606716760
transform 1 0 40020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1606716760
transform 1 0 39652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_425
timestamp 1606716760
transform 1 0 39468 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_428
timestamp 1606716760
transform 1 0 39744 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[171\]
timestamp 1606716760
transform 1 0 38456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_417
timestamp 1606716760
transform 1 0 38732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[97\]_TE
timestamp 1606716760
transform 1 0 37904 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_406
timestamp 1606716760
transform 1 0 37720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_410
timestamp 1606716760
transform 1 0 38088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[79\]
timestamp 1606716760
transform 1 0 36064 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[121\]_B
timestamp 1606716760
transform 1 0 35512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_380
timestamp 1606716760
transform 1 0 35328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_384
timestamp 1606716760
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[97\]_A
timestamp 1606716760
transform 1 0 39468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_423
timestamp 1606716760
transform 1 0 39284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_427
timestamp 1606716760
transform 1 0 39652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[97\]
timestamp 1606716760
transform 1 0 37628 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_17_404
timestamp 1606716760
transform 1 0 37536 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1606716760
transform 1 0 36892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[79\]_A
timestamp 1606716760
transform 1 0 37352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_398
timestamp 1606716760
transform 1 0 36984 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[121\]_A
timestamp 1606716760
transform 1 0 35788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[79\]_TE
timestamp 1606716760
transform 1 0 36156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_387
timestamp 1606716760
transform 1 0 35972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_391
timestamp 1606716760
transform 1 0 36340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_383
timestamp 1606716760
transform 1 0 35604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1606716760
transform 1 0 39652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[93\]_A
timestamp 1606716760
transform 1 0 38916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_421
timestamp 1606716760
transform 1 0 39100 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_428
timestamp 1606716760
transform 1 0 39744 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_417
timestamp 1606716760
transform 1 0 38732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[8\]
timestamp 1606716760
transform 1 0 37904 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_400
timestamp 1606716760
transform 1 0 37168 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[84\]
timestamp 1606716760
transform 1 0 36340 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_388
timestamp 1606716760
transform 1 0 36064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_376
timestamp 1606716760
transform 1 0 34960 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[15\]
timestamp 1606716760
transform 1 0 39744 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1606716760
transform 1 0 39652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[8\]_A
timestamp 1606716760
transform 1 0 39100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_419
timestamp 1606716760
transform 1 0 38916 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_419
timestamp 1606716760
transform 1 0 38916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_423
timestamp 1606716760
transform 1 0 39284 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[345\]
timestamp 1606716760
transform 1 0 38640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_415
timestamp 1606716760
transform 1 0 38548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[93\]
timestamp 1606716760
transform 1 0 38088 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[124\]_A
timestamp 1606716760
transform 1 0 37628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_403
timestamp 1606716760
transform 1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_407
timestamp 1606716760
transform 1 0 37812 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_409
timestamp 1606716760
transform 1 0 37996 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[153\]
timestamp 1606716760
transform 1 0 36984 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1606716760
transform 1 0 36892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[84\]_A
timestamp 1606716760
transform 1 0 36708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_401
timestamp 1606716760
transform 1 0 37260 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[124\]
timestamp 1606716760
transform 1 0 36616 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_391
timestamp 1606716760
transform 1 0 36340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_391
timestamp 1606716760
transform 1 0 36340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[451\]
timestamp 1606716760
transform 1 0 34960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_383
timestamp 1606716760
transform 1 0 35604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1606716760
transform 1 0 35236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[18\]_A
timestamp 1606716760
transform 1 0 38916 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[12\]_B
timestamp 1606716760
transform 1 0 39652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[15\]_B
timestamp 1606716760
transform 1 0 39284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_421
timestamp 1606716760
transform 1 0 39100 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_425
timestamp 1606716760
transform 1 0 39468 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_417
timestamp 1606716760
transform 1 0 38732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[18\]
timestamp 1606716760
transform 1 0 37076 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1606716760
transform 1 0 36892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[124\]_B
timestamp 1606716760
transform 1 0 36708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_398
timestamp 1606716760
transform 1 0 36984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[454\]
timestamp 1606716760
transform 1 0 35880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[18\]_TE
timestamp 1606716760
transform 1 0 36340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_389
timestamp 1606716760
transform 1 0 36156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1606716760
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[125\]_A
timestamp 1606716760
transform 1 0 35420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_378
timestamp 1606716760
transform 1 0 35144 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_383
timestamp 1606716760
transform 1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[10\]
timestamp 1606716760
transform 1 0 39744 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1606716760
transform 1 0 39652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_425
timestamp 1606716760
transform 1 0 39468 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[127\]_B
timestamp 1606716760
transform 1 0 38548 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_417
timestamp 1606716760
transform 1 0 38732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[127\]
timestamp 1606716760
transform 1 0 37536 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_413
timestamp 1606716760
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[113\]_B
timestamp 1606716760
transform 1 0 37168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_396
timestamp 1606716760
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_402
timestamp 1606716760
transform 1 0 37352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[112\]
timestamp 1606716760
transform 1 0 35972 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_386
timestamp 1606716760
transform 1 0 35880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_382
timestamp 1606716760
transform 1 0 35512 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[84\]
timestamp 1606716760
transform 1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[42\]_TE
timestamp 1606716760
transform 1 0 39652 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[10\]_TE
timestamp 1606716760
transform 1 0 39284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_421
timestamp 1606716760
transform 1 0 39100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_425
timestamp 1606716760
transform 1 0 39468 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_415
timestamp 1606716760
transform 1 0 38548 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[113\]_A
timestamp 1606716760
transform 1 0 37996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[127\]_A
timestamp 1606716760
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_407
timestamp 1606716760
transform 1 0 37812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_411
timestamp 1606716760
transform 1 0 38180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[113\]
timestamp 1606716760
transform 1 0 36984 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1606716760
transform 1 0 36892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_396
timestamp 1606716760
transform 1 0 36800 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[112\]_A
timestamp 1606716760
transform 1 0 36616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[112\]_B
timestamp 1606716760
transform 1 0 36156 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_388
timestamp 1606716760
transform 1 0 36064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_391
timestamp 1606716760
transform 1 0 36340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[441\]
timestamp 1606716760
transform 1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_382
timestamp 1606716760
transform 1 0 35512 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[116\]
timestamp 1606716760
transform 1 0 39744 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1606716760
transform 1 0 39652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_419
timestamp 1606716760
transform 1 0 38916 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[457\]
timestamp 1606716760
transform 1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_407
timestamp 1606716760
transform 1 0 37812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_396
timestamp 1606716760
transform 1 0 36800 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[442\]
timestamp 1606716760
transform 1 0 36524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[116\]_A
timestamp 1606716760
transform 1 0 35972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_385
timestamp 1606716760
transform 1 0 35788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_389
timestamp 1606716760
transform 1 0 36156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[80\]
timestamp 1606716760
transform 1 0 34500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1606716760
transform 1 0 34040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_367
timestamp 1606716760
transform 1 0 34132 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_365
timestamp 1606716760
transform 1 0 33948 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_353
timestamp 1606716760
transform 1 0 32844 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[120\]_B
timestamp 1606716760
transform 1 0 32660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_349
timestamp 1606716760
transform 1 0 32476 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[75\]
timestamp 1606716760
transform 1 0 31648 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_332
timestamp 1606716760
transform 1 0 30912 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[6\]
timestamp 1606716760
transform 1 0 30084 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[121\]
timestamp 1606716760
transform 1 0 34776 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[80\]_A
timestamp 1606716760
transform 1 0 34592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_360
timestamp 1606716760
transform 1 0 33488 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[120\]_A
timestamp 1606716760
transform 1 0 33304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_356
timestamp 1606716760
transform 1 0 33120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[120\]
timestamp 1606716760
transform 1 0 32292 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[75\]_A
timestamp 1606716760
transform 1 0 32016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_343
timestamp 1606716760
transform 1 0 31924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_346
timestamp 1606716760
transform 1 0 32200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1606716760
transform 1 0 31280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[6\]_A
timestamp 1606716760
transform 1 0 30728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_328
timestamp 1606716760
transform 1 0 30544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1606716760
transform 1 0 30912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_337
timestamp 1606716760
transform 1 0 31372 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[452\]
timestamp 1606716760
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_323
timestamp 1606716760
transform 1 0 30084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[173\]
timestamp 1606716760
transform 1 0 34684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1606716760
transform 1 0 34040 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_367
timestamp 1606716760
transform 1 0 34132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_362
timestamp 1606716760
transform 1 0 33672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[450\]
timestamp 1606716760
transform 1 0 32292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_350
timestamp 1606716760
transform 1 0 32568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_339
timestamp 1606716760
transform 1 0 31556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[122\]
timestamp 1606716760
transform 1 0 30728 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_329
timestamp 1606716760
transform 1 0 30636 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[125\]
timestamp 1606716760
transform 1 0 34776 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1606716760
transform 1 0 34040 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_367
timestamp 1606716760
transform 1 0 34132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_373
timestamp 1606716760
transform 1 0 34684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_368
timestamp 1606716760
transform 1 0 34224 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[455\]
timestamp 1606716760
transform 1 0 33948 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_354
timestamp 1606716760
transform 1 0 32936 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_353
timestamp 1606716760
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_342
timestamp 1606716760
transform 1 0 31832 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_341
timestamp 1606716760
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[122\]_A
timestamp 1606716760
transform 1 0 31556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1606716760
transform 1 0 31280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[122\]_B
timestamp 1606716760
transform 1 0 30912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_330
timestamp 1606716760
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_326
timestamp 1606716760
transform 1 0 30360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1606716760
transform 1 0 31096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1606716760
transform 1 0 31372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[92\]
timestamp 1606716760
transform 1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[125\]_B
timestamp 1606716760
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1606716760
transform 1 0 33580 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1606716760
transform 1 0 32476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1606716760
transform 1 0 31280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1606716760
transform 1 0 30912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1606716760
transform 1 0 31372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[189\]
timestamp 1606716760
transform 1 0 34132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1606716760
transform 1 0 34040 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_370
timestamp 1606716760
transform 1 0 34408 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[111\]_B
timestamp 1606716760
transform 1 0 33856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1606716760
transform 1 0 33672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_354
timestamp 1606716760
transform 1 0 32936 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_342
timestamp 1606716760
transform 1 0 31832 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_330
timestamp 1606716760
transform 1 0 30728 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[111\]_A
timestamp 1606716760
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_371
timestamp 1606716760
transform 1 0 34500 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_375
timestamp 1606716760
transform 1 0 34868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[111\]
timestamp 1606716760
transform 1 0 33672 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_361
timestamp 1606716760
transform 1 0 33580 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1606716760
transform 1 0 32476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1606716760
transform 1 0 31280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1606716760
transform 1 0 30728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1606716760
transform 1 0 31372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[116\]
timestamp 1606716760
transform 1 0 34132 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1606716760
transform 1 0 34040 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_365
timestamp 1606716760
transform 1 0 33948 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_353
timestamp 1606716760
transform 1 0 32844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_341
timestamp 1606716760
transform 1 0 31740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_329
timestamp 1606716760
transform 1 0 30636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_315
timestamp 1606716760
transform 1 0 29348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[64\]
timestamp 1606716760
transform 1 0 28520 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1606716760
transform 1 0 28428 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[119\]_B
timestamp 1606716760
transform 1 0 27876 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_301
timestamp 1606716760
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[62\]
timestamp 1606716760
transform 1 0 26864 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1606716760
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_280
timestamp 1606716760
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[59\]
timestamp 1606716760
transform 1 0 25300 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_315
timestamp 1606716760
transform 1 0 29348 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[151\]
timestamp 1606716760
transform 1 0 29072 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[119\]_A
timestamp 1606716760
transform 1 0 28520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[64\]_A
timestamp 1606716760
transform 1 0 28888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_308
timestamp 1606716760
transform 1 0 28704 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_304
timestamp 1606716760
transform 1 0 28336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[119\]
timestamp 1606716760
transform 1 0 27508 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[60\]_A
timestamp 1606716760
transform 1 0 26956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[62\]_A
timestamp 1606716760
transform 1 0 27324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_287
timestamp 1606716760
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_291
timestamp 1606716760
transform 1 0 27140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[60\]
timestamp 1606716760
transform 1 0 25944 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1606716760
transform 1 0 25668 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[59\]_A
timestamp 1606716760
transform 1 0 25484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_272
timestamp 1606716760
transform 1 0 25392 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_276
timestamp 1606716760
transform 1 0 25760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_321
timestamp 1606716760
transform 1 0 29900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[449\]
timestamp 1606716760
transform 1 0 28520 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1606716760
transform 1 0 28796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1606716760
transform 1 0 28428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_304
timestamp 1606716760
transform 1 0 28336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[118\]_B
timestamp 1606716760
transform 1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[123\]_B
timestamp 1606716760
transform 1 0 27600 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_289
timestamp 1606716760
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_293
timestamp 1606716760
transform 1 0 27324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_298
timestamp 1606716760
transform 1 0 27784 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[118\]
timestamp 1606716760
transform 1 0 26128 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[114\]_B
timestamp 1606716760
transform 1 0 25944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_272
timestamp 1606716760
transform 1 0 25392 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_318
timestamp 1606716760
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_314
timestamp 1606716760
transform 1 0 29256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[453\]
timestamp 1606716760
transform 1 0 28980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_306
timestamp 1606716760
transform 1 0 28520 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_307
timestamp 1606716760
transform 1 0 28612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[123\]
timestamp 1606716760
transform 1 0 27416 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_297
timestamp 1606716760
transform 1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_303
timestamp 1606716760
transform 1 0 28244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[123\]_A
timestamp 1606716760
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1606716760
transform 1 0 28428 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[114\]_A
timestamp 1606716760
transform 1 0 26772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_289
timestamp 1606716760
transform 1 0 26956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[444\]
timestamp 1606716760
transform 1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[118\]_A
timestamp 1606716760
transform 1 0 27140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_293
timestamp 1606716760
transform 1 0 27324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[114\]
timestamp 1606716760
transform 1 0 25760 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[117\]_B
timestamp 1606716760
transform 1 0 25944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[440\]
timestamp 1606716760
transform 1 0 26404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_280
timestamp 1606716760
transform 1 0 26128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_286
timestamp 1606716760
transform 1 0 26680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_285
timestamp 1606716760
transform 1 0 26588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[11\]_A
timestamp 1606716760
transform 1 0 25208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1606716760
transform 1 0 25668 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_275
timestamp 1606716760
transform 1 0 25668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_272
timestamp 1606716760
transform 1 0 25392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_320
timestamp 1606716760
transform 1 0 29808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_308
timestamp 1606716760
transform 1 0 28704 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[447\]
timestamp 1606716760
transform 1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[117\]_A
timestamp 1606716760
transform 1 0 26772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_289
timestamp 1606716760
transform 1 0 26956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_296
timestamp 1606716760
transform 1 0 27600 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_285
timestamp 1606716760
transform 1 0 26588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[117\]
timestamp 1606716760
transform 1 0 25760 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1606716760
transform 1 0 25668 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[110\]_A
timestamp 1606716760
transform 1 0 25484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_270
timestamp 1606716760
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_318
timestamp 1606716760
transform 1 0 29624 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_306
timestamp 1606716760
transform 1 0 28520 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1606716760
transform 1 0 28428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_299
timestamp 1606716760
transform 1 0 27876 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_287
timestamp 1606716760
transform 1 0 26772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[181\]
timestamp 1606716760
transform 1 0 26496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_283
timestamp 1606716760
transform 1 0 26404 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_271
timestamp 1606716760
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_318
timestamp 1606716760
transform 1 0 29624 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_306
timestamp 1606716760
transform 1 0 28520 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[107\]_A
timestamp 1606716760
transform 1 0 28336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_302
timestamp 1606716760
transform 1 0 28152 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[107\]
timestamp 1606716760
transform 1 0 26496 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[107\]_TE
timestamp 1606716760
transform 1 0 26312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1606716760
transform 1 0 25668 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_269
timestamp 1606716760
transform 1 0 25116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_276
timestamp 1606716760
transform 1 0 25760 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[122\]
timestamp 1606716760
transform 1 0 29808 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_318
timestamp 1606716760
transform 1 0 29624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_306
timestamp 1606716760
transform 1 0 28520 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1606716760
transform 1 0 28428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_304
timestamp 1606716760
transform 1 0 28336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[445\]
timestamp 1606716760
transform 1 0 27324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_296
timestamp 1606716760
transform 1 0 27600 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_285
timestamp 1606716760
transform 1 0 26588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[115\]
timestamp 1606716760
transform 1 0 25760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1606716760
transform 1 0 25300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_275
timestamp 1606716760
transform 1 0 25668 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_263
timestamp 1606716760
transform 1 0 24564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[55\]
timestamp 1606716760
transform 1 0 23736 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_253
timestamp 1606716760
transform 1 0 23644 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[116\]_B
timestamp 1606716760
transform 1 0 23460 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1606716760
transform 1 0 22816 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1606716760
transform 1 0 22908 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[59\]_A
timestamp 1606716760
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_228
timestamp 1606716760
transform 1 0 21344 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_232
timestamp 1606716760
transform 1 0 21712 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[55\]_A
timestamp 1606716760
transform 1 0 24656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_262
timestamp 1606716760
transform 1 0 24472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_266
timestamp 1606716760
transform 1 0 24840 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[116\]_A
timestamp 1606716760
transform 1 0 24288 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1606716760
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[116\]
timestamp 1606716760
transform 1 0 23276 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[62\]_A
timestamp 1606716760
transform 1 0 21988 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1606716760
transform 1 0 22172 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_233
timestamp 1606716760
transform 1 0 21804 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[62\]
timestamp 1606716760
transform 1 0 20148 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[11\]
timestamp 1606716760
transform 1 0 24564 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_260
timestamp 1606716760
transform 1 0 24288 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_248
timestamp 1606716760
transform 1 0 23184 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[340\]
timestamp 1606716760
transform 1 0 22908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1606716760
transform 1 0 22816 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_235
timestamp 1606716760
transform 1 0 21988 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_243
timestamp 1606716760
transform 1 0 22724 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[142\]
timestamp 1606716760
transform 1 0 21344 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[24\]_TE
timestamp 1606716760
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_231
timestamp 1606716760
transform 1 0 21620 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[62\]_TE
timestamp 1606716760
transform 1 0 20792 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_220
timestamp 1606716760
transform 1 0 20608 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1606716760
transform 1 0 20976 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[110\]
timestamp 1606716760
transform 1 0 24840 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[11\]_B
timestamp 1606716760
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_262
timestamp 1606716760
transform 1 0 24472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_267
timestamp 1606716760
transform 1 0 24932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_255
timestamp 1606716760
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1606716760
transform 1 0 24104 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_254
timestamp 1606716760
transform 1 0 23736 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[24\]_A
timestamp 1606716760
transform 1 0 23644 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[118\]_A
timestamp 1606716760
transform 1 0 23920 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[438\]
timestamp 1606716760
transform 1 0 24196 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_251
timestamp 1606716760
transform 1 0 23460 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[10\]
timestamp 1606716760
transform 1 0 22908 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1606716760
transform 1 0 22816 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[118\]_TE
timestamp 1606716760
transform 1 0 22080 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_234
timestamp 1606716760
transform 1 0 21896 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_238
timestamp 1606716760
transform 1 0 22264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[103\]
timestamp 1606716760
transform 1 0 21068 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[106\]
timestamp 1606716760
transform 1 0 20148 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  la_buf\[24\]
timestamp 1606716760
transform 1 0 21804 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[0\]_A
timestamp 1606716760
transform 1 0 21160 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_224
timestamp 1606716760
transform 1 0 20976 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_232
timestamp 1606716760
transform 1 0 21712 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_228
timestamp 1606716760
transform 1 0 21344 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[106\]_A
timestamp 1606716760
transform 1 0 21528 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1606716760
transform 1 0 20332 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[104\]_A
timestamp 1606716760
transform 1 0 20516 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[103\]_B
timestamp 1606716760
transform 1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1606716760
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[192\]
timestamp 1606716760
transform 1 0 24472 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[110\]_B
timestamp 1606716760
transform 1 0 25024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_265
timestamp 1606716760
transform 1 0 24748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[10\]_A
timestamp 1606716760
transform 1 0 23920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_254
timestamp 1606716760
transform 1 0 23736 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_258
timestamp 1606716760
transform 1 0 24104 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[118\]
timestamp 1606716760
transform 1 0 22080 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_13_234
timestamp 1606716760
transform 1 0 21896 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[103\]_A
timestamp 1606716760
transform 1 0 21712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_231
timestamp 1606716760
transform 1 0 21620 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[107\]
timestamp 1606716760
transform 1 0 20424 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_215
timestamp 1606716760
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_227
timestamp 1606716760
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[37\]
timestamp 1606716760
transform 1 0 23644 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[10\]_B
timestamp 1606716760
transform 1 0 23092 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_249
timestamp 1606716760
transform 1 0 23276 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1606716760
transform 1 0 22816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[108\]_A
timestamp 1606716760
transform 1 0 22264 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_236
timestamp 1606716760
transform 1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_240
timestamp 1606716760
transform 1 0 22448 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_245
timestamp 1606716760
transform 1 0 22908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[108\]
timestamp 1606716760
transform 1 0 21252 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[107\]_A
timestamp 1606716760
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[107\]_B
timestamp 1606716760
transform 1 0 20700 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_219
timestamp 1606716760
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_223
timestamp 1606716760
transform 1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[37\]_A
timestamp 1606716760
transform 1 0 24932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_266
timestamp 1606716760
transform 1 0 24840 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[111\]
timestamp 1606716760
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[37\]_TE
timestamp 1606716760
transform 1 0 23644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_258
timestamp 1606716760
transform 1 0 24104 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[119\]_A
timestamp 1606716760
transform 1 0 23276 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_247
timestamp 1606716760
transform 1 0 23092 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_251
timestamp 1606716760
transform 1 0 23460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[119\]
timestamp 1606716760
transform 1 0 21436 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[433\]
timestamp 1606716760
transform 1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[109\]_A
timestamp 1606716760
transform 1 0 20884 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[119\]_TE
timestamp 1606716760
transform 1 0 21252 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_215
timestamp 1606716760
transform 1 0 20148 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1606716760
transform 1 0 20700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1606716760
transform 1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_259
timestamp 1606716760
transform 1 0 24196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[11\]
timestamp 1606716760
transform 1 0 23368 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_249
timestamp 1606716760
transform 1 0 23276 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1606716760
transform 1 0 22816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_234
timestamp 1606716760
transform 1 0 21896 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_242
timestamp 1606716760
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_245
timestamp 1606716760
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[114\]_TE
timestamp 1606716760
transform 1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[108\]_B
timestamp 1606716760
transform 1 0 21712 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_230
timestamp 1606716760
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_226
timestamp 1606716760
transform 1 0 21160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[59\]
timestamp 1606716760
transform 1 0 19688 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_202
timestamp 1606716760
transform 1 0 18952 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[57\]
timestamp 1606716760
transform 1 0 17296 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1606716760
transform 1 0 17204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[131\]
timestamp 1606716760
transform 1 0 16192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1606716760
transform 1 0 15364 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_171
timestamp 1606716760
transform 1 0 16100 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_175
timestamp 1606716760
transform 1 0 16468 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1606716760
transform 1 0 20056 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[59\]_TE
timestamp 1606716760
transform 1 0 19688 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1606716760
transform 1 0 19872 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[134\]
timestamp 1606716760
transform 1 0 19044 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_200
timestamp 1606716760
transform 1 0 18768 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1606716760
transform 1 0 19320 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[57\]_A
timestamp 1606716760
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[57\]_TE
timestamp 1606716760
transform 1 0 17296 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_183
timestamp 1606716760
transform 1 0 17204 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_186
timestamp 1606716760
transform 1 0 17480 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_177
timestamp 1606716760
transform 1 0 16652 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[431\]
timestamp 1606716760
transform 1 0 16376 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_166
timestamp 1606716760
transform 1 0 15640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[0\]
timestamp 1606716760
transform 1 0 19780 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[330\]
timestamp 1606716760
transform 1 0 18768 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_203
timestamp 1606716760
transform 1 0 19044 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[435\]
timestamp 1606716760
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1606716760
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_180
timestamp 1606716760
transform 1 0 16928 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_184
timestamp 1606716760
transform 1 0 17296 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_188
timestamp 1606716760
transform 1 0 17664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1606716760
transform 1 0 18032 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[430\]
timestamp 1606716760
transform 1 0 15548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[11\]_TE
timestamp 1606716760
transform 1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_164
timestamp 1606716760
transform 1 0 15456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1606716760
transform 1 0 15824 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[104\]
timestamp 1606716760
transform 1 0 19504 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[106\]_B
timestamp 1606716760
transform 1 0 19504 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1606716760
transform 1 0 20056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[0\]_B
timestamp 1606716760
transform 1 0 19872 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_210
timestamp 1606716760
transform 1 0 19688 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_207
timestamp 1606716760
transform 1 0 19412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_201
timestamp 1606716760
transform 1 0 18860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_207
timestamp 1606716760
transform 1 0 19412 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_201
timestamp 1606716760
transform 1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[105\]_B
timestamp 1606716760
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[100\]_A
timestamp 1606716760
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1606716760
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[100\]
timestamp 1606716760
transform 1 0 17664 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[101\]
timestamp 1606716760
transform 1 0 17296 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1606716760
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[11\]_A
timestamp 1606716760
transform 1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[100\]_B
timestamp 1606716760
transform 1 0 17480 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_193
timestamp 1606716760
transform 1 0 18124 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_180
timestamp 1606716760
transform 1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1606716760
transform 1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[11\]
timestamp 1606716760
transform 1 0 15272 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[102\]
timestamp 1606716760
transform 1 0 15640 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_175
timestamp 1606716760
transform 1 0 16468 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1606716760
transform 1 0 20056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[104\]_B
timestamp 1606716760
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_210
timestamp 1606716760
transform 1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[105\]_A
timestamp 1606716760
transform 1 0 19504 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_206
timestamp 1606716760
transform 1 0 19320 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[105\]
timestamp 1606716760
transform 1 0 18492 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[101\]_B
timestamp 1606716760
transform 1 0 18308 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[437\]
timestamp 1606716760
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[101\]_A
timestamp 1606716760
transform 1 0 17940 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_189
timestamp 1606716760
transform 1 0 17756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1606716760
transform 1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[102\]_A
timestamp 1606716760
transform 1 0 16560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_178
timestamp 1606716760
transform 1 0 16744 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[85\]
timestamp 1606716760
transform 1 0 16100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[102\]_B
timestamp 1606716760
transform 1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1606716760
transform 1 0 15364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1606716760
transform 1 0 15732 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_170
timestamp 1606716760
transform 1 0 16008 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_174
timestamp 1606716760
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[109\]
timestamp 1606716760
transform 1 0 19688 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[434\]
timestamp 1606716760
transform 1 0 18676 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_202
timestamp 1606716760
transform 1 0 18952 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[439\]
timestamp 1606716760
transform 1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1606716760
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_184
timestamp 1606716760
transform 1 0 17296 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_191
timestamp 1606716760
transform 1 0 17940 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[13\]_A
timestamp 1606716760
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1606716760
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_171
timestamp 1606716760
transform 1 0 16100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1606716760
transform 1 0 20056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[109\]_B
timestamp 1606716760
transform 1 0 19872 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[436\]
timestamp 1606716760
transform 1 0 19044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_206
timestamp 1606716760
transform 1 0 19320 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_195
timestamp 1606716760
transform 1 0 18308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[98\]
timestamp 1606716760
transform 1 0 18032 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1606716760
transform 1 0 17664 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_176
timestamp 1606716760
transform 1 0 16560 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[121\]_A
timestamp 1606716760
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1606716760
transform 1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[1\]
timestamp 1606716760
transform 1 0 19504 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_10_196
timestamp 1606716760
transform 1 0 18400 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1606716760
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1606716760
transform 1 0 17020 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1606716760
transform 1 0 17296 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[186\]
timestamp 1606716760
transform 1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_167
timestamp 1606716760
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_173
timestamp 1606716760
transform 1 0 16284 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_151
timestamp 1606716760
transform 1 0 14260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[55\]
timestamp 1606716760
transform 1 0 12604 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_18_131
timestamp 1606716760
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1606716760
transform 1 0 11592 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1606716760
transform 1 0 10396 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1606716760
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_123
timestamp 1606716760
transform 1 0 11684 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1606716760
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[55\]_A
timestamp 1606716760
transform 1 0 13892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_149
timestamp 1606716760
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_154
timestamp 1606716760
transform 1 0 14536 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[55\]_TE
timestamp 1606716760
transform 1 0 12604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1606716760
transform 1 0 12788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_109
timestamp 1606716760
transform 1 0 10396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_121
timestamp 1606716760
transform 1 0 11500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_159
timestamp 1606716760
transform 1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_147
timestamp 1606716760
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_135
timestamp 1606716760
transform 1 0 12788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1606716760
transform 1 0 11592 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_112
timestamp 1606716760
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1606716760
transform 1 0 11408 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1606716760
transform 1 0 11684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_158
timestamp 1606716760
transform 1 0 14904 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1606716760
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_154
timestamp 1606716760
transform 1 0 14536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[22\]
timestamp 1606716760
transform 1 0 13248 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1606716760
transform 1 0 12788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1606716760
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_129
timestamp 1606716760
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_141
timestamp 1606716760
transform 1 0 13340 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1606716760
transform 1 0 11592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_116
timestamp 1606716760
transform 1 0 11040 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1606716760
transform 1 0 11684 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_117
timestamp 1606716760
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[432\]
timestamp 1606716760
transform 1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1606716760
transform 1 0 14904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1606716760
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[22\]_A
timestamp 1606716760
transform 1 0 14720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_145
timestamp 1606716760
transform 1 0 13708 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_154
timestamp 1606716760
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[87\]
timestamp 1606716760
transform 1 0 13432 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[22\]_TE
timestamp 1606716760
transform 1 0 13248 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_132
timestamp 1606716760
transform 1 0 12512 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_108
timestamp 1606716760
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_120
timestamp 1606716760
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[13\]
timestamp 1606716760
transform 1 0 14076 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[195\]
timestamp 1606716760
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_135
timestamp 1606716760
transform 1 0 12788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1606716760
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1606716760
transform 1 0 11592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_116
timestamp 1606716760
transform 1 0 11040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1606716760
transform 1 0 11684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[121\]
timestamp 1606716760
transform 1 0 14536 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1606716760
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[121\]_TE
timestamp 1606716760
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[13\]_TE
timestamp 1606716760
transform 1 0 13892 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_145
timestamp 1606716760
transform 1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1606716760
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[96\]
timestamp 1606716760
transform 1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1606716760
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_139
timestamp 1606716760
transform 1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[20\]_A
timestamp 1606716760
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_111
timestamp 1606716760
transform 1 0 10580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1606716760
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_159
timestamp 1606716760
transform 1 0 14996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_147
timestamp 1606716760
transform 1 0 13892 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_135
timestamp 1606716760
transform 1 0 12788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1606716760
transform 1 0 11592 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[39\]_TE
timestamp 1606716760
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_111
timestamp 1606716760
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_119
timestamp 1606716760
transform 1 0 11316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1606716760
transform 1 0 11684 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[78\]
timestamp 1606716760
transform 1 0 10120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_98
timestamp 1606716760
transform 1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[48\]
timestamp 1606716760
transform 1 0 7728 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_72
timestamp 1606716760
transform 1 0 6992 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[122\]
timestamp 1606716760
transform 1 0 6716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1606716760
transform 1 0 5980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[53\]_TE
timestamp 1606716760
transform 1 0 6256 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_60
timestamp 1606716760
transform 1 0 5888 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_62
timestamp 1606716760
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_66
timestamp 1606716760
transform 1 0 6440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1606716760
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[48\]_A
timestamp 1606716760
transform 1 0 9108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1606716760
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_97
timestamp 1606716760
transform 1 0 9292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[109\]_A
timestamp 1606716760
transform 1 0 7912 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[48\]_TE
timestamp 1606716760
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1606716760
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1606716760
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1606716760
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[109\]
timestamp 1606716760
transform 1 0 6072 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[109\]_TE
timestamp 1606716760
transform 1 0 5888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[48\]_B
timestamp 1606716760
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1606716760
transform 1 0 5520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_100
timestamp 1606716760
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[183\]
timestamp 1606716760
transform 1 0 7084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_76
timestamp 1606716760
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_88
timestamp 1606716760
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[125\]
timestamp 1606716760
transform 1 0 6072 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1606716760
transform 1 0 5980 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[104\]_TE
timestamp 1606716760
transform 1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_58
timestamp 1606716760
transform 1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1606716760
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_69
timestamp 1606716760
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_105
timestamp 1606716760
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1606716760
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_92
timestamp 1606716760
transform 1 0 8832 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_104
timestamp 1606716760
transform 1 0 9936 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1606716760
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_91
timestamp 1606716760
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[104\]_A
timestamp 1606716760
transform 1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1606716760
transform 1 0 7728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_83
timestamp 1606716760
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1606716760
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[104\]
timestamp 1606716760
transform 1 0 6348 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1606716760
transform 1 0 6624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[178\]
timestamp 1606716760
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1606716760
transform 1 0 5980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[101\]_A
timestamp 1606716760
transform 1 0 5796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[106\]_A
timestamp 1606716760
transform 1 0 5428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 1606716760
transform 1 0 5612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1606716760
transform 1 0 5612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_61
timestamp 1606716760
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_62
timestamp 1606716760
transform 1 0 6072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[94\]
timestamp 1606716760
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1606716760
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_96
timestamp 1606716760
transform 1 0 9200 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_76
timestamp 1606716760
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_88
timestamp 1606716760
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[180\]
timestamp 1606716760
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[103\]_A
timestamp 1606716760
transform 1 0 5428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1606716760
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_64
timestamp 1606716760
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[0\]_A
timestamp 1606716760
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_100
timestamp 1606716760
transform 1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_104
timestamp 1606716760
transform 1 0 9936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[0\]
timestamp 1606716760
transform 1 0 7912 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 1606716760
transform 1 0 7176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1606716760
transform 1 0 5980 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[110\]_A
timestamp 1606716760
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1606716760
transform 1 0 5612 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1606716760
transform 1 0 6072 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[20\]
timestamp 1606716760
transform 1 0 8924 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1606716760
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[20\]_TE
timestamp 1606716760
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[74\]
timestamp 1606716760
transform 1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[0\]_TE
timestamp 1606716760
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_78
timestamp 1606716760
transform 1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1606716760
transform 1 0 8096 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp 1606716760
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[100\]_A
timestamp 1606716760
transform 1 0 6256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1606716760
transform 1 0 6072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_66
timestamp 1606716760
transform 1 0 6440 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_106
timestamp 1606716760
transform 1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[113\]
timestamp 1606716760
transform 1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_95
timestamp 1606716760
transform 1 0 9108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[102\]
timestamp 1606716760
transform 1 0 7452 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[182\]
timestamp 1606716760
transform 1 0 6072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1606716760
transform 1 0 5980 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[108\]_TE
timestamp 1606716760
transform 1 0 5796 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_57
timestamp 1606716760
transform 1 0 5612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1606716760
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[48\]
timestamp 1606716760
transform 1 0 4324 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[4\]_B
timestamp 1606716760
transform 1 0 3956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1606716760
transform 1 0 4140 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_52
timestamp 1606716760
transform 1 0 5152 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[334\]
timestamp 1606716760
transform 1 0 3312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606716760
transform 1 0 2852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_31
timestamp 1606716760
transform 1 0 3220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_35
timestamp 1606716760
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606716760
transform 1 0 368 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606716760
transform 1 0 644 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606716760
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[48\]_A
timestamp 1606716760
transform 1 0 4968 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_46
timestamp 1606716760
transform 1 0 4600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_52
timestamp 1606716760
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[4\]
timestamp 1606716760
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1606716760
transform 1 0 3220 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1606716760
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_32
timestamp 1606716760
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_36
timestamp 1606716760
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606716760
transform 1 0 368 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606716760
transform 1 0 644 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606716760
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[175\]
timestamp 1606716760
transform 1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[4\]_A
timestamp 1606716760
transform 1 0 4416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_42
timestamp 1606716760
transform 1 0 4232 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_46
timestamp 1606716760
transform 1 0 4600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1606716760
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606716760
transform 1 0 368 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606716760
transform 1 0 644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606716760
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_53
timestamp 1606716760
transform 1 0 5244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[101\]
timestamp 1606716760
transform 1 0 3956 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[106\]
timestamp 1606716760
transform 1 0 3588 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1606716760
transform 1 0 3220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[101\]_TE
timestamp 1606716760
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_27
timestamp 1606716760
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1606716760
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1606716760
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_36
timestamp 1606716760
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606716760
transform 1 0 368 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606716760
transform 1 0 368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606716760
transform 1 0 644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606716760
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606716760
transform 1 0 644 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606716760
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1606716760
transform 1 0 5244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[103\]
timestamp 1606716760
transform 1 0 3588 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[177\]
timestamp 1606716760
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1606716760
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[103\]_TE
timestamp 1606716760
transform 1 0 3036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[106\]_TE
timestamp 1606716760
transform 1 0 2668 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_19
timestamp 1606716760
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_23
timestamp 1606716760
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1606716760
transform 1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_32
timestamp 1606716760
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606716760
transform 1 0 368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606716760
transform 1 0 644 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1606716760
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_53
timestamp 1606716760
transform 1 0 5244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[110\]
timestamp 1606716760
transform 1 0 3588 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_27
timestamp 1606716760
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606716760
transform 1 0 368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606716760
transform 1 0 644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606716760
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[100\]
timestamp 1606716760
transform 1 0 4416 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[100\]_TE
timestamp 1606716760
transform 1 0 4232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[110\]_TE
timestamp 1606716760
transform 1 0 3864 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_40
timestamp 1606716760
transform 1 0 4048 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[184\]
timestamp 1606716760
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1606716760
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1606716760
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_32
timestamp 1606716760
transform 1 0 3312 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_36
timestamp 1606716760
transform 1 0 3680 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606716760
transform 1 0 368 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606716760
transform 1 0 644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606716760
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[174\]
timestamp 1606716760
transform 1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_38
timestamp 1606716760
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_45
timestamp 1606716760
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[179\]
timestamp 1606716760
transform 1 0 3220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[120\]_TE
timestamp 1606716760
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606716760
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_34
timestamp 1606716760
transform 1 0 3496 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606716760
transform 1 0 368 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606716760
transform 1 0 644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606716760
transform 1 0 1748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606716760
transform -1 0 169556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606716760
transform -1 0 169556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606716760
transform -1 0 169556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1832
timestamp 1606716760
transform 1 0 168912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1832
timestamp 1606716760
transform 1 0 168912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1824
timestamp 1606716760
transform 1 0 168176 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606716760
transform -1 0 169556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606716760
transform -1 0 169556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1832
timestamp 1606716760
transform 1 0 168912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1834
timestamp 1606716760
transform 1 0 169096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606716760
transform -1 0 169556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606716760
transform -1 0 169556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1832
timestamp 1606716760
transform 1 0 168912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1832
timestamp 1606716760
transform 1 0 168912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606716760
transform -1 0 169556 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606716760
transform -1 0 169556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606716760
transform -1 0 169556 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1834
timestamp 1606716760
transform 1 0 169096 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1834
timestamp 1606716760
transform 1 0 169096 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1832
timestamp 1606716760
transform 1 0 168912 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1820
timestamp 1606716760
transform 1 0 167808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1808
timestamp 1606716760
transform 1 0 166704 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1606716760
transform 1 0 166612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_we_buf_A
timestamp 1606716760
transform 1 0 165416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_sel_buf\[2\]_A
timestamp 1606716760
transform 1 0 165784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1796
timestamp 1606716760
transform 1 0 165600 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1800
timestamp 1606716760
transform 1 0 165968 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1806
timestamp 1606716760
transform 1 0 166520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1792
timestamp 1606716760
transform 1 0 165232 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_we_buf
timestamp 1606716760
transform 1 0 163576 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_sel_buf\[2\]_TE
timestamp 1606716760
transform 1 0 163392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1812
timestamp 1606716760
transform 1 0 167072 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1800
timestamp 1606716760
transform 1 0 165968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1606716760
transform 1 0 164588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1606716760
transform 1 0 163760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1777
timestamp 1606716760
transform 1 0 163852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1788
timestamp 1606716760
transform 1 0 164864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1770
timestamp 1606716760
transform 1 0 163208 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1822
timestamp 1606716760
transform 1 0 167992 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1820
timestamp 1606716760
transform 1 0 167808 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1810
timestamp 1606716760
transform 1 0 166888 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1808
timestamp 1606716760
transform 1 0 166704 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1606716760
transform 1 0 165508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1606716760
transform 1 0 166612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1798
timestamp 1606716760
transform 1 0 165784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1799
timestamp 1606716760
transform 1 0 165876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1789
timestamp 1606716760
transform 1 0 164956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1606716760
transform 1 0 163760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1606716760
transform 1 0 164588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1777
timestamp 1606716760
transform 1 0 163852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1776
timestamp 1606716760
transform 1 0 163760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1784
timestamp 1606716760
transform 1 0 164496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1787
timestamp 1606716760
transform 1 0 164772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1606716760
transform 1 0 163576 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1774
timestamp 1606716760
transform 1 0 163576 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1772
timestamp 1606716760
transform 1 0 163392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1820
timestamp 1606716760
transform 1 0 167808 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1808
timestamp 1606716760
transform 1 0 166704 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1606716760
transform 1 0 166612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1606716760
transform 1 0 165508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1797
timestamp 1606716760
transform 1 0 165692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1805
timestamp 1606716760
transform 1 0 166428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1606716760
transform 1 0 164128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1606716760
transform 1 0 164588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1779
timestamp 1606716760
transform 1 0 164036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1783
timestamp 1606716760
transform 1 0 164404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1787
timestamp 1606716760
transform 1 0 164772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1773
timestamp 1606716760
transform 1 0 163484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1820
timestamp 1606716760
transform 1 0 167808 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1808
timestamp 1606716760
transform 1 0 166704 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1606716760
transform 1 0 165416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1796
timestamp 1606716760
transform 1 0 165600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1606716760
transform 1 0 164956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1792
timestamp 1606716760
transform 1 0 165232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1606716760
transform 1 0 163944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1606716760
transform 1 0 163760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_vdd_pwrgood_A
timestamp 1606716760
transform 1 0 164680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1777
timestamp 1606716760
transform 1 0 163852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1781
timestamp 1606716760
transform 1 0 164220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1785
timestamp 1606716760
transform 1 0 164588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1788
timestamp 1606716760
transform 1 0 164864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1772
timestamp 1606716760
transform 1 0 163392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1820
timestamp 1606716760
transform 1 0 167808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1808
timestamp 1606716760
transform 1 0 166704 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1606716760
transform 1 0 166612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1797
timestamp 1606716760
transform 1 0 165692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1805
timestamp 1606716760
transform 1 0 166428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  mprj_vdd_pwrgood
timestamp 1606716760
transform 1 0 164588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1606716760
transform 1 0 163944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1777
timestamp 1606716760
transform 1 0 163852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1780
timestamp 1606716760
transform 1 0 164128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1784
timestamp 1606716760
transform 1 0 164496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1771
timestamp 1606716760
transform 1 0 163300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1820
timestamp 1606716760
transform 1 0 167808 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  mprj2_vdd_pwrgood
timestamp 1606716760
transform 1 0 166704 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1800
timestamp 1606716760
transform 1 0 165968 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1606716760
transform 1 0 163852 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  mprj2_pwrgood
timestamp 1606716760
transform 1 0 164864 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1606716760
transform 1 0 163760 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1775
timestamp 1606716760
transform 1 0 163668 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1780
timestamp 1606716760
transform 1 0 164128 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1771
timestamp 1606716760
transform 1 0 163300 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1822
timestamp 1606716760
transform 1 0 167992 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1822
timestamp 1606716760
transform 1 0 167992 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1817
timestamp 1606716760
transform 1 0 167532 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj2_vdd_pwrgood_A
timestamp 1606716760
transform 1 0 167532 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1606716760
transform 1 0 167624 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[458\]
timestamp 1606716760
transform 1 0 167716 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[294\]
timestamp 1606716760
transform 1 0 167716 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1606716760
transform 1 0 166704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[92\]_A
timestamp 1606716760
transform 1 0 166796 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1811
timestamp 1606716760
transform 1 0 166980 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1811
timestamp 1606716760
transform 1 0 166980 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1815
timestamp 1606716760
transform 1 0 167348 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1606716760
transform 1 0 167164 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1807
timestamp 1606716760
transform 1 0 166612 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1606716760
transform 1 0 166612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1803
timestamp 1606716760
transform 1 0 166244 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_pwrgood_A
timestamp 1606716760
transform 1 0 166428 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj2_pwrgood_A
timestamp 1606716760
transform 1 0 166060 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1799
timestamp 1606716760
transform 1 0 165876 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[92\]
timestamp 1606716760
transform 1 0 164956 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_8  mprj_pwrgood
timestamp 1606716760
transform 1 0 164772 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A
timestamp 1606716760
transform 1 0 164036 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1606716760
transform 1 0 164404 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1779
timestamp 1606716760
transform 1 0 164036 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1781
timestamp 1606716760
transform 1 0 164220 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1606716760
transform 1 0 164772 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[92\]_TE
timestamp 1606716760
transform 1 0 164588 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1788
timestamp 1606716760
transform 1 0 164864 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1785
timestamp 1606716760
transform 1 0 164588 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1606716760
transform 1 0 163576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[9\]_A
timestamp 1606716760
transform 1 0 163852 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1775
timestamp 1606716760
transform 1 0 163668 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1777
timestamp 1606716760
transform 1 0 163852 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[5\]
timestamp 1606716760
transform 1 0 162564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1766
timestamp 1606716760
transform 1 0 162840 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1759
timestamp 1606716760
transform 1 0 162196 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1606716760
transform 1 0 161000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1745
timestamp 1606716760
transform 1 0 160908 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1747
timestamp 1606716760
transform 1 0 161092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1606716760
transform 1 0 159160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__A
timestamp 1606716760
transform 1 0 159620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1729
timestamp 1606716760
transform 1 0 159436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1733
timestamp 1606716760
transform 1 0 159804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__A
timestamp 1606716760
transform 1 0 158608 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1718
timestamp 1606716760
transform 1 0 158424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1722
timestamp 1606716760
transform 1 0 158792 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1758
timestamp 1606716760
transform 1 0 162104 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1746
timestamp 1606716760
transform 1 0 161000 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1734
timestamp 1606716760
transform 1 0 159896 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[27\]
timestamp 1606716760
transform 1 0 158240 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1606716760
transform 1 0 163116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1762
timestamp 1606716760
transform 1 0 162472 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1767
timestamp 1606716760
transform 1 0 162932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _447_
timestamp 1606716760
transform 1 0 162196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1759
timestamp 1606716760
transform 1 0 162196 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1606716760
transform 1 0 161184 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1606716760
transform 1 0 161000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1751
timestamp 1606716760
transform 1 0 161460 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1744
timestamp 1606716760
transform 1 0 160816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1747
timestamp 1606716760
transform 1 0 161092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1606716760
transform 1 0 160172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1740
timestamp 1606716760
transform 1 0 160448 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[27\]_A
timestamp 1606716760
transform 1 0 159528 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1733
timestamp 1606716760
transform 1 0 159804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1732
timestamp 1606716760
transform 1 0 159712 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1606716760
transform 1 0 158424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[27\]_TE
timestamp 1606716760
transform 1 0 158240 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1716
timestamp 1606716760
transform 1 0 158240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1721
timestamp 1606716760
transform 1 0 158700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1718
timestamp 1606716760
transform 1 0 158424 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1761
timestamp 1606716760
transform 1 0 162380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A
timestamp 1606716760
transform 1 0 162196 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1606716760
transform 1 0 161000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__A
timestamp 1606716760
transform 1 0 161276 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1745
timestamp 1606716760
transform 1 0 160908 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1747
timestamp 1606716760
transform 1 0 161092 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1751
timestamp 1606716760
transform 1 0 161460 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__A
timestamp 1606716760
transform 1 0 160172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1739
timestamp 1606716760
transform 1 0 160356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[300\]
timestamp 1606716760
transform 1 0 159620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1728
timestamp 1606716760
transform 1 0 159344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1734
timestamp 1606716760
transform 1 0 159896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__A
timestamp 1606716760
transform 1 0 158424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1720
timestamp 1606716760
transform 1 0 158608 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1760
timestamp 1606716760
transform 1 0 162288 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[211\]
timestamp 1606716760
transform 1 0 162012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1606716760
transform 1 0 160632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1745
timestamp 1606716760
transform 1 0 160908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1740
timestamp 1606716760
transform 1 0 160448 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _467_
timestamp 1606716760
transform 1 0 159436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1727
timestamp 1606716760
transform 1 0 159252 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1732
timestamp 1606716760
transform 1 0 159712 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[298\]
timestamp 1606716760
transform 1 0 158240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1719
timestamp 1606716760
transform 1 0 158516 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1606716760
transform 1 0 162656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1606716760
transform 1 0 163116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1760
timestamp 1606716760
transform 1 0 162288 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1767
timestamp 1606716760
transform 1 0 162932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__A
timestamp 1606716760
transform 1 0 162104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1756
timestamp 1606716760
transform 1 0 161920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1606716760
transform 1 0 161644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1606716760
transform 1 0 161000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__A
timestamp 1606716760
transform 1 0 160632 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1744
timestamp 1606716760
transform 1 0 160816 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1747
timestamp 1606716760
transform 1 0 161092 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__A
timestamp 1606716760
transform 1 0 160172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1735
timestamp 1606716760
transform 1 0 159988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1739
timestamp 1606716760
transform 1 0 160356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1606716760
transform 1 0 159344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1606716760
transform 1 0 159804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1724
timestamp 1606716760
transform 1 0 158976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1731
timestamp 1606716760
transform 1 0 159620 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1606716760
transform 1 0 158332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1606716760
transform 1 0 158792 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1716
timestamp 1606716760
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1720
timestamp 1606716760
transform 1 0 158608 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1606716760
transform 1 0 161920 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1755
timestamp 1606716760
transform 1 0 161828 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1759
timestamp 1606716760
transform 1 0 162196 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1606716760
transform 1 0 160816 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1747
timestamp 1606716760
transform 1 0 161092 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1736
timestamp 1606716760
transform 1 0 160080 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1606716760
transform 1 0 159804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[90\]_A
timestamp 1606716760
transform 1 0 159528 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1723
timestamp 1606716760
transform 1 0 158884 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1729
timestamp 1606716760
transform 1 0 159436 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1732
timestamp 1606716760
transform 1 0 159712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1606716760
transform 1 0 158240 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[90\]_TE
timestamp 1606716760
transform 1 0 158700 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1719
timestamp 1606716760
transform 1 0 158516 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[9\]
timestamp 1606716760
transform 1 0 162012 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1768
timestamp 1606716760
transform 1 0 163024 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1764
timestamp 1606716760
transform 1 0 162656 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__608__A
timestamp 1606716760
transform 1 0 162840 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1606716760
transform 1 0 161920 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1606716760
transform 1 0 161920 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[9\]_TE
timestamp 1606716760
transform 1 0 161736 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1754
timestamp 1606716760
transform 1 0 161736 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1758
timestamp 1606716760
transform 1 0 162104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _608_
timestamp 1606716760
transform 1 0 162380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[98\]_A
timestamp 1606716760
transform 1 0 161276 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1750
timestamp 1606716760
transform 1 0 161368 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1606716760
transform 1 0 161552 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1751
timestamp 1606716760
transform 1 0 161460 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1606716760
transform 1 0 161092 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1606716760
transform 1 0 161000 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__A
timestamp 1606716760
transform 1 0 160816 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1747
timestamp 1606716760
transform 1 0 161092 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1738
timestamp 1606716760
transform 1 0 160264 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1606716760
transform 1 0 160080 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[98\]
timestamp 1606716760
transform 1 0 159436 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1606716760
transform 1 0 159068 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[98\]_TE
timestamp 1606716760
transform 1 0 158884 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1726
timestamp 1606716760
transform 1 0 159160 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1734
timestamp 1606716760
transform 1 0 159896 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[90\]
timestamp 1606716760
transform 1 0 158240 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[96\]_A
timestamp 1606716760
transform 1 0 158516 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1717
timestamp 1606716760
transform 1 0 158332 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1721
timestamp 1606716760
transform 1 0 158700 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp 1606716760
transform 1 0 158148 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[25\]_A
timestamp 1606716760
transform 1 0 157596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1711
timestamp 1606716760
transform 1 0 157780 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1707
timestamp 1606716760
transform 1 0 157412 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[25\]
timestamp 1606716760
transform 1 0 155756 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1606716760
transform 1 0 155388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[20\]_A
timestamp 1606716760
transform 1 0 155204 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1686
timestamp 1606716760
transform 1 0 155480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[0\]_A
timestamp 1606716760
transform 1 0 154836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1677
timestamp 1606716760
transform 1 0 154652 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1681
timestamp 1606716760
transform 1 0 155020 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1606716760
transform 1 0 158148 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1714
timestamp 1606716760
transform 1 0 158056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1702
timestamp 1606716760
transform 1 0 156952 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[21\]
timestamp 1606716760
transform 1 0 155296 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1676
timestamp 1606716760
transform 1 0 154560 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1606716760
transform 1 0 158148 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1715
timestamp 1606716760
transform 1 0 158148 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1703
timestamp 1606716760
transform 1 0 157044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1707
timestamp 1606716760
transform 1 0 157412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[67\]
timestamp 1606716760
transform 1 0 156768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1695
timestamp 1606716760
transform 1 0 156308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1606716760
transform 1 0 156032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__A
timestamp 1606716760
transform 1 0 156216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[21\]_A
timestamp 1606716760
transform 1 0 156584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1692
timestamp 1606716760
transform 1 0 156032 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1696
timestamp 1606716760
transform 1 0 156400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1606716760
transform 1 0 155388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[21\]_TE
timestamp 1606716760
transform 1 0 155204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1684
timestamp 1606716760
transform 1 0 155296 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1686
timestamp 1606716760
transform 1 0 155480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1606716760
transform 1 0 155756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1667
timestamp 1606716760
transform 1 0 153732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__A
timestamp 1606716760
transform 1 0 154376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[16\]_A
timestamp 1606716760
transform 1 0 154744 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1672
timestamp 1606716760
transform 1 0 154192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1676
timestamp 1606716760
transform 1 0 154560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1606716760
transform 1 0 155020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1679
timestamp 1606716760
transform 1 0 154836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1680
timestamp 1606716760
transform 1 0 154928 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1665
timestamp 1606716760
transform 1 0 153548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1663
timestamp 1606716760
transform 1 0 153364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[16\]_TE
timestamp 1606716760
transform 1 0 153364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[62\]
timestamp 1606716760
transform 1 0 153456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1606716760
transform 1 0 153916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1706
timestamp 1606716760
transform 1 0 157320 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__A
timestamp 1606716760
transform 1 0 156032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1694
timestamp 1606716760
transform 1 0 156216 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1606716760
transform 1 0 155388 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1683
timestamp 1606716760
transform 1 0 155204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1686
timestamp 1606716760
transform 1 0 155480 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__A
timestamp 1606716760
transform 1 0 155020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1674
timestamp 1606716760
transform 1 0 154376 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1680
timestamp 1606716760
transform 1 0 154928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1606716760
transform 1 0 158148 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1709
timestamp 1606716760
transform 1 0 157596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1606716760
transform 1 0 156216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1697
timestamp 1606716760
transform 1 0 156492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1606716760
transform 1 0 155204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1686
timestamp 1606716760
transform 1 0 155480 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1606716760
transform 1 0 154192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1671
timestamp 1606716760
transform 1 0 154100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1675
timestamp 1606716760
transform 1 0 154468 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1667
timestamp 1606716760
transform 1 0 153732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__A
timestamp 1606716760
transform 1 0 157688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1708
timestamp 1606716760
transform 1 0 157504 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1712
timestamp 1606716760
transform 1 0 157872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 1606716760
transform 1 0 157228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1700
timestamp 1606716760
transform 1 0 156768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1704
timestamp 1606716760
transform 1 0 157136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1606716760
transform 1 0 155756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A
timestamp 1606716760
transform 1 0 156216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__A
timestamp 1606716760
transform 1 0 156584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1692
timestamp 1606716760
transform 1 0 156032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1696
timestamp 1606716760
transform 1 0 156400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1606716760
transform 1 0 155388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__A
timestamp 1606716760
transform 1 0 155204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1682
timestamp 1606716760
transform 1 0 155112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1686
timestamp 1606716760
transform 1 0 155480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__A
timestamp 1606716760
transform 1 0 154192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1674
timestamp 1606716760
transform 1 0 154376 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1666
timestamp 1606716760
transform 1 0 153640 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1606716760
transform 1 0 158148 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1714
timestamp 1606716760
transform 1 0 158056 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1606716760
transform 1 0 157136 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1702
timestamp 1606716760
transform 1 0 156952 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1706
timestamp 1606716760
transform 1 0 157320 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1606716760
transform 1 0 156676 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__A
timestamp 1606716760
transform 1 0 156124 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1691
timestamp 1606716760
transform 1 0 155940 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1695
timestamp 1606716760
transform 1 0 156308 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1606716760
transform 1 0 155664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1606716760
transform 1 0 154652 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1680
timestamp 1606716760
transform 1 0 154928 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1606716760
transform 1 0 153640 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1669
timestamp 1606716760
transform 1 0 153916 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1606716760
transform 1 0 158056 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[94\]_A
timestamp 1606716760
transform 1 0 157596 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1711
timestamp 1606716760
transform 1 0 157780 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1707
timestamp 1606716760
transform 1 0 157412 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[96\]
timestamp 1606716760
transform 1 0 156676 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[94\]
timestamp 1606716760
transform 1 0 155756 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1695
timestamp 1606716760
transform 1 0 156308 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1691
timestamp 1606716760
transform 1 0 155940 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[96\]_TE
timestamp 1606716760
transform 1 0 156492 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1606716760
transform 1 0 156216 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[292\]
timestamp 1606716760
transform 1 0 155204 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1682
timestamp 1606716760
transform 1 0 155112 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1606716760
transform 1 0 155388 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1686
timestamp 1606716760
transform 1 0 155480 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1686
timestamp 1606716760
transform 1 0 155480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[94\]_TE
timestamp 1606716760
transform 1 0 155756 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1664
timestamp 1606716760
transform 1 0 153456 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[296\]
timestamp 1606716760
transform 1 0 154376 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1676
timestamp 1606716760
transform 1 0 154560 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__A
timestamp 1606716760
transform 1 0 154836 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1677
timestamp 1606716760
transform 1 0 154652 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1681
timestamp 1606716760
transform 1 0 155020 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1668
timestamp 1606716760
transform 1 0 153824 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1665
timestamp 1606716760
transform 1 0 153548 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__A
timestamp 1606716760
transform 1 0 153640 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1606716760
transform 1 0 153364 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[20\]
timestamp 1606716760
transform 1 0 152996 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_dat_buf\[0\]_TE
timestamp 1606716760
transform 1 0 152812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[58\]
timestamp 1606716760
transform 1 0 151984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1651
timestamp 1606716760
transform 1 0 152260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[66\]
timestamp 1606716760
transform 1 0 150972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1640
timestamp 1606716760
transform 1 0 151248 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1629
timestamp 1606716760
transform 1 0 150236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1606716760
transform 1 0 149776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[29\]_A
timestamp 1606716760
transform 1 0 150052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1625
timestamp 1606716760
transform 1 0 149868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[39\]
timestamp 1606716760
transform 1 0 148764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_adr_buf\[29\]_TE
timestamp 1606716760
transform 1 0 148396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1611
timestamp 1606716760
transform 1 0 148580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1616
timestamp 1606716760
transform 1 0 149040 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[16\]
timestamp 1606716760
transform 1 0 152904 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1606716760
transform 1 0 152536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1655
timestamp 1606716760
transform 1 0 152628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1642
timestamp 1606716760
transform 1 0 151432 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1630
timestamp 1606716760
transform 1 0 150328 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1618
timestamp 1606716760
transform 1 0 149224 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[63\]
timestamp 1606716760
transform 1 0 152904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1657
timestamp 1606716760
transform 1 0 152812 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1661
timestamp 1606716760
transform 1 0 153180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1606716760
transform 1 0 152536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__A
timestamp 1606716760
transform 1 0 152076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1655
timestamp 1606716760
transform 1 0 152628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1647
timestamp 1606716760
transform 1 0 151892 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1651
timestamp 1606716760
transform 1 0 152260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1606716760
transform 1 0 151616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1642
timestamp 1606716760
transform 1 0 151432 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1642
timestamp 1606716760
transform 1 0 151432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1630
timestamp 1606716760
transform 1 0 150328 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1634
timestamp 1606716760
transform 1 0 150696 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1630
timestamp 1606716760
transform 1 0 150328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A
timestamp 1606716760
transform 1 0 150512 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1625
timestamp 1606716760
transform 1 0 149868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1623
timestamp 1606716760
transform 1 0 149684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1621
timestamp 1606716760
transform 1 0 149500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1606716760
transform 1 0 149776 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1606716760
transform 1 0 150052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1606716760
transform 1 0 150052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1609
timestamp 1606716760
transform 1 0 148396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1615
timestamp 1606716760
transform 1 0 148948 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1662
timestamp 1606716760
transform 1 0 153272 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A
timestamp 1606716760
transform 1 0 151984 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1650
timestamp 1606716760
transform 1 0 152168 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1606716760
transform 1 0 151524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1642
timestamp 1606716760
transform 1 0 151432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1646
timestamp 1606716760
transform 1 0 151800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1606716760
transform 1 0 150328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A
timestamp 1606716760
transform 1 0 150696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1628
timestamp 1606716760
transform 1 0 150144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1632
timestamp 1606716760
transform 1 0 150512 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1636
timestamp 1606716760
transform 1 0 150880 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1606716760
transform 1 0 149868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1606716760
transform 1 0 149776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1620
timestamp 1606716760
transform 1 0 149408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1606716760
transform 1 0 152536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1651
timestamp 1606716760
transform 1 0 152260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1655
timestamp 1606716760
transform 1 0 152628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1643
timestamp 1606716760
transform 1 0 151524 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1631
timestamp 1606716760
transform 1 0 150420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1619
timestamp 1606716760
transform 1 0 149316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1606716760
transform 1 0 149040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1614
timestamp 1606716760
transform 1 0 148856 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1606716760
transform 1 0 151892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__A
timestamp 1606716760
transform 1 0 152352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1650
timestamp 1606716760
transform 1 0 152168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1654
timestamp 1606716760
transform 1 0 152536 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__A
timestamp 1606716760
transform 1 0 151340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1639
timestamp 1606716760
transform 1 0 151156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1643
timestamp 1606716760
transform 1 0 151524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1606716760
transform 1 0 150880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1606716760
transform 1 0 150328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1628
timestamp 1606716760
transform 1 0 150144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1632
timestamp 1606716760
transform 1 0 150512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1606716760
transform 1 0 149868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1606716760
transform 1 0 149776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1606716760
transform 1 0 149500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1619
timestamp 1606716760
transform 1 0 149316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1623
timestamp 1606716760
transform 1 0 149684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1606716760
transform 1 0 148672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1606716760
transform 1 0 149132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1615
timestamp 1606716760
transform 1 0 148948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1658
timestamp 1606716760
transform 1 0 152904 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1606716760
transform 1 0 152628 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1606716760
transform 1 0 152536 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1652
timestamp 1606716760
transform 1 0 152352 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1644
timestamp 1606716760
transform 1 0 151616 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1606716760
transform 1 0 150236 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1632
timestamp 1606716760
transform 1 0 150512 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1621
timestamp 1606716760
transform 1 0 149500 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1657
timestamp 1606716760
transform 1 0 152812 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1655
timestamp 1606716760
transform 1 0 152628 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__A
timestamp 1606716760
transform 1 0 152628 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1654
timestamp 1606716760
transform 1 0 152536 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1648
timestamp 1606716760
transform 1 0 151984 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1651
timestamp 1606716760
transform 1 0 152260 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[89\]_A
timestamp 1606716760
transform 1 0 152444 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[89\]
timestamp 1606716760
transform 1 0 150604 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1606716760
transform 1 0 151340 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1640
timestamp 1606716760
transform 1 0 151248 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1644
timestamp 1606716760
transform 1 0 151616 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1606716760
transform 1 0 151800 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1606716760
transform 1 0 150512 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1606716760
transform 1 0 150328 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A
timestamp 1606716760
transform 1 0 150696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[89\]_TE
timestamp 1606716760
transform 1 0 150328 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1628
timestamp 1606716760
transform 1 0 150144 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1632
timestamp 1606716760
transform 1 0 150512 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1636
timestamp 1606716760
transform 1 0 150880 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1606716760
transform 1 0 149868 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1606716760
transform 1 0 149776 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1624
timestamp 1606716760
transform 1 0 149776 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1623
timestamp 1606716760
transform 1 0 149684 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1616
timestamp 1606716760
transform 1 0 149040 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1617
timestamp 1606716760
transform 1 0 149132 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[69\]_A
timestamp 1606716760
transform 1 0 149132 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[291\]
timestamp 1606716760
transform 1 0 149500 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1619
timestamp 1606716760
transform 1 0 149316 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1610
timestamp 1606716760
transform 1 0 148488 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1608
timestamp 1606716760
transform 1 0 148304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1600
timestamp 1606716760
transform 1 0 147568 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1588
timestamp 1606716760
transform 1 0 146464 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1576
timestamp 1606716760
transform 1 0 145360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1606716760
transform 1 0 144164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1564
timestamp 1606716760
transform 1 0 144256 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1606
timestamp 1606716760
transform 1 0 148120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1606716760
transform 1 0 146924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1594
timestamp 1606716760
transform 1 0 147016 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1591
timestamp 1606716760
transform 1 0 146740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1606716760
transform 1 0 145728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1577
timestamp 1606716760
transform 1 0 145452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1583
timestamp 1606716760
transform 1 0 146004 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1569
timestamp 1606716760
transform 1 0 144716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1557
timestamp 1606716760
transform 1 0 143612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1606716760
transform 1 0 148120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1606716760
transform 1 0 147200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1606716760
transform 1 0 146924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1606716760
transform 1 0 147660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1594
timestamp 1606716760
transform 1 0 147016 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1594
timestamp 1606716760
transform 1 0 147016 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1599
timestamp 1606716760
transform 1 0 147476 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1603
timestamp 1606716760
transform 1 0 147844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1606716760
transform 1 0 145728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1581
timestamp 1606716760
transform 1 0 145820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1576
timestamp 1606716760
transform 1 0 145360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1582
timestamp 1606716760
transform 1 0 145912 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1569
timestamp 1606716760
transform 1 0 144716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1606716760
transform 1 0 144164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1557
timestamp 1606716760
transform 1 0 143612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1564
timestamp 1606716760
transform 1 0 144256 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1606716760
transform 1 0 148120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1605
timestamp 1606716760
transform 1 0 148028 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1608
timestamp 1606716760
transform 1 0 148304 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1601
timestamp 1606716760
transform 1 0 147660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1606716760
transform 1 0 146372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1585
timestamp 1606716760
transform 1 0 146188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1589
timestamp 1606716760
transform 1 0 146556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1606716760
transform 1 0 145912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1576
timestamp 1606716760
transform 1 0 145360 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1606716760
transform 1 0 144164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1558
timestamp 1606716760
transform 1 0 143704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1562
timestamp 1606716760
transform 1 0 144072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1564
timestamp 1606716760
transform 1 0 144256 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1606
timestamp 1606716760
transform 1 0 148120 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1606716760
transform 1 0 146924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1594
timestamp 1606716760
transform 1 0 147016 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1590
timestamp 1606716760
transform 1 0 146648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1606716760
transform 1 0 145268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1578
timestamp 1606716760
transform 1 0 145544 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1567
timestamp 1606716760
transform 1 0 144532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1555
timestamp 1606716760
transform 1 0 143428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1606716760
transform 1 0 148120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1604
timestamp 1606716760
transform 1 0 147936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1608
timestamp 1606716760
transform 1 0 148304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1606716760
transform 1 0 147660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1593
timestamp 1606716760
transform 1 0 146924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1606716760
transform 1 0 146280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1606716760
transform 1 0 146740 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1589
timestamp 1606716760
transform 1 0 146556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1606716760
transform 1 0 145268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1606716760
transform 1 0 145728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1606716760
transform 1 0 146096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1578
timestamp 1606716760
transform 1 0 145544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1582
timestamp 1606716760
transform 1 0 145912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1572
timestamp 1606716760
transform 1 0 144992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1606716760
transform 1 0 144164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1555
timestamp 1606716760
transform 1 0 143428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1564
timestamp 1606716760
transform 1 0 144256 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[69\]
timestamp 1606716760
transform 1 0 147844 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1606716760
transform 1 0 146924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1594
timestamp 1606716760
transform 1 0 147016 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1602
timestamp 1606716760
transform 1 0 147752 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1585
timestamp 1606716760
transform 1 0 146188 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1606716760
transform 1 0 145912 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1570
timestamp 1606716760
transform 1 0 144808 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1605
timestamp 1606716760
transform 1 0 148028 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[271\]
timestamp 1606716760
transform 1 0 147844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1606
timestamp 1606716760
transform 1 0 148120 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[69\]_TE
timestamp 1606716760
transform 1 0 148304 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1593
timestamp 1606716760
transform 1 0 146924 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[289\]
timestamp 1606716760
transform 1 0 147752 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1606716760
transform 1 0 147660 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[87\]_A
timestamp 1606716760
transform 1 0 147016 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1596
timestamp 1606716760
transform 1 0 147200 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1600
timestamp 1606716760
transform 1 0 147568 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1601
timestamp 1606716760
transform 1 0 147660 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[87\]
timestamp 1606716760
transform 1 0 145176 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1606716760
transform 1 0 146372 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A
timestamp 1606716760
transform 1 0 146740 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1592
timestamp 1606716760
transform 1 0 146832 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1585
timestamp 1606716760
transform 1 0 146188 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1589
timestamp 1606716760
transform 1 0 146556 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1574
timestamp 1606716760
transform 1 0 145176 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1606716760
transform 1 0 145912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1606716760
transform 1 0 145360 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1578
timestamp 1606716760
transform 1 0 145544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1564
timestamp 1606716760
transform 1 0 144256 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1606716760
transform 1 0 144900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1606716760
transform 1 0 144808 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[67\]_A
timestamp 1606716760
transform 1 0 144440 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[87\]_TE
timestamp 1606716760
transform 1 0 144624 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1566
timestamp 1606716760
transform 1 0 144440 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1571
timestamp 1606716760
transform 1 0 144900 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1568
timestamp 1606716760
transform 1 0 144624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1562
timestamp 1606716760
transform 1 0 144072 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1556
timestamp 1606716760
transform 1 0 143520 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1558
timestamp 1606716760
transform 1 0 143704 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1606716760
transform 1 0 143520 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1606716760
transform 1 0 144164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1551
timestamp 1606716760
transform 1 0 143060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1539
timestamp 1606716760
transform 1 0 141956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1527
timestamp 1606716760
transform 1 0 140852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1515
timestamp 1606716760
transform 1 0 139748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1606716760
transform 1 0 138552 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1503
timestamp 1606716760
transform 1 0 138644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1545
timestamp 1606716760
transform 1 0 142508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1533
timestamp 1606716760
transform 1 0 141404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1606716760
transform 1 0 141312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1520
timestamp 1606716760
transform 1 0 140208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1508
timestamp 1606716760
transform 1 0 139104 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1545
timestamp 1606716760
transform 1 0 142508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1551
timestamp 1606716760
transform 1 0 143060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1533
timestamp 1606716760
transform 1 0 141404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1539
timestamp 1606716760
transform 1 0 141956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1606716760
transform 1 0 141312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1522
timestamp 1606716760
transform 1 0 140392 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1530
timestamp 1606716760
transform 1 0 141128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1527
timestamp 1606716760
transform 1 0 140852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1515
timestamp 1606716760
transform 1 0 139748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1606716760
transform 1 0 138552 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1510
timestamp 1606716760
transform 1 0 139288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1503
timestamp 1606716760
transform 1 0 138644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1546
timestamp 1606716760
transform 1 0 142600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1534
timestamp 1606716760
transform 1 0 141496 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1522
timestamp 1606716760
transform 1 0 140392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _660_
timestamp 1606716760
transform 1 0 138644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1606716760
transform 1 0 138552 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__660__A
timestamp 1606716760
transform 1 0 139104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1506
timestamp 1606716760
transform 1 0 138920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1510
timestamp 1606716760
transform 1 0 139288 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[269\]
timestamp 1606716760
transform 1 0 143152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1548
timestamp 1606716760
transform 1 0 142784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[287\]
timestamp 1606716760
transform 1 0 141404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1536
timestamp 1606716760
transform 1 0 141680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1606716760
transform 1 0 141312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1530
timestamp 1606716760
transform 1 0 141128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[207\]
timestamp 1606716760
transform 1 0 139748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1518
timestamp 1606716760
transform 1 0 140024 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1606716760
transform 1 0 138736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1606716760
transform 1 0 139196 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1507
timestamp 1606716760
transform 1 0 139012 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1511
timestamp 1606716760
transform 1 0 139380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1606716760
transform 1 0 143244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1606716760
transform 1 0 142784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1544
timestamp 1606716760
transform 1 0 142416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1551
timestamp 1606716760
transform 1 0 143060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[285\]
timestamp 1606716760
transform 1 0 141036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[65\]_A
timestamp 1606716760
transform 1 0 140484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1521
timestamp 1606716760
transform 1 0 140300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1525
timestamp 1606716760
transform 1 0 140668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1532
timestamp 1606716760
transform 1 0 141312 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[65\]
timestamp 1606716760
transform 1 0 138644 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1606716760
transform 1 0 138552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[67\]
timestamp 1606716760
transform 1 0 143152 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1540
timestamp 1606716760
transform 1 0 142048 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1606716760
transform 1 0 141404 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A
timestamp 1606716760
transform 1 0 141864 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1536
timestamp 1606716760
transform 1 0 141680 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1606716760
transform 1 0 141312 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[85\]_TE
timestamp 1606716760
transform 1 0 141128 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1527
timestamp 1606716760
transform 1 0 140852 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1606716760
transform 1 0 139932 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1515
timestamp 1606716760
transform 1 0 139748 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1519
timestamp 1606716760
transform 1 0 140116 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1606716760
transform 1 0 139472 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[5\]_TE
timestamp 1606716760
transform 1 0 138920 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[65\]_TE
timestamp 1606716760
transform 1 0 139288 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1504
timestamp 1606716760
transform 1 0 138736 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1508
timestamp 1606716760
transform 1 0 139104 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1554
timestamp 1606716760
transform 1 0 143336 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[67\]_TE
timestamp 1606716760
transform 1 0 143336 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[85\]_A
timestamp 1606716760
transform 1 0 142968 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1606716760
transform 1 0 143060 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1552
timestamp 1606716760
transform 1 0 143152 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1548
timestamp 1606716760
transform 1 0 142784 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1547
timestamp 1606716760
transform 1 0 142692 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1606716760
transform 1 0 142508 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1543
timestamp 1606716760
transform 1 0 142324 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1606716760
transform 1 0 142048 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1606716760
transform 1 0 141956 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[85\]
timestamp 1606716760
transform 1 0 141128 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[5\]_A
timestamp 1606716760
transform 1 0 140484 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[83\]_A
timestamp 1606716760
transform 1 0 141036 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1527
timestamp 1606716760
transform 1 0 140852 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1531
timestamp 1606716760
transform 1 0 141220 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1521
timestamp 1606716760
transform 1 0 140300 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1525
timestamp 1606716760
transform 1 0 140668 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1529
timestamp 1606716760
transform 1 0 141036 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[83\]
timestamp 1606716760
transform 1 0 139196 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[5\]
timestamp 1606716760
transform 1 0 138644 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1505
timestamp 1606716760
transform 1 0 138828 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[83\]_TE
timestamp 1606716760
transform 1 0 138920 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1606716760
transform 1 0 138552 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1606716760
transform 1 0 139104 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1490
timestamp 1606716760
transform 1 0 137448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1478
timestamp 1606716760
transform 1 0 136344 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1466
timestamp 1606716760
transform 1 0 135240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1454
timestamp 1606716760
transform 1 0 134136 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1496
timestamp 1606716760
transform 1 0 138000 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1484
timestamp 1606716760
transform 1 0 136896 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1606716760
transform 1 0 135700 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1472
timestamp 1606716760
transform 1 0 135792 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1459
timestamp 1606716760
transform 1 0 134596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[267\]
timestamp 1606716760
transform 1 0 137908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1492
timestamp 1606716760
transform 1 0 137632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1498
timestamp 1606716760
transform 1 0 138184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1490
timestamp 1606716760
transform 1 0 137448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1484
timestamp 1606716760
transform 1 0 136896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1606716760
transform 1 0 135700 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1470
timestamp 1606716760
transform 1 0 135608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1472
timestamp 1606716760
transform 1 0 135792 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1478
timestamp 1606716760
transform 1 0 136344 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1462
timestamp 1606716760
transform 1 0 134872 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1466
timestamp 1606716760
transform 1 0 135240 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1450
timestamp 1606716760
transform 1 0 133768 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1454
timestamp 1606716760
transform 1 0 134136 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1499
timestamp 1606716760
transform 1 0 138276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[263\]
timestamp 1606716760
transform 1 0 137264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1491
timestamp 1606716760
transform 1 0 137540 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1485
timestamp 1606716760
transform 1 0 136988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1477
timestamp 1606716760
transform 1 0 136252 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1465
timestamp 1606716760
transform 1 0 135148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__A
timestamp 1606716760
transform 1 0 133860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1449
timestamp 1606716760
transform 1 0 133676 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1453
timestamp 1606716760
transform 1 0 134044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _604_
timestamp 1606716760
transform 1 0 137724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1492
timestamp 1606716760
transform 1 0 137632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1496
timestamp 1606716760
transform 1 0 138000 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _657_
timestamp 1606716760
transform 1 0 136620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1484
timestamp 1606716760
transform 1 0 136896 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1606716760
transform 1 0 135700 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1469
timestamp 1606716760
transform 1 0 135516 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1472
timestamp 1606716760
transform 1 0 135792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1480
timestamp 1606716760
transform 1 0 136528 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _644_
timestamp 1606716760
transform 1 0 134136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1457
timestamp 1606716760
transform 1 0 134412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1606716760
transform 1 0 138368 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1606716760
transform 1 0 137540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__A
timestamp 1606716760
transform 1 0 138000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__A
timestamp 1606716760
transform 1 0 137172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1489
timestamp 1606716760
transform 1 0 137356 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1494
timestamp 1606716760
transform 1 0 137816 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1498
timestamp 1606716760
transform 1 0 138184 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__657__A
timestamp 1606716760
transform 1 0 136804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1481
timestamp 1606716760
transform 1 0 136620 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1485
timestamp 1606716760
transform 1 0 136988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _606_
timestamp 1606716760
transform 1 0 136344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__A
timestamp 1606716760
transform 1 0 135424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1470
timestamp 1606716760
transform 1 0 135608 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _646_
timestamp 1606716760
transform 1 0 134964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1462
timestamp 1606716760
transform 1 0 134872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1466
timestamp 1606716760
transform 1 0 135240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__A
timestamp 1606716760
transform 1 0 134136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1456
timestamp 1606716760
transform 1 0 134320 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[61\]
timestamp 1606716760
transform 1 0 137080 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1485
timestamp 1606716760
transform 1 0 136988 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1606716760
transform 1 0 135792 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1606716760
transform 1 0 135700 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1606716760
transform 1 0 136252 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[58\]_TE
timestamp 1606716760
transform 1 0 135332 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1469
timestamp 1606716760
transform 1 0 135516 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1475
timestamp 1606716760
transform 1 0 136068 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1479
timestamp 1606716760
transform 1 0 136436 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1463
timestamp 1606716760
transform 1 0 134964 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[260\]
timestamp 1606716760
transform 1 0 134688 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[283\]
timestamp 1606716760
transform 1 0 133676 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1448
timestamp 1606716760
transform 1 0 133584 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1452
timestamp 1606716760
transform 1 0 133952 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1499
timestamp 1606716760
transform 1 0 138276 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1501
timestamp 1606716760
transform 1 0 138460 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[63\]_A
timestamp 1606716760
transform 1 0 138276 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[61\]_A
timestamp 1606716760
transform 1 0 138368 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[58\]_A
timestamp 1606716760
transform 1 0 137172 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[61\]_TE
timestamp 1606716760
transform 1 0 137540 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1497
timestamp 1606716760
transform 1 0 138092 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1489
timestamp 1606716760
transform 1 0 137356 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1493
timestamp 1606716760
transform 1 0 137724 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1485
timestamp 1606716760
transform 1 0 136988 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[58\]
timestamp 1606716760
transform 1 0 135332 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[63\]
timestamp 1606716760
transform 1 0 136436 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1606716760
transform 1 0 136252 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[81\]_A
timestamp 1606716760
transform 1 0 135700 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[63\]_TE
timestamp 1606716760
transform 1 0 136068 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1469
timestamp 1606716760
transform 1 0 135516 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1473
timestamp 1606716760
transform 1 0 135884 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1478
timestamp 1606716760
transform 1 0 136344 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[265\]
timestamp 1606716760
transform 1 0 134320 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[81\]
timestamp 1606716760
transform 1 0 133860 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1606716760
transform 1 0 133584 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[81\]_TE
timestamp 1606716760
transform 1 0 133676 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1450
timestamp 1606716760
transform 1 0 133768 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1459
timestamp 1606716760
transform 1 0 134596 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1606716760
transform 1 0 132940 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1432
timestamp 1606716760
transform 1 0 132112 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1440
timestamp 1606716760
transform 1 0 132848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1442
timestamp 1606716760
transform 1 0 133032 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[3\]_A
timestamp 1606716760
transform 1 0 130824 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1416
timestamp 1606716760
transform 1 0 130640 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1420
timestamp 1606716760
transform 1 0 131008 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[3\]
timestamp 1606716760
transform 1 0 128984 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[3\]_TE
timestamp 1606716760
transform 1 0 128800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1447
timestamp 1606716760
transform 1 0 133492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1435
timestamp 1606716760
transform 1 0 132388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1423
timestamp 1606716760
transform 1 0 131284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1606716760
transform 1 0 130088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1411
timestamp 1606716760
transform 1 0 130180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1399
timestamp 1606716760
transform 1 0 129076 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1407
timestamp 1606716760
transform 1 0 129812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1606716760
transform 1 0 132940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1438
timestamp 1606716760
transform 1 0 132664 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1440
timestamp 1606716760
transform 1 0 132848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1442
timestamp 1606716760
transform 1 0 133032 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1426
timestamp 1606716760
transform 1 0 131560 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1428
timestamp 1606716760
transform 1 0 131744 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _641_
timestamp 1606716760
transform 1 0 131284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__A
timestamp 1606716760
transform 1 0 131560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1424
timestamp 1606716760
transform 1 0 131376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__A
timestamp 1606716760
transform 1 0 130548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1414
timestamp 1606716760
transform 1 0 130456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1413
timestamp 1606716760
transform 1 0 130364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1417
timestamp 1606716760
transform 1 0 130732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1606716760
transform 1 0 131100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1422
timestamp 1606716760
transform 1 0 131192 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1606716760
transform 1 0 130088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1606716760
transform 1 0 130180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _638_
timestamp 1606716760
transform 1 0 130088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1606716760
transform 1 0 129076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__637__A
timestamp 1606716760
transform 1 0 129536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1402
timestamp 1606716760
transform 1 0 129352 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1398
timestamp 1606716760
transform 1 0 128984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1402
timestamp 1606716760
transform 1 0 129352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1406
timestamp 1606716760
transform 1 0 129720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _645_
timestamp 1606716760
transform 1 0 133400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1606716760
transform 1 0 132940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1440
timestamp 1606716760
transform 1 0 132848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1442
timestamp 1606716760
transform 1 0 133032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1428
timestamp 1606716760
transform 1 0 131744 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1606716760
transform 1 0 130732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__A
timestamp 1606716760
transform 1 0 131192 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__A
timestamp 1606716760
transform 1 0 131560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1413
timestamp 1606716760
transform 1 0 130364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1420
timestamp 1606716760
transform 1 0 131008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1424
timestamp 1606716760
transform 1 0 131376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__A
timestamp 1606716760
transform 1 0 130180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1405
timestamp 1606716760
transform 1 0 129628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _643_
timestamp 1606716760
transform 1 0 133124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1435
timestamp 1606716760
transform 1 0 132388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1446
timestamp 1606716760
transform 1 0 133400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1423
timestamp 1606716760
transform 1 0 131284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1606716760
transform 1 0 130088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1409
timestamp 1606716760
transform 1 0 129996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1411
timestamp 1606716760
transform 1 0 130180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1401
timestamp 1606716760
transform 1 0 129260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1606716760
transform 1 0 132940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__A
timestamp 1606716760
transform 1 0 133216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1438
timestamp 1606716760
transform 1 0 132664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1442
timestamp 1606716760
transform 1 0 133032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1446
timestamp 1606716760
transform 1 0 133400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1430
timestamp 1606716760
transform 1 0 131928 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__A
timestamp 1606716760
transform 1 0 130640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1414
timestamp 1606716760
transform 1 0 130456 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1418
timestamp 1606716760
transform 1 0 130824 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _636_
timestamp 1606716760
transform 1 0 130180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1410
timestamp 1606716760
transform 1 0 130088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1404
timestamp 1606716760
transform 1 0 129536 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1432
timestamp 1606716760
transform 1 0 132112 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1444
timestamp 1606716760
transform 1 0 133216 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _602_
timestamp 1606716760
transform 1 0 130732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[7\]_A
timestamp 1606716760
transform 1 0 130456 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1416
timestamp 1606716760
transform 1 0 130640 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1420
timestamp 1606716760
transform 1 0 131008 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1606716760
transform 1 0 130088 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1411
timestamp 1606716760
transform 1 0 130180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[7\]_TE
timestamp 1606716760
transform 1 0 129168 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1402
timestamp 1606716760
transform 1 0 129352 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1447
timestamp 1606716760
transform 1 0 133492 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1606716760
transform 1 0 133124 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1606716760
transform 1 0 133400 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1442
timestamp 1606716760
transform 1 0 133032 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1442
timestamp 1606716760
transform 1 0 133032 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1446
timestamp 1606716760
transform 1 0 133400 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1606716760
transform 1 0 132940 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A
timestamp 1606716760
transform 1 0 132848 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1438
timestamp 1606716760
transform 1 0 132664 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1437
timestamp 1606716760
transform 1 0 132572 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1434
timestamp 1606716760
transform 1 0 132296 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1433
timestamp 1606716760
transform 1 0 132204 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1606716760
transform 1 0 132388 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1606716760
transform 1 0 132388 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1606716760
transform 1 0 131560 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1424
timestamp 1606716760
transform 1 0 131376 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1422
timestamp 1606716760
transform 1 0 131192 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1606716760
transform 1 0 131928 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1428
timestamp 1606716760
transform 1 0 131744 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1606716760
transform 1 0 130548 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1416
timestamp 1606716760
transform 1 0 130640 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1606716760
transform 1 0 131100 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__A
timestamp 1606716760
transform 1 0 131008 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1420
timestamp 1606716760
transform 1 0 131008 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1418
timestamp 1606716760
transform 1 0 130824 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1412
timestamp 1606716760
transform 1 0 130272 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[209\]
timestamp 1606716760
transform 1 0 129260 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[7\]
timestamp 1606716760
transform 1 0 129168 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__655__A
timestamp 1606716760
transform 1 0 128708 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1397
timestamp 1606716760
transform 1 0 128892 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1404
timestamp 1606716760
transform 1 0 129536 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1606716760
transform 1 0 129076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1606716760
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1381
timestamp 1606716760
transform 1 0 127420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1393
timestamp 1606716760
transform 1 0 128524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1377
timestamp 1606716760
transform 1 0 127052 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1365
timestamp 1606716760
transform 1 0 125948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[2\]_A
timestamp 1606716760
transform 1 0 124660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1349
timestamp 1606716760
transform 1 0 124476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1353
timestamp 1606716760
transform 1 0 124844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _634_
timestamp 1606716760
transform 1 0 127696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1382
timestamp 1606716760
transform 1 0 127512 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1387
timestamp 1606716760
transform 1 0 127972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1362
timestamp 1606716760
transform 1 0 125672 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1374
timestamp 1606716760
transform 1 0 126776 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1606716760
transform 1 0 124476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1350
timestamp 1606716760
transform 1 0 124568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1606716760
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__634__A
timestamp 1606716760
transform 1 0 127696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1390
timestamp 1606716760
transform 1 0 128248 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1379
timestamp 1606716760
transform 1 0 127236 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1381
timestamp 1606716760
transform 1 0 127420 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1386
timestamp 1606716760
transform 1 0 127880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1378
timestamp 1606716760
transform 1 0 127144 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _627_
timestamp 1606716760
transform 1 0 125580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1606716760
transform 1 0 126868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__A
timestamp 1606716760
transform 1 0 126316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1364
timestamp 1606716760
transform 1 0 125856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1368
timestamp 1606716760
transform 1 0 126224 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1371
timestamp 1606716760
transform 1 0 126500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1363
timestamp 1606716760
transform 1 0 125764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1375
timestamp 1606716760
transform 1 0 126868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _622_
timestamp 1606716760
transform 1 0 124568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1606716760
transform 1 0 124476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1344
timestamp 1606716760
transform 1 0 124016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1348
timestamp 1606716760
transform 1 0 124384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1353
timestamp 1606716760
transform 1 0 124844 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1351
timestamp 1606716760
transform 1 0 124660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1606716760
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1381
timestamp 1606716760
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1393
timestamp 1606716760
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1377
timestamp 1606716760
transform 1 0 127052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _635_
timestamp 1606716760
transform 1 0 126316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__A
timestamp 1606716760
transform 1 0 125672 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__632__A
timestamp 1606716760
transform 1 0 126868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1360
timestamp 1606716760
transform 1 0 125488 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1364
timestamp 1606716760
transform 1 0 125856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1368
timestamp 1606716760
transform 1 0 126224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1372
timestamp 1606716760
transform 1 0 126592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__A
timestamp 1606716760
transform 1 0 125304 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _623_
timestamp 1606716760
transform 1 0 124844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__A
timestamp 1606716760
transform 1 0 124568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1347
timestamp 1606716760
transform 1 0 124292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1352
timestamp 1606716760
transform 1 0 124752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1356
timestamp 1606716760
transform 1 0 125120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _633_
timestamp 1606716760
transform 1 0 127880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1384
timestamp 1606716760
transform 1 0 127696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1389
timestamp 1606716760
transform 1 0 128156 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1606716760
transform 1 0 126316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1362
timestamp 1606716760
transform 1 0 125672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1368
timestamp 1606716760
transform 1 0 126224 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1372
timestamp 1606716760
transform 1 0 126592 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1606716760
transform 1 0 124476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1350
timestamp 1606716760
transform 1 0 124568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1341
timestamp 1606716760
transform 1 0 123740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _629_
timestamp 1606716760
transform 1 0 127420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1606716760
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__A
timestamp 1606716760
transform 1 0 127880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__A
timestamp 1606716760
transform 1 0 128248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1384
timestamp 1606716760
transform 1 0 127696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1388
timestamp 1606716760
transform 1 0 128064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1392
timestamp 1606716760
transform 1 0 128432 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1376
timestamp 1606716760
transform 1 0 126960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _601_
timestamp 1606716760
transform 1 0 125948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__A
timestamp 1606716760
transform 1 0 126408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__A
timestamp 1606716760
transform 1 0 126776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1360
timestamp 1606716760
transform 1 0 125488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1364
timestamp 1606716760
transform 1 0 125856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1368
timestamp 1606716760
transform 1 0 126224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1372
timestamp 1606716760
transform 1 0 126592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__A
timestamp 1606716760
transform 1 0 125304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _628_
timestamp 1606716760
transform 1 0 124844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A
timestamp 1606716760
transform 1 0 124108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1343
timestamp 1606716760
transform 1 0 123924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1347
timestamp 1606716760
transform 1 0 124292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1356
timestamp 1606716760
transform 1 0 125120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1606716760
transform 1 0 128156 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1379
timestamp 1606716760
transform 1 0 127236 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1387
timestamp 1606716760
transform 1 0 127972 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1392
timestamp 1606716760
transform 1 0 128432 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[56\]
timestamp 1606716760
transform 1 0 125580 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1357
timestamp 1606716760
transform 1 0 125212 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1606716760
transform 1 0 124568 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1606716760
transform 1 0 124476 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__A
timestamp 1606716760
transform 1 0 125028 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[54\]_TE
timestamp 1606716760
transform 1 0 123924 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1345
timestamp 1606716760
transform 1 0 124108 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1353
timestamp 1606716760
transform 1 0 124844 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1342
timestamp 1606716760
transform 1 0 123832 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _655_
timestamp 1606716760
transform 1 0 128248 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__A
timestamp 1606716760
transform 1 0 128156 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1389
timestamp 1606716760
transform 1 0 128156 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1393
timestamp 1606716760
transform 1 0 128524 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1391
timestamp 1606716760
transform 1 0 128340 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1606716760
transform 1 0 127696 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1606716760
transform 1 0 127328 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1380
timestamp 1606716760
transform 1 0 127328 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1381
timestamp 1606716760
transform 1 0 127420 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1385
timestamp 1606716760
transform 1 0 127788 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1368
timestamp 1606716760
transform 1 0 126224 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[258\]
timestamp 1606716760
transform 1 0 126316 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[56\]_A
timestamp 1606716760
transform 1 0 126868 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1372
timestamp 1606716760
transform 1 0 126592 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1377
timestamp 1606716760
transform 1 0 127052 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _653_
timestamp 1606716760
transform 1 0 125580 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__A
timestamp 1606716760
transform 1 0 126040 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[54\]_A
timestamp 1606716760
transform 1 0 125764 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1360
timestamp 1606716760
transform 1 0 125488 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1364
timestamp 1606716760
transform 1 0 125856 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1361
timestamp 1606716760
transform 1 0 125580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1365
timestamp 1606716760
transform 1 0 125948 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[56\]_TE
timestamp 1606716760
transform 1 0 126132 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[54\]
timestamp 1606716760
transform 1 0 123924 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1606716760
transform 1 0 124844 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1344
timestamp 1606716760
transform 1 0 124016 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1352
timestamp 1606716760
transform 1 0 124752 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1354
timestamp 1606716760
transform 1 0 124936 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1341
timestamp 1606716760
transform 1 0 123740 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[256\]
timestamp 1606716760
transform 1 0 123740 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[2\]
timestamp 1606716760
transform 1 0 122820 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[25\]_A
timestamp 1606716760
transform 1 0 122268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1327
timestamp 1606716760
transform 1 0 122452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[231\]
timestamp 1606716760
transform 1 0 121808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1606716760
transform 1 0 121716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[25\]_TE
timestamp 1606716760
transform 1 0 120888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1312
timestamp 1606716760
transform 1 0 121072 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1318
timestamp 1606716760
transform 1 0 121624 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1323
timestamp 1606716760
transform 1 0 122084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1302
timestamp 1606716760
transform 1 0 120152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1290
timestamp 1606716760
transform 1 0 119048 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1325
timestamp 1606716760
transform 1 0 122268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1337
timestamp 1606716760
transform 1 0 123372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1313
timestamp 1606716760
transform 1 0 121164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1301
timestamp 1606716760
transform 1 0 120060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1606716760
transform 1 0 118864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1289
timestamp 1606716760
transform 1 0 118956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__A
timestamp 1606716760
transform 1 0 122268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1332
timestamp 1606716760
transform 1 0 122912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1327
timestamp 1606716760
transform 1 0 122452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1339
timestamp 1606716760
transform 1 0 123556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _615_
timestamp 1606716760
transform 1 0 121532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _618_
timestamp 1606716760
transform 1 0 121808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1606716760
transform 1 0 121716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1310
timestamp 1606716760
transform 1 0 120888 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1316
timestamp 1606716760
transform 1 0 121440 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1320
timestamp 1606716760
transform 1 0 121808 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1307
timestamp 1606716760
transform 1 0 120612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1323
timestamp 1606716760
transform 1 0 122084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _614_
timestamp 1606716760
transform 1 0 119508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1298
timestamp 1606716760
transform 1 0 119784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1295
timestamp 1606716760
transform 1 0 119508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1606716760
transform 1 0 118864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1289
timestamp 1606716760
transform 1 0 118956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__A
timestamp 1606716760
transform 1 0 122268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1327
timestamp 1606716760
transform 1 0 122452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1339
timestamp 1606716760
transform 1 0 123556 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _619_
timestamp 1606716760
transform 1 0 121808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1606716760
transform 1 0 121716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__615__A
timestamp 1606716760
transform 1 0 121532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1309
timestamp 1606716760
transform 1 0 120796 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1323
timestamp 1606716760
transform 1 0 122084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__614__A
timestamp 1606716760
transform 1 0 119508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1297
timestamp 1606716760
transform 1 0 119692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _620_
timestamp 1606716760
transform 1 0 122360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1325
timestamp 1606716760
transform 1 0 122268 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1329
timestamp 1606716760
transform 1 0 122636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1313
timestamp 1606716760
transform 1 0 121164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1301
timestamp 1606716760
transform 1 0 120060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1606716760
transform 1 0 118864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1289
timestamp 1606716760
transform 1 0 118956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _624_
timestamp 1606716760
transform 1 0 123648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__A
timestamp 1606716760
transform 1 0 122360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1328
timestamp 1606716760
transform 1 0 122544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _613_
timestamp 1606716760
transform 1 0 120704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1606716760
transform 1 0 121716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__A
timestamp 1606716760
transform 1 0 121164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1311
timestamp 1606716760
transform 1 0 120980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1315
timestamp 1606716760
transform 1 0 121348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1320
timestamp 1606716760
transform 1 0 121808 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[280\]
timestamp 1606716760
transform 1 0 119324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1296
timestamp 1606716760
transform 1 0 119600 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A
timestamp 1606716760
transform 1 0 118772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1289
timestamp 1606716760
transform 1 0 118956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _621_
timestamp 1606716760
transform 1 0 122820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1326
timestamp 1606716760
transform 1 0 122360 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1330
timestamp 1606716760
transform 1 0 122728 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1334
timestamp 1606716760
transform 1 0 123096 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _617_
timestamp 1606716760
transform 1 0 120980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1314
timestamp 1606716760
transform 1 0 121256 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _651_
timestamp 1606716760
transform 1 0 119968 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__A
timestamp 1606716760
transform 1 0 119416 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[52\]_A
timestamp 1606716760
transform 1 0 119784 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1292
timestamp 1606716760
transform 1 0 119232 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1296
timestamp 1606716760
transform 1 0 119600 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1303
timestamp 1606716760
transform 1 0 120244 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _616_
timestamp 1606716760
transform 1 0 118956 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1606716760
transform 1 0 118864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1333
timestamp 1606716760
transform 1 0 123004 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1338
timestamp 1606716760
transform 1 0 123464 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1327
timestamp 1606716760
transform 1 0 122452 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1330
timestamp 1606716760
transform 1 0 122728 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1326
timestamp 1606716760
transform 1 0 122360 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__649__A
timestamp 1606716760
transform 1 0 122268 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__A
timestamp 1606716760
transform 1 0 122544 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A
timestamp 1606716760
transform 1 0 122820 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _649_
timestamp 1606716760
transform 1 0 121808 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1606716760
transform 1 0 121992 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1606716760
transform 1 0 121716 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _648_
timestamp 1606716760
transform 1 0 122084 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1323
timestamp 1606716760
transform 1 0 122084 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__617__A
timestamp 1606716760
transform 1 0 120980 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[78\]_A
timestamp 1606716760
transform 1 0 121072 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1310
timestamp 1606716760
transform 1 0 120888 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1313
timestamp 1606716760
transform 1 0 121164 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1314
timestamp 1606716760
transform 1 0 121256 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1305
timestamp 1606716760
transform 1 0 120428 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[78\]
timestamp 1606716760
transform 1 0 119232 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1606716760
transform 1 0 119140 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__651__A
timestamp 1606716760
transform 1 0 120244 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1301
timestamp 1606716760
transform 1 0 120060 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[78\]_TE
timestamp 1606716760
transform 1 0 118956 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1278
timestamp 1606716760
transform 1 0 117944 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _600_
timestamp 1606716760
transform 1 0 116196 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1606716760
transform 1 0 116104 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__A
timestamp 1606716760
transform 1 0 116656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1257
timestamp 1606716760
transform 1 0 116012 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1262
timestamp 1606716760
transform 1 0 116472 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1266
timestamp 1606716760
transform 1 0 116840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp 1606716760
transform 1 0 114632 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1606716760
transform 1 0 115092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1240
timestamp 1606716760
transform 1 0 114448 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1245
timestamp 1606716760
transform 1 0 114908 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1249
timestamp 1606716760
transform 1 0 115276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1276
timestamp 1606716760
transform 1 0 117760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1264
timestamp 1606716760
transform 1 0 116656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _625_
timestamp 1606716760
transform 1 0 115276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1240
timestamp 1606716760
transform 1 0 114448 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1248
timestamp 1606716760
transform 1 0 115184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1252
timestamp 1606716760
transform 1 0 115552 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1282
timestamp 1606716760
transform 1 0 118312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1283
timestamp 1606716760
transform 1 0 118404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1271
timestamp 1606716760
transform 1 0 117300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1606716760
transform 1 0 115828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1606716760
transform 1 0 116104 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1254
timestamp 1606716760
transform 1 0 115736 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1258
timestamp 1606716760
transform 1 0 116104 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1270
timestamp 1606716760
transform 1 0 117208 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1257
timestamp 1606716760
transform 1 0 116012 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1259
timestamp 1606716760
transform 1 0 116196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1606716760
transform 1 0 114724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__A
timestamp 1606716760
transform 1 0 115276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1246
timestamp 1606716760
transform 1 0 115000 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1246
timestamp 1606716760
transform 1 0 115000 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1251
timestamp 1606716760
transform 1 0 115460 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1235
timestamp 1606716760
transform 1 0 113988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1234
timestamp 1606716760
transform 1 0 113896 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1283
timestamp 1606716760
transform 1 0 118404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1271
timestamp 1606716760
transform 1 0 117300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1606716760
transform 1 0 116104 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1606716760
transform 1 0 115828 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1253
timestamp 1606716760
transform 1 0 115644 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1257
timestamp 1606716760
transform 1 0 116012 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1259
timestamp 1606716760
transform 1 0 116196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1606716760
transform 1 0 114724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1242
timestamp 1606716760
transform 1 0 114632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1245
timestamp 1606716760
transform 1 0 114908 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1234
timestamp 1606716760
transform 1 0 113896 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1272
timestamp 1606716760
transform 1 0 117392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1284
timestamp 1606716760
transform 1 0 118496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1606716760
transform 1 0 117116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1258
timestamp 1606716760
transform 1 0 116104 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1266
timestamp 1606716760
transform 1 0 116840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1246
timestamp 1606716760
transform 1 0 115000 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1234
timestamp 1606716760
transform 1 0 113896 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _611_
timestamp 1606716760
transform 1 0 118312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1606716760
transform 1 0 117760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1274
timestamp 1606716760
transform 1 0 117576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1278
timestamp 1606716760
transform 1 0 117944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1285
timestamp 1606716760
transform 1 0 118588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1606716760
transform 1 0 117300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _612_
timestamp 1606716760
transform 1 0 116196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1606716760
transform 1 0 116104 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1606716760
transform 1 0 117116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__A
timestamp 1606716760
transform 1 0 116656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1254
timestamp 1606716760
transform 1 0 115736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1262
timestamp 1606716760
transform 1 0 116472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1266
timestamp 1606716760
transform 1 0 116840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A
timestamp 1606716760
transform 1 0 114448 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1238
timestamp 1606716760
transform 1 0 114264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1242
timestamp 1606716760
transform 1 0 114632 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1606716760
transform 1 0 114080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1234
timestamp 1606716760
transform 1 0 113896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1606716760
transform 1 0 117668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[52\]_TE
timestamp 1606716760
transform 1 0 118404 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1274
timestamp 1606716760
transform 1 0 117576 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1278
timestamp 1606716760
transform 1 0 117944 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1282
timestamp 1606716760
transform 1 0 118312 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1285
timestamp 1606716760
transform 1 0 118588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1606716760
transform 1 0 116196 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1262
timestamp 1606716760
transform 1 0 116472 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1251
timestamp 1606716760
transform 1 0 115460 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[254\]
timestamp 1606716760
transform 1 0 117392 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[52\]
timestamp 1606716760
transform 1 0 118404 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1606716760
transform 1 0 117852 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[76\]_A
timestamp 1606716760
transform 1 0 118220 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1279
timestamp 1606716760
transform 1 0 118036 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1283
timestamp 1606716760
transform 1 0 118404 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1275
timestamp 1606716760
transform 1 0 117668 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1279
timestamp 1606716760
transform 1 0 118036 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[76\]
timestamp 1606716760
transform 1 0 116380 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1606716760
transform 1 0 116656 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1262
timestamp 1606716760
transform 1 0 116472 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1266
timestamp 1606716760
transform 1 0 116840 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[278\]
timestamp 1606716760
transform 1 0 116196 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1606716760
transform 1 0 116288 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1606716760
transform 1 0 116104 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[50\]_A
timestamp 1606716760
transform 1 0 115736 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[76\]_TE
timestamp 1606716760
transform 1 0 116104 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1256
timestamp 1606716760
transform 1 0 115920 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1253
timestamp 1606716760
transform 1 0 115644 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1257
timestamp 1606716760
transform 1 0 116012 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[252\]
timestamp 1606716760
transform 1 0 115000 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[49\]_A
timestamp 1606716760
transform 1 0 115460 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1252
timestamp 1606716760
transform 1 0 115552 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1238
timestamp 1606716760
transform 1 0 114264 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1249
timestamp 1606716760
transform 1 0 115276 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[50\]
timestamp 1606716760
transform 1 0 113896 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[251\]
timestamp 1606716760
transform 1 0 113988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1220
timestamp 1606716760
transform 1 0 112608 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1232
timestamp 1606716760
transform 1 0 113712 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1606716760
transform 1 0 110860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1606716760
transform 1 0 111320 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1204
timestamp 1606716760
transform 1 0 111136 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1208
timestamp 1606716760
transform 1 0 111504 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1606716760
transform 1 0 110492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1198
timestamp 1606716760
transform 1 0 110584 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1185
timestamp 1606716760
transform 1 0 109388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1606716760
transform 1 0 113252 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1221
timestamp 1606716760
transform 1 0 112700 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1228
timestamp 1606716760
transform 1 0 113344 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1209
timestamp 1606716760
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1606716760
transform 1 0 110216 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1191
timestamp 1606716760
transform 1 0 109940 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1197
timestamp 1606716760
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1606716760
transform 1 0 113712 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1606716760
transform 1 0 113252 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1226
timestamp 1606716760
transform 1 0 113160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1228
timestamp 1606716760
transform 1 0 113344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1222
timestamp 1606716760
transform 1 0 112792 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1218
timestamp 1606716760
transform 1 0 112424 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1206
timestamp 1606716760
transform 1 0 111320 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1210
timestamp 1606716760
transform 1 0 111688 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1606716760
transform 1 0 110492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1606716760
transform 1 0 110216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1194
timestamp 1606716760
transform 1 0 110216 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1192
timestamp 1606716760
transform 1 0 110032 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1196
timestamp 1606716760
transform 1 0 110400 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1198
timestamp 1606716760
transform 1 0 110584 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1182
timestamp 1606716760
transform 1 0 109112 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1184
timestamp 1606716760
transform 1 0 109296 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1606716760
transform 1 0 113712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1222
timestamp 1606716760
transform 1 0 112792 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1230
timestamp 1606716760
transform 1 0 113528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1210
timestamp 1606716760
transform 1 0 111688 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1606716760
transform 1 0 110492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1193
timestamp 1606716760
transform 1 0 110124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1198
timestamp 1606716760
transform 1 0 110584 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1181
timestamp 1606716760
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1606716760
transform 1 0 113620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1606716760
transform 1 0 113252 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1224
timestamp 1606716760
transform 1 0 112976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1228
timestamp 1606716760
transform 1 0 113344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _609_
timestamp 1606716760
transform 1 0 110860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1204
timestamp 1606716760
transform 1 0 111136 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1216
timestamp 1606716760
transform 1 0 112240 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1606716760
transform 1 0 109572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1186
timestamp 1606716760
transform 1 0 109480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1190
timestamp 1606716760
transform 1 0 109848 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1198
timestamp 1606716760
transform 1 0 110584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1182
timestamp 1606716760
transform 1 0 109112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1606716760
transform 1 0 112608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1606716760
transform 1 0 113620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1606716760
transform 1 0 113068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1223
timestamp 1606716760
transform 1 0 112884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1227
timestamp 1606716760
transform 1 0 113252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1606716760
transform 1 0 111596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1606716760
transform 1 0 111044 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__A
timestamp 1606716760
transform 1 0 111412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1606716760
transform 1 0 112056 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1201
timestamp 1606716760
transform 1 0 110860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1205
timestamp 1606716760
transform 1 0 111228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1212
timestamp 1606716760
transform 1 0 111872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1216
timestamp 1606716760
transform 1 0 112240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1606716760
transform 1 0 110584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1606716760
transform 1 0 110492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1606716760
transform 1 0 109848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1606716760
transform 1 0 110216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1188
timestamp 1606716760
transform 1 0 109664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1192
timestamp 1606716760
transform 1 0 110032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1196
timestamp 1606716760
transform 1 0 110400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1606716760
transform 1 0 109388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1181
timestamp 1606716760
transform 1 0 109020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[49\]
timestamp 1606716760
transform 1 0 113804 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1606716760
transform 1 0 113252 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__A
timestamp 1606716760
transform 1 0 112608 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1222
timestamp 1606716760
transform 1 0 112792 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1226
timestamp 1606716760
transform 1 0 113160 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1228
timestamp 1606716760
transform 1 0 113344 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1232
timestamp 1606716760
transform 1 0 113712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1218
timestamp 1606716760
transform 1 0 112424 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _556_
timestamp 1606716760
transform 1 0 112148 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[85\]_TE
timestamp 1606716760
transform 1 0 111596 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1207
timestamp 1606716760
transform 1 0 111412 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1211
timestamp 1606716760
transform 1 0 111780 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[74\]
timestamp 1606716760
transform 1 0 109756 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1181
timestamp 1606716760
transform 1 0 109020 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[49\]_TE
timestamp 1606716760
transform 1 0 113804 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[50\]_TE
timestamp 1606716760
transform 1 0 113712 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1231
timestamp 1606716760
transform 1 0 113620 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1227
timestamp 1606716760
transform 1 0 113252 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1606716760
transform 1 0 113436 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[85\]_A
timestamp 1606716760
transform 1 0 113436 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1230
timestamp 1606716760
transform 1 0 113528 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1219
timestamp 1606716760
transform 1 0 112516 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[87\]_A
timestamp 1606716760
transform 1 0 112700 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1223
timestamp 1606716760
transform 1 0 112884 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  la_buf\[85\]
timestamp 1606716760
transform 1 0 111596 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[87\]
timestamp 1606716760
transform 1 0 110860 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1606716760
transform 1 0 111044 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[74\]_A
timestamp 1606716760
transform 1 0 111412 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1201
timestamp 1606716760
transform 1 0 110860 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1205
timestamp 1606716760
transform 1 0 111228 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1199
timestamp 1606716760
transform 1 0 110676 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _558_
timestamp 1606716760
transform 1 0 110584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1606716760
transform 1 0 110584 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1606716760
transform 1 0 110492 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[87\]_TE
timestamp 1606716760
transform 1 0 110400 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[159\]
timestamp 1606716760
transform 1 0 109572 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[74\]_TE
timestamp 1606716760
transform 1 0 109940 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1190
timestamp 1606716760
transform 1 0 109848 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1189
timestamp 1606716760
transform 1 0 109756 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1193
timestamp 1606716760
transform 1 0 110124 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1606716760
transform 1 0 108928 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1183
timestamp 1606716760
transform 1 0 109204 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1182
timestamp 1606716760
transform 1 0 109112 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[161\]
timestamp 1606716760
transform 1 0 109480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1173
timestamp 1606716760
transform 1 0 108284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1149
timestamp 1606716760
transform 1 0 106076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1161
timestamp 1606716760
transform 1 0 107180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1606716760
transform 1 0 104880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1135
timestamp 1606716760
transform 1 0 104788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1137
timestamp 1606716760
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1127
timestamp 1606716760
transform 1 0 104052 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1167
timestamp 1606716760
transform 1 0 107732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1179
timestamp 1606716760
transform 1 0 108836 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1606716760
transform 1 0 107640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1165
timestamp 1606716760
transform 1 0 107548 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1149
timestamp 1606716760
transform 1 0 106076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1161
timestamp 1606716760
transform 1 0 107180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1606716760
transform 1 0 105800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1134
timestamp 1606716760
transform 1 0 104696 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1606716760
transform 1 0 107732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1170
timestamp 1606716760
transform 1 0 108008 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1172
timestamp 1606716760
transform 1 0 108192 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1606716760
transform 1 0 107640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1165
timestamp 1606716760
transform 1 0 107548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1606716760
transform 1 0 106536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1153
timestamp 1606716760
transform 1 0 106444 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1157
timestamp 1606716760
transform 1 0 106812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1160
timestamp 1606716760
transform 1 0 107088 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1606716760
transform 1 0 105800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1147
timestamp 1606716760
transform 1 0 105892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1145
timestamp 1606716760
transform 1 0 105708 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1148
timestamp 1606716760
transform 1 0 105984 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1606716760
transform 1 0 104880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1135
timestamp 1606716760
transform 1 0 104788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1137
timestamp 1606716760
transform 1 0 104972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[115\]_A
timestamp 1606716760
transform 1 0 104328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1129
timestamp 1606716760
transform 1 0 104236 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1132
timestamp 1606716760
transform 1 0 104512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1606716760
transform 1 0 107732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1169
timestamp 1606716760
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1164
timestamp 1606716760
transform 1 0 107456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1606716760
transform 1 0 106536 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1149
timestamp 1606716760
transform 1 0 106076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1153
timestamp 1606716760
transform 1 0 106444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1156
timestamp 1606716760
transform 1 0 106720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1606716760
transform 1 0 104880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1134
timestamp 1606716760
transform 1 0 104696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1137
timestamp 1606716760
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1606716760
transform 1 0 107732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1170
timestamp 1606716760
transform 1 0 108008 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1606716760
transform 1 0 107640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1165
timestamp 1606716760
transform 1 0 107548 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1157
timestamp 1606716760
transform 1 0 106812 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1145
timestamp 1606716760
transform 1 0 105708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[163\]
timestamp 1606716760
transform 1 0 104328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1133
timestamp 1606716760
transform 1 0 104604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1606716760
transform 1 0 108376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1606716760
transform 1 0 107732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1606716760
transform 1 0 108836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1169
timestamp 1606716760
transform 1 0 107916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1173
timestamp 1606716760
transform 1 0 108284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1177
timestamp 1606716760
transform 1 0 108652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1164
timestamp 1606716760
transform 1 0 107456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1152
timestamp 1606716760
transform 1 0 106352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[272\]
timestamp 1606716760
transform 1 0 104972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1606716760
transform 1 0 104880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1140
timestamp 1606716760
transform 1 0 105248 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1606716760
transform 1 0 104144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1130
timestamp 1606716760
transform 1 0 104328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1606716760
transform 1 0 107732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1606716760
transform 1 0 108744 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1170
timestamp 1606716760
transform 1 0 108008 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1606716760
transform 1 0 107640 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1164
timestamp 1606716760
transform 1 0 107456 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1606716760
transform 1 0 106444 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1156
timestamp 1606716760
transform 1 0 106720 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1141
timestamp 1606716760
transform 1 0 105340 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1171
timestamp 1606716760
transform 1 0 108100 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1178
timestamp 1606716760
transform 1 0 108744 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1606716760
transform 1 0 107916 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1606716760
transform 1 0 107732 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1606716760
transform 1 0 107732 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[276\]
timestamp 1606716760
transform 1 0 108468 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[274\]
timestamp 1606716760
transform 1 0 107824 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1166
timestamp 1606716760
transform 1 0 107640 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[83\]_A
timestamp 1606716760
transform 1 0 107180 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1162
timestamp 1606716760
transform 1 0 107272 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1163
timestamp 1606716760
transform 1 0 107364 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1606716760
transform 1 0 106812 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1155
timestamp 1606716760
transform 1 0 106628 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[157\]
timestamp 1606716760
transform 1 0 106996 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1159
timestamp 1606716760
transform 1 0 106996 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1151
timestamp 1606716760
transform 1 0 106260 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A
timestamp 1606716760
transform 1 0 106444 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _554_
timestamp 1606716760
transform 1 0 105984 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[89\]_A
timestamp 1606716760
transform 1 0 105800 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[83\]
timestamp 1606716760
transform 1 0 105340 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _552_
timestamp 1606716760
transform 1 0 104972 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1606716760
transform 1 0 104880 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1606716760
transform 1 0 104880 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A
timestamp 1606716760
transform 1 0 105432 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[83\]_TE
timestamp 1606716760
transform 1 0 105156 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1137
timestamp 1606716760
transform 1 0 104972 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1140
timestamp 1606716760
transform 1 0 105248 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1144
timestamp 1606716760
transform 1 0 105616 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1130
timestamp 1606716760
transform 1 0 104328 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1130
timestamp 1606716760
transform 1 0 104328 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[70\]_TE
timestamp 1606716760
transform 1 0 104512 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[89\]_TE
timestamp 1606716760
transform 1 0 104512 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[70\]_A
timestamp 1606716760
transform 1 0 104144 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[81\]_A
timestamp 1606716760
transform 1 0 104144 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1134
timestamp 1606716760
transform 1 0 104696 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1134
timestamp 1606716760
transform 1 0 104696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1115
timestamp 1606716760
transform 1 0 102948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__A
timestamp 1606716760
transform 1 0 102764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1111
timestamp 1606716760
transform 1 0 102580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _599_
timestamp 1606716760
transform 1 0 102304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606716760
transform 1 0 102028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[115\]
timestamp 1606716760
transform 1 0 103040 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606716760
transform 1 0 102028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1108
timestamp 1606716760
transform 1 0 102304 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[115\]_TE
timestamp 1606716760
transform 1 0 103316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1123
timestamp 1606716760
transform 1 0 103684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1117
timestamp 1606716760
transform 1 0 103132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1121
timestamp 1606716760
transform 1 0 103500 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[317\]
timestamp 1606716760
transform 1 0 102856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1111
timestamp 1606716760
transform 1 0 102580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp 1606716760
transform 1 0 102304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606716760
transform 1 0 102028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606716760
transform 1 0 102028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1108
timestamp 1606716760
transform 1 0 102304 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[155\]
timestamp 1606716760
transform 1 0 103316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__A
timestamp 1606716760
transform 1 0 103132 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1115
timestamp 1606716760
transform 1 0 102948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1122
timestamp 1606716760
transform 1 0 103592 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__563__A
timestamp 1606716760
transform 1 0 102764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1111
timestamp 1606716760
transform 1 0 102580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _563_
timestamp 1606716760
transform 1 0 102304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606716760
transform 1 0 102028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _560_
timestamp 1606716760
transform 1 0 103316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[72\]_A
timestamp 1606716760
transform 1 0 103776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[72\]_TE
timestamp 1606716760
transform 1 0 103132 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1115
timestamp 1606716760
transform 1 0 102948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1122
timestamp 1606716760
transform 1 0 103592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1126
timestamp 1606716760
transform 1 0 103960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A
timestamp 1606716760
transform 1 0 102764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1111
timestamp 1606716760
transform 1 0 102580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _547_
timestamp 1606716760
transform 1 0 102304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606716760
transform 1 0 102028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1126
timestamp 1606716760
transform 1 0 103960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[72\]
timestamp 1606716760
transform 1 0 102304 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606716760
transform 1 0 102028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[89\]
timestamp 1606716760
transform 1 0 103684 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[81\]_TE
timestamp 1606716760
transform 1 0 103132 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1115
timestamp 1606716760
transform 1 0 102948 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1119
timestamp 1606716760
transform 1 0 103316 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__A
timestamp 1606716760
transform 1 0 102764 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1111
timestamp 1606716760
transform 1 0 102580 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1606716760
transform 1 0 102304 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606716760
transform 1 0 102028 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1126
timestamp 1606716760
transform 1 0 103960 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1126
timestamp 1606716760
transform 1 0 103960 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[81\]
timestamp 1606716760
transform 1 0 102304 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[70\]
timestamp 1606716760
transform 1 0 102304 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606716760
transform 1 0 102028 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606716760
transform 1 0 102028 0 1 1088
box -38 -48 314 592
use mgmt_protect_hv  powergood_check
timestamp 1606716760
transform 1 0 95062 0 1 1121
box 0 0 4932 5000
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606716760
transform -1 0 93012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_996
timestamp 1606716760
transform 1 0 92000 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[150\]
timestamp 1606716760
transform 1 0 91724 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[112\]_A
timestamp 1606716760
transform 1 0 91540 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_985
timestamp 1606716760
transform 1 0 90988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[164\]
timestamp 1606716760
transform 1 0 90712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[112\]_TE
timestamp 1606716760
transform 1 0 90252 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_979
timestamp 1606716760
transform 1 0 90436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[109\]_A
timestamp 1606716760
transform 1 0 89332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_969
timestamp 1606716760
transform 1 0 89516 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606716760
transform -1 0 93012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_996
timestamp 1606716760
transform 1 0 92000 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _561_
timestamp 1606716760
transform 1 0 91724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_985
timestamp 1606716760
transform 1 0 90988 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _543_
timestamp 1606716760
transform 1 0 90712 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[113\]_A
timestamp 1606716760
transform 1 0 90436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_977
timestamp 1606716760
transform 1 0 90252 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_981
timestamp 1606716760
transform 1 0 90620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1606716760
transform 1 0 90160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[110\]_A
timestamp 1606716760
transform 1 0 89608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_968
timestamp 1606716760
transform 1 0 89424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_972
timestamp 1606716760
transform 1 0 89792 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606716760
transform -1 0 93012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606716760
transform -1 0 93012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1606716760
transform 1 0 92552 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1606716760
transform 1 0 91724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_996
timestamp 1606716760
transform 1 0 92000 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1606716760
transform 1 0 91724 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A
timestamp 1606716760
transform 1 0 92184 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_996
timestamp 1606716760
transform 1 0 92000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1000
timestamp 1606716760
transform 1 0 92368 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_984
timestamp 1606716760
transform 1 0 90896 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_992
timestamp 1606716760
transform 1 0 91632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_992
timestamp 1606716760
transform 1 0 91632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _541_
timestamp 1606716760
transform 1 0 90252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1606716760
transform 1 0 90712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_980
timestamp 1606716760
transform 1 0 90528 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_979
timestamp 1606716760
transform 1 0 90436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606716760
transform 1 0 90160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_968
timestamp 1606716760
transform 1 0 89424 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606716760
transform -1 0 93012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1606716760
transform 1 0 92552 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1000
timestamp 1606716760
transform 1 0 92368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_996
timestamp 1606716760
transform 1 0 92000 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1606716760
transform 1 0 92184 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1606716760
transform 1 0 91724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_985
timestamp 1606716760
transform 1 0 90988 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _540_
timestamp 1606716760
transform 1 0 90344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__A
timestamp 1606716760
transform 1 0 90804 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_981
timestamp 1606716760
transform 1 0 90620 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _538_
timestamp 1606716760
transform 1 0 89332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__538__A
timestamp 1606716760
transform 1 0 89792 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__A
timestamp 1606716760
transform 1 0 90160 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_970
timestamp 1606716760
transform 1 0 89608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_974
timestamp 1606716760
transform 1 0 89976 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606716760
transform -1 0 93012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1000
timestamp 1606716760
transform 1 0 92368 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_996
timestamp 1606716760
transform 1 0 92000 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[90\]_A
timestamp 1606716760
transform 1 0 92184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[90\]
timestamp 1606716760
transform 1 0 90344 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_4_977
timestamp 1606716760
transform 1 0 90252 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606716760
transform 1 0 90160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_971
timestamp 1606716760
transform 1 0 89700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_975
timestamp 1606716760
transform 1 0 90068 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606716760
transform -1 0 93012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1000
timestamp 1606716760
transform 1 0 92368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_996
timestamp 1606716760
transform 1 0 92000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[7\]_A
timestamp 1606716760
transform 1 0 92184 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[7\]
timestamp 1606716760
transform 1 0 90344 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[90\]_TE
timestamp 1606716760
transform 1 0 90160 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[7\]_TE
timestamp 1606716760
transform 1 0 89792 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_971
timestamp 1606716760
transform 1 0 89700 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_974
timestamp 1606716760
transform 1 0 89976 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606716760
transform -1 0 93012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_996
timestamp 1606716760
transform 1 0 92000 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[76\]
timestamp 1606716760
transform 1 0 90344 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_2_977
timestamp 1606716760
transform 1 0 90252 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606716760
transform 1 0 90160 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1003
timestamp 1606716760
transform 1 0 92644 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606716760
transform -1 0 93012 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606716760
transform -1 0 93012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1000
timestamp 1606716760
transform 1 0 92368 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_999
timestamp 1606716760
transform 1 0 92276 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__A
timestamp 1606716760
transform 1 0 92184 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[76\]_A
timestamp 1606716760
transform 1 0 92092 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_996
timestamp 1606716760
transform 1 0 92000 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_995
timestamp 1606716760
transform 1 0 91908 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_991
timestamp 1606716760
transform 1 0 91540 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _478_
timestamp 1606716760
transform 1 0 91724 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1606716760
transform 1 0 91632 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__536__A
timestamp 1606716760
transform 1 0 91724 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_984
timestamp 1606716760
transform 1 0 90896 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[76\]_TE
timestamp 1606716760
transform 1 0 91080 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _536_
timestamp 1606716760
transform 1 0 91264 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__A
timestamp 1606716760
transform 1 0 90344 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[58\]_A
timestamp 1606716760
transform 1 0 90712 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_980
timestamp 1606716760
transform 1 0 90528 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_980
timestamp 1606716760
transform 1 0 90528 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _529_
timestamp 1606716760
transform 1 0 89884 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__A
timestamp 1606716760
transform 1 0 89332 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_969
timestamp 1606716760
transform 1 0 89516 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_976
timestamp 1606716760
transform 1 0 90160 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_965
timestamp 1606716760
transform 1 0 89148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[109\]
timestamp 1606716760
transform 1 0 87492 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1606716760
transform 1 0 87400 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_934
timestamp 1606716760
transform 1 0 86296 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_922
timestamp 1606716760
transform 1 0 85192 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[110\]
timestamp 1606716760
transform 1 0 87768 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_942
timestamp 1606716760
transform 1 0 87032 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[315\]
timestamp 1606716760
transform 1 0 86756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_936
timestamp 1606716760
transform 1 0 86480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_928
timestamp 1606716760
transform 1 0 85744 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1606716760
transform 1 0 84548 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_916
timestamp 1606716760
transform 1 0 84640 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[113\]
timestamp 1606716760
transform 1 0 88780 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[113\]_TE
timestamp 1606716760
transform 1 0 88596 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _545_
timestamp 1606716760
transform 1 0 89148 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[132\]
timestamp 1606716760
transform 1 0 88136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[312\]
timestamp 1606716760
transform 1 0 87768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_oen_buffers\[110\]_TE
timestamp 1606716760
transform 1 0 88228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_952
timestamp 1606716760
transform 1 0 87952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_957
timestamp 1606716760
transform 1 0 88412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_953
timestamp 1606716760
transform 1 0 88044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_957
timestamp 1606716760
transform 1 0 88412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_940
timestamp 1606716760
transform 1 0 86848 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_947
timestamp 1606716760
transform 1 0 87492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606716760
transform 1 0 87400 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_934
timestamp 1606716760
transform 1 0 86296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_928
timestamp 1606716760
transform 1 0 85744 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606716760
transform 1 0 84548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_916
timestamp 1606716760
transform 1 0 84640 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_922
timestamp 1606716760
transform 1 0 85192 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__A
timestamp 1606716760
transform 1 0 89148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__A
timestamp 1606716760
transform 1 0 88688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_962
timestamp 1606716760
transform 1 0 88872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _549_
timestamp 1606716760
transform 1 0 88228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_958
timestamp 1606716760
transform 1 0 88504 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606716760
transform 1 0 87400 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_947
timestamp 1606716760
transform 1 0 87492 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_934
timestamp 1606716760
transform 1 0 86296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_922
timestamp 1606716760
transform 1 0 85192 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_959
timestamp 1606716760
transform 1 0 88596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _534_
timestamp 1606716760
transform 1 0 88320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _565_
timestamp 1606716760
transform 1 0 87308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_948
timestamp 1606716760
transform 1 0 87584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[148\]
timestamp 1606716760
transform 1 0 86296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_937
timestamp 1606716760
transform 1 0 86572 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_928
timestamp 1606716760
transform 1 0 85744 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606716760
transform 1 0 84548 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_914
timestamp 1606716760
transform 1 0 84456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_916
timestamp 1606716760
transform 1 0 84640 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__A
timestamp 1606716760
transform 1 0 88964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_961
timestamp 1606716760
transform 1 0 88780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_965
timestamp 1606716760
transform 1 0 89148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__A
timestamp 1606716760
transform 1 0 88320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _532_
timestamp 1606716760
transform 1 0 88504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_954
timestamp 1606716760
transform 1 0 88136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__A
timestamp 1606716760
transform 1 0 87952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_950
timestamp 1606716760
transform 1 0 87768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _527_
timestamp 1606716760
transform 1 0 87492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1606716760
transform 1 0 87216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606716760
transform 1 0 87400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_942
timestamp 1606716760
transform 1 0 87032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A
timestamp 1606716760
transform 1 0 86848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _567_
timestamp 1606716760
transform 1 0 86388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_938
timestamp 1606716760
transform 1 0 86664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_927
timestamp 1606716760
transform 1 0 85652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[81\]
timestamp 1606716760
transform 1 0 85376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_921
timestamp 1606716760
transform 1 0 85100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[58\]_TE
timestamp 1606716760
transform 1 0 88872 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_964
timestamp 1606716760
transform 1 0 89056 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_958
timestamp 1606716760
transform 1 0 88504 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[74\]
timestamp 1606716760
transform 1 0 86848 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_2_938
timestamp 1606716760
transform 1 0 86664 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _520_
timestamp 1606716760
transform 1 0 85652 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_930
timestamp 1606716760
transform 1 0 85928 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _487_
timestamp 1606716760
transform 1 0 84640 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606716760
transform 1 0 84548 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[92\]_A
timestamp 1606716760
transform 1 0 84272 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_914
timestamp 1606716760
transform 1 0 84456 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_919
timestamp 1606716760
transform 1 0 84916 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[58\]
timestamp 1606716760
transform 1 0 88872 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_0_965
timestamp 1606716760
transform 1 0 89148 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1606716760
transform 1 0 88780 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _525_
timestamp 1606716760
transform 1 0 88872 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__A
timestamp 1606716760
transform 1 0 87952 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__A
timestamp 1606716760
transform 1 0 87860 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[74\]_A
timestamp 1606716760
transform 1 0 88320 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_953
timestamp 1606716760
transform 1 0 88044 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_950
timestamp 1606716760
transform 1 0 87768 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_954
timestamp 1606716760
transform 1 0 88136 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_958
timestamp 1606716760
transform 1 0 88504 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_949
timestamp 1606716760
transform 1 0 87676 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1606716760
transform 1 0 87400 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _523_
timestamp 1606716760
transform 1 0 87492 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606716760
transform 1 0 87400 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__A
timestamp 1606716760
transform 1 0 86848 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[74\]_TE
timestamp 1606716760
transform 1 0 87216 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_942
timestamp 1606716760
transform 1 0 87032 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _516_
timestamp 1606716760
transform 1 0 86020 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__A
timestamp 1606716760
transform 1 0 86204 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_931
timestamp 1606716760
transform 1 0 86020 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _521_
timestamp 1606716760
transform 1 0 86388 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__A
timestamp 1606716760
transform 1 0 86480 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_934
timestamp 1606716760
transform 1 0 86296 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_938
timestamp 1606716760
transform 1 0 86664 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_938
timestamp 1606716760
transform 1 0 86664 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_918
timestamp 1606716760
transform 1 0 84824 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _518_
timestamp 1606716760
transform 1 0 85376 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1606716760
transform 1 0 85928 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__A
timestamp 1606716760
transform 1 0 85836 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_927
timestamp 1606716760
transform 1 0 85652 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_920
timestamp 1606716760
transform 1 0 85008 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_916
timestamp 1606716760
transform 1 0 84640 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_914
timestamp 1606716760
transform 1 0 84456 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__A
timestamp 1606716760
transform 1 0 84640 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__A
timestamp 1606716760
transform 1 0 84824 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_910
timestamp 1606716760
transform 1 0 84088 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_898
timestamp 1606716760
transform 1 0 82984 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1606716760
transform 1 0 81788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_886
timestamp 1606716760
transform 1 0 81880 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_861
timestamp 1606716760
transform 1 0 79580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_873
timestamp 1606716760
transform 1 0 80684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_903
timestamp 1606716760
transform 1 0 83444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_891
timestamp 1606716760
transform 1 0 82340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_879
timestamp 1606716760
transform 1 0 81236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_867
timestamp 1606716760
transform 1 0 80132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_910
timestamp 1606716760
transform 1 0 84088 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_903
timestamp 1606716760
transform 1 0 83444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_898
timestamp 1606716760
transform 1 0 82984 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_891
timestamp 1606716760
transform 1 0 82340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606716760
transform 1 0 81788 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_879
timestamp 1606716760
transform 1 0 81236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_886
timestamp 1606716760
transform 1 0 81880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_867
timestamp 1606716760
transform 1 0 80132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_861
timestamp 1606716760
transform 1 0 79580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_873
timestamp 1606716760
transform 1 0 80684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_910
timestamp 1606716760
transform 1 0 84088 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_898
timestamp 1606716760
transform 1 0 82984 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606716760
transform 1 0 81788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_886
timestamp 1606716760
transform 1 0 81880 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_861
timestamp 1606716760
transform 1 0 79580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_873
timestamp 1606716760
transform 1 0 80684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[166\]
timestamp 1606716760
transform 1 0 83076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_898
timestamp 1606716760
transform 1 0 82984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_902
timestamp 1606716760
transform 1 0 83352 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_890
timestamp 1606716760
transform 1 0 82248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_878
timestamp 1606716760
transform 1 0 81144 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[339\]
timestamp 1606716760
transform 1 0 80868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_867
timestamp 1606716760
transform 1 0 80132 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__A
timestamp 1606716760
transform 1 0 83812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_909
timestamp 1606716760
transform 1 0 83996 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _511_
timestamp 1606716760
transform 1 0 83352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_901
timestamp 1606716760
transform 1 0 83260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_905
timestamp 1606716760
transform 1 0 83628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__A
timestamp 1606716760
transform 1 0 82340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_889
timestamp 1606716760
transform 1 0 82156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_893
timestamp 1606716760
transform 1 0 82524 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 1606716760
transform 1 0 81880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606716760
transform 1 0 81788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__A
timestamp 1606716760
transform 1 0 81144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_880
timestamp 1606716760
transform 1 0 81328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_884
timestamp 1606716760
transform 1 0 81696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_876
timestamp 1606716760
transform 1 0 80960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _501_
timestamp 1606716760
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_861
timestamp 1606716760
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[428\]
timestamp 1606716760
transform 1 0 79304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__A
timestamp 1606716760
transform 1 0 83812 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_909
timestamp 1606716760
transform 1 0 83996 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _514_
timestamp 1606716760
transform 1 0 83352 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[92\]_TE
timestamp 1606716760
transform 1 0 82984 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_900
timestamp 1606716760
transform 1 0 83168 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_905
timestamp 1606716760
transform 1 0 83628 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _504_
timestamp 1606716760
transform 1 0 82156 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_892
timestamp 1606716760
transform 1 0 82432 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_881
timestamp 1606716760
transform 1 0 81420 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[9\]
timestamp 1606716760
transform 1 0 80592 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_862
timestamp 1606716760
transform 1 0 79672 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_870
timestamp 1606716760
transform 1 0 80408 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[98\]_B
timestamp 1606716760
transform 1 0 79488 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_858
timestamp 1606716760
transform 1 0 79304 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _512_
timestamp 1606716760
transform 1 0 84180 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_907
timestamp 1606716760
transform 1 0 83812 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[92\]
timestamp 1606716760
transform 1 0 82984 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_1_897
timestamp 1606716760
transform 1 0 82892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_903
timestamp 1606716760
transform 1 0 83444 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__A
timestamp 1606716760
transform 1 0 83628 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1606716760
transform 1 0 83076 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _509_
timestamp 1606716760
transform 1 0 83168 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__A
timestamp 1606716760
transform 1 0 82708 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__A
timestamp 1606716760
transform 1 0 82524 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_895
timestamp 1606716760
transform 1 0 82708 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_893
timestamp 1606716760
transform 1 0 82524 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1606716760
transform 1 0 82064 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__A
timestamp 1606716760
transform 1 0 82340 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_891
timestamp 1606716760
transform 1 0 82340 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_889
timestamp 1606716760
transform 1 0 82156 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_884
timestamp 1606716760
transform 1 0 81696 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[9\]_B
timestamp 1606716760
transform 1 0 81604 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[9\]_A
timestamp 1606716760
transform 1 0 81512 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606716760
transform 1 0 81788 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 1606716760
transform 1 0 81880 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_881
timestamp 1606716760
transform 1 0 81420 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_880
timestamp 1606716760
transform 1 0 81328 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[9\]_A
timestamp 1606716760
transform 1 0 81236 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[9\]
timestamp 1606716760
transform 1 0 80500 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _503_
timestamp 1606716760
transform 1 0 80592 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1606716760
transform 1 0 80224 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__A
timestamp 1606716760
transform 1 0 80408 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_869
timestamp 1606716760
transform 1 0 80316 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_868
timestamp 1606716760
transform 1 0 80224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_875
timestamp 1606716760
transform 1 0 80868 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_860
timestamp 1606716760
transform 1 0 79488 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[98\]_A
timestamp 1606716760
transform 1 0 80040 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[98\]_A
timestamp 1606716760
transform 1 0 79672 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_864
timestamp 1606716760
transform 1 0 79856 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_864
timestamp 1606716760
transform 1 0 79856 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_849
timestamp 1606716760
transform 1 0 78476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_837
timestamp 1606716760
transform 1 0 77372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1606716760
transform 1 0 76176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_825
timestamp 1606716760
transform 1 0 76268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_808
timestamp 1606716760
transform 1 0 74704 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_820
timestamp 1606716760
transform 1 0 75808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1606716760
transform 1 0 78936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_855
timestamp 1606716760
transform 1 0 79028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_842
timestamp 1606716760
transform 1 0 77832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_830
timestamp 1606716760
transform 1 0 76728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_806
timestamp 1606716760
transform 1 0 74520 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_818
timestamp 1606716760
transform 1 0 75624 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606716760
transform 1 0 78936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_855
timestamp 1606716760
transform 1 0 79028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_849
timestamp 1606716760
transform 1 0 78476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_842
timestamp 1606716760
transform 1 0 77832 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_837
timestamp 1606716760
transform 1 0 77372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606716760
transform 1 0 76176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_830
timestamp 1606716760
transform 1 0 76728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_825
timestamp 1606716760
transform 1 0 76268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_806
timestamp 1606716760
transform 1 0 74520 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_818
timestamp 1606716760
transform 1 0 75624 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_812
timestamp 1606716760
transform 1 0 75072 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_849
timestamp 1606716760
transform 1 0 78476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_837
timestamp 1606716760
transform 1 0 77372 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606716760
transform 1 0 76176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_825
timestamp 1606716760
transform 1 0 76268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_812
timestamp 1606716760
transform 1 0 75072 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606716760
transform 1 0 78936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_850
timestamp 1606716760
transform 1 0 78568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_855
timestamp 1606716760
transform 1 0 79028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[426\]
timestamp 1606716760
transform 1 0 77188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_838
timestamp 1606716760
transform 1 0 77464 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[168\]
timestamp 1606716760
transform 1 0 76176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[96\]_B
timestamp 1606716760
transform 1 0 76636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_827
timestamp 1606716760
transform 1 0 76452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_831
timestamp 1606716760
transform 1 0 76820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[424\]
timestamp 1606716760
transform 1 0 74428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_808
timestamp 1606716760
transform 1 0 74704 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_820
timestamp 1606716760
transform 1 0 75808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_850
timestamp 1606716760
transform 1 0 78568 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[96\]_A
timestamp 1606716760
transform 1 0 77280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_838
timestamp 1606716760
transform 1 0 77464 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[96\]
timestamp 1606716760
transform 1 0 76268 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606716760
transform 1 0 76176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_834
timestamp 1606716760
transform 1 0 77096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_821
timestamp 1606716760
transform 1 0 75900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _500_
timestamp 1606716760
transform 1 0 74520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__A
timestamp 1606716760
transform 1 0 74980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_805
timestamp 1606716760
transform 1 0 74428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_809
timestamp 1606716760
transform 1 0 74796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_813
timestamp 1606716760
transform 1 0 75164 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _473_
timestamp 1606716760
transform 1 0 79028 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606716760
transform 1 0 78936 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_853
timestamp 1606716760
transform 1 0 78844 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[94\]_A
timestamp 1606716760
transform 1 0 77924 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_845
timestamp 1606716760
transform 1 0 78108 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _497_
timestamp 1606716760
transform 1 0 77464 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_841
timestamp 1606716760
transform 1 0 77740 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[78\]_A
timestamp 1606716760
transform 1 0 76912 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_830
timestamp 1606716760
transform 1 0 76728 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_834
timestamp 1606716760
transform 1 0 77096 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[78\]
timestamp 1606716760
transform 1 0 75072 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_2_809
timestamp 1606716760
transform 1 0 74796 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[98\]
timestamp 1606716760
transform 1 0 78660 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[98\]
timestamp 1606716760
transform 1 0 79028 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__A
timestamp 1606716760
transform 1 0 78844 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A
timestamp 1606716760
transform 1 0 78108 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__A
timestamp 1606716760
transform 1 0 77924 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_845
timestamp 1606716760
transform 1 0 78108 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_843
timestamp 1606716760
transform 1 0 77924 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_847
timestamp 1606716760
transform 1 0 78292 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _499_
timestamp 1606716760
transform 1 0 77464 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1606716760
transform 1 0 77372 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_841
timestamp 1606716760
transform 1 0 77740 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[94\]
timestamp 1606716760
transform 1 0 76268 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606716760
transform 1 0 76176 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[96\]_A
timestamp 1606716760
transform 1 0 76820 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_829
timestamp 1606716760
transform 1 0 76636 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_833
timestamp 1606716760
transform 1 0 77004 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[96\]
timestamp 1606716760
transform 1 0 75808 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_1_815
timestamp 1606716760
transform 1 0 75348 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_821
timestamp 1606716760
transform 1 0 75900 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[94\]_TE
timestamp 1606716760
transform 1 0 75992 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[152\]
timestamp 1606716760
transform 1 0 74796 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1606716760
transform 1 0 74520 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[5\]_A
timestamp 1606716760
transform 1 0 74796 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_805
timestamp 1606716760
transform 1 0 74428 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_807
timestamp 1606716760
transform 1 0 74612 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_807
timestamp 1606716760
transform 1 0 74612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_811
timestamp 1606716760
transform 1 0 74980 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[78\]_TE
timestamp 1606716760
transform 1 0 75164 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_812
timestamp 1606716760
transform 1 0 75072 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_796
timestamp 1606716760
transform 1 0 73600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_784
timestamp 1606716760
transform 1 0 72496 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[27\]_A
timestamp 1606716760
transform 1 0 71208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_772
timestamp 1606716760
transform 1 0 71392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1606716760
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_758
timestamp 1606716760
transform 1 0 70104 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_762
timestamp 1606716760
transform 1 0 70472 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_764
timestamp 1606716760
transform 1 0 70656 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[27\]_TE
timestamp 1606716760
transform 1 0 69920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_755
timestamp 1606716760
transform 1 0 69828 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1606716760
transform 1 0 73324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_794
timestamp 1606716760
transform 1 0 73416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_781
timestamp 1606716760
transform 1 0 72220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_757
timestamp 1606716760
transform 1 0 70012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_769
timestamp 1606716760
transform 1 0 71116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606716760
transform 1 0 73324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_794
timestamp 1606716760
transform 1 0 73416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_800
timestamp 1606716760
transform 1 0 73968 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_788
timestamp 1606716760
transform 1 0 72864 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _598_
timestamp 1606716760
transform 1 0 71944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_770
timestamp 1606716760
transform 1 0 71208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_781
timestamp 1606716760
transform 1 0 72220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_776
timestamp 1606716760
transform 1 0 71760 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _595_
timestamp 1606716760
transform 1 0 70932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606716760
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_759
timestamp 1606716760
transform 1 0 70196 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_764
timestamp 1606716760
transform 1 0 70656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _594_
timestamp 1606716760
transform 1 0 69920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_754
timestamp 1606716760
transform 1 0 69736 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_751
timestamp 1606716760
transform 1 0 69460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[79\]
timestamp 1606716760
transform 1 0 73692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__597__A
timestamp 1606716760
transform 1 0 73140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_789
timestamp 1606716760
transform 1 0 72956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_793
timestamp 1606716760
transform 1 0 73324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_800
timestamp 1606716760
transform 1 0 73968 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _597_
timestamp 1606716760
transform 1 0 72680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__A
timestamp 1606716760
transform 1 0 72496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_782
timestamp 1606716760
transform 1 0 72312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _498_
timestamp 1606716760
transform 1 0 71668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__A
timestamp 1606716760
transform 1 0 72128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__A
timestamp 1606716760
transform 1 0 71484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_771
timestamp 1606716760
transform 1 0 71300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_778
timestamp 1606716760
transform 1 0 71944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _517_
timestamp 1606716760
transform 1 0 70656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606716760
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__595__A
timestamp 1606716760
transform 1 0 71116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_758
timestamp 1606716760
transform 1 0 70104 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_762
timestamp 1606716760
transform 1 0 70472 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_767
timestamp 1606716760
transform 1 0 70932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__594__A
timestamp 1606716760
transform 1 0 69920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_752
timestamp 1606716760
transform 1 0 69552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _494_
timestamp 1606716760
transform 1 0 73416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606716760
transform 1 0 73324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_792
timestamp 1606716760
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_797
timestamp 1606716760
transform 1 0 73692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_788
timestamp 1606716760
transform 1 0 72864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _489_
timestamp 1606716760
transform 1 0 71484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_776
timestamp 1606716760
transform 1 0 71760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _496_
timestamp 1606716760
transform 1 0 70472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_765
timestamp 1606716760
transform 1 0 70748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _491_
timestamp 1606716760
transform 1 0 69460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_754
timestamp 1606716760
transform 1 0 69736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1606716760
transform 1 0 74244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _490_
timestamp 1606716760
transform 1 0 73416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__A
timestamp 1606716760
transform 1 0 73876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_791
timestamp 1606716760
transform 1 0 73140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_797
timestamp 1606716760
transform 1 0 73692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_801
timestamp 1606716760
transform 1 0 74060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_783
timestamp 1606716760
transform 1 0 72404 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _484_
timestamp 1606716760
transform 1 0 71760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__A
timestamp 1606716760
transform 1 0 72220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__A
timestamp 1606716760
transform 1 0 71484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_771
timestamp 1606716760
transform 1 0 71300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_775
timestamp 1606716760
transform 1 0 71668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_779
timestamp 1606716760
transform 1 0 72036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_767
timestamp 1606716760
transform 1 0 70932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1606716760
transform 1 0 71116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606716760
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _493_
timestamp 1606716760
transform 1 0 70656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_759
timestamp 1606716760
transform 1 0 70196 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__A
timestamp 1606716760
transform 1 0 70380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_755
timestamp 1606716760
transform 1 0 69828 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__A
timestamp 1606716760
transform 1 0 70012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_751
timestamp 1606716760
transform 1 0 69460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__A
timestamp 1606716760
transform 1 0 69644 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1606716760
transform 1 0 73416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606716760
transform 1 0 73324 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__A
timestamp 1606716760
transform 1 0 73876 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[5\]_TE
timestamp 1606716760
transform 1 0 72956 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_791
timestamp 1606716760
transform 1 0 73140 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_797
timestamp 1606716760
transform 1 0 73692 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_801
timestamp 1606716760
transform 1 0 74060 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_785
timestamp 1606716760
transform 1 0 72588 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1606716760
transform 1 0 72312 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[94\]_B
timestamp 1606716760
transform 1 0 71576 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_770
timestamp 1606716760
transform 1 0 71208 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_776
timestamp 1606716760
transform 1 0 71760 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 1606716760
transform 1 0 70932 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_759
timestamp 1606716760
transform 1 0 70196 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1606716760
transform 1 0 69920 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_754
timestamp 1606716760
transform 1 0 69736 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[5\]
timestamp 1606716760
transform 1 0 72956 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[422\]
timestamp 1606716760
transform 1 0 73416 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_790
timestamp 1606716760
transform 1 0 73048 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_797
timestamp 1606716760
transform 1 0 73692 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[94\]
timestamp 1606716760
transform 1 0 71392 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[94\]
timestamp 1606716760
transform 1 0 71852 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_781
timestamp 1606716760
transform 1 0 72220 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_785
timestamp 1606716760
transform 1 0 72588 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_786
timestamp 1606716760
transform 1 0 72680 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[94\]_A
timestamp 1606716760
transform 1 0 72864 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__A
timestamp 1606716760
transform 1 0 72772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[94\]_A
timestamp 1606716760
transform 1 0 72404 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_776
timestamp 1606716760
transform 1 0 71760 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1606716760
transform 1 0 71668 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__A
timestamp 1606716760
transform 1 0 70932 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__A
timestamp 1606716760
transform 1 0 70932 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_765
timestamp 1606716760
transform 1 0 70748 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_769
timestamp 1606716760
transform 1 0 71116 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_769
timestamp 1606716760
transform 1 0 71116 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _593_
timestamp 1606716760
transform 1 0 70472 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_758
timestamp 1606716760
transform 1 0 70104 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_758
timestamp 1606716760
transform 1 0 70104 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_762
timestamp 1606716760
transform 1 0 70472 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606716760
transform 1 0 70564 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_764
timestamp 1606716760
transform 1 0 70656 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_752
timestamp 1606716760
transform 1 0 69552 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_754
timestamp 1606716760
transform 1 0 69736 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[92\]_A
timestamp 1606716760
transform 1 0 69920 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__A
timestamp 1606716760
transform 1 0 69920 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_749
timestamp 1606716760
transform 1 0 69276 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_737
timestamp 1606716760
transform 1 0 68172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_725
timestamp 1606716760
transform 1 0 67068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1606716760
transform 1 0 64952 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[124\]_A
timestamp 1606716760
transform 1 0 65780 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_699
timestamp 1606716760
transform 1 0 64676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_703
timestamp 1606716760
transform 1 0 65044 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_713
timestamp 1606716760
transform 1 0 65964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_745
timestamp 1606716760
transform 1 0 68908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1606716760
transform 1 0 67712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_733
timestamp 1606716760
transform 1 0 67804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_720
timestamp 1606716760
transform 1 0 66608 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_708
timestamp 1606716760
transform 1 0 65504 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _592_
timestamp 1606716760
transform 1 0 68356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_742
timestamp 1606716760
transform 1 0 68632 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_739
timestamp 1606716760
transform 1 0 68356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606716760
transform 1 0 67712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_733
timestamp 1606716760
transform 1 0 67804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_722
timestamp 1606716760
transform 1 0 66792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_730
timestamp 1606716760
transform 1 0 67528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_727
timestamp 1606716760
transform 1 0 67252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606716760
transform 1 0 64952 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_698
timestamp 1606716760
transform 1 0 64584 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_710
timestamp 1606716760
transform 1 0 65688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_703
timestamp 1606716760
transform 1 0 65044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_715
timestamp 1606716760
transform 1 0 66148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _515_
timestamp 1606716760
transform 1 0 68908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__A
timestamp 1606716760
transform 1 0 69368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_748
timestamp 1606716760
transform 1 0 69184 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__A
timestamp 1606716760
transform 1 0 67988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__592__A
timestamp 1606716760
transform 1 0 68356 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_737
timestamp 1606716760
transform 1 0 68172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_741
timestamp 1606716760
transform 1 0 68540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_733
timestamp 1606716760
transform 1 0 67804 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _589_
timestamp 1606716760
transform 1 0 67528 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[170\]
timestamp 1606716760
transform 1 0 66516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_722
timestamp 1606716760
transform 1 0 66792 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606716760
transform 1 0 64952 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_703
timestamp 1606716760
transform 1 0 65044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_715
timestamp 1606716760
transform 1 0 66148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _495_
timestamp 1606716760
transform 1 0 68448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_739
timestamp 1606716760
transform 1 0 68356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_743
timestamp 1606716760
transform 1 0 68724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606716760
transform 1 0 67712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_733
timestamp 1606716760
transform 1 0 67804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[135\]
timestamp 1606716760
transform 1 0 66700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_724
timestamp 1606716760
transform 1 0 66976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[420\]
timestamp 1606716760
transform 1 0 65320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_698
timestamp 1606716760
transform 1 0 64584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_709
timestamp 1606716760
transform 1 0 65596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _483_
timestamp 1606716760
transform 1 0 69184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__A
timestamp 1606716760
transform 1 0 68448 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_736
timestamp 1606716760
transform 1 0 68080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_742
timestamp 1606716760
transform 1 0 68632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__A
timestamp 1606716760
transform 1 0 67896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_732
timestamp 1606716760
transform 1 0 67712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _482_
timestamp 1606716760
transform 1 0 67436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1606716760
transform 1 0 66424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__A
timestamp 1606716760
transform 1 0 66884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_721
timestamp 1606716760
transform 1 0 66700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_725
timestamp 1606716760
transform 1 0 67068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[419\]
timestamp 1606716760
transform 1 0 65044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606716760
transform 1 0 64952 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_698
timestamp 1606716760
transform 1 0 64584 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_706
timestamp 1606716760
transform 1 0 65320 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[92\]_A
timestamp 1606716760
transform 1 0 68816 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_746
timestamp 1606716760
transform 1 0 69000 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_742
timestamp 1606716760
transform 1 0 68632 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[92\]
timestamp 1606716760
transform 1 0 67804 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606716760
transform 1 0 67712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 1606716760
transform 1 0 66700 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[61\]_TE
timestamp 1606716760
transform 1 0 67528 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_718
timestamp 1606716760
transform 1 0 66424 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_724
timestamp 1606716760
transform 1 0 66976 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1606716760
transform 1 0 65044 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_702
timestamp 1606716760
transform 1 0 64952 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_706
timestamp 1606716760
transform 1 0 65320 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[92\]
timestamp 1606716760
transform 1 0 68908 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1606716760
transform 1 0 68816 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[61\]_A
timestamp 1606716760
transform 1 0 69368 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_748
timestamp 1606716760
transform 1 0 69184 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[96\]_A
timestamp 1606716760
transform 1 0 68264 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[92\]_B
timestamp 1606716760
transform 1 0 68632 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_736
timestamp 1606716760
transform 1 0 68080 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_740
timestamp 1606716760
transform 1 0 68448 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1606716760
transform 1 0 66516 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[61\]
timestamp 1606716760
transform 1 0 67528 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[96\]
timestamp 1606716760
transform 1 0 66424 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__A
timestamp 1606716760
transform 1 0 66976 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__A
timestamp 1606716760
transform 1 0 67344 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_718
timestamp 1606716760
transform 1 0 66424 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_722
timestamp 1606716760
transform 1 0 66792 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_726
timestamp 1606716760
transform 1 0 67160 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[96\]_TE
timestamp 1606716760
transform 1 0 66240 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_699
timestamp 1606716760
transform 1 0 64676 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1606716760
transform 1 0 65964 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A
timestamp 1606716760
transform 1 0 65504 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__A
timestamp 1606716760
transform 1 0 65872 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_711
timestamp 1606716760
transform 1 0 65780 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_714
timestamp 1606716760
transform 1 0 66056 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_710
timestamp 1606716760
transform 1 0 65688 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_714
timestamp 1606716760
transform 1 0 66056 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _485_
timestamp 1606716760
transform 1 0 65044 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606716760
transform 1 0 64952 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_698
timestamp 1606716760
transform 1 0 64584 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_706
timestamp 1606716760
transform 1 0 65320 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[124\]_TE
timestamp 1606716760
transform 1 0 64492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_696
timestamp 1606716760
transform 1 0 64400 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_690
timestamp 1606716760
transform 1 0 63848 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_678
timestamp 1606716760
transform 1 0 62744 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_666
timestamp 1606716760
transform 1 0 61640 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_654
timestamp 1606716760
transform 1 0 60536 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_696
timestamp 1606716760
transform 1 0 64400 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_684
timestamp 1606716760
transform 1 0 63296 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1606716760
transform 1 0 62100 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_672
timestamp 1606716760
transform 1 0 62192 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_668
timestamp 1606716760
transform 1 0 61824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_656
timestamp 1606716760
transform 1 0 60720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_644
timestamp 1606716760
transform 1 0 59616 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1606716760
transform 1 0 63204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_686
timestamp 1606716760
transform 1 0 63480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_690
timestamp 1606716760
transform 1 0 63848 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_679
timestamp 1606716760
transform 1 0 62836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1606716760
transform 1 0 62192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606716760
transform 1 0 62100 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[47\]_A
timestamp 1606716760
transform 1 0 62652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_675
timestamp 1606716760
transform 1 0 62468 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_678
timestamp 1606716760
transform 1 0 62744 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_666
timestamp 1606716760
transform 1 0 61640 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1606716760
transform 1 0 61088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_659
timestamp 1606716760
transform 1 0 60996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_663
timestamp 1606716760
transform 1 0 61364 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_647
timestamp 1606716760
transform 1 0 59892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_654
timestamp 1606716760
transform 1 0 60536 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_696
timestamp 1606716760
transform 1 0 64400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1606716760
transform 1 0 63756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__A
timestamp 1606716760
transform 1 0 63204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__581__A
timestamp 1606716760
transform 1 0 64216 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_685
timestamp 1606716760
transform 1 0 63388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_692
timestamp 1606716760
transform 1 0 64032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_681
timestamp 1606716760
transform 1 0 63020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[47\]
timestamp 1606716760
transform 1 0 62192 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__A
timestamp 1606716760
transform 1 0 62008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A
timestamp 1606716760
transform 1 0 61640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_664
timestamp 1606716760
transform 1 0 61456 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_668
timestamp 1606716760
transform 1 0 61824 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _591_
timestamp 1606716760
transform 1 0 61180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__A
timestamp 1606716760
transform 1 0 60996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_657
timestamp 1606716760
transform 1 0 60812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_645
timestamp 1606716760
transform 1 0 59708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _596_
timestamp 1606716760
transform 1 0 64308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1606716760
transform 1 0 63296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_683
timestamp 1606716760
transform 1 0 63204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_687
timestamp 1606716760
transform 1 0 63572 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _572_
timestamp 1606716760
transform 1 0 62192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606716760
transform 1 0 62100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_675
timestamp 1606716760
transform 1 0 62468 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_665
timestamp 1606716760
transform 1 0 61548 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[39\]_A
timestamp 1606716760
transform 1 0 61364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_661
timestamp 1606716760
transform 1 0 61180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[87\]
timestamp 1606716760
transform 1 0 60352 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[87\]_B
timestamp 1606716760
transform 1 0 60168 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_648
timestamp 1606716760
transform 1 0 59984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__596__A
timestamp 1606716760
transform 1 0 64400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _579_
timestamp 1606716760
transform 1 0 63572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__A
timestamp 1606716760
transform 1 0 64032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__A
timestamp 1606716760
transform 1 0 63388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_683
timestamp 1606716760
transform 1 0 63204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_690
timestamp 1606716760
transform 1 0 63848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_694
timestamp 1606716760
transform 1 0 64216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__A
timestamp 1606716760
transform 1 0 63020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_679
timestamp 1606716760
transform 1 0 62836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 1606716760
transform 1 0 62560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1606716760
transform 1 0 62192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_674
timestamp 1606716760
transform 1 0 62376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_668
timestamp 1606716760
transform 1 0 61824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[39\]
timestamp 1606716760
transform 1 0 60996 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[87\]_A
timestamp 1606716760
transform 1 0 60812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[37\]_A
timestamp 1606716760
transform 1 0 60444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_651
timestamp 1606716760
transform 1 0 60260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_655
timestamp 1606716760
transform 1 0 60628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_696
timestamp 1606716760
transform 1 0 64400 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _574_
timestamp 1606716760
transform 1 0 63756 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1606716760
transform 1 0 64216 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[90\]_B
timestamp 1606716760
transform 1 0 63572 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_692
timestamp 1606716760
transform 1 0 64032 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_681
timestamp 1606716760
transform 1 0 63020 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[89\]
timestamp 1606716760
transform 1 0 62192 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606716760
transform 1 0 62100 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[63\]_A
timestamp 1606716760
transform 1 0 61548 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_667
timestamp 1606716760
transform 1 0 61732 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_663
timestamp 1606716760
transform 1 0 61364 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[85\]
timestamp 1606716760
transform 1 0 60536 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[83\]_A
timestamp 1606716760
transform 1 0 59984 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[85\]_B
timestamp 1606716760
transform 1 0 60352 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_646
timestamp 1606716760
transform 1 0 59800 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_650
timestamp 1606716760
transform 1 0 60168 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_695
timestamp 1606716760
transform 1 0 64308 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[90\]_A
timestamp 1606716760
transform 1 0 64492 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[90\]_A
timestamp 1606716760
transform 1 0 64400 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[90\]
timestamp 1606716760
transform 1 0 63388 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[90\]
timestamp 1606716760
transform 1 0 63480 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_694
timestamp 1606716760
transform 1 0 64216 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_683
timestamp 1606716760
transform 1 0 63204 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[89\]_B
timestamp 1606716760
transform 1 0 63204 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1606716760
transform 1 0 63112 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_681
timestamp 1606716760
transform 1 0 63020 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_680
timestamp 1606716760
transform 1 0 62928 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[89\]_A
timestamp 1606716760
transform 1 0 62836 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_672
timestamp 1606716760
transform 1 0 62192 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_677
timestamp 1606716760
transform 1 0 62652 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[417\]
timestamp 1606716760
transform 1 0 61916 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[89\]
timestamp 1606716760
transform 1 0 61824 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[89\]_A
timestamp 1606716760
transform 1 0 61640 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_665
timestamp 1606716760
transform 1 0 61548 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_664
timestamp 1606716760
transform 1 0 61456 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[85\]_A
timestamp 1606716760
transform 1 0 61272 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[87\]_A
timestamp 1606716760
transform 1 0 61364 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_661
timestamp 1606716760
transform 1 0 61180 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_660
timestamp 1606716760
transform 1 0 61088 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[87\]
timestamp 1606716760
transform 1 0 60352 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1606716760
transform 1 0 60260 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_645
timestamp 1606716760
transform 1 0 59708 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1606716760
transform 1 0 59340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[122\]_A
timestamp 1606716760
transform 1 0 58972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[46\]_A
timestamp 1606716760
transform 1 0 58604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_631
timestamp 1606716760
transform 1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_635
timestamp 1606716760
transform 1 0 58788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_639
timestamp 1606716760
transform 1 0 59156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_642
timestamp 1606716760
transform 1 0 59432 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[46\]
timestamp 1606716760
transform 1 0 57592 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[45\]_A
timestamp 1606716760
transform 1 0 57040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[122\]_TE
timestamp 1606716760
transform 1 0 57408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1606716760
transform 1 0 56856 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_618
timestamp 1606716760
transform 1 0 57224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[45\]
timestamp 1606716760
transform 1 0 56028 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_601
timestamp 1606716760
transform 1 0 55660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[36\]_A
timestamp 1606716760
transform 1 0 55476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_597
timestamp 1606716760
transform 1 0 55292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_632
timestamp 1606716760
transform 1 0 58512 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_620
timestamp 1606716760
transform 1 0 57408 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[44\]
timestamp 1606716760
transform 1 0 56580 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1606716760
transform 1 0 56488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_598
timestamp 1606716760
transform 1 0 55384 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606716760
transform 1 0 59340 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_635
timestamp 1606716760
transform 1 0 58788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_630
timestamp 1606716760
transform 1 0 58328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_638
timestamp 1606716760
transform 1 0 59064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_642
timestamp 1606716760
transform 1 0 59432 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[44\]_A
timestamp 1606716760
transform 1 0 57040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_623
timestamp 1606716760
transform 1 0 57684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_614
timestamp 1606716760
transform 1 0 56856 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_618
timestamp 1606716760
transform 1 0 57224 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606716760
transform 1 0 56488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[43\]_A
timestamp 1606716760
transform 1 0 56672 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_611
timestamp 1606716760
transform 1 0 56580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_610
timestamp 1606716760
transform 1 0 56488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[43\]
timestamp 1606716760
transform 1 0 55660 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_607
timestamp 1606716760
transform 1 0 56212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_600
timestamp 1606716760
transform 1 0 55568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[38\]
timestamp 1606716760
transform 1 0 54648 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[32\]_A
timestamp 1606716760
transform 1 0 54832 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_599
timestamp 1606716760
transform 1 0 55476 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_590
timestamp 1606716760
transform 1 0 54648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_594
timestamp 1606716760
transform 1 0 55016 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _576_
timestamp 1606716760
transform 1 0 58144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[415\]
timestamp 1606716760
transform 1 0 59432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606716760
transform 1 0 59340 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__A
timestamp 1606716760
transform 1 0 58604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_631
timestamp 1606716760
transform 1 0 58420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_635
timestamp 1606716760
transform 1 0 58788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_626
timestamp 1606716760
transform 1 0 57960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[411\]
timestamp 1606716760
transform 1 0 56948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_618
timestamp 1606716760
transform 1 0 57224 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A
timestamp 1606716760
transform 1 0 56396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_611
timestamp 1606716760
transform 1 0 56580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _578_
timestamp 1606716760
transform 1 0 55936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_600
timestamp 1606716760
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_607
timestamp 1606716760
transform 1 0 56212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[38\]_A
timestamp 1606716760
transform 1 0 55384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_596
timestamp 1606716760
transform 1 0 55200 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _573_
timestamp 1606716760
transform 1 0 58604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_636
timestamp 1606716760
transform 1 0 58880 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[413\]
timestamp 1606716760
transform 1 0 57592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[81\]_B
timestamp 1606716760
transform 1 0 57316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_614
timestamp 1606716760
transform 1 0 56856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_618
timestamp 1606716760
transform 1 0 57224 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_621
timestamp 1606716760
transform 1 0 57500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_625
timestamp 1606716760
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _571_
timestamp 1606716760
transform 1 0 56580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606716760
transform 1 0 56488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[42\]_A
timestamp 1606716760
transform 1 0 55936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_606
timestamp 1606716760
transform 1 0 56120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _510_
timestamp 1606716760
transform 1 0 55108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_591
timestamp 1606716760
transform 1 0 54740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_598
timestamp 1606716760
transform 1 0 55384 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[37\]
timestamp 1606716760
transform 1 0 59432 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606716760
transform 1 0 59340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[81\]_A
timestamp 1606716760
transform 1 0 58144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1606716760
transform 1 0 58604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_630
timestamp 1606716760
transform 1 0 58328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_635
timestamp 1606716760
transform 1 0 58788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_626
timestamp 1606716760
transform 1 0 57960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[81\]
timestamp 1606716760
transform 1 0 57132 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_613
timestamp 1606716760
transform 1 0 56764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__A
timestamp 1606716760
transform 1 0 56580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_609
timestamp 1606716760
transform 1 0 56396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[42\]
timestamp 1606716760
transform 1 0 55568 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__A
timestamp 1606716760
transform 1 0 55108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_592
timestamp 1606716760
transform 1 0 54832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_597
timestamp 1606716760
transform 1 0 55292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[83\]
timestamp 1606716760
transform 1 0 58972 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_629
timestamp 1606716760
transform 1 0 58236 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[34\]
timestamp 1606716760
transform 1 0 57408 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[7\]_B
timestamp 1606716760
transform 1 0 57132 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_619
timestamp 1606716760
transform 1 0 57316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606716760
transform 1 0 56488 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_611
timestamp 1606716760
transform 1 0 56580 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[78\]_B
timestamp 1606716760
transform 1 0 55568 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_602
timestamp 1606716760
transform 1 0 55752 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_598
timestamp 1606716760
transform 1 0 55384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[63\]
timestamp 1606716760
transform 1 0 59432 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[85\]
timestamp 1606716760
transform 1 0 58512 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606716760
transform 1 0 59340 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[85\]_A
timestamp 1606716760
transform 1 0 59524 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[63\]_TE
timestamp 1606716760
transform 1 0 59156 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_641
timestamp 1606716760
transform 1 0 59340 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_637
timestamp 1606716760
transform 1 0 58972 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[34\]_A
timestamp 1606716760
transform 1 0 58328 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[83\]_B
timestamp 1606716760
transform 1 0 58788 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_628
timestamp 1606716760
transform 1 0 58144 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_632
timestamp 1606716760
transform 1 0 58512 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[7\]
timestamp 1606716760
transform 1 0 56948 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_624
timestamp 1606716760
transform 1 0 57776 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_624
timestamp 1606716760
transform 1 0 57776 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1606716760
transform 1 0 57408 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[137\]
timestamp 1606716760
transform 1 0 57500 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[7\]_A
timestamp 1606716760
transform 1 0 57960 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_611
timestamp 1606716760
transform 1 0 56580 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_612
timestamp 1606716760
transform 1 0 56672 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[78\]_A
timestamp 1606716760
transform 1 0 56396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_616
timestamp 1606716760
transform 1 0 57040 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[83\]_A
timestamp 1606716760
transform 1 0 56856 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[78\]
timestamp 1606716760
transform 1 0 55384 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[83\]
timestamp 1606716760
transform 1 0 55844 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_607
timestamp 1606716760
transform 1 0 56212 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[337\]
timestamp 1606716760
transform 1 0 54832 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[76\]_A
timestamp 1606716760
transform 1 0 54832 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_590
timestamp 1606716760
transform 1 0 54648 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_590
timestamp 1606716760
transform 1 0 54648 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[41\]_A
timestamp 1606716760
transform 1 0 55200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_594
timestamp 1606716760
transform 1 0 55016 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_595
timestamp 1606716760
transform 1 0 55108 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[36\]
timestamp 1606716760
transform 1 0 54464 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_587
timestamp 1606716760
transform 1 0 54372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1606716760
transform 1 0 53728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_577
timestamp 1606716760
transform 1 0 53452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_581
timestamp 1606716760
transform 1 0 53820 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[15\]_A
timestamp 1606716760
transform 1 0 52532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_569
timestamp 1606716760
transform 1 0 52716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[15\]_TE
timestamp 1606716760
transform 1 0 51612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_559
timestamp 1606716760
transform 1 0 51796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[89\]
timestamp 1606716760
transform 1 0 51152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[24\]_A
timestamp 1606716760
transform 1 0 50600 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_544
timestamp 1606716760
transform 1 0 50416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_548
timestamp 1606716760
transform 1 0 50784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_555
timestamp 1606716760
transform 1 0 51428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[33\]
timestamp 1606716760
transform 1 0 53452 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_586
timestamp 1606716760
transform 1 0 54280 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_574
timestamp 1606716760
transform 1 0 53176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_562
timestamp 1606716760
transform 1 0 52072 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1606716760
transform 1 0 50876 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_548
timestamp 1606716760
transform 1 0 50784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_550
timestamp 1606716760
transform 1 0 50968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_540
timestamp 1606716760
transform 1 0 50048 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[408\]
timestamp 1606716760
transform 1 0 53636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[32\]
timestamp 1606716760
transform 1 0 53820 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606716760
transform 1 0 53728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[33\]_A
timestamp 1606716760
transform 1 0 53544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_578
timestamp 1606716760
transform 1 0 53544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_582
timestamp 1606716760
transform 1 0 53912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_577
timestamp 1606716760
transform 1 0 53452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[31\]
timestamp 1606716760
transform 1 0 51980 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_570
timestamp 1606716760
transform 1 0 52808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1606716760
transform 1 0 51980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_573
timestamp 1606716760
transform 1 0 53084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_558
timestamp 1606716760
transform 1 0 51704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606716760
transform 1 0 50876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_548
timestamp 1606716760
transform 1 0 50784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_550
timestamp 1606716760
transform 1 0 50968 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_549
timestamp 1606716760
transform 1 0 50876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_540
timestamp 1606716760
transform 1 0 50048 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_537
timestamp 1606716760
transform 1 0 49772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[40\]
timestamp 1606716760
transform 1 0 54372 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606716760
transform 1 0 53728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[40\]_A
timestamp 1606716760
transform 1 0 54188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_579
timestamp 1606716760
transform 1 0 53636 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_581
timestamp 1606716760
transform 1 0 53820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[31\]_A
timestamp 1606716760
transform 1 0 52348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_561
timestamp 1606716760
transform 1 0 51980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_567
timestamp 1606716760
transform 1 0 52532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[27\]_A
timestamp 1606716760
transform 1 0 51796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_557
timestamp 1606716760
transform 1 0 51612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[27\]
timestamp 1606716760
transform 1 0 50784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_545
timestamp 1606716760
transform 1 0 50508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_537
timestamp 1606716760
transform 1 0 49772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[35\]_A
timestamp 1606716760
transform 1 0 54556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_587
timestamp 1606716760
transform 1 0 54372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[3\]
timestamp 1606716760
transform 1 0 53544 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_574
timestamp 1606716760
transform 1 0 53176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_562
timestamp 1606716760
transform 1 0 52072 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606716760
transform 1 0 50876 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_545
timestamp 1606716760
transform 1 0 50508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_550
timestamp 1606716760
transform 1 0 50968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[35\]
timestamp 1606716760
transform 1 0 54004 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606716760
transform 1 0 53728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[3\]_A
timestamp 1606716760
transform 1 0 53544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_576
timestamp 1606716760
transform 1 0 53360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_581
timestamp 1606716760
transform 1 0 53820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__A
timestamp 1606716760
transform 1 0 53176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _481_
timestamp 1606716760
transform 1 0 52716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_563
timestamp 1606716760
transform 1 0 52164 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_572
timestamp 1606716760
transform 1 0 52992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[30\]_A
timestamp 1606716760
transform 1 0 50876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_547
timestamp 1606716760
transform 1 0 50692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_551
timestamp 1606716760
transform 1 0 51060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[30\]
timestamp 1606716760
transform 1 0 49864 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[41\]
timestamp 1606716760
transform 1 0 54556 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[76\]_B
timestamp 1606716760
transform 1 0 54004 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_581
timestamp 1606716760
transform 1 0 53820 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_585
timestamp 1606716760
transform 1 0 54188 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[98\]
timestamp 1606716760
transform 1 0 52164 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[406\]
timestamp 1606716760
transform 1 0 51152 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606716760
transform 1 0 50876 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_546
timestamp 1606716760
transform 1 0 50600 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_550
timestamp 1606716760
transform 1 0 50968 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_555
timestamp 1606716760
transform 1 0 51428 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[76\]
timestamp 1606716760
transform 1 0 53820 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 1606716760
transform 1 0 54096 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1606716760
transform 1 0 54556 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_588
timestamp 1606716760
transform 1 0 54464 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _508_
timestamp 1606716760
transform 1 0 53452 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606716760
transform 1 0 53728 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[98\]_A
timestamp 1606716760
transform 1 0 53452 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_576
timestamp 1606716760
transform 1 0 53360 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_580
timestamp 1606716760
transform 1 0 53728 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_576
timestamp 1606716760
transform 1 0 53360 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_579
timestamp 1606716760
transform 1 0 53636 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__A
timestamp 1606716760
transform 1 0 53912 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[74\]
timestamp 1606716760
transform 1 0 51796 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_568
timestamp 1606716760
transform 1 0 52624 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_572
timestamp 1606716760
transform 1 0 52992 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_568
timestamp 1606716760
transform 1 0 52624 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[98\]_TE
timestamp 1606716760
transform 1 0 52440 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[74\]_A
timestamp 1606716760
transform 1 0 52808 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1606716760
transform 1 0 51704 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[74\]_B
timestamp 1606716760
transform 1 0 51520 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_558
timestamp 1606716760
transform 1 0 51704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_564
timestamp 1606716760
transform 1 0 52256 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[172\]
timestamp 1606716760
transform 1 0 51980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1606716760
transform 1 0 50968 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_546
timestamp 1606716760
transform 1 0 50600 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_548
timestamp 1606716760
transform 1 0 50784 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_541
timestamp 1606716760
transform 1 0 50140 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[81\]_A
timestamp 1606716760
transform 1 0 50784 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[404\]
timestamp 1606716760
transform 1 0 50508 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[81\]
timestamp 1606716760
transform 1 0 49772 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_537
timestamp 1606716760
transform 1 0 49772 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[78\]_A
timestamp 1606716760
transform 1 0 49956 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[24\]
timestamp 1606716760
transform 1 0 49588 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_532
timestamp 1606716760
transform 1 0 49312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1606716760
transform 1 0 48116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_516
timestamp 1606716760
transform 1 0 47840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_520
timestamp 1606716760
transform 1 0 48208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[117\]_A
timestamp 1606716760
transform 1 0 46920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[16\]_A
timestamp 1606716760
transform 1 0 46276 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_497
timestamp 1606716760
transform 1 0 46092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_501
timestamp 1606716760
transform 1 0 46460 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_505
timestamp 1606716760
transform 1 0 46828 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1606716760
transform 1 0 47104 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[16\]
timestamp 1606716760
transform 1 0 45264 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_485
timestamp 1606716760
transform 1 0 44988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[28\]
timestamp 1606716760
transform 1 0 49220 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_523
timestamp 1606716760
transform 1 0 48484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[20\]
timestamp 1606716760
transform 1 0 47656 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[21\]
timestamp 1606716760
transform 1 0 46092 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_506
timestamp 1606716760
transform 1 0 46920 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1606716760
transform 1 0 45264 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[117\]_TE
timestamp 1606716760
transform 1 0 45632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_489
timestamp 1606716760
transform 1 0 45356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_494
timestamp 1606716760
transform 1 0 45816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[28\]_A
timestamp 1606716760
transform 1 0 49588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[26\]
timestamp 1606716760
transform 1 0 49220 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[25\]_A
timestamp 1606716760
transform 1 0 49220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_523
timestamp 1606716760
transform 1 0 48484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_529
timestamp 1606716760
transform 1 0 49036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_533
timestamp 1606716760
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[22\]
timestamp 1606716760
transform 1 0 47656 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[25\]
timestamp 1606716760
transform 1 0 48208 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606716760
transform 1 0 48116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[20\]_A
timestamp 1606716760
transform 1 0 47932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_509
timestamp 1606716760
transform 1 0 47196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_513
timestamp 1606716760
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_515
timestamp 1606716760
transform 1 0 47748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[21\]_A
timestamp 1606716760
transform 1 0 46460 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_497
timestamp 1606716760
transform 1 0 46092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_503
timestamp 1606716760
transform 1 0 46644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606716760
transform 1 0 45264 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[72\]_B
timestamp 1606716760
transform 1 0 45908 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_487
timestamp 1606716760
transform 1 0 45172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_489
timestamp 1606716760
transform 1 0 45356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_483
timestamp 1606716760
transform 1 0 44804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_495
timestamp 1606716760
transform 1 0 45908 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[26\]_A
timestamp 1606716760
transform 1 0 49588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[14\]_A
timestamp 1606716760
transform 1 0 49220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_529
timestamp 1606716760
transform 1 0 49036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_533
timestamp 1606716760
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[14\]
timestamp 1606716760
transform 1 0 48208 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606716760
transform 1 0 48116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[22\]_A
timestamp 1606716760
transform 1 0 47932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_514
timestamp 1606716760
transform 1 0 47656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[72\]_A
timestamp 1606716760
transform 1 0 46736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1606716760
transform 1 0 46552 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_506
timestamp 1606716760
transform 1 0 46920 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[72\]
timestamp 1606716760
transform 1 0 45724 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_492
timestamp 1606716760
transform 1 0 45632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[23\]
timestamp 1606716760
transform 1 0 48576 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_523
timestamp 1606716760
transform 1 0 48484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1606716760
transform 1 0 49404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 1606716760
transform 1 0 47472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_510
timestamp 1606716760
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_515
timestamp 1606716760
transform 1 0 47748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[70\]_B
timestamp 1606716760
transform 1 0 46368 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_498
timestamp 1606716760
transform 1 0 46184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_502
timestamp 1606716760
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[2\]
timestamp 1606716760
transform 1 0 45356 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606716760
transform 1 0 45264 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_484
timestamp 1606716760
transform 1 0 44896 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[23\]_A
timestamp 1606716760
transform 1 0 48944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_530
timestamp 1606716760
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606716760
transform 1 0 48116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__A
timestamp 1606716760
transform 1 0 47472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_511
timestamp 1606716760
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_514
timestamp 1606716760
transform 1 0 47656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_518
timestamp 1606716760
transform 1 0 48024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_520
timestamp 1606716760
transform 1 0 48208 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[70\]_A
timestamp 1606716760
transform 1 0 46644 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_501
timestamp 1606716760
transform 1 0 46460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_505
timestamp 1606716760
transform 1 0 46828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[70\]
timestamp 1606716760
transform 1 0 45632 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[65\]_A
timestamp 1606716760
transform 1 0 45080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[2\]_A
timestamp 1606716760
transform 1 0 45448 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_484
timestamp 1606716760
transform 1 0 44896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_488
timestamp 1606716760
transform 1 0 45264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_534
timestamp 1606716760
transform 1 0 49496 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[7\]
timestamp 1606716760
transform 1 0 48668 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_517
timestamp 1606716760
transform 1 0 47932 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[74\]
timestamp 1606716760
transform 1 0 47104 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_500
timestamp 1606716760
transform 1 0 46368 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[72\]
timestamp 1606716760
transform 1 0 45540 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606716760
transform 1 0 45264 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_487
timestamp 1606716760
transform 1 0 45172 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_489
timestamp 1606716760
transform 1 0 45356 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[7\]_A
timestamp 1606716760
transform 1 0 49588 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[78\]
timestamp 1606716760
transform 1 0 48944 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_533
timestamp 1606716760
transform 1 0 49404 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_529
timestamp 1606716760
transform 1 0 49036 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1606716760
transform 1 0 48668 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[76\]_A
timestamp 1606716760
transform 1 0 49220 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1606716760
transform 1 0 48852 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[402\]
timestamp 1606716760
transform 1 0 47656 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[76\]
timestamp 1606716760
transform 1 0 48208 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606716760
transform 1 0 48116 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[74\]_A
timestamp 1606716760
transform 1 0 47472 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_510
timestamp 1606716760
transform 1 0 47288 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1606716760
transform 1 0 47932 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_514
timestamp 1606716760
transform 1 0 47656 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_518
timestamp 1606716760
transform 1 0 48024 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[400\]
timestamp 1606716760
transform 1 0 46644 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[70\]
timestamp 1606716760
transform 1 0 46092 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1606716760
transform 1 0 46000 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[69\]_A
timestamp 1606716760
transform 1 0 46092 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[70\]_A
timestamp 1606716760
transform 1 0 47104 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[72\]_A
timestamp 1606716760
transform 1 0 46460 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_506
timestamp 1606716760
transform 1 0 46920 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_499
timestamp 1606716760
transform 1 0 46276 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_506
timestamp 1606716760
transform 1 0 46920 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[395\]
timestamp 1606716760
transform 1 0 44804 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[69\]
timestamp 1606716760
transform 1 0 45080 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_486
timestamp 1606716760
transform 1 0 45080 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_494
timestamp 1606716760
transform 1 0 45816 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_495
timestamp 1606716760
transform 1 0 45908 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_477
timestamp 1606716760
transform 1 0 44252 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1606716760
transform 1 0 42504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[25\]_A
timestamp 1606716760
transform 1 0 42964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_459
timestamp 1606716760
transform 1 0 42596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_465
timestamp 1606716760
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[25\]_TE
timestamp 1606716760
transform 1 0 41952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_450
timestamp 1606716760
transform 1 0 41768 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_454
timestamp 1606716760
transform 1 0 42136 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[99\]
timestamp 1606716760
transform 1 0 41492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_437
timestamp 1606716760
transform 1 0 40572 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_445
timestamp 1606716760
transform 1 0 41308 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_476
timestamp 1606716760
transform 1 0 44160 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_464
timestamp 1606716760
transform 1 0 43056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_452
timestamp 1606716760
transform 1 0 41952 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_440
timestamp 1606716760
transform 1 0 40848 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_475
timestamp 1606716760
transform 1 0 44068 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_471
timestamp 1606716760
transform 1 0 43700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606716760
transform 1 0 42504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_463
timestamp 1606716760
transform 1 0 42964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_457
timestamp 1606716760
transform 1 0 42412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_459
timestamp 1606716760
transform 1 0 42596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_451
timestamp 1606716760
transform 1 0 41860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_453
timestamp 1606716760
transform 1 0 42044 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[1\]
timestamp 1606716760
transform 1 0 41032 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[19\]_A
timestamp 1606716760
transform 1 0 40756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_440
timestamp 1606716760
transform 1 0 40848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_437
timestamp 1606716760
transform 1 0 40572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_441
timestamp 1606716760
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[17\]_A
timestamp 1606716760
transform 1 0 44344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_476
timestamp 1606716760
transform 1 0 44160 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_480
timestamp 1606716760
transform 1 0 44528 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[17\]
timestamp 1606716760
transform 1 0 43332 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606716760
transform 1 0 42504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_456
timestamp 1606716760
transform 1 0 42320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_459
timestamp 1606716760
transform 1 0 42596 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_448
timestamp 1606716760
transform 1 0 41584 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[1\]_A
timestamp 1606716760
transform 1 0 41400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_443
timestamp 1606716760
transform 1 0 41124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_435
timestamp 1606716760
transform 1 0 40388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[69\]
timestamp 1606716760
transform 1 0 43700 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[69\]_A
timestamp 1606716760
transform 1 0 44712 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_480
timestamp 1606716760
transform 1 0 44528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[83\]
timestamp 1606716760
transform 1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_463
timestamp 1606716760
transform 1 0 42964 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_448
timestamp 1606716760
transform 1 0 41584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _587_
timestamp 1606716760
transform 1 0 41308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_437
timestamp 1606716760
transform 1 0 40572 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[65\]
timestamp 1606716760
transform 1 0 44068 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[65\]_B
timestamp 1606716760
transform 1 0 43884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_471
timestamp 1606716760
transform 1 0 43700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__A
timestamp 1606716760
transform 1 0 43516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_467
timestamp 1606716760
transform 1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _513_
timestamp 1606716760
transform 1 0 43056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606716760
transform 1 0 42504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_459
timestamp 1606716760
transform 1 0 42596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_463
timestamp 1606716760
transform 1 0 42964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_455
timestamp 1606716760
transform 1 0 42228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__587__A
timestamp 1606716760
transform 1 0 41308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_442
timestamp 1606716760
transform 1 0 41032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_447
timestamp 1606716760
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[126\]_A
timestamp 1606716760
transform 1 0 40112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_430
timestamp 1606716760
transform 1 0 39928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_434
timestamp 1606716760
transform 1 0 40296 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[65\]_A
timestamp 1606716760
transform 1 0 44068 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[69\]_B
timestamp 1606716760
transform 1 0 44436 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_473
timestamp 1606716760
transform 1 0 43884 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1606716760
transform 1 0 44252 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_481
timestamp 1606716760
transform 1 0 44620 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[65\]
timestamp 1606716760
transform 1 0 43056 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[9\]_TE
timestamp 1606716760
transform 1 0 42688 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_456
timestamp 1606716760
transform 1 0 42320 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_462
timestamp 1606716760
transform 1 0 42872 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[399\]
timestamp 1606716760
transform 1 0 42044 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_452
timestamp 1606716760
transform 1 0 41952 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_440
timestamp 1606716760
transform 1 0 40848 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[9\]_A
timestamp 1606716760
transform 1 0 44528 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[67\]_A
timestamp 1606716760
transform 1 0 44252 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_475
timestamp 1606716760
transform 1 0 44068 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_479
timestamp 1606716760
transform 1 0 44436 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_478
timestamp 1606716760
transform 1 0 44344 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1606716760
transform 1 0 44712 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[67\]
timestamp 1606716760
transform 1 0 41584 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[67\]
timestamp 1606716760
transform 1 0 43240 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  la_buf\[9\]
timestamp 1606716760
transform 1 0 42688 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_1_459
timestamp 1606716760
transform 1 0 42596 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1606716760
transform 1 0 42780 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[67\]_A
timestamp 1606716760
transform 1 0 42596 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1606716760
transform 1 0 43148 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606716760
transform 1 0 42504 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_450
timestamp 1606716760
transform 1 0 41768 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_457
timestamp 1606716760
transform 1 0 42412 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_434
timestamp 1606716760
transform 1 0 40296 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_446
timestamp 1606716760
transform 1 0 41400 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_443
timestamp 1606716760
transform 1 0 41124 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[67\]_B
timestamp 1606716760
transform 1 0 41400 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[397\]
timestamp 1606716760
transform 1 0 41492 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1606716760
transform 1 0 40296 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[63\]_A
timestamp 1606716760
transform 1 0 40112 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_432
timestamp 1606716760
transform 1 0 40112 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_435
timestamp 1606716760
transform 1 0 40388 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_430
timestamp 1606716760
transform 1 0 39928 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_425
timestamp 1606716760
transform 1 0 39468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_413
timestamp 1606716760
transform 1 0 38364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[443\]
timestamp 1606716760
transform 1 0 36984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1606716760
transform 1 0 36892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_389
timestamp 1606716760
transform 1 0 36156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_401
timestamp 1606716760
transform 1 0 37260 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[115\]_A
timestamp 1606716760
transform 1 0 35972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_385
timestamp 1606716760
transform 1 0 35788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1606716760
transform 1 0 39652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_428
timestamp 1606716760
transform 1 0 39744 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_424
timestamp 1606716760
transform 1 0 39376 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_412
timestamp 1606716760
transform 1 0 38272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_400
timestamp 1606716760
transform 1 0 37168 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_388
timestamp 1606716760
transform 1 0 36064 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_376
timestamp 1606716760
transform 1 0 34960 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[19\]
timestamp 1606716760
transform 1 0 39744 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606716760
transform 1 0 39652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_428
timestamp 1606716760
transform 1 0 39744 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_422
timestamp 1606716760
transform 1 0 39192 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_415
timestamp 1606716760
transform 1 0 38548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_403
timestamp 1606716760
transform 1 0 37444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_410
timestamp 1606716760
transform 1 0 38088 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606716760
transform 1 0 36892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_391
timestamp 1606716760
transform 1 0 36340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_398
timestamp 1606716760
transform 1 0 36984 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_385
timestamp 1606716760
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_379
timestamp 1606716760
transform 1 0 35236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_423
timestamp 1606716760
transform 1 0 39284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[124\]_A
timestamp 1606716760
transform 1 0 37996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_407
timestamp 1606716760
transform 1 0 37812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_411
timestamp 1606716760
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[124\]
timestamp 1606716760
transform 1 0 36984 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606716760
transform 1 0 36892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_389
timestamp 1606716760
transform 1 0 36156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_377
timestamp 1606716760
transform 1 0 35052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[126\]
timestamp 1606716760
transform 1 0 39744 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606716760
transform 1 0 39652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[63\]_B
timestamp 1606716760
transform 1 0 38916 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_418
timestamp 1606716760
transform 1 0 38824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_421
timestamp 1606716760
transform 1 0 39100 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_410
timestamp 1606716760
transform 1 0 38088 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[29\]
timestamp 1606716760
transform 1 0 36156 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_398
timestamp 1606716760
transform 1 0 36984 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_387
timestamp 1606716760
transform 1 0 35972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_379
timestamp 1606716760
transform 1 0 35236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[63\]_A
timestamp 1606716760
transform 1 0 39744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_426
timestamp 1606716760
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[63\]
timestamp 1606716760
transform 1 0 38732 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_416
timestamp 1606716760
transform 1 0 38640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_410
timestamp 1606716760
transform 1 0 38088 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606716760
transform 1 0 36892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[29\]_A
timestamp 1606716760
transform 1 0 36524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_395
timestamp 1606716760
transform 1 0 36708 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_398
timestamp 1606716760
transform 1 0 36984 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_385
timestamp 1606716760
transform 1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606716760
transform 1 0 39652 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_428
timestamp 1606716760
transform 1 0 39744 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_426
timestamp 1606716760
transform 1 0 39560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_414
timestamp 1606716760
transform 1 0 38456 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_402
timestamp 1606716760
transform 1 0 37352 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[61\]_B
timestamp 1606716760
transform 1 0 37168 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_389
timestamp 1606716760
transform 1 0 36156 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_397
timestamp 1606716760
transform 1 0 36892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[391\]
timestamp 1606716760
transform 1 0 35880 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[5\]_B
timestamp 1606716760
transform 1 0 35512 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_384
timestamp 1606716760
transform 1 0 35696 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[63\]
timestamp 1606716760
transform 1 0 39100 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_419
timestamp 1606716760
transform 1 0 38916 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_424
timestamp 1606716760
transform 1 0 39376 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[393\]
timestamp 1606716760
transform 1 0 39100 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[61\]_A
timestamp 1606716760
transform 1 0 38548 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_417
timestamp 1606716760
transform 1 0 38732 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[61\]
timestamp 1606716760
transform 1 0 37536 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1606716760
transform 1 0 37444 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[61\]_A
timestamp 1606716760
transform 1 0 37996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_413
timestamp 1606716760
transform 1 0 38364 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_407
timestamp 1606716760
transform 1 0 37812 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_411
timestamp 1606716760
transform 1 0 38180 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[61\]
timestamp 1606716760
transform 1 0 36984 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606716760
transform 1 0 36892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[5\]_A
timestamp 1606716760
transform 1 0 36340 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[5\]_A
timestamp 1606716760
transform 1 0 36248 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_392
timestamp 1606716760
transform 1 0 36432 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_400
timestamp 1606716760
transform 1 0 37168 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_389
timestamp 1606716760
transform 1 0 36156 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1606716760
transform 1 0 36524 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_388
timestamp 1606716760
transform 1 0 36064 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[5\]
timestamp 1606716760
transform 1 0 35236 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[5\]
timestamp 1606716760
transform 1 0 35328 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_376
timestamp 1606716760
transform 1 0 34960 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[115\]
timestamp 1606716760
transform 1 0 34132 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[115\]_TE
timestamp 1606716760
transform 1 0 33948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[116\]_TE
timestamp 1606716760
transform 1 0 33580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_363
timestamp 1606716760
transform 1 0 33764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[190\]
timestamp 1606716760
transform 1 0 33120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_355
timestamp 1606716760
transform 1 0 33028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_359
timestamp 1606716760
transform 1 0 33396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_349
timestamp 1606716760
transform 1 0 32476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1606716760
transform 1 0 31280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1606716760
transform 1 0 31096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1606716760
transform 1 0 31372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[122\]_A
timestamp 1606716760
transform 1 0 30176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_326
timestamp 1606716760
transform 1 0 30360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[125\]
timestamp 1606716760
transform 1 0 34132 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606716760
transform 1 0 34040 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_354
timestamp 1606716760
transform 1 0 32936 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_342
timestamp 1606716760
transform 1 0 31832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_330
timestamp 1606716760
transform 1 0 30728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606716760
transform 1 0 34040 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[125\]_A
timestamp 1606716760
transform 1 0 34500 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_367
timestamp 1606716760
transform 1 0 34132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_368
timestamp 1606716760
transform 1 0 34224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1606716760
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_364
timestamp 1606716760
transform 1 0 33856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_360
timestamp 1606716760
transform 1 0 33488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[121\]_A
timestamp 1606716760
transform 1 0 33304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_356
timestamp 1606716760
transform 1 0 33120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_356
timestamp 1606716760
transform 1 0 33120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[120\]
timestamp 1606716760
transform 1 0 32292 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[121\]
timestamp 1606716760
transform 1 0 32292 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_342
timestamp 1606716760
transform 1 0 31832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_346
timestamp 1606716760
transform 1 0 32200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_345
timestamp 1606716760
transform 1 0 32108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606716760
transform 1 0 31280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1606716760
transform 1 0 31188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_337
timestamp 1606716760
transform 1 0 31372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[13\]_A
timestamp 1606716760
transform 1 0 30452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_330
timestamp 1606716760
transform 1 0 30728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_325
timestamp 1606716760
transform 1 0 30268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1606716760
transform 1 0 30636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_365
timestamp 1606716760
transform 1 0 33948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[120\]_A
timestamp 1606716760
transform 1 0 32660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_353
timestamp 1606716760
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_349
timestamp 1606716760
transform 1 0 32476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606716760
transform 1 0 31280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1606716760
transform 1 0 31188 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1606716760
transform 1 0 31372 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1606716760
transform 1 0 30820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606716760
transform 1 0 34040 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_367
timestamp 1606716760
transform 1 0 34132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_361
timestamp 1606716760
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_365
timestamp 1606716760
transform 1 0 33948 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_349
timestamp 1606716760
transform 1 0 32476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_337
timestamp 1606716760
transform 1 0 31372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[18\]
timestamp 1606716760
transform 1 0 30544 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_327
timestamp 1606716760
transform 1 0 30452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1606716760
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1606716760
transform 1 0 33580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1606716760
transform 1 0 32476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606716760
transform 1 0 31280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[18\]_A
timestamp 1606716760
transform 1 0 30912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1606716760
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1606716760
transform 1 0 31372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[144\]
timestamp 1606716760
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_328
timestamp 1606716760
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[335\]
timestamp 1606716760
transform 1 0 34500 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606716760
transform 1 0 34040 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_367
timestamp 1606716760
transform 1 0 34132 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_374
timestamp 1606716760
transform 1 0 34776 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_362
timestamp 1606716760
transform 1 0 33672 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[388\]
timestamp 1606716760
transform 1 0 32292 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_350
timestamp 1606716760
transform 1 0 32568 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[386\]
timestamp 1606716760
transform 1 0 31280 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_332
timestamp 1606716760
transform 1 0 30912 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_339
timestamp 1606716760
transform 1 0 31556 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[56\]_B
timestamp 1606716760
transform 1 0 30728 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_328
timestamp 1606716760
transform 1 0 30544 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1606716760
transform 1 0 34592 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[58\]_A
timestamp 1606716760
transform 1 0 34776 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_366
timestamp 1606716760
transform 1 0 34040 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_373
timestamp 1606716760
transform 1 0 34684 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_372
timestamp 1606716760
transform 1 0 34592 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[58\]
timestamp 1606716760
transform 1 0 33764 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[58\]_A
timestamp 1606716760
transform 1 0 33856 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[58\]_B
timestamp 1606716760
transform 1 0 33580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1606716760
transform 1 0 33672 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[58\]
timestamp 1606716760
transform 1 0 32844 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[70\]_A
timestamp 1606716760
transform 1 0 33212 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_355
timestamp 1606716760
transform 1 0 33028 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_359
timestamp 1606716760
transform 1 0 33396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[384\]
timestamp 1606716760
transform 1 0 31832 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1606716760
transform 1 0 31740 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_345
timestamp 1606716760
transform 1 0 32108 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[70\]
timestamp 1606716760
transform 1 0 31372 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_1_332
timestamp 1606716760
transform 1 0 30912 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_340
timestamp 1606716760
transform 1 0 31648 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_332
timestamp 1606716760
transform 1 0 30912 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[70\]_TE
timestamp 1606716760
transform 1 0 31096 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606716760
transform 1 0 31280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_328
timestamp 1606716760
transform 1 0 30544 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_322
timestamp 1606716760
transform 1 0 29992 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_328
timestamp 1606716760
transform 1 0 30544 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[56\]_A
timestamp 1606716760
transform 1 0 30728 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[65\]_A
timestamp 1606716760
transform 1 0 30728 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[56\]_A
timestamp 1606716760
transform 1 0 30360 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_321
timestamp 1606716760
transform 1 0 29900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_313
timestamp 1606716760
transform 1 0 29164 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_301
timestamp 1606716760
transform 1 0 28060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[115\]_A
timestamp 1606716760
transform 1 0 26772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_289
timestamp 1606716760
transform 1 0 26956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_285
timestamp 1606716760
transform 1 0 26588 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[123\]
timestamp 1606716760
transform 1 0 25760 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1606716760
transform 1 0 25668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[115\]_B
timestamp 1606716760
transform 1 0 25484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_272
timestamp 1606716760
transform 1 0 25392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_318
timestamp 1606716760
transform 1 0 29624 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_306
timestamp 1606716760
transform 1 0 28520 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606716760
transform 1 0 28428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_302
timestamp 1606716760
transform 1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_294
timestamp 1606716760
transform 1 0 27416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[123\]_A
timestamp 1606716760
transform 1 0 26128 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_282
timestamp 1606716760
transform 1 0 26312 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[185\]
timestamp 1606716760
transform 1 0 25300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_274
timestamp 1606716760
transform 1 0 25576 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[13\]
timestamp 1606716760
transform 1 0 29440 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_318
timestamp 1606716760
transform 1 0 29624 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_306
timestamp 1606716760
transform 1 0 28520 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_313
timestamp 1606716760
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606716760
transform 1 0 28428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_303
timestamp 1606716760
transform 1 0 28244 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_301
timestamp 1606716760
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[119\]_A
timestamp 1606716760
transform 1 0 26772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_295
timestamp 1606716760
transform 1 0 27508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_289
timestamp 1606716760
transform 1 0 26956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_283
timestamp 1606716760
transform 1 0 26404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_285
timestamp 1606716760
transform 1 0 26588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[119\]
timestamp 1606716760
transform 1 0 25760 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[118\]
timestamp 1606716760
transform 1 0 25576 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_274
timestamp 1606716760
transform 1 0 25576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606716760
transform 1 0 25668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1606716760
transform 1 0 25208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[15\]_A
timestamp 1606716760
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_315
timestamp 1606716760
transform 1 0 29348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_319
timestamp 1606716760
transform 1 0 29716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[15\]
timestamp 1606716760
transform 1 0 28520 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[127\]_A
timestamp 1606716760
transform 1 0 27876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1606716760
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_305
timestamp 1606716760
transform 1 0 28428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[127\]
timestamp 1606716760
transform 1 0 26864 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1606716760
transform 1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[118\]_A
timestamp 1606716760
transform 1 0 26312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_280
timestamp 1606716760
transform 1 0 26128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_284
timestamp 1606716760
transform 1 0 26496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[146\]
timestamp 1606716760
transform 1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606716760
transform 1 0 25668 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_269
timestamp 1606716760
transform 1 0 25116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1606716760
transform 1 0 25760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_315
timestamp 1606716760
transform 1 0 29348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[12\]
timestamp 1606716760
transform 1 0 28520 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606716760
transform 1 0 28428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[67\]_TE
timestamp 1606716760
transform 1 0 27876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_301
timestamp 1606716760
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _585_
timestamp 1606716760
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_292
timestamp 1606716760
transform 1 0 27232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1606716760
transform 1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1606716760
transform 1 0 26128 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[54\]_B
timestamp 1606716760
transform 1 0 25944 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_276
timestamp 1606716760
transform 1 0 25760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[12\]_A
timestamp 1606716760
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_315
timestamp 1606716760
transform 1 0 29348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_319
timestamp 1606716760
transform 1 0 29716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[67\]_A
timestamp 1606716760
transform 1 0 29164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_311
timestamp 1606716760
transform 1 0 28980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[67\]
timestamp 1606716760
transform 1 0 27324 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[54\]_A
timestamp 1606716760
transform 1 0 26772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__585__A
timestamp 1606716760
transform 1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_289
timestamp 1606716760
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_285
timestamp 1606716760
transform 1 0 26588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[54\]
timestamp 1606716760
transform 1 0 25760 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606716760
transform 1 0 25668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[113\]_A
timestamp 1606716760
transform 1 0 25300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_273
timestamp 1606716760
transform 1 0 25484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[56\]
timestamp 1606716760
transform 1 0 29716 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_317
timestamp 1606716760
transform 1 0 29532 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[139\]
timestamp 1606716760
transform 1 0 28520 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1606716760
transform 1 0 28796 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606716760
transform 1 0 28428 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_300
timestamp 1606716760
transform 1 0 27968 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_304
timestamp 1606716760
transform 1 0 28336 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_288
timestamp 1606716760
transform 1 0 26864 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[115\]
timestamp 1606716760
transform 1 0 26036 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_271
timestamp 1606716760
transform 1 0 25300 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[56\]
timestamp 1606716760
transform 1 0 29716 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1606716760
transform 1 0 28888 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_306
timestamp 1606716760
transform 1 0 28520 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_311
timestamp 1606716760
transform 1 0 28980 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[65\]
timestamp 1606716760
transform 1 0 28336 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[72\]_A
timestamp 1606716760
transform 1 0 28336 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[65\]_TE
timestamp 1606716760
transform 1 0 28152 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_302
timestamp 1606716760
transform 1 0 28152 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[141\]
timestamp 1606716760
transform 1 0 27324 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[115\]_A
timestamp 1606716760
transform 1 0 26772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1606716760
transform 1 0 26956 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_296
timestamp 1606716760
transform 1 0 27600 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[54\]
timestamp 1606716760
transform 1 0 25760 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  la_buf\[72\]
timestamp 1606716760
transform 1 0 26496 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1606716760
transform 1 0 26036 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_285
timestamp 1606716760
transform 1 0 26588 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_280
timestamp 1606716760
transform 1 0 26128 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[54\]_A
timestamp 1606716760
transform 1 0 26312 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_269
timestamp 1606716760
transform 1 0 25116 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_269
timestamp 1606716760
transform 1 0 25116 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606716760
transform 1 0 25668 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__A
timestamp 1606716760
transform 1 0 25300 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[69\]_TE
timestamp 1606716760
transform 1 0 25300 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[72\]_TE
timestamp 1606716760
transform 1 0 25852 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1606716760
transform 1 0 25484 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_273
timestamp 1606716760
transform 1 0 25484 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[116\]_A
timestamp 1606716760
transform 1 0 24472 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_264
timestamp 1606716760
transform 1 0 24656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_260
timestamp 1606716760
transform 1 0 24288 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[116\]
timestamp 1606716760
transform 1 0 23460 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[11\]_A
timestamp 1606716760
transform 1 0 23276 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_247
timestamp 1606716760
transform 1 0 23092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[114\]_A
timestamp 1606716760
transform 1 0 22908 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_243
timestamp 1606716760
transform 1 0 22724 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[114\]
timestamp 1606716760
transform 1 0 21068 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[1\]_A
timestamp 1606716760
transform 1 0 20792 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_215
timestamp 1606716760
transform 1 0 20148 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_221
timestamp 1606716760
transform 1 0 20700 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_224
timestamp 1606716760
transform 1 0 20976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[113\]_A
timestamp 1606716760
transform 1 0 24748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_263
timestamp 1606716760
transform 1 0 24564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_267
timestamp 1606716760
transform 1 0 24932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[113\]
timestamp 1606716760
transform 1 0 22908 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606716760
transform 1 0 22816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_236
timestamp 1606716760
transform 1 0 22080 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[193\]
timestamp 1606716760
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[103\]
timestamp 1606716760
transform 1 0 21252 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_219
timestamp 1606716760
transform 1 0 20516 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_268
timestamp 1606716760
transform 1 0 25024 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1606716760
transform 1 0 24656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_266
timestamp 1606716760
transform 1 0 24840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[114\]_A
timestamp 1606716760
transform 1 0 25024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[111\]_A
timestamp 1606716760
transform 1 0 24840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[114\]
timestamp 1606716760
transform 1 0 24012 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_245
timestamp 1606716760
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[111\]
timestamp 1606716760
transform 1 0 23000 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_7_242
timestamp 1606716760
transform 1 0 22632 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_238
timestamp 1606716760
transform 1 0 22264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_241
timestamp 1606716760
transform 1 0 22540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[113\]_TE
timestamp 1606716760
transform 1 0 22448 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[111\]_TE
timestamp 1606716760
transform 1 0 22816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606716760
transform 1 0 22816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[187\]
timestamp 1606716760
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1606716760
transform 1 0 21436 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_227
timestamp 1606716760
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[52\]_B
timestamp 1606716760
transform 1 0 20976 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[382\]
timestamp 1606716760
transform 1 0 21160 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[188\]
timestamp 1606716760
transform 1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[103\]_A
timestamp 1606716760
transform 1 0 21620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_233
timestamp 1606716760
transform 1 0 21804 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1606716760
transform 1 0 20884 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1606716760
transform 1 0 20148 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_223
timestamp 1606716760
transform 1 0 20884 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1606716760
transform 1 0 20148 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[112\]_A
timestamp 1606716760
transform 1 0 24932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_265
timestamp 1606716760
transform 1 0 24748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[112\]
timestamp 1606716760
transform 1 0 23920 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[117\]_A
timestamp 1606716760
transform 1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_248
timestamp 1606716760
transform 1 0 23184 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_252
timestamp 1606716760
transform 1 0 23552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[117\]
timestamp 1606716760
transform 1 0 22356 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_235
timestamp 1606716760
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[52\]_A
timestamp 1606716760
transform 1 0 21804 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_231
timestamp 1606716760
transform 1 0 21620 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[52\]
timestamp 1606716760
transform 1 0 20792 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_215
timestamp 1606716760
transform 1 0 20148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_221
timestamp 1606716760
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[113\]
timestamp 1606716760
transform 1 0 24932 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_259
timestamp 1606716760
transform 1 0 24196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[110\]
timestamp 1606716760
transform 1 0 23368 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_249
timestamp 1606716760
transform 1 0 23276 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606716760
transform 1 0 22816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_236
timestamp 1606716760
transform 1 0 22080 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_245
timestamp 1606716760
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _590_
timestamp 1606716760
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1606716760
transform 1 0 20700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[111\]_A
timestamp 1606716760
transform 1 0 24840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1606716760
transform 1 0 24656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_268
timestamp 1606716760
transform 1 0 25024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[111\]
timestamp 1606716760
transform 1 0 23828 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[110\]_A
timestamp 1606716760
transform 1 0 23644 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[10\]_A
timestamp 1606716760
transform 1 0 22724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_241
timestamp 1606716760
transform 1 0 22540 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1606716760
transform 1 0 22908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[10\]
timestamp 1606716760
transform 1 0 21712 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__A
timestamp 1606716760
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_228
timestamp 1606716760
transform 1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[107\]
timestamp 1606716760
transform 1 0 20148 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[107\]_A
timestamp 1606716760
transform 1 0 21160 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_224
timestamp 1606716760
transform 1 0 20976 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[69\]
timestamp 1606716760
transform 1 0 23644 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606716760
transform 1 0 22816 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[45\]_TE
timestamp 1606716760
transform 1 0 22540 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_235
timestamp 1606716760
transform 1 0 21988 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_243
timestamp 1606716760
transform 1 0 22724 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_245
timestamp 1606716760
transform 1 0 22908 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[119\]
timestamp 1606716760
transform 1 0 21712 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1606716760
transform 1 0 21344 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[38\]_A
timestamp 1606716760
transform 1 0 21160 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_224
timestamp 1606716760
transform 1 0 20976 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_263
timestamp 1606716760
transform 1 0 24564 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1606716760
transform 1 0 24472 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[69\]_A
timestamp 1606716760
transform 1 0 24932 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[45\]_A
timestamp 1606716760
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1606716760
transform 1 0 24840 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[52\]_A
timestamp 1606716760
transform 1 0 24288 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1606716760
transform 1 0 24104 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_259
timestamp 1606716760
transform 1 0 24196 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[52\]
timestamp 1606716760
transform 1 0 23276 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1606716760
transform 1 0 23184 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  la_buf\[45\]
timestamp 1606716760
transform 1 0 22540 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[143\]
timestamp 1606716760
transform 1 0 22172 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[36\]_A
timestamp 1606716760
transform 1 0 21988 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240
timestamp 1606716760
transform 1 0 22448 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1606716760
transform 1 0 22172 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[109\]_A
timestamp 1606716760
transform 1 0 21436 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_231
timestamp 1606716760
transform 1 0 21620 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_233
timestamp 1606716760
transform 1 0 21804 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[109\]
timestamp 1606716760
transform 1 0 20424 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  la_buf\[36\]
timestamp 1606716760
transform 1 0 20148 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_0_227
timestamp 1606716760
transform 1 0 21252 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1606716760
transform 1 0 20332 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1606716760
transform 1 0 20056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_210
timestamp 1606716760
transform 1 0 19688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[75\]
timestamp 1606716760
transform 1 0 19044 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[1\]_TE
timestamp 1606716760
transform 1 0 19504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_200
timestamp 1606716760
transform 1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_206
timestamp 1606716760
transform 1 0 19320 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[112\]_A
timestamp 1606716760
transform 1 0 17848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1606716760
transform 1 0 17664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_192
timestamp 1606716760
transform 1 0 18032 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[112\]
timestamp 1606716760
transform 1 0 16008 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[112\]_TE
timestamp 1606716760
transform 1 0 15824 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1606716760
transform 1 0 15640 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_214
timestamp 1606716760
transform 1 0 20056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[105\]_A
timestamp 1606716760
transform 1 0 18768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1606716760
transform 1 0 18952 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_198
timestamp 1606716760
transform 1 0 18584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[105\]
timestamp 1606716760
transform 1 0 17756 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606716760
transform 1 0 17204 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_182
timestamp 1606716760
transform 1 0 17112 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1606716760
transform 1 0 17296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_188
timestamp 1606716760
transform 1 0 17664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[100\]
timestamp 1606716760
transform 1 0 15548 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_174
timestamp 1606716760
transform 1 0 16376 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606716760
transform 1 0 20056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[102\]_A
timestamp 1606716760
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_203
timestamp 1606716760
transform 1 0 19044 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1606716760
transform 1 0 18952 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1606716760
transform 1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[102\]
timestamp 1606716760
transform 1 0 17756 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[104\]
timestamp 1606716760
transform 1 0 18216 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606716760
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[101\]_A
timestamp 1606716760
transform 1 0 17204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_184
timestamp 1606716760
transform 1 0 17296 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_192
timestamp 1606716760
transform 1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606716760
transform 1 0 17020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1606716760
transform 1 0 17388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[101\]
timestamp 1606716760
transform 1 0 16192 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[100\]_A
timestamp 1606716760
transform 1 0 15916 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1606716760
transform 1 0 16100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_166
timestamp 1606716760
transform 1 0 15640 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_171
timestamp 1606716760
transform 1 0 16100 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606716760
transform 1 0 20056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_212
timestamp 1606716760
transform 1 0 19872 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_200
timestamp 1606716760
transform 1 0 18768 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[104\]_A
timestamp 1606716760
transform 1 0 18584 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_195
timestamp 1606716760
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[0\]
timestamp 1606716760
transform 1 0 17112 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[0\]_A
timestamp 1606716760
transform 1 0 18124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_191
timestamp 1606716760
transform 1 0 17940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1606716760
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1606716760
transform 1 0 15640 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[108\]
timestamp 1606716760
transform 1 0 19872 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_211
timestamp 1606716760
transform 1 0 19780 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[50\]_B
timestamp 1606716760
transform 1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1606716760
transform 1 0 18860 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_205
timestamp 1606716760
transform 1 0 19228 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[106\]
timestamp 1606716760
transform 1 0 18032 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606716760
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_184
timestamp 1606716760
transform 1 0 17296 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_177
timestamp 1606716760
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1606716760
transform 1 0 15548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606716760
transform 1 0 20056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[108\]_A
timestamp 1606716760
transform 1 0 19872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1606716760
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[50\]_A
timestamp 1606716760
transform 1 0 19504 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_206
timestamp 1606716760
transform 1 0 19320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[50\]
timestamp 1606716760
transform 1 0 18492 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[106\]_A
timestamp 1606716760
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1606716760
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_194
timestamp 1606716760
transform 1 0 18216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1606716760
transform 1 0 16744 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1606716760
transform 1 0 15640 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[38\]
timestamp 1606716760
transform 1 0 19320 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[112\]
timestamp 1606716760
transform 1 0 18308 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_198
timestamp 1606716760
transform 1 0 18584 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[380\]
timestamp 1606716760
transform 1 0 17296 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606716760
transform 1 0 17204 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1606716760
transform 1 0 17572 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_163
timestamp 1606716760
transform 1 0 15364 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_175
timestamp 1606716760
transform 1 0 16468 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606716760
transform 1 0 20056 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1606716760
transform 1 0 19964 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_206
timestamp 1606716760
transform 1 0 19320 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[50\]_A
timestamp 1606716760
transform 1 0 19504 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[110\]
timestamp 1606716760
transform 1 0 19320 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[36\]_TE
timestamp 1606716760
transform 1 0 19872 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[38\]_TE
timestamp 1606716760
transform 1 0 19780 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1606716760
transform 1 0 19596 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_210
timestamp 1606716760
transform 1 0 19688 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_200
timestamp 1606716760
transform 1 0 18768 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_183
timestamp 1606716760
transform 1 0 17204 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[49\]
timestamp 1606716760
transform 1 0 17572 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[50\]
timestamp 1606716760
transform 1 0 18492 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_195
timestamp 1606716760
transform 1 0 18308 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1606716760
transform 1 0 18400 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_buffers\[49\]_A
timestamp 1606716760
transform 1 0 18584 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1606716760
transform 1 0 17112 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[3\]_A
timestamp 1606716760
transform 1 0 17020 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[49\]_A
timestamp 1606716760
transform 1 0 16928 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1606716760
transform 1 0 17480 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1606716760
transform 1 0 16744 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1606716760
transform 1 0 16836 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[3\]
timestamp 1606716760
transform 1 0 15180 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[49\]
timestamp 1606716760
transform 1 0 15916 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_user_to_mprj_in_gates\[49\]_B
timestamp 1606716760
transform 1 0 15732 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1606716760
transform 1 0 15180 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1606716760
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1606716760
transform 1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1606716760
transform 1 0 14536 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_143
timestamp 1606716760
transform 1 0 13524 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[39\]_A
timestamp 1606716760
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1606716760
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_131
timestamp 1606716760
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[39\]
timestamp 1606716760
transform 1 0 10396 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_8_159
timestamp 1606716760
transform 1 0 14996 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_147
timestamp 1606716760
transform 1 0 13892 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_135
timestamp 1606716760
transform 1 0 12788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606716760
transform 1 0 11592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_114
timestamp 1606716760
transform 1 0 10856 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1606716760
transform 1 0 11684 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1606716760
transform 1 0 14996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606716760
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1606716760
transform 1 0 13892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1606716760
transform 1 0 14536 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1606716760
transform 1 0 12788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_129
timestamp 1606716760
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_141
timestamp 1606716760
transform 1 0 13340 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606716760
transform 1 0 11592 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_115
timestamp 1606716760
transform 1 0 10948 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_121
timestamp 1606716760
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1606716760
transform 1 0 11684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1606716760
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606716760
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_154
timestamp 1606716760
transform 1 0 14536 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1606716760
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1606716760
transform 1 0 13340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[95\]
timestamp 1606716760
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[19\]_A
timestamp 1606716760
transform 1 0 11408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1606716760
transform 1 0 11224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_122
timestamp 1606716760
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1606716760
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1606716760
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[21\]
timestamp 1606716760
transform 1 0 11684 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606716760
transform 1 0 11592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1606716760
transform 1 0 11224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606716760
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1606716760
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1606716760
transform 1 0 14536 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[97\]
timestamp 1606716760
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[21\]_A
timestamp 1606716760
transform 1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_130
timestamp 1606716760
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_136
timestamp 1606716760
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1606716760
transform 1 0 13156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[21\]_TE
timestamp 1606716760
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[23\]_A
timestamp 1606716760
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_119
timestamp 1606716760
transform 1 0 11316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1606716760
transform 1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[77\]
timestamp 1606716760
transform 1 0 15088 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1606716760
transform 1 0 14904 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_150
timestamp 1606716760
transform 1 0 14168 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_138
timestamp 1606716760
transform 1 0 13064 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_126
timestamp 1606716760
transform 1 0 11960 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[123\]
timestamp 1606716760
transform 1 0 11684 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606716760
transform 1 0 11592 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[49\]_TE
timestamp 1606716760
transform 1 0 11040 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_114
timestamp 1606716760
transform 1 0 10856 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1606716760
transform 1 0 11224 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1606716760
transform 1 0 14720 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1606716760
transform 1 0 14628 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1606716760
transform 1 0 14904 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[3\]_TE
timestamp 1606716760
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[379\]
timestamp 1606716760
transform 1 0 14904 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_154
timestamp 1606716760
transform 1 0 14536 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_152
timestamp 1606716760
transform 1 0 14352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1606716760
transform 1 0 14260 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606716760
transform 1 0 14444 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1606716760
transform 1 0 13892 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[47\]_A
timestamp 1606716760
transform 1 0 14076 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[47\]
timestamp 1606716760
transform 1 0 12236 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[121\]
timestamp 1606716760
transform 1 0 12972 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[49\]_A
timestamp 1606716760
transform 1 0 12420 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[47\]_TE
timestamp 1606716760
transform 1 0 12052 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1606716760
transform 1 0 12236 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1606716760
transform 1 0 12604 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_140
timestamp 1606716760
transform 1 0 13248 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1606716760
transform 1 0 11776 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1606716760
transform 1 0 11868 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[49\]
timestamp 1606716760
transform 1 0 10580 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[26\]_A
timestamp 1606716760
transform 1 0 10396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[54\]_A
timestamp 1606716760
transform 1 0 10856 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_112
timestamp 1606716760
transform 1 0 10672 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116
timestamp 1606716760
transform 1 0 11040 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_108
timestamp 1606716760
transform 1 0 10304 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1606716760
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[102\]_A
timestamp 1606716760
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1606716760
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_97
timestamp 1606716760
transform 1 0 9292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_91
timestamp 1606716760
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[108\]_A
timestamp 1606716760
transform 1 0 7636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[102\]_TE
timestamp 1606716760
transform 1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1606716760
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_81
timestamp 1606716760
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_85
timestamp 1606716760
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  la_buf\[108\]
timestamp 1606716760
transform 1 0 5796 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_9_55
timestamp 1606716760
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1606716760
transform 1 0 9752 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_90
timestamp 1606716760
transform 1 0 8648 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[176\]
timestamp 1606716760
transform 1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1606716760
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_78
timestamp 1606716760
transform 1 0 7544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606716760
transform 1 0 5980 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_55
timestamp 1606716760
transform 1 0 5428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1606716760
transform 1 0 6072 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1606716760
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[93\]
timestamp 1606716760
transform 1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606716760
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_92
timestamp 1606716760
transform 1 0 8832 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_103
timestamp 1606716760
transform 1 0 9844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1606716760
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[91\]
timestamp 1606716760
transform 1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606716760
transform 1 0 7728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_73
timestamp 1606716760
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_77
timestamp 1606716760
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_89
timestamp 1606716760
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[56\]
timestamp 1606716760
transform 1 0 6072 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606716760
transform 1 0 5980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[123\]_A
timestamp 1606716760
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 1606716760
transform 1 0 5888 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1606716760
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_61
timestamp 1606716760
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[19\]
timestamp 1606716760
transform 1 0 9568 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606716760
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[19\]_TE
timestamp 1606716760
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1606716760
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1606716760
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1606716760
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1606716760
transform 1 0 7544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[56\]_A
timestamp 1606716760
transform 1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_76
timestamp 1606716760
transform 1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_80
timestamp 1606716760
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_84
timestamp 1606716760
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[125\]_A
timestamp 1606716760
transform 1 0 6532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[56\]_TE
timestamp 1606716760
transform 1 0 6900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_65
timestamp 1606716760
transform 1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_69
timestamp 1606716760
transform 1 0 6716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_106
timestamp 1606716760
transform 1 0 10120 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[17\]
timestamp 1606716760
transform 1 0 8464 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_4_80
timestamp 1606716760
transform 1 0 7728 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[14\]
timestamp 1606716760
transform 1 0 6072 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606716760
transform 1 0 5980 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[12\]_TE
timestamp 1606716760
transform 1 0 5428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1606716760
transform 1 0 5612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[23\]
timestamp 1606716760
transform 1 0 9660 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606716760
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[17\]_A
timestamp 1606716760
transform 1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[23\]_TE
timestamp 1606716760
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp 1606716760
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_97
timestamp 1606716760
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1606716760
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[102\]
timestamp 1606716760
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[14\]_A
timestamp 1606716760
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[17\]_TE
timestamp 1606716760
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1606716760
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_81
timestamp 1606716760
transform 1 0 7820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_87
timestamp 1606716760
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[12\]_A
timestamp 1606716760
transform 1 0 6624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1606716760
transform 1 0 6440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1606716760
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[26\]
timestamp 1606716760
transform 1 0 9200 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_2_94
timestamp 1606716760
transform 1 0 9016 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_86
timestamp 1606716760
transform 1 0 8280 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[28\]
timestamp 1606716760
transform 1 0 6624 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606716760
transform 1 0 5980 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[14\]_TE
timestamp 1606716760
transform 1 0 6256 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_62
timestamp 1606716760
transform 1 0 6072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1606716760
transform 1 0 6440 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[54\]
timestamp 1606716760
transform 1 0 9016 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_1_102
timestamp 1606716760
transform 1 0 9752 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_98
timestamp 1606716760
transform 1 0 9384 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_93
timestamp 1606716760
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[26\]_TE
timestamp 1606716760
transform 1 0 9200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1606716760
transform 1 0 8924 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606716760
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[100\]
timestamp 1606716760
transform 1 0 9476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1606716760
transform 1 0 8372 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[54\]_TE
timestamp 1606716760
transform 1 0 8740 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_91
timestamp 1606716760
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[130\]
timestamp 1606716760
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[52\]_A
timestamp 1606716760
transform 1 0 8004 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_81
timestamp 1606716760
transform 1 0 7820 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1606716760
transform 1 0 8004 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[28\]_A
timestamp 1606716760
transform 1 0 8188 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1606716760
transform 1 0 8188 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[28\]_TE
timestamp 1606716760
transform 1 0 7176 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1606716760
transform 1 0 7360 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[52\]
timestamp 1606716760
transform 1 0 6164 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[124\]
timestamp 1606716760
transform 1 0 6716 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1606716760
transform 1 0 6348 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1606716760
transform 1 0 6992 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[50\]_A
timestamp 1606716760
transform 1 0 5520 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[52\]_TE
timestamp 1606716760
transform 1 0 5888 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1606716760
transform 1 0 5336 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1606716760
transform 1 0 5704 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_61
timestamp 1606716760
transform 1 0 5980 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1606716760
transform 1 0 6072 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[41\]_A
timestamp 1606716760
transform 1 0 6164 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[120\]_A
timestamp 1606716760
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_51
timestamp 1606716760
transform 1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[120\]
timestamp 1606716760
transform 1 0 3404 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[194\]
timestamp 1606716760
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1606716760
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1606716760
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_23
timestamp 1606716760
transform 1 0 2484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_32
timestamp 1606716760
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606716760
transform 1 0 368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606716760
transform 1 0 644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1606716760
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[105\]_A
timestamp 1606716760
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_51
timestamp 1606716760
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[105\]
timestamp 1606716760
transform 1 0 3404 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_8_27
timestamp 1606716760
transform 1 0 2852 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606716760
transform 1 0 368 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606716760
transform 1 0 644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606716760
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[123\]
timestamp 1606716760
transform 1 0 3956 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[0\]
timestamp 1606716760
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[123\]_TE
timestamp 1606716760
transform 1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1606716760
transform 1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_48
timestamp 1606716760
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[197\]
timestamp 1606716760
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606716760
transform 1 0 3220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[105\]_TE
timestamp 1606716760
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_27
timestamp 1606716760
transform 1 0 2852 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp 1606716760
transform 1 0 3404 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1606716760
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1606716760
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_32
timestamp 1606716760
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp 1606716760
transform 1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606716760
transform 1 0 368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606716760
transform 1 0 368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606716760
transform 1 0 644 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606716760
transform 1 0 1748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606716760
transform 1 0 644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606716760
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[125\]
timestamp 1606716760
transform 1 0 4692 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[125\]_TE
timestamp 1606716760
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_39
timestamp 1606716760
transform 1 0 3956 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[199\]
timestamp 1606716760
transform 1 0 3680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606716760
transform 1 0 3220 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1606716760
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1606716760
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606716760
transform 1 0 368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606716760
transform 1 0 644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606716760
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_53
timestamp 1606716760
transform 1 0 5244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[88\]
timestamp 1606716760
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  mprj_rstn_buf
timestamp 1606716760
transform 1 0 3588 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_4_23
timestamp 1606716760
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_27
timestamp 1606716760
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606716760
transform 1 0 368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606716760
transform 1 0 644 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_15
timestamp 1606716760
transform 1 0 1748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[12\]
timestamp 1606716760
transform 1 0 4784 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1606716760
transform 1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_rstn_buf_A
timestamp 1606716760
transform 1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_40
timestamp 1606716760
transform 1 0 4048 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1606716760
transform 1 0 4416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1606716760
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[86\]
timestamp 1606716760
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606716760
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mprj_rstn_buf_TE
timestamp 1606716760
transform 1 0 3588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1606716760
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_23
timestamp 1606716760
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_32
timestamp 1606716760
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606716760
transform 1 0 368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606716760
transform 1 0 644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1606716760
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_53
timestamp 1606716760
transform 1 0 5244 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[43\]_A
timestamp 1606716760
transform 1 0 5060 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1606716760
transform 1 0 4876 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[43\]
timestamp 1606716760
transform 1 0 3220 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[117\]
timestamp 1606716760
transform 1 0 2208 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_19
timestamp 1606716760
transform 1 0 2116 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1606716760
transform 1 0 2484 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606716760
transform 1 0 368 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606716760
transform 1 0 644 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1606716760
transform 1 0 1748 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[41\]
timestamp 1606716760
transform 1 0 4324 0 1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[41\]_TE
timestamp 1606716760
transform 1 0 4140 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1606716760
transform 1 0 3956 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[50\]
timestamp 1606716760
transform 1 0 3680 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[115\]
timestamp 1606716760
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606716760
transform 1 0 3220 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1606716760
transform 1 0 3220 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[43\]_TE
timestamp 1606716760
transform 1 0 3772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_la_buf\[50\]_TE
timestamp 1606716760
transform 1 0 3496 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1606716760
transform 1 0 3312 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1606716760
transform 1 0 3588 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[126\]
timestamp 1606716760
transform 1 0 2208 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[128\]
timestamp 1606716760
transform 1 0 2208 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19
timestamp 1606716760
transform 1 0 2116 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23
timestamp 1606716760
transform 1 0 2484 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19
timestamp 1606716760
transform 1 0 2116 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_23
timestamp 1606716760
transform 1 0 2484 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606716760
transform 1 0 368 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606716760
transform 1 0 368 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1606716760
transform 1 0 644 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1606716760
transform 1 0 1748 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606716760
transform 1 0 644 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1606716760
transform 1 0 1748 0 1 1088
box -38 -48 406 592
<< labels >>
rlabel metal2 s 570 0 626 800 4 caravel_clk
port 1 nsew
rlabel metal2 s 938 0 994 800 4 caravel_clk2
port 2 nsew
rlabel metal3 s 0 1096 800 1216 4 caravel_rstn
port 3 nsew
rlabel metal2 s 754 12200 810 13000 4 la_data_in_core[0]
port 4 nsew
rlabel metal3 s 0 11976 800 12096 4 la_data_in_core[100]
port 5 nsew
rlabel metal2 s 1122 12200 1178 13000 4 la_data_in_core[101]
port 6 nsew
rlabel metal3 s 0 11432 800 11552 4 la_data_in_core[102]
port 7 nsew
rlabel metal2 s 1490 12200 1546 13000 4 la_data_in_core[103]
port 8 nsew
rlabel metal2 s 1858 12200 1914 13000 4 la_data_in_core[104]
port 9 nsew
rlabel metal3 s 0 10888 800 11008 4 la_data_in_core[105]
port 10 nsew
rlabel metal2 s 2226 12200 2282 13000 4 la_data_in_core[106]
port 11 nsew
rlabel metal3 s 0 10344 800 10464 4 la_data_in_core[107]
port 12 nsew
rlabel metal2 s 2594 12200 2650 13000 4 la_data_in_core[108]
port 13 nsew
rlabel metal2 s 2962 12200 3018 13000 4 la_data_in_core[109]
port 14 nsew
rlabel metal3 s 0 9800 800 9920 4 la_data_in_core[10]
port 15 nsew
rlabel metal2 s 3330 12200 3386 13000 4 la_data_in_core[110]
port 16 nsew
rlabel metal3 s 0 9256 800 9376 4 la_data_in_core[111]
port 17 nsew
rlabel metal2 s 3698 12200 3754 13000 4 la_data_in_core[112]
port 18 nsew
rlabel metal2 s 4066 12200 4122 13000 4 la_data_in_core[113]
port 19 nsew
rlabel metal3 s 0 8712 800 8832 4 la_data_in_core[114]
port 20 nsew
rlabel metal2 s 4434 12200 4490 13000 4 la_data_in_core[115]
port 21 nsew
rlabel metal3 s 0 8168 800 8288 4 la_data_in_core[116]
port 22 nsew
rlabel metal2 s 4802 12200 4858 13000 4 la_data_in_core[117]
port 23 nsew
rlabel metal2 s 5170 12200 5226 13000 4 la_data_in_core[118]
port 24 nsew
rlabel metal3 s 0 7624 800 7744 4 la_data_in_core[119]
port 25 nsew
rlabel metal2 s 5538 12200 5594 13000 4 la_data_in_core[11]
port 26 nsew
rlabel metal3 s 0 7080 800 7200 4 la_data_in_core[120]
port 27 nsew
rlabel metal2 s 5906 12200 5962 13000 4 la_data_in_core[121]
port 28 nsew
rlabel metal2 s 6274 12200 6330 13000 4 la_data_in_core[122]
port 29 nsew
rlabel metal3 s 0 6536 800 6656 4 la_data_in_core[123]
port 30 nsew
rlabel metal2 s 6642 12200 6698 13000 4 la_data_in_core[124]
port 31 nsew
rlabel metal3 s 0 5992 800 6112 4 la_data_in_core[125]
port 32 nsew
rlabel metal2 s 7010 12200 7066 13000 4 la_data_in_core[126]
port 33 nsew
rlabel metal2 s 7378 12200 7434 13000 4 la_data_in_core[127]
port 34 nsew
rlabel metal3 s 0 5448 800 5568 4 la_data_in_core[12]
port 35 nsew
rlabel metal2 s 7746 12200 7802 13000 4 la_data_in_core[13]
port 36 nsew
rlabel metal3 s 0 4904 800 5024 4 la_data_in_core[14]
port 37 nsew
rlabel metal2 s 8114 12200 8170 13000 4 la_data_in_core[15]
port 38 nsew
rlabel metal2 s 8482 12200 8538 13000 4 la_data_in_core[16]
port 39 nsew
rlabel metal3 s 0 4360 800 4480 4 la_data_in_core[17]
port 40 nsew
rlabel metal2 s 8850 12200 8906 13000 4 la_data_in_core[18]
port 41 nsew
rlabel metal3 s 0 3816 800 3936 4 la_data_in_core[19]
port 42 nsew
rlabel metal2 s 9218 12200 9274 13000 4 la_data_in_core[1]
port 43 nsew
rlabel metal2 s 9586 12200 9642 13000 4 la_data_in_core[20]
port 44 nsew
rlabel metal3 s 0 3272 800 3392 4 la_data_in_core[21]
port 45 nsew
rlabel metal2 s 9954 12200 10010 13000 4 la_data_in_core[22]
port 46 nsew
rlabel metal3 s 0 2728 800 2848 4 la_data_in_core[23]
port 47 nsew
rlabel metal2 s 10322 12200 10378 13000 4 la_data_in_core[24]
port 48 nsew
rlabel metal2 s 10690 12200 10746 13000 4 la_data_in_core[25]
port 49 nsew
rlabel metal3 s 0 2184 800 2304 4 la_data_in_core[26]
port 50 nsew
rlabel metal2 s 11058 12200 11114 13000 4 la_data_in_core[27]
port 51 nsew
rlabel metal3 s 0 1640 800 1760 4 la_data_in_core[28]
port 52 nsew
rlabel metal2 s 11426 12200 11482 13000 4 la_data_in_core[29]
port 53 nsew
rlabel metal2 s 11794 12200 11850 13000 4 la_data_in_core[2]
port 54 nsew
rlabel metal2 s 12162 12200 12218 13000 4 la_data_in_core[30]
port 55 nsew
rlabel metal2 s 12530 12200 12586 13000 4 la_data_in_core[31]
port 56 nsew
rlabel metal2 s 12898 12200 12954 13000 4 la_data_in_core[32]
port 57 nsew
rlabel metal2 s 13266 12200 13322 13000 4 la_data_in_core[33]
port 58 nsew
rlabel metal2 s 13634 12200 13690 13000 4 la_data_in_core[34]
port 59 nsew
rlabel metal2 s 14002 12200 14058 13000 4 la_data_in_core[35]
port 60 nsew
rlabel metal2 s 1306 0 1362 800 4 la_data_in_core[36]
port 61 nsew
rlabel metal2 s 14370 12200 14426 13000 4 la_data_in_core[37]
port 62 nsew
rlabel metal2 s 1674 0 1730 800 4 la_data_in_core[38]
port 63 nsew
rlabel metal2 s 14738 12200 14794 13000 4 la_data_in_core[39]
port 64 nsew
rlabel metal2 s 2042 0 2098 800 4 la_data_in_core[3]
port 65 nsew
rlabel metal2 s 15106 12200 15162 13000 4 la_data_in_core[40]
port 66 nsew
rlabel metal2 s 2410 0 2466 800 4 la_data_in_core[41]
port 67 nsew
rlabel metal2 s 15474 12200 15530 13000 4 la_data_in_core[42]
port 68 nsew
rlabel metal2 s 2778 0 2834 800 4 la_data_in_core[43]
port 69 nsew
rlabel metal2 s 15842 12200 15898 13000 4 la_data_in_core[44]
port 70 nsew
rlabel metal2 s 3146 0 3202 800 4 la_data_in_core[45]
port 71 nsew
rlabel metal2 s 16210 12200 16266 13000 4 la_data_in_core[46]
port 72 nsew
rlabel metal2 s 3514 0 3570 800 4 la_data_in_core[47]
port 73 nsew
rlabel metal2 s 16578 12200 16634 13000 4 la_data_in_core[48]
port 74 nsew
rlabel metal2 s 3882 0 3938 800 4 la_data_in_core[49]
port 75 nsew
rlabel metal2 s 16946 12200 17002 13000 4 la_data_in_core[4]
port 76 nsew
rlabel metal2 s 4250 0 4306 800 4 la_data_in_core[50]
port 77 nsew
rlabel metal2 s 17314 12200 17370 13000 4 la_data_in_core[51]
port 78 nsew
rlabel metal2 s 4618 0 4674 800 4 la_data_in_core[52]
port 79 nsew
rlabel metal2 s 17682 12200 17738 13000 4 la_data_in_core[53]
port 80 nsew
rlabel metal2 s 4986 0 5042 800 4 la_data_in_core[54]
port 81 nsew
rlabel metal2 s 18050 12200 18106 13000 4 la_data_in_core[55]
port 82 nsew
rlabel metal2 s 5354 0 5410 800 4 la_data_in_core[56]
port 83 nsew
rlabel metal2 s 18418 12200 18474 13000 4 la_data_in_core[57]
port 84 nsew
rlabel metal2 s 5722 0 5778 800 4 la_data_in_core[58]
port 85 nsew
rlabel metal2 s 18786 12200 18842 13000 4 la_data_in_core[59]
port 86 nsew
rlabel metal2 s 6090 0 6146 800 4 la_data_in_core[5]
port 87 nsew
rlabel metal2 s 19154 12200 19210 13000 4 la_data_in_core[60]
port 88 nsew
rlabel metal2 s 6458 0 6514 800 4 la_data_in_core[61]
port 89 nsew
rlabel metal2 s 19522 12200 19578 13000 4 la_data_in_core[62]
port 90 nsew
rlabel metal2 s 6826 0 6882 800 4 la_data_in_core[63]
port 91 nsew
rlabel metal2 s 19890 12200 19946 13000 4 la_data_in_core[64]
port 92 nsew
rlabel metal2 s 7194 0 7250 800 4 la_data_in_core[65]
port 93 nsew
rlabel metal2 s 20258 12200 20314 13000 4 la_data_in_core[66]
port 94 nsew
rlabel metal2 s 7562 0 7618 800 4 la_data_in_core[67]
port 95 nsew
rlabel metal2 s 20626 12200 20682 13000 4 la_data_in_core[68]
port 96 nsew
rlabel metal2 s 7930 0 7986 800 4 la_data_in_core[69]
port 97 nsew
rlabel metal2 s 20994 12200 21050 13000 4 la_data_in_core[6]
port 98 nsew
rlabel metal2 s 8298 0 8354 800 4 la_data_in_core[70]
port 99 nsew
rlabel metal2 s 21362 12200 21418 13000 4 la_data_in_core[71]
port 100 nsew
rlabel metal2 s 8666 0 8722 800 4 la_data_in_core[72]
port 101 nsew
rlabel metal2 s 21730 12200 21786 13000 4 la_data_in_core[73]
port 102 nsew
rlabel metal2 s 9034 0 9090 800 4 la_data_in_core[74]
port 103 nsew
rlabel metal2 s 22098 12200 22154 13000 4 la_data_in_core[75]
port 104 nsew
rlabel metal2 s 9402 0 9458 800 4 la_data_in_core[76]
port 105 nsew
rlabel metal2 s 22466 12200 22522 13000 4 la_data_in_core[77]
port 106 nsew
rlabel metal2 s 9770 0 9826 800 4 la_data_in_core[78]
port 107 nsew
rlabel metal2 s 22834 12200 22890 13000 4 la_data_in_core[79]
port 108 nsew
rlabel metal2 s 10138 0 10194 800 4 la_data_in_core[7]
port 109 nsew
rlabel metal2 s 23202 12200 23258 13000 4 la_data_in_core[80]
port 110 nsew
rlabel metal2 s 10506 0 10562 800 4 la_data_in_core[81]
port 111 nsew
rlabel metal2 s 23570 12200 23626 13000 4 la_data_in_core[82]
port 112 nsew
rlabel metal2 s 10874 0 10930 800 4 la_data_in_core[83]
port 113 nsew
rlabel metal2 s 23938 12200 23994 13000 4 la_data_in_core[84]
port 114 nsew
rlabel metal2 s 11242 0 11298 800 4 la_data_in_core[85]
port 115 nsew
rlabel metal2 s 24306 12200 24362 13000 4 la_data_in_core[86]
port 116 nsew
rlabel metal2 s 11610 0 11666 800 4 la_data_in_core[87]
port 117 nsew
rlabel metal2 s 24674 12200 24730 13000 4 la_data_in_core[88]
port 118 nsew
rlabel metal2 s 11978 0 12034 800 4 la_data_in_core[89]
port 119 nsew
rlabel metal2 s 25042 12200 25098 13000 4 la_data_in_core[8]
port 120 nsew
rlabel metal2 s 12346 0 12402 800 4 la_data_in_core[90]
port 121 nsew
rlabel metal2 s 25410 12200 25466 13000 4 la_data_in_core[91]
port 122 nsew
rlabel metal2 s 12714 0 12770 800 4 la_data_in_core[92]
port 123 nsew
rlabel metal2 s 25778 12200 25834 13000 4 la_data_in_core[93]
port 124 nsew
rlabel metal2 s 13082 0 13138 800 4 la_data_in_core[94]
port 125 nsew
rlabel metal2 s 26146 12200 26202 13000 4 la_data_in_core[95]
port 126 nsew
rlabel metal2 s 13450 0 13506 800 4 la_data_in_core[96]
port 127 nsew
rlabel metal2 s 26514 12200 26570 13000 4 la_data_in_core[97]
port 128 nsew
rlabel metal2 s 13818 0 13874 800 4 la_data_in_core[98]
port 129 nsew
rlabel metal2 s 26882 12200 26938 13000 4 la_data_in_core[99]
port 130 nsew
rlabel metal2 s 14186 0 14242 800 4 la_data_in_core[9]
port 131 nsew
rlabel metal2 s 14554 0 14610 800 4 la_data_in_mprj[0]
port 132 nsew
rlabel metal2 s 14922 0 14978 800 4 la_data_in_mprj[100]
port 133 nsew
rlabel metal2 s 15290 0 15346 800 4 la_data_in_mprj[101]
port 134 nsew
rlabel metal2 s 15658 0 15714 800 4 la_data_in_mprj[102]
port 135 nsew
rlabel metal2 s 16026 0 16082 800 4 la_data_in_mprj[103]
port 136 nsew
rlabel metal2 s 16394 0 16450 800 4 la_data_in_mprj[104]
port 137 nsew
rlabel metal2 s 16762 0 16818 800 4 la_data_in_mprj[105]
port 138 nsew
rlabel metal2 s 17130 0 17186 800 4 la_data_in_mprj[106]
port 139 nsew
rlabel metal2 s 17498 0 17554 800 4 la_data_in_mprj[107]
port 140 nsew
rlabel metal2 s 17866 0 17922 800 4 la_data_in_mprj[108]
port 141 nsew
rlabel metal2 s 18234 0 18290 800 4 la_data_in_mprj[109]
port 142 nsew
rlabel metal2 s 18602 0 18658 800 4 la_data_in_mprj[10]
port 143 nsew
rlabel metal2 s 18970 0 19026 800 4 la_data_in_mprj[110]
port 144 nsew
rlabel metal2 s 19338 0 19394 800 4 la_data_in_mprj[111]
port 145 nsew
rlabel metal2 s 19706 0 19762 800 4 la_data_in_mprj[112]
port 146 nsew
rlabel metal2 s 20074 0 20130 800 4 la_data_in_mprj[113]
port 147 nsew
rlabel metal2 s 20442 0 20498 800 4 la_data_in_mprj[114]
port 148 nsew
rlabel metal2 s 20810 0 20866 800 4 la_data_in_mprj[115]
port 149 nsew
rlabel metal2 s 21178 0 21234 800 4 la_data_in_mprj[116]
port 150 nsew
rlabel metal2 s 21546 0 21602 800 4 la_data_in_mprj[117]
port 151 nsew
rlabel metal2 s 21914 0 21970 800 4 la_data_in_mprj[118]
port 152 nsew
rlabel metal2 s 22282 0 22338 800 4 la_data_in_mprj[119]
port 153 nsew
rlabel metal2 s 22650 0 22706 800 4 la_data_in_mprj[11]
port 154 nsew
rlabel metal2 s 23018 0 23074 800 4 la_data_in_mprj[120]
port 155 nsew
rlabel metal2 s 23386 0 23442 800 4 la_data_in_mprj[121]
port 156 nsew
rlabel metal2 s 23754 0 23810 800 4 la_data_in_mprj[122]
port 157 nsew
rlabel metal2 s 24122 0 24178 800 4 la_data_in_mprj[123]
port 158 nsew
rlabel metal2 s 24490 0 24546 800 4 la_data_in_mprj[124]
port 159 nsew
rlabel metal2 s 24858 0 24914 800 4 la_data_in_mprj[125]
port 160 nsew
rlabel metal2 s 25226 0 25282 800 4 la_data_in_mprj[126]
port 161 nsew
rlabel metal2 s 25594 0 25650 800 4 la_data_in_mprj[127]
port 162 nsew
rlabel metal2 s 25962 0 26018 800 4 la_data_in_mprj[12]
port 163 nsew
rlabel metal2 s 26330 0 26386 800 4 la_data_in_mprj[13]
port 164 nsew
rlabel metal2 s 26698 0 26754 800 4 la_data_in_mprj[14]
port 165 nsew
rlabel metal2 s 27066 0 27122 800 4 la_data_in_mprj[15]
port 166 nsew
rlabel metal2 s 27434 0 27490 800 4 la_data_in_mprj[16]
port 167 nsew
rlabel metal2 s 27802 0 27858 800 4 la_data_in_mprj[17]
port 168 nsew
rlabel metal2 s 28170 0 28226 800 4 la_data_in_mprj[18]
port 169 nsew
rlabel metal2 s 28538 0 28594 800 4 la_data_in_mprj[19]
port 170 nsew
rlabel metal2 s 28906 0 28962 800 4 la_data_in_mprj[1]
port 171 nsew
rlabel metal2 s 29274 0 29330 800 4 la_data_in_mprj[20]
port 172 nsew
rlabel metal2 s 29642 0 29698 800 4 la_data_in_mprj[21]
port 173 nsew
rlabel metal2 s 30010 0 30066 800 4 la_data_in_mprj[22]
port 174 nsew
rlabel metal2 s 30378 0 30434 800 4 la_data_in_mprj[23]
port 175 nsew
rlabel metal2 s 30746 0 30802 800 4 la_data_in_mprj[24]
port 176 nsew
rlabel metal2 s 31114 0 31170 800 4 la_data_in_mprj[25]
port 177 nsew
rlabel metal2 s 31482 0 31538 800 4 la_data_in_mprj[26]
port 178 nsew
rlabel metal2 s 31850 0 31906 800 4 la_data_in_mprj[27]
port 179 nsew
rlabel metal2 s 32218 0 32274 800 4 la_data_in_mprj[28]
port 180 nsew
rlabel metal2 s 32586 0 32642 800 4 la_data_in_mprj[29]
port 181 nsew
rlabel metal2 s 32954 0 33010 800 4 la_data_in_mprj[2]
port 182 nsew
rlabel metal2 s 33322 0 33378 800 4 la_data_in_mprj[30]
port 183 nsew
rlabel metal2 s 33690 0 33746 800 4 la_data_in_mprj[31]
port 184 nsew
rlabel metal2 s 34058 0 34114 800 4 la_data_in_mprj[32]
port 185 nsew
rlabel metal2 s 34426 0 34482 800 4 la_data_in_mprj[33]
port 186 nsew
rlabel metal2 s 34794 0 34850 800 4 la_data_in_mprj[34]
port 187 nsew
rlabel metal2 s 35162 0 35218 800 4 la_data_in_mprj[35]
port 188 nsew
rlabel metal2 s 35530 0 35586 800 4 la_data_in_mprj[36]
port 189 nsew
rlabel metal2 s 35898 0 35954 800 4 la_data_in_mprj[37]
port 190 nsew
rlabel metal2 s 36266 0 36322 800 4 la_data_in_mprj[38]
port 191 nsew
rlabel metal2 s 36634 0 36690 800 4 la_data_in_mprj[39]
port 192 nsew
rlabel metal2 s 37002 0 37058 800 4 la_data_in_mprj[3]
port 193 nsew
rlabel metal2 s 37370 0 37426 800 4 la_data_in_mprj[40]
port 194 nsew
rlabel metal2 s 37738 0 37794 800 4 la_data_in_mprj[41]
port 195 nsew
rlabel metal2 s 38106 0 38162 800 4 la_data_in_mprj[42]
port 196 nsew
rlabel metal2 s 38474 0 38530 800 4 la_data_in_mprj[43]
port 197 nsew
rlabel metal2 s 38842 0 38898 800 4 la_data_in_mprj[44]
port 198 nsew
rlabel metal2 s 39210 0 39266 800 4 la_data_in_mprj[45]
port 199 nsew
rlabel metal2 s 39578 0 39634 800 4 la_data_in_mprj[46]
port 200 nsew
rlabel metal2 s 39946 0 40002 800 4 la_data_in_mprj[47]
port 201 nsew
rlabel metal2 s 27250 12200 27306 13000 4 la_data_in_mprj[48]
port 202 nsew
rlabel metal2 s 40314 0 40370 800 4 la_data_in_mprj[49]
port 203 nsew
rlabel metal2 s 27618 12200 27674 13000 4 la_data_in_mprj[4]
port 204 nsew
rlabel metal2 s 40682 0 40738 800 4 la_data_in_mprj[50]
port 205 nsew
rlabel metal2 s 27986 12200 28042 13000 4 la_data_in_mprj[51]
port 206 nsew
rlabel metal2 s 41050 0 41106 800 4 la_data_in_mprj[52]
port 207 nsew
rlabel metal2 s 28354 12200 28410 13000 4 la_data_in_mprj[53]
port 208 nsew
rlabel metal2 s 41418 0 41474 800 4 la_data_in_mprj[54]
port 209 nsew
rlabel metal2 s 28722 12200 28778 13000 4 la_data_in_mprj[55]
port 210 nsew
rlabel metal2 s 41786 0 41842 800 4 la_data_in_mprj[56]
port 211 nsew
rlabel metal2 s 29090 12200 29146 13000 4 la_data_in_mprj[57]
port 212 nsew
rlabel metal2 s 42154 0 42210 800 4 la_data_in_mprj[58]
port 213 nsew
rlabel metal2 s 29458 12200 29514 13000 4 la_data_in_mprj[59]
port 214 nsew
rlabel metal2 s 42522 0 42578 800 4 la_data_in_mprj[5]
port 215 nsew
rlabel metal2 s 29826 12200 29882 13000 4 la_data_in_mprj[60]
port 216 nsew
rlabel metal2 s 42890 0 42946 800 4 la_data_in_mprj[61]
port 217 nsew
rlabel metal2 s 30194 12200 30250 13000 4 la_data_in_mprj[62]
port 218 nsew
rlabel metal2 s 43258 0 43314 800 4 la_data_in_mprj[63]
port 219 nsew
rlabel metal2 s 30562 12200 30618 13000 4 la_data_in_mprj[64]
port 220 nsew
rlabel metal2 s 43626 0 43682 800 4 la_data_in_mprj[65]
port 221 nsew
rlabel metal2 s 30930 12200 30986 13000 4 la_data_in_mprj[66]
port 222 nsew
rlabel metal2 s 43994 0 44050 800 4 la_data_in_mprj[67]
port 223 nsew
rlabel metal2 s 31298 12200 31354 13000 4 la_data_in_mprj[68]
port 224 nsew
rlabel metal2 s 44362 0 44418 800 4 la_data_in_mprj[69]
port 225 nsew
rlabel metal2 s 31666 12200 31722 13000 4 la_data_in_mprj[6]
port 226 nsew
rlabel metal2 s 44730 0 44786 800 4 la_data_in_mprj[70]
port 227 nsew
rlabel metal2 s 32034 12200 32090 13000 4 la_data_in_mprj[71]
port 228 nsew
rlabel metal2 s 45098 0 45154 800 4 la_data_in_mprj[72]
port 229 nsew
rlabel metal2 s 32402 12200 32458 13000 4 la_data_in_mprj[73]
port 230 nsew
rlabel metal2 s 45466 0 45522 800 4 la_data_in_mprj[74]
port 231 nsew
rlabel metal2 s 32770 12200 32826 13000 4 la_data_in_mprj[75]
port 232 nsew
rlabel metal2 s 45834 0 45890 800 4 la_data_in_mprj[76]
port 233 nsew
rlabel metal2 s 33138 12200 33194 13000 4 la_data_in_mprj[77]
port 234 nsew
rlabel metal2 s 46202 0 46258 800 4 la_data_in_mprj[78]
port 235 nsew
rlabel metal2 s 33506 12200 33562 13000 4 la_data_in_mprj[79]
port 236 nsew
rlabel metal2 s 46570 0 46626 800 4 la_data_in_mprj[7]
port 237 nsew
rlabel metal2 s 33874 12200 33930 13000 4 la_data_in_mprj[80]
port 238 nsew
rlabel metal2 s 46938 0 46994 800 4 la_data_in_mprj[81]
port 239 nsew
rlabel metal2 s 34242 12200 34298 13000 4 la_data_in_mprj[82]
port 240 nsew
rlabel metal2 s 47306 0 47362 800 4 la_data_in_mprj[83]
port 241 nsew
rlabel metal2 s 34610 12200 34666 13000 4 la_data_in_mprj[84]
port 242 nsew
rlabel metal2 s 47674 0 47730 800 4 la_data_in_mprj[85]
port 243 nsew
rlabel metal2 s 34978 12200 35034 13000 4 la_data_in_mprj[86]
port 244 nsew
rlabel metal2 s 48042 0 48098 800 4 la_data_in_mprj[87]
port 245 nsew
rlabel metal2 s 35346 12200 35402 13000 4 la_data_in_mprj[88]
port 246 nsew
rlabel metal2 s 48410 0 48466 800 4 la_data_in_mprj[89]
port 247 nsew
rlabel metal2 s 35714 12200 35770 13000 4 la_data_in_mprj[8]
port 248 nsew
rlabel metal2 s 48778 0 48834 800 4 la_data_in_mprj[90]
port 249 nsew
rlabel metal2 s 36082 12200 36138 13000 4 la_data_in_mprj[91]
port 250 nsew
rlabel metal2 s 49146 0 49202 800 4 la_data_in_mprj[92]
port 251 nsew
rlabel metal2 s 36450 12200 36506 13000 4 la_data_in_mprj[93]
port 252 nsew
rlabel metal2 s 49514 0 49570 800 4 la_data_in_mprj[94]
port 253 nsew
rlabel metal2 s 36818 12200 36874 13000 4 la_data_in_mprj[95]
port 254 nsew
rlabel metal2 s 49882 0 49938 800 4 la_data_in_mprj[96]
port 255 nsew
rlabel metal2 s 37186 12200 37242 13000 4 la_data_in_mprj[97]
port 256 nsew
rlabel metal2 s 50250 0 50306 800 4 la_data_in_mprj[98]
port 257 nsew
rlabel metal2 s 37554 12200 37610 13000 4 la_data_in_mprj[99]
port 258 nsew
rlabel metal2 s 50618 0 50674 800 4 la_data_in_mprj[9]
port 259 nsew
rlabel metal2 s 37922 12200 37978 13000 4 la_data_out_core[0]
port 260 nsew
rlabel metal2 s 38290 12200 38346 13000 4 la_data_out_core[100]
port 261 nsew
rlabel metal2 s 38658 12200 38714 13000 4 la_data_out_core[101]
port 262 nsew
rlabel metal2 s 39026 12200 39082 13000 4 la_data_out_core[102]
port 263 nsew
rlabel metal2 s 39394 12200 39450 13000 4 la_data_out_core[103]
port 264 nsew
rlabel metal2 s 39762 12200 39818 13000 4 la_data_out_core[104]
port 265 nsew
rlabel metal2 s 40130 12200 40186 13000 4 la_data_out_core[105]
port 266 nsew
rlabel metal2 s 40498 12200 40554 13000 4 la_data_out_core[106]
port 267 nsew
rlabel metal2 s 40866 12200 40922 13000 4 la_data_out_core[107]
port 268 nsew
rlabel metal2 s 41234 12200 41290 13000 4 la_data_out_core[108]
port 269 nsew
rlabel metal2 s 41602 12200 41658 13000 4 la_data_out_core[109]
port 270 nsew
rlabel metal2 s 41970 12200 42026 13000 4 la_data_out_core[10]
port 271 nsew
rlabel metal2 s 42338 12200 42394 13000 4 la_data_out_core[110]
port 272 nsew
rlabel metal2 s 42706 12200 42762 13000 4 la_data_out_core[111]
port 273 nsew
rlabel metal2 s 43074 12200 43130 13000 4 la_data_out_core[112]
port 274 nsew
rlabel metal2 s 43442 12200 43498 13000 4 la_data_out_core[113]
port 275 nsew
rlabel metal2 s 43810 12200 43866 13000 4 la_data_out_core[114]
port 276 nsew
rlabel metal2 s 44178 12200 44234 13000 4 la_data_out_core[115]
port 277 nsew
rlabel metal2 s 44546 12200 44602 13000 4 la_data_out_core[116]
port 278 nsew
rlabel metal2 s 44914 12200 44970 13000 4 la_data_out_core[117]
port 279 nsew
rlabel metal2 s 45282 12200 45338 13000 4 la_data_out_core[118]
port 280 nsew
rlabel metal2 s 45650 12200 45706 13000 4 la_data_out_core[119]
port 281 nsew
rlabel metal2 s 46018 12200 46074 13000 4 la_data_out_core[11]
port 282 nsew
rlabel metal2 s 46386 12200 46442 13000 4 la_data_out_core[120]
port 283 nsew
rlabel metal2 s 46754 12200 46810 13000 4 la_data_out_core[121]
port 284 nsew
rlabel metal2 s 47122 12200 47178 13000 4 la_data_out_core[122]
port 285 nsew
rlabel metal2 s 47490 12200 47546 13000 4 la_data_out_core[123]
port 286 nsew
rlabel metal2 s 47858 12200 47914 13000 4 la_data_out_core[124]
port 287 nsew
rlabel metal2 s 48226 12200 48282 13000 4 la_data_out_core[125]
port 288 nsew
rlabel metal2 s 48594 12200 48650 13000 4 la_data_out_core[126]
port 289 nsew
rlabel metal2 s 48962 12200 49018 13000 4 la_data_out_core[127]
port 290 nsew
rlabel metal2 s 49330 12200 49386 13000 4 la_data_out_core[12]
port 291 nsew
rlabel metal2 s 49698 12200 49754 13000 4 la_data_out_core[13]
port 292 nsew
rlabel metal2 s 50066 12200 50122 13000 4 la_data_out_core[14]
port 293 nsew
rlabel metal2 s 50434 12200 50490 13000 4 la_data_out_core[15]
port 294 nsew
rlabel metal2 s 50802 12200 50858 13000 4 la_data_out_core[16]
port 295 nsew
rlabel metal2 s 51170 12200 51226 13000 4 la_data_out_core[17]
port 296 nsew
rlabel metal2 s 51538 12200 51594 13000 4 la_data_out_core[18]
port 297 nsew
rlabel metal2 s 51906 12200 51962 13000 4 la_data_out_core[19]
port 298 nsew
rlabel metal2 s 52274 12200 52330 13000 4 la_data_out_core[1]
port 299 nsew
rlabel metal2 s 52642 12200 52698 13000 4 la_data_out_core[20]
port 300 nsew
rlabel metal2 s 53010 12200 53066 13000 4 la_data_out_core[21]
port 301 nsew
rlabel metal2 s 53378 12200 53434 13000 4 la_data_out_core[22]
port 302 nsew
rlabel metal2 s 53746 12200 53802 13000 4 la_data_out_core[23]
port 303 nsew
rlabel metal2 s 54114 12200 54170 13000 4 la_data_out_core[24]
port 304 nsew
rlabel metal2 s 54482 12200 54538 13000 4 la_data_out_core[25]
port 305 nsew
rlabel metal2 s 54850 12200 54906 13000 4 la_data_out_core[26]
port 306 nsew
rlabel metal2 s 55218 12200 55274 13000 4 la_data_out_core[27]
port 307 nsew
rlabel metal2 s 55586 12200 55642 13000 4 la_data_out_core[28]
port 308 nsew
rlabel metal2 s 55954 12200 56010 13000 4 la_data_out_core[29]
port 309 nsew
rlabel metal2 s 56322 12200 56378 13000 4 la_data_out_core[2]
port 310 nsew
rlabel metal2 s 56690 12200 56746 13000 4 la_data_out_core[30]
port 311 nsew
rlabel metal2 s 57058 12200 57114 13000 4 la_data_out_core[31]
port 312 nsew
rlabel metal2 s 57426 12200 57482 13000 4 la_data_out_core[32]
port 313 nsew
rlabel metal2 s 57794 12200 57850 13000 4 la_data_out_core[33]
port 314 nsew
rlabel metal2 s 58162 12200 58218 13000 4 la_data_out_core[34]
port 315 nsew
rlabel metal2 s 58530 12200 58586 13000 4 la_data_out_core[35]
port 316 nsew
rlabel metal2 s 58898 12200 58954 13000 4 la_data_out_core[36]
port 317 nsew
rlabel metal2 s 59266 12200 59322 13000 4 la_data_out_core[37]
port 318 nsew
rlabel metal2 s 59634 12200 59690 13000 4 la_data_out_core[38]
port 319 nsew
rlabel metal2 s 60002 12200 60058 13000 4 la_data_out_core[39]
port 320 nsew
rlabel metal2 s 60370 12200 60426 13000 4 la_data_out_core[3]
port 321 nsew
rlabel metal2 s 60738 12200 60794 13000 4 la_data_out_core[40]
port 322 nsew
rlabel metal2 s 61106 12200 61162 13000 4 la_data_out_core[41]
port 323 nsew
rlabel metal2 s 61474 12200 61530 13000 4 la_data_out_core[42]
port 324 nsew
rlabel metal2 s 61842 12200 61898 13000 4 la_data_out_core[43]
port 325 nsew
rlabel metal2 s 62210 12200 62266 13000 4 la_data_out_core[44]
port 326 nsew
rlabel metal2 s 62578 12200 62634 13000 4 la_data_out_core[45]
port 327 nsew
rlabel metal2 s 62946 12200 63002 13000 4 la_data_out_core[46]
port 328 nsew
rlabel metal2 s 63314 12200 63370 13000 4 la_data_out_core[47]
port 329 nsew
rlabel metal2 s 63682 12200 63738 13000 4 la_data_out_core[48]
port 330 nsew
rlabel metal2 s 50986 0 51042 800 4 la_data_out_core[49]
port 331 nsew
rlabel metal2 s 64050 12200 64106 13000 4 la_data_out_core[4]
port 332 nsew
rlabel metal2 s 51354 0 51410 800 4 la_data_out_core[50]
port 333 nsew
rlabel metal2 s 64418 12200 64474 13000 4 la_data_out_core[51]
port 334 nsew
rlabel metal2 s 51722 0 51778 800 4 la_data_out_core[52]
port 335 nsew
rlabel metal2 s 64786 12200 64842 13000 4 la_data_out_core[53]
port 336 nsew
rlabel metal2 s 52090 0 52146 800 4 la_data_out_core[54]
port 337 nsew
rlabel metal2 s 65154 12200 65210 13000 4 la_data_out_core[55]
port 338 nsew
rlabel metal2 s 52458 0 52514 800 4 la_data_out_core[56]
port 339 nsew
rlabel metal2 s 65522 12200 65578 13000 4 la_data_out_core[57]
port 340 nsew
rlabel metal2 s 52826 0 52882 800 4 la_data_out_core[58]
port 341 nsew
rlabel metal2 s 65890 12200 65946 13000 4 la_data_out_core[59]
port 342 nsew
rlabel metal2 s 53194 0 53250 800 4 la_data_out_core[5]
port 343 nsew
rlabel metal2 s 66258 12200 66314 13000 4 la_data_out_core[60]
port 344 nsew
rlabel metal2 s 53562 0 53618 800 4 la_data_out_core[61]
port 345 nsew
rlabel metal2 s 66626 12200 66682 13000 4 la_data_out_core[62]
port 346 nsew
rlabel metal2 s 53930 0 53986 800 4 la_data_out_core[63]
port 347 nsew
rlabel metal2 s 66994 12200 67050 13000 4 la_data_out_core[64]
port 348 nsew
rlabel metal2 s 54298 0 54354 800 4 la_data_out_core[65]
port 349 nsew
rlabel metal2 s 67362 12200 67418 13000 4 la_data_out_core[66]
port 350 nsew
rlabel metal2 s 54666 0 54722 800 4 la_data_out_core[67]
port 351 nsew
rlabel metal2 s 67730 12200 67786 13000 4 la_data_out_core[68]
port 352 nsew
rlabel metal2 s 55034 0 55090 800 4 la_data_out_core[69]
port 353 nsew
rlabel metal2 s 68098 12200 68154 13000 4 la_data_out_core[6]
port 354 nsew
rlabel metal2 s 55402 0 55458 800 4 la_data_out_core[70]
port 355 nsew
rlabel metal2 s 68466 12200 68522 13000 4 la_data_out_core[71]
port 356 nsew
rlabel metal2 s 55770 0 55826 800 4 la_data_out_core[72]
port 357 nsew
rlabel metal2 s 68834 12200 68890 13000 4 la_data_out_core[73]
port 358 nsew
rlabel metal2 s 56138 0 56194 800 4 la_data_out_core[74]
port 359 nsew
rlabel metal2 s 69202 12200 69258 13000 4 la_data_out_core[75]
port 360 nsew
rlabel metal2 s 56506 0 56562 800 4 la_data_out_core[76]
port 361 nsew
rlabel metal2 s 69570 12200 69626 13000 4 la_data_out_core[77]
port 362 nsew
rlabel metal2 s 56874 0 56930 800 4 la_data_out_core[78]
port 363 nsew
rlabel metal2 s 69938 12200 69994 13000 4 la_data_out_core[79]
port 364 nsew
rlabel metal2 s 57242 0 57298 800 4 la_data_out_core[7]
port 365 nsew
rlabel metal2 s 70306 12200 70362 13000 4 la_data_out_core[80]
port 366 nsew
rlabel metal2 s 57610 0 57666 800 4 la_data_out_core[81]
port 367 nsew
rlabel metal2 s 70674 12200 70730 13000 4 la_data_out_core[82]
port 368 nsew
rlabel metal2 s 57978 0 58034 800 4 la_data_out_core[83]
port 369 nsew
rlabel metal2 s 71042 12200 71098 13000 4 la_data_out_core[84]
port 370 nsew
rlabel metal2 s 58346 0 58402 800 4 la_data_out_core[85]
port 371 nsew
rlabel metal2 s 71410 12200 71466 13000 4 la_data_out_core[86]
port 372 nsew
rlabel metal2 s 58714 0 58770 800 4 la_data_out_core[87]
port 373 nsew
rlabel metal2 s 71778 12200 71834 13000 4 la_data_out_core[88]
port 374 nsew
rlabel metal2 s 59082 0 59138 800 4 la_data_out_core[89]
port 375 nsew
rlabel metal2 s 72146 12200 72202 13000 4 la_data_out_core[8]
port 376 nsew
rlabel metal2 s 59450 0 59506 800 4 la_data_out_core[90]
port 377 nsew
rlabel metal2 s 72514 12200 72570 13000 4 la_data_out_core[91]
port 378 nsew
rlabel metal2 s 59818 0 59874 800 4 la_data_out_core[92]
port 379 nsew
rlabel metal2 s 72882 12200 72938 13000 4 la_data_out_core[93]
port 380 nsew
rlabel metal2 s 60186 0 60242 800 4 la_data_out_core[94]
port 381 nsew
rlabel metal2 s 73250 12200 73306 13000 4 la_data_out_core[95]
port 382 nsew
rlabel metal2 s 60554 0 60610 800 4 la_data_out_core[96]
port 383 nsew
rlabel metal2 s 73618 12200 73674 13000 4 la_data_out_core[97]
port 384 nsew
rlabel metal2 s 60922 0 60978 800 4 la_data_out_core[98]
port 385 nsew
rlabel metal2 s 73986 12200 74042 13000 4 la_data_out_core[99]
port 386 nsew
rlabel metal2 s 61290 0 61346 800 4 la_data_out_core[9]
port 387 nsew
rlabel metal2 s 61658 0 61714 800 4 la_data_out_mprj[0]
port 388 nsew
rlabel metal2 s 62026 0 62082 800 4 la_data_out_mprj[100]
port 389 nsew
rlabel metal2 s 62394 0 62450 800 4 la_data_out_mprj[101]
port 390 nsew
rlabel metal2 s 62762 0 62818 800 4 la_data_out_mprj[102]
port 391 nsew
rlabel metal2 s 63130 0 63186 800 4 la_data_out_mprj[103]
port 392 nsew
rlabel metal2 s 63498 0 63554 800 4 la_data_out_mprj[104]
port 393 nsew
rlabel metal2 s 63866 0 63922 800 4 la_data_out_mprj[105]
port 394 nsew
rlabel metal2 s 64234 0 64290 800 4 la_data_out_mprj[106]
port 395 nsew
rlabel metal2 s 64602 0 64658 800 4 la_data_out_mprj[107]
port 396 nsew
rlabel metal2 s 64970 0 65026 800 4 la_data_out_mprj[108]
port 397 nsew
rlabel metal2 s 65338 0 65394 800 4 la_data_out_mprj[109]
port 398 nsew
rlabel metal2 s 65706 0 65762 800 4 la_data_out_mprj[10]
port 399 nsew
rlabel metal2 s 66074 0 66130 800 4 la_data_out_mprj[110]
port 400 nsew
rlabel metal2 s 66442 0 66498 800 4 la_data_out_mprj[111]
port 401 nsew
rlabel metal2 s 66810 0 66866 800 4 la_data_out_mprj[112]
port 402 nsew
rlabel metal2 s 67178 0 67234 800 4 la_data_out_mprj[113]
port 403 nsew
rlabel metal2 s 67546 0 67602 800 4 la_data_out_mprj[114]
port 404 nsew
rlabel metal2 s 67914 0 67970 800 4 la_data_out_mprj[115]
port 405 nsew
rlabel metal2 s 68282 0 68338 800 4 la_data_out_mprj[116]
port 406 nsew
rlabel metal2 s 68650 0 68706 800 4 la_data_out_mprj[117]
port 407 nsew
rlabel metal2 s 69018 0 69074 800 4 la_data_out_mprj[118]
port 408 nsew
rlabel metal2 s 69386 0 69442 800 4 la_data_out_mprj[119]
port 409 nsew
rlabel metal2 s 69754 0 69810 800 4 la_data_out_mprj[11]
port 410 nsew
rlabel metal2 s 70122 0 70178 800 4 la_data_out_mprj[120]
port 411 nsew
rlabel metal2 s 70490 0 70546 800 4 la_data_out_mprj[121]
port 412 nsew
rlabel metal2 s 70858 0 70914 800 4 la_data_out_mprj[122]
port 413 nsew
rlabel metal2 s 71226 0 71282 800 4 la_data_out_mprj[123]
port 414 nsew
rlabel metal2 s 71594 0 71650 800 4 la_data_out_mprj[124]
port 415 nsew
rlabel metal2 s 71962 0 72018 800 4 la_data_out_mprj[125]
port 416 nsew
rlabel metal2 s 72330 0 72386 800 4 la_data_out_mprj[126]
port 417 nsew
rlabel metal2 s 72698 0 72754 800 4 la_data_out_mprj[127]
port 418 nsew
rlabel metal2 s 73066 0 73122 800 4 la_data_out_mprj[12]
port 419 nsew
rlabel metal2 s 73434 0 73490 800 4 la_data_out_mprj[13]
port 420 nsew
rlabel metal2 s 73802 0 73858 800 4 la_data_out_mprj[14]
port 421 nsew
rlabel metal2 s 74170 0 74226 800 4 la_data_out_mprj[15]
port 422 nsew
rlabel metal2 s 74538 0 74594 800 4 la_data_out_mprj[16]
port 423 nsew
rlabel metal2 s 74906 0 74962 800 4 la_data_out_mprj[17]
port 424 nsew
rlabel metal2 s 75274 0 75330 800 4 la_data_out_mprj[18]
port 425 nsew
rlabel metal2 s 75642 0 75698 800 4 la_data_out_mprj[19]
port 426 nsew
rlabel metal2 s 76010 0 76066 800 4 la_data_out_mprj[1]
port 427 nsew
rlabel metal2 s 76378 0 76434 800 4 la_data_out_mprj[20]
port 428 nsew
rlabel metal2 s 76746 0 76802 800 4 la_data_out_mprj[21]
port 429 nsew
rlabel metal2 s 77114 0 77170 800 4 la_data_out_mprj[22]
port 430 nsew
rlabel metal2 s 77482 0 77538 800 4 la_data_out_mprj[23]
port 431 nsew
rlabel metal2 s 77850 0 77906 800 4 la_data_out_mprj[24]
port 432 nsew
rlabel metal2 s 78218 0 78274 800 4 la_data_out_mprj[25]
port 433 nsew
rlabel metal2 s 78586 0 78642 800 4 la_data_out_mprj[26]
port 434 nsew
rlabel metal2 s 78954 0 79010 800 4 la_data_out_mprj[27]
port 435 nsew
rlabel metal2 s 79322 0 79378 800 4 la_data_out_mprj[28]
port 436 nsew
rlabel metal2 s 79690 0 79746 800 4 la_data_out_mprj[29]
port 437 nsew
rlabel metal2 s 80058 0 80114 800 4 la_data_out_mprj[2]
port 438 nsew
rlabel metal2 s 80426 0 80482 800 4 la_data_out_mprj[30]
port 439 nsew
rlabel metal2 s 80794 0 80850 800 4 la_data_out_mprj[31]
port 440 nsew
rlabel metal2 s 81162 0 81218 800 4 la_data_out_mprj[32]
port 441 nsew
rlabel metal2 s 81530 0 81586 800 4 la_data_out_mprj[33]
port 442 nsew
rlabel metal2 s 81898 0 81954 800 4 la_data_out_mprj[34]
port 443 nsew
rlabel metal2 s 82266 0 82322 800 4 la_data_out_mprj[35]
port 444 nsew
rlabel metal2 s 82634 0 82690 800 4 la_data_out_mprj[36]
port 445 nsew
rlabel metal2 s 83002 0 83058 800 4 la_data_out_mprj[37]
port 446 nsew
rlabel metal2 s 83370 0 83426 800 4 la_data_out_mprj[38]
port 447 nsew
rlabel metal2 s 83738 0 83794 800 4 la_data_out_mprj[39]
port 448 nsew
rlabel metal2 s 84106 0 84162 800 4 la_data_out_mprj[3]
port 449 nsew
rlabel metal2 s 84474 0 84530 800 4 la_data_out_mprj[40]
port 450 nsew
rlabel metal2 s 84842 0 84898 800 4 la_data_out_mprj[41]
port 451 nsew
rlabel metal2 s 85210 0 85266 800 4 la_data_out_mprj[42]
port 452 nsew
rlabel metal2 s 85578 0 85634 800 4 la_data_out_mprj[43]
port 453 nsew
rlabel metal2 s 85946 0 86002 800 4 la_data_out_mprj[44]
port 454 nsew
rlabel metal2 s 86314 0 86370 800 4 la_data_out_mprj[45]
port 455 nsew
rlabel metal2 s 86682 0 86738 800 4 la_data_out_mprj[46]
port 456 nsew
rlabel metal2 s 87050 0 87106 800 4 la_data_out_mprj[47]
port 457 nsew
rlabel metal2 s 74354 12200 74410 13000 4 la_data_out_mprj[48]
port 458 nsew
rlabel metal2 s 87418 0 87474 800 4 la_data_out_mprj[49]
port 459 nsew
rlabel metal2 s 74722 12200 74778 13000 4 la_data_out_mprj[4]
port 460 nsew
rlabel metal2 s 87786 0 87842 800 4 la_data_out_mprj[50]
port 461 nsew
rlabel metal2 s 75090 12200 75146 13000 4 la_data_out_mprj[51]
port 462 nsew
rlabel metal2 s 88154 0 88210 800 4 la_data_out_mprj[52]
port 463 nsew
rlabel metal2 s 75458 12200 75514 13000 4 la_data_out_mprj[53]
port 464 nsew
rlabel metal2 s 88522 0 88578 800 4 la_data_out_mprj[54]
port 465 nsew
rlabel metal2 s 75826 12200 75882 13000 4 la_data_out_mprj[55]
port 466 nsew
rlabel metal2 s 88890 0 88946 800 4 la_data_out_mprj[56]
port 467 nsew
rlabel metal2 s 76194 12200 76250 13000 4 la_data_out_mprj[57]
port 468 nsew
rlabel metal2 s 89258 0 89314 800 4 la_data_out_mprj[58]
port 469 nsew
rlabel metal2 s 76562 12200 76618 13000 4 la_data_out_mprj[59]
port 470 nsew
rlabel metal2 s 89626 0 89682 800 4 la_data_out_mprj[5]
port 471 nsew
rlabel metal2 s 76930 12200 76986 13000 4 la_data_out_mprj[60]
port 472 nsew
rlabel metal2 s 89994 0 90050 800 4 la_data_out_mprj[61]
port 473 nsew
rlabel metal2 s 77298 12200 77354 13000 4 la_data_out_mprj[62]
port 474 nsew
rlabel metal2 s 90362 0 90418 800 4 la_data_out_mprj[63]
port 475 nsew
rlabel metal2 s 77666 12200 77722 13000 4 la_data_out_mprj[64]
port 476 nsew
rlabel metal2 s 90730 0 90786 800 4 la_data_out_mprj[65]
port 477 nsew
rlabel metal2 s 78034 12200 78090 13000 4 la_data_out_mprj[66]
port 478 nsew
rlabel metal2 s 91098 0 91154 800 4 la_data_out_mprj[67]
port 479 nsew
rlabel metal2 s 78402 12200 78458 13000 4 la_data_out_mprj[68]
port 480 nsew
rlabel metal2 s 91466 0 91522 800 4 la_data_out_mprj[69]
port 481 nsew
rlabel metal2 s 78770 12200 78826 13000 4 la_data_out_mprj[6]
port 482 nsew
rlabel metal2 s 91834 0 91890 800 4 la_data_out_mprj[70]
port 483 nsew
rlabel metal2 s 79138 12200 79194 13000 4 la_data_out_mprj[71]
port 484 nsew
rlabel metal2 s 92202 0 92258 800 4 la_data_out_mprj[72]
port 485 nsew
rlabel metal2 s 79506 12200 79562 13000 4 la_data_out_mprj[73]
port 486 nsew
rlabel metal2 s 92570 0 92626 800 4 la_data_out_mprj[74]
port 487 nsew
rlabel metal2 s 79874 12200 79930 13000 4 la_data_out_mprj[75]
port 488 nsew
rlabel metal2 s 92938 0 92994 800 4 la_data_out_mprj[76]
port 489 nsew
rlabel metal2 s 80242 12200 80298 13000 4 la_data_out_mprj[77]
port 490 nsew
rlabel metal2 s 93306 0 93362 800 4 la_data_out_mprj[78]
port 491 nsew
rlabel metal2 s 80610 12200 80666 13000 4 la_data_out_mprj[79]
port 492 nsew
rlabel metal2 s 93674 0 93730 800 4 la_data_out_mprj[7]
port 493 nsew
rlabel metal2 s 80978 12200 81034 13000 4 la_data_out_mprj[80]
port 494 nsew
rlabel metal2 s 94042 0 94098 800 4 la_data_out_mprj[81]
port 495 nsew
rlabel metal2 s 81346 12200 81402 13000 4 la_data_out_mprj[82]
port 496 nsew
rlabel metal2 s 94410 0 94466 800 4 la_data_out_mprj[83]
port 497 nsew
rlabel metal2 s 81714 12200 81770 13000 4 la_data_out_mprj[84]
port 498 nsew
rlabel metal2 s 94778 0 94834 800 4 la_data_out_mprj[85]
port 499 nsew
rlabel metal2 s 82082 12200 82138 13000 4 la_data_out_mprj[86]
port 500 nsew
rlabel metal2 s 95146 0 95202 800 4 la_data_out_mprj[87]
port 501 nsew
rlabel metal2 s 82450 12200 82506 13000 4 la_data_out_mprj[88]
port 502 nsew
rlabel metal2 s 95514 0 95570 800 4 la_data_out_mprj[89]
port 503 nsew
rlabel metal2 s 82818 12200 82874 13000 4 la_data_out_mprj[8]
port 504 nsew
rlabel metal2 s 95882 0 95938 800 4 la_data_out_mprj[90]
port 505 nsew
rlabel metal2 s 83186 12200 83242 13000 4 la_data_out_mprj[91]
port 506 nsew
rlabel metal2 s 96250 0 96306 800 4 la_data_out_mprj[92]
port 507 nsew
rlabel metal2 s 83554 12200 83610 13000 4 la_data_out_mprj[93]
port 508 nsew
rlabel metal2 s 96618 0 96674 800 4 la_data_out_mprj[94]
port 509 nsew
rlabel metal2 s 83922 12200 83978 13000 4 la_data_out_mprj[95]
port 510 nsew
rlabel metal2 s 96986 0 97042 800 4 la_data_out_mprj[96]
port 511 nsew
rlabel metal2 s 84290 12200 84346 13000 4 la_data_out_mprj[97]
port 512 nsew
rlabel metal2 s 97354 0 97410 800 4 la_data_out_mprj[98]
port 513 nsew
rlabel metal2 s 84658 12200 84714 13000 4 la_data_out_mprj[99]
port 514 nsew
rlabel metal2 s 97722 0 97778 800 4 la_data_out_mprj[9]
port 515 nsew
rlabel metal2 s 85026 12200 85082 13000 4 la_oen_core[0]
port 516 nsew
rlabel metal2 s 85394 12200 85450 13000 4 la_oen_core[100]
port 517 nsew
rlabel metal2 s 85762 12200 85818 13000 4 la_oen_core[101]
port 518 nsew
rlabel metal2 s 86130 12200 86186 13000 4 la_oen_core[102]
port 519 nsew
rlabel metal2 s 86498 12200 86554 13000 4 la_oen_core[103]
port 520 nsew
rlabel metal2 s 86866 12200 86922 13000 4 la_oen_core[104]
port 521 nsew
rlabel metal2 s 87234 12200 87290 13000 4 la_oen_core[105]
port 522 nsew
rlabel metal2 s 87602 12200 87658 13000 4 la_oen_core[106]
port 523 nsew
rlabel metal2 s 87970 12200 88026 13000 4 la_oen_core[107]
port 524 nsew
rlabel metal2 s 88338 12200 88394 13000 4 la_oen_core[108]
port 525 nsew
rlabel metal2 s 88706 12200 88762 13000 4 la_oen_core[109]
port 526 nsew
rlabel metal2 s 89074 12200 89130 13000 4 la_oen_core[10]
port 527 nsew
rlabel metal2 s 89442 12200 89498 13000 4 la_oen_core[110]
port 528 nsew
rlabel metal2 s 89810 12200 89866 13000 4 la_oen_core[111]
port 529 nsew
rlabel metal2 s 90178 12200 90234 13000 4 la_oen_core[112]
port 530 nsew
rlabel metal2 s 90546 12200 90602 13000 4 la_oen_core[113]
port 531 nsew
rlabel metal2 s 90914 12200 90970 13000 4 la_oen_core[114]
port 532 nsew
rlabel metal2 s 91282 12200 91338 13000 4 la_oen_core[115]
port 533 nsew
rlabel metal2 s 91650 12200 91706 13000 4 la_oen_core[116]
port 534 nsew
rlabel metal2 s 92018 12200 92074 13000 4 la_oen_core[117]
port 535 nsew
rlabel metal2 s 92386 12200 92442 13000 4 la_oen_core[118]
port 536 nsew
rlabel metal2 s 92754 12200 92810 13000 4 la_oen_core[119]
port 537 nsew
rlabel metal2 s 93122 12200 93178 13000 4 la_oen_core[11]
port 538 nsew
rlabel metal2 s 93490 12200 93546 13000 4 la_oen_core[120]
port 539 nsew
rlabel metal2 s 93858 12200 93914 13000 4 la_oen_core[121]
port 540 nsew
rlabel metal2 s 94226 12200 94282 13000 4 la_oen_core[122]
port 541 nsew
rlabel metal2 s 94594 12200 94650 13000 4 la_oen_core[123]
port 542 nsew
rlabel metal2 s 94962 12200 95018 13000 4 la_oen_core[124]
port 543 nsew
rlabel metal2 s 95330 12200 95386 13000 4 la_oen_core[125]
port 544 nsew
rlabel metal2 s 95698 12200 95754 13000 4 la_oen_core[126]
port 545 nsew
rlabel metal2 s 96066 12200 96122 13000 4 la_oen_core[127]
port 546 nsew
rlabel metal2 s 96434 12200 96490 13000 4 la_oen_core[12]
port 547 nsew
rlabel metal2 s 96802 12200 96858 13000 4 la_oen_core[13]
port 548 nsew
rlabel metal2 s 97170 12200 97226 13000 4 la_oen_core[14]
port 549 nsew
rlabel metal2 s 97538 12200 97594 13000 4 la_oen_core[15]
port 550 nsew
rlabel metal2 s 97906 12200 97962 13000 4 la_oen_core[16]
port 551 nsew
rlabel metal2 s 98274 12200 98330 13000 4 la_oen_core[17]
port 552 nsew
rlabel metal2 s 98642 12200 98698 13000 4 la_oen_core[18]
port 553 nsew
rlabel metal2 s 99010 12200 99066 13000 4 la_oen_core[19]
port 554 nsew
rlabel metal2 s 99378 12200 99434 13000 4 la_oen_core[1]
port 555 nsew
rlabel metal2 s 99746 12200 99802 13000 4 la_oen_core[20]
port 556 nsew
rlabel metal2 s 100114 12200 100170 13000 4 la_oen_core[21]
port 557 nsew
rlabel metal2 s 100482 12200 100538 13000 4 la_oen_core[22]
port 558 nsew
rlabel metal2 s 100850 12200 100906 13000 4 la_oen_core[23]
port 559 nsew
rlabel metal2 s 101218 12200 101274 13000 4 la_oen_core[24]
port 560 nsew
rlabel metal2 s 101586 12200 101642 13000 4 la_oen_core[25]
port 561 nsew
rlabel metal2 s 101954 12200 102010 13000 4 la_oen_core[26]
port 562 nsew
rlabel metal2 s 102322 12200 102378 13000 4 la_oen_core[27]
port 563 nsew
rlabel metal2 s 102690 12200 102746 13000 4 la_oen_core[28]
port 564 nsew
rlabel metal2 s 103058 12200 103114 13000 4 la_oen_core[29]
port 565 nsew
rlabel metal2 s 103426 12200 103482 13000 4 la_oen_core[2]
port 566 nsew
rlabel metal2 s 103794 12200 103850 13000 4 la_oen_core[30]
port 567 nsew
rlabel metal2 s 104162 12200 104218 13000 4 la_oen_core[31]
port 568 nsew
rlabel metal2 s 104530 12200 104586 13000 4 la_oen_core[32]
port 569 nsew
rlabel metal2 s 104898 12200 104954 13000 4 la_oen_core[33]
port 570 nsew
rlabel metal2 s 105266 12200 105322 13000 4 la_oen_core[34]
port 571 nsew
rlabel metal2 s 105634 12200 105690 13000 4 la_oen_core[35]
port 572 nsew
rlabel metal2 s 106002 12200 106058 13000 4 la_oen_core[36]
port 573 nsew
rlabel metal2 s 106370 12200 106426 13000 4 la_oen_core[37]
port 574 nsew
rlabel metal2 s 106738 12200 106794 13000 4 la_oen_core[38]
port 575 nsew
rlabel metal2 s 107106 12200 107162 13000 4 la_oen_core[39]
port 576 nsew
rlabel metal2 s 107474 12200 107530 13000 4 la_oen_core[3]
port 577 nsew
rlabel metal2 s 107842 12200 107898 13000 4 la_oen_core[40]
port 578 nsew
rlabel metal2 s 108210 12200 108266 13000 4 la_oen_core[41]
port 579 nsew
rlabel metal2 s 108578 12200 108634 13000 4 la_oen_core[42]
port 580 nsew
rlabel metal2 s 108946 12200 109002 13000 4 la_oen_core[43]
port 581 nsew
rlabel metal2 s 109314 12200 109370 13000 4 la_oen_core[44]
port 582 nsew
rlabel metal2 s 109682 12200 109738 13000 4 la_oen_core[45]
port 583 nsew
rlabel metal2 s 110050 12200 110106 13000 4 la_oen_core[46]
port 584 nsew
rlabel metal2 s 110418 12200 110474 13000 4 la_oen_core[47]
port 585 nsew
rlabel metal2 s 110786 12200 110842 13000 4 la_oen_core[48]
port 586 nsew
rlabel metal2 s 98090 0 98146 800 4 la_oen_core[49]
port 587 nsew
rlabel metal2 s 111154 12200 111210 13000 4 la_oen_core[4]
port 588 nsew
rlabel metal2 s 98458 0 98514 800 4 la_oen_core[50]
port 589 nsew
rlabel metal2 s 111522 12200 111578 13000 4 la_oen_core[51]
port 590 nsew
rlabel metal2 s 98826 0 98882 800 4 la_oen_core[52]
port 591 nsew
rlabel metal2 s 111890 12200 111946 13000 4 la_oen_core[53]
port 592 nsew
rlabel metal2 s 99194 0 99250 800 4 la_oen_core[54]
port 593 nsew
rlabel metal2 s 112258 12200 112314 13000 4 la_oen_core[55]
port 594 nsew
rlabel metal2 s 99562 0 99618 800 4 la_oen_core[56]
port 595 nsew
rlabel metal2 s 112626 12200 112682 13000 4 la_oen_core[57]
port 596 nsew
rlabel metal2 s 99930 0 99986 800 4 la_oen_core[58]
port 597 nsew
rlabel metal2 s 112994 12200 113050 13000 4 la_oen_core[59]
port 598 nsew
rlabel metal2 s 100298 0 100354 800 4 la_oen_core[5]
port 599 nsew
rlabel metal2 s 113362 12200 113418 13000 4 la_oen_core[60]
port 600 nsew
rlabel metal2 s 100666 0 100722 800 4 la_oen_core[61]
port 601 nsew
rlabel metal2 s 113730 12200 113786 13000 4 la_oen_core[62]
port 602 nsew
rlabel metal2 s 101034 0 101090 800 4 la_oen_core[63]
port 603 nsew
rlabel metal2 s 114098 12200 114154 13000 4 la_oen_core[64]
port 604 nsew
rlabel metal2 s 101402 0 101458 800 4 la_oen_core[65]
port 605 nsew
rlabel metal2 s 114466 12200 114522 13000 4 la_oen_core[66]
port 606 nsew
rlabel metal2 s 101770 0 101826 800 4 la_oen_core[67]
port 607 nsew
rlabel metal2 s 114834 12200 114890 13000 4 la_oen_core[68]
port 608 nsew
rlabel metal2 s 102138 0 102194 800 4 la_oen_core[69]
port 609 nsew
rlabel metal2 s 115202 12200 115258 13000 4 la_oen_core[6]
port 610 nsew
rlabel metal2 s 102506 0 102562 800 4 la_oen_core[70]
port 611 nsew
rlabel metal2 s 115570 12200 115626 13000 4 la_oen_core[71]
port 612 nsew
rlabel metal2 s 102874 0 102930 800 4 la_oen_core[72]
port 613 nsew
rlabel metal2 s 115938 12200 115994 13000 4 la_oen_core[73]
port 614 nsew
rlabel metal2 s 103242 0 103298 800 4 la_oen_core[74]
port 615 nsew
rlabel metal2 s 116306 12200 116362 13000 4 la_oen_core[75]
port 616 nsew
rlabel metal2 s 103610 0 103666 800 4 la_oen_core[76]
port 617 nsew
rlabel metal2 s 116674 12200 116730 13000 4 la_oen_core[77]
port 618 nsew
rlabel metal2 s 103978 0 104034 800 4 la_oen_core[78]
port 619 nsew
rlabel metal2 s 117042 12200 117098 13000 4 la_oen_core[79]
port 620 nsew
rlabel metal2 s 104346 0 104402 800 4 la_oen_core[7]
port 621 nsew
rlabel metal2 s 117410 12200 117466 13000 4 la_oen_core[80]
port 622 nsew
rlabel metal2 s 104714 0 104770 800 4 la_oen_core[81]
port 623 nsew
rlabel metal2 s 117778 12200 117834 13000 4 la_oen_core[82]
port 624 nsew
rlabel metal2 s 105082 0 105138 800 4 la_oen_core[83]
port 625 nsew
rlabel metal2 s 118146 12200 118202 13000 4 la_oen_core[84]
port 626 nsew
rlabel metal2 s 105450 0 105506 800 4 la_oen_core[85]
port 627 nsew
rlabel metal2 s 118514 12200 118570 13000 4 la_oen_core[86]
port 628 nsew
rlabel metal2 s 105818 0 105874 800 4 la_oen_core[87]
port 629 nsew
rlabel metal2 s 118882 12200 118938 13000 4 la_oen_core[88]
port 630 nsew
rlabel metal2 s 106186 0 106242 800 4 la_oen_core[89]
port 631 nsew
rlabel metal2 s 119250 12200 119306 13000 4 la_oen_core[8]
port 632 nsew
rlabel metal2 s 106554 0 106610 800 4 la_oen_core[90]
port 633 nsew
rlabel metal2 s 119618 12200 119674 13000 4 la_oen_core[91]
port 634 nsew
rlabel metal2 s 106922 0 106978 800 4 la_oen_core[92]
port 635 nsew
rlabel metal2 s 119986 12200 120042 13000 4 la_oen_core[93]
port 636 nsew
rlabel metal2 s 107290 0 107346 800 4 la_oen_core[94]
port 637 nsew
rlabel metal2 s 120354 12200 120410 13000 4 la_oen_core[95]
port 638 nsew
rlabel metal2 s 107658 0 107714 800 4 la_oen_core[96]
port 639 nsew
rlabel metal2 s 120722 12200 120778 13000 4 la_oen_core[97]
port 640 nsew
rlabel metal2 s 108026 0 108082 800 4 la_oen_core[98]
port 641 nsew
rlabel metal2 s 121090 12200 121146 13000 4 la_oen_core[99]
port 642 nsew
rlabel metal2 s 108394 0 108450 800 4 la_oen_core[9]
port 643 nsew
rlabel metal2 s 108762 0 108818 800 4 la_oen_mprj[0]
port 644 nsew
rlabel metal2 s 109130 0 109186 800 4 la_oen_mprj[100]
port 645 nsew
rlabel metal2 s 109498 0 109554 800 4 la_oen_mprj[101]
port 646 nsew
rlabel metal2 s 109866 0 109922 800 4 la_oen_mprj[102]
port 647 nsew
rlabel metal2 s 110234 0 110290 800 4 la_oen_mprj[103]
port 648 nsew
rlabel metal2 s 110602 0 110658 800 4 la_oen_mprj[104]
port 649 nsew
rlabel metal2 s 110970 0 111026 800 4 la_oen_mprj[105]
port 650 nsew
rlabel metal2 s 111338 0 111394 800 4 la_oen_mprj[106]
port 651 nsew
rlabel metal2 s 111706 0 111762 800 4 la_oen_mprj[107]
port 652 nsew
rlabel metal2 s 112074 0 112130 800 4 la_oen_mprj[108]
port 653 nsew
rlabel metal2 s 112442 0 112498 800 4 la_oen_mprj[109]
port 654 nsew
rlabel metal2 s 112810 0 112866 800 4 la_oen_mprj[10]
port 655 nsew
rlabel metal2 s 113178 0 113234 800 4 la_oen_mprj[110]
port 656 nsew
rlabel metal2 s 113546 0 113602 800 4 la_oen_mprj[111]
port 657 nsew
rlabel metal2 s 113914 0 113970 800 4 la_oen_mprj[112]
port 658 nsew
rlabel metal2 s 114282 0 114338 800 4 la_oen_mprj[113]
port 659 nsew
rlabel metal2 s 114650 0 114706 800 4 la_oen_mprj[114]
port 660 nsew
rlabel metal2 s 115018 0 115074 800 4 la_oen_mprj[115]
port 661 nsew
rlabel metal2 s 115386 0 115442 800 4 la_oen_mprj[116]
port 662 nsew
rlabel metal2 s 115754 0 115810 800 4 la_oen_mprj[117]
port 663 nsew
rlabel metal2 s 116122 0 116178 800 4 la_oen_mprj[118]
port 664 nsew
rlabel metal2 s 116490 0 116546 800 4 la_oen_mprj[119]
port 665 nsew
rlabel metal2 s 116858 0 116914 800 4 la_oen_mprj[11]
port 666 nsew
rlabel metal2 s 117226 0 117282 800 4 la_oen_mprj[120]
port 667 nsew
rlabel metal2 s 117594 0 117650 800 4 la_oen_mprj[121]
port 668 nsew
rlabel metal2 s 117962 0 118018 800 4 la_oen_mprj[122]
port 669 nsew
rlabel metal2 s 118330 0 118386 800 4 la_oen_mprj[123]
port 670 nsew
rlabel metal2 s 118698 0 118754 800 4 la_oen_mprj[124]
port 671 nsew
rlabel metal2 s 119066 0 119122 800 4 la_oen_mprj[125]
port 672 nsew
rlabel metal2 s 119434 0 119490 800 4 la_oen_mprj[126]
port 673 nsew
rlabel metal2 s 119802 0 119858 800 4 la_oen_mprj[127]
port 674 nsew
rlabel metal2 s 120170 0 120226 800 4 la_oen_mprj[12]
port 675 nsew
rlabel metal2 s 120538 0 120594 800 4 la_oen_mprj[13]
port 676 nsew
rlabel metal2 s 120906 0 120962 800 4 la_oen_mprj[14]
port 677 nsew
rlabel metal2 s 121274 0 121330 800 4 la_oen_mprj[15]
port 678 nsew
rlabel metal2 s 121642 0 121698 800 4 la_oen_mprj[16]
port 679 nsew
rlabel metal2 s 122010 0 122066 800 4 la_oen_mprj[17]
port 680 nsew
rlabel metal2 s 122378 0 122434 800 4 la_oen_mprj[18]
port 681 nsew
rlabel metal2 s 122746 0 122802 800 4 la_oen_mprj[19]
port 682 nsew
rlabel metal2 s 123114 0 123170 800 4 la_oen_mprj[1]
port 683 nsew
rlabel metal2 s 123482 0 123538 800 4 la_oen_mprj[20]
port 684 nsew
rlabel metal2 s 123850 0 123906 800 4 la_oen_mprj[21]
port 685 nsew
rlabel metal2 s 124218 0 124274 800 4 la_oen_mprj[22]
port 686 nsew
rlabel metal2 s 124586 0 124642 800 4 la_oen_mprj[23]
port 687 nsew
rlabel metal2 s 124954 0 125010 800 4 la_oen_mprj[24]
port 688 nsew
rlabel metal2 s 125322 0 125378 800 4 la_oen_mprj[25]
port 689 nsew
rlabel metal2 s 125690 0 125746 800 4 la_oen_mprj[26]
port 690 nsew
rlabel metal2 s 126058 0 126114 800 4 la_oen_mprj[27]
port 691 nsew
rlabel metal2 s 126426 0 126482 800 4 la_oen_mprj[28]
port 692 nsew
rlabel metal2 s 126794 0 126850 800 4 la_oen_mprj[29]
port 693 nsew
rlabel metal2 s 127162 0 127218 800 4 la_oen_mprj[2]
port 694 nsew
rlabel metal2 s 127530 0 127586 800 4 la_oen_mprj[30]
port 695 nsew
rlabel metal2 s 127898 0 127954 800 4 la_oen_mprj[31]
port 696 nsew
rlabel metal2 s 128266 0 128322 800 4 la_oen_mprj[32]
port 697 nsew
rlabel metal2 s 128634 0 128690 800 4 la_oen_mprj[33]
port 698 nsew
rlabel metal2 s 129002 0 129058 800 4 la_oen_mprj[34]
port 699 nsew
rlabel metal2 s 129370 0 129426 800 4 la_oen_mprj[35]
port 700 nsew
rlabel metal2 s 129738 0 129794 800 4 la_oen_mprj[36]
port 701 nsew
rlabel metal2 s 130106 0 130162 800 4 la_oen_mprj[37]
port 702 nsew
rlabel metal2 s 130474 0 130530 800 4 la_oen_mprj[38]
port 703 nsew
rlabel metal2 s 130842 0 130898 800 4 la_oen_mprj[39]
port 704 nsew
rlabel metal2 s 131210 0 131266 800 4 la_oen_mprj[3]
port 705 nsew
rlabel metal2 s 131578 0 131634 800 4 la_oen_mprj[40]
port 706 nsew
rlabel metal2 s 131946 0 132002 800 4 la_oen_mprj[41]
port 707 nsew
rlabel metal2 s 132314 0 132370 800 4 la_oen_mprj[42]
port 708 nsew
rlabel metal2 s 132682 0 132738 800 4 la_oen_mprj[43]
port 709 nsew
rlabel metal2 s 133050 0 133106 800 4 la_oen_mprj[44]
port 710 nsew
rlabel metal2 s 133418 0 133474 800 4 la_oen_mprj[45]
port 711 nsew
rlabel metal2 s 133786 0 133842 800 4 la_oen_mprj[46]
port 712 nsew
rlabel metal2 s 134154 0 134210 800 4 la_oen_mprj[47]
port 713 nsew
rlabel metal2 s 121458 12200 121514 13000 4 la_oen_mprj[48]
port 714 nsew
rlabel metal2 s 134522 0 134578 800 4 la_oen_mprj[49]
port 715 nsew
rlabel metal2 s 121826 12200 121882 13000 4 la_oen_mprj[4]
port 716 nsew
rlabel metal2 s 134890 0 134946 800 4 la_oen_mprj[50]
port 717 nsew
rlabel metal2 s 122194 12200 122250 13000 4 la_oen_mprj[51]
port 718 nsew
rlabel metal2 s 135258 0 135314 800 4 la_oen_mprj[52]
port 719 nsew
rlabel metal2 s 122562 12200 122618 13000 4 la_oen_mprj[53]
port 720 nsew
rlabel metal2 s 135626 0 135682 800 4 la_oen_mprj[54]
port 721 nsew
rlabel metal2 s 122930 12200 122986 13000 4 la_oen_mprj[55]
port 722 nsew
rlabel metal2 s 135994 0 136050 800 4 la_oen_mprj[56]
port 723 nsew
rlabel metal2 s 123298 12200 123354 13000 4 la_oen_mprj[57]
port 724 nsew
rlabel metal2 s 136362 0 136418 800 4 la_oen_mprj[58]
port 725 nsew
rlabel metal2 s 123666 12200 123722 13000 4 la_oen_mprj[59]
port 726 nsew
rlabel metal2 s 136730 0 136786 800 4 la_oen_mprj[5]
port 727 nsew
rlabel metal2 s 124034 12200 124090 13000 4 la_oen_mprj[60]
port 728 nsew
rlabel metal2 s 137098 0 137154 800 4 la_oen_mprj[61]
port 729 nsew
rlabel metal2 s 124402 12200 124458 13000 4 la_oen_mprj[62]
port 730 nsew
rlabel metal2 s 137466 0 137522 800 4 la_oen_mprj[63]
port 731 nsew
rlabel metal2 s 124770 12200 124826 13000 4 la_oen_mprj[64]
port 732 nsew
rlabel metal2 s 137834 0 137890 800 4 la_oen_mprj[65]
port 733 nsew
rlabel metal2 s 125138 12200 125194 13000 4 la_oen_mprj[66]
port 734 nsew
rlabel metal2 s 138202 0 138258 800 4 la_oen_mprj[67]
port 735 nsew
rlabel metal2 s 125506 12200 125562 13000 4 la_oen_mprj[68]
port 736 nsew
rlabel metal2 s 138570 0 138626 800 4 la_oen_mprj[69]
port 737 nsew
rlabel metal2 s 125874 12200 125930 13000 4 la_oen_mprj[6]
port 738 nsew
rlabel metal2 s 138938 0 138994 800 4 la_oen_mprj[70]
port 739 nsew
rlabel metal2 s 126242 12200 126298 13000 4 la_oen_mprj[71]
port 740 nsew
rlabel metal2 s 139306 0 139362 800 4 la_oen_mprj[72]
port 741 nsew
rlabel metal2 s 126610 12200 126666 13000 4 la_oen_mprj[73]
port 742 nsew
rlabel metal2 s 139674 0 139730 800 4 la_oen_mprj[74]
port 743 nsew
rlabel metal2 s 126978 12200 127034 13000 4 la_oen_mprj[75]
port 744 nsew
rlabel metal2 s 140042 0 140098 800 4 la_oen_mprj[76]
port 745 nsew
rlabel metal2 s 127346 12200 127402 13000 4 la_oen_mprj[77]
port 746 nsew
rlabel metal2 s 140410 0 140466 800 4 la_oen_mprj[78]
port 747 nsew
rlabel metal2 s 127714 12200 127770 13000 4 la_oen_mprj[79]
port 748 nsew
rlabel metal2 s 140778 0 140834 800 4 la_oen_mprj[7]
port 749 nsew
rlabel metal2 s 128082 12200 128138 13000 4 la_oen_mprj[80]
port 750 nsew
rlabel metal2 s 141146 0 141202 800 4 la_oen_mprj[81]
port 751 nsew
rlabel metal2 s 128450 12200 128506 13000 4 la_oen_mprj[82]
port 752 nsew
rlabel metal2 s 141514 0 141570 800 4 la_oen_mprj[83]
port 753 nsew
rlabel metal2 s 128818 12200 128874 13000 4 la_oen_mprj[84]
port 754 nsew
rlabel metal2 s 141882 0 141938 800 4 la_oen_mprj[85]
port 755 nsew
rlabel metal2 s 129186 12200 129242 13000 4 la_oen_mprj[86]
port 756 nsew
rlabel metal2 s 142250 0 142306 800 4 la_oen_mprj[87]
port 757 nsew
rlabel metal2 s 129554 12200 129610 13000 4 la_oen_mprj[88]
port 758 nsew
rlabel metal2 s 142618 0 142674 800 4 la_oen_mprj[89]
port 759 nsew
rlabel metal2 s 129922 12200 129978 13000 4 la_oen_mprj[8]
port 760 nsew
rlabel metal2 s 142986 0 143042 800 4 la_oen_mprj[90]
port 761 nsew
rlabel metal2 s 130290 12200 130346 13000 4 la_oen_mprj[91]
port 762 nsew
rlabel metal2 s 143354 0 143410 800 4 la_oen_mprj[92]
port 763 nsew
rlabel metal2 s 130658 12200 130714 13000 4 la_oen_mprj[93]
port 764 nsew
rlabel metal2 s 143722 0 143778 800 4 la_oen_mprj[94]
port 765 nsew
rlabel metal2 s 131026 12200 131082 13000 4 la_oen_mprj[95]
port 766 nsew
rlabel metal2 s 144090 0 144146 800 4 la_oen_mprj[96]
port 767 nsew
rlabel metal2 s 131394 12200 131450 13000 4 la_oen_mprj[97]
port 768 nsew
rlabel metal2 s 144458 0 144514 800 4 la_oen_mprj[98]
port 769 nsew
rlabel metal2 s 131762 12200 131818 13000 4 la_oen_mprj[99]
port 770 nsew
rlabel metal2 s 144826 0 144882 800 4 la_oen_mprj[9]
port 771 nsew
rlabel metal2 s 132130 12200 132186 13000 4 mprj_adr_o_core[0]
port 772 nsew
rlabel metal2 s 145194 0 145250 800 4 mprj_adr_o_core[10]
port 773 nsew
rlabel metal2 s 132498 12200 132554 13000 4 mprj_adr_o_core[11]
port 774 nsew
rlabel metal2 s 145562 0 145618 800 4 mprj_adr_o_core[12]
port 775 nsew
rlabel metal2 s 132866 12200 132922 13000 4 mprj_adr_o_core[13]
port 776 nsew
rlabel metal2 s 145930 0 145986 800 4 mprj_adr_o_core[14]
port 777 nsew
rlabel metal2 s 133234 12200 133290 13000 4 mprj_adr_o_core[15]
port 778 nsew
rlabel metal2 s 146298 0 146354 800 4 mprj_adr_o_core[16]
port 779 nsew
rlabel metal2 s 133602 12200 133658 13000 4 mprj_adr_o_core[17]
port 780 nsew
rlabel metal2 s 146666 0 146722 800 4 mprj_adr_o_core[18]
port 781 nsew
rlabel metal2 s 133970 12200 134026 13000 4 mprj_adr_o_core[19]
port 782 nsew
rlabel metal2 s 147034 0 147090 800 4 mprj_adr_o_core[1]
port 783 nsew
rlabel metal2 s 134338 12200 134394 13000 4 mprj_adr_o_core[20]
port 784 nsew
rlabel metal2 s 147402 0 147458 800 4 mprj_adr_o_core[21]
port 785 nsew
rlabel metal2 s 134706 12200 134762 13000 4 mprj_adr_o_core[22]
port 786 nsew
rlabel metal2 s 147770 0 147826 800 4 mprj_adr_o_core[23]
port 787 nsew
rlabel metal2 s 135074 12200 135130 13000 4 mprj_adr_o_core[24]
port 788 nsew
rlabel metal2 s 148138 0 148194 800 4 mprj_adr_o_core[25]
port 789 nsew
rlabel metal2 s 135442 12200 135498 13000 4 mprj_adr_o_core[26]
port 790 nsew
rlabel metal2 s 148506 0 148562 800 4 mprj_adr_o_core[27]
port 791 nsew
rlabel metal2 s 135810 12200 135866 13000 4 mprj_adr_o_core[28]
port 792 nsew
rlabel metal2 s 148874 0 148930 800 4 mprj_adr_o_core[29]
port 793 nsew
rlabel metal2 s 136178 12200 136234 13000 4 mprj_adr_o_core[2]
port 794 nsew
rlabel metal2 s 149242 0 149298 800 4 mprj_adr_o_core[30]
port 795 nsew
rlabel metal2 s 136546 12200 136602 13000 4 mprj_adr_o_core[31]
port 796 nsew
rlabel metal2 s 149610 0 149666 800 4 mprj_adr_o_core[3]
port 797 nsew
rlabel metal2 s 136914 12200 136970 13000 4 mprj_adr_o_core[4]
port 798 nsew
rlabel metal2 s 149978 0 150034 800 4 mprj_adr_o_core[5]
port 799 nsew
rlabel metal2 s 137282 12200 137338 13000 4 mprj_adr_o_core[6]
port 800 nsew
rlabel metal2 s 150346 0 150402 800 4 mprj_adr_o_core[7]
port 801 nsew
rlabel metal2 s 137650 12200 137706 13000 4 mprj_adr_o_core[8]
port 802 nsew
rlabel metal2 s 150714 0 150770 800 4 mprj_adr_o_core[9]
port 803 nsew
rlabel metal2 s 138018 12200 138074 13000 4 mprj_adr_o_user[0]
port 804 nsew
rlabel metal2 s 138386 12200 138442 13000 4 mprj_adr_o_user[10]
port 805 nsew
rlabel metal2 s 138754 12200 138810 13000 4 mprj_adr_o_user[11]
port 806 nsew
rlabel metal2 s 139122 12200 139178 13000 4 mprj_adr_o_user[12]
port 807 nsew
rlabel metal2 s 139490 12200 139546 13000 4 mprj_adr_o_user[13]
port 808 nsew
rlabel metal2 s 139858 12200 139914 13000 4 mprj_adr_o_user[14]
port 809 nsew
rlabel metal2 s 140226 12200 140282 13000 4 mprj_adr_o_user[15]
port 810 nsew
rlabel metal2 s 140594 12200 140650 13000 4 mprj_adr_o_user[16]
port 811 nsew
rlabel metal2 s 140962 12200 141018 13000 4 mprj_adr_o_user[17]
port 812 nsew
rlabel metal2 s 141330 12200 141386 13000 4 mprj_adr_o_user[18]
port 813 nsew
rlabel metal2 s 141698 12200 141754 13000 4 mprj_adr_o_user[19]
port 814 nsew
rlabel metal2 s 142066 12200 142122 13000 4 mprj_adr_o_user[1]
port 815 nsew
rlabel metal2 s 142434 12200 142490 13000 4 mprj_adr_o_user[20]
port 816 nsew
rlabel metal2 s 142802 12200 142858 13000 4 mprj_adr_o_user[21]
port 817 nsew
rlabel metal2 s 143170 12200 143226 13000 4 mprj_adr_o_user[22]
port 818 nsew
rlabel metal2 s 143538 12200 143594 13000 4 mprj_adr_o_user[23]
port 819 nsew
rlabel metal2 s 143906 12200 143962 13000 4 mprj_adr_o_user[24]
port 820 nsew
rlabel metal2 s 144274 12200 144330 13000 4 mprj_adr_o_user[25]
port 821 nsew
rlabel metal2 s 144642 12200 144698 13000 4 mprj_adr_o_user[26]
port 822 nsew
rlabel metal2 s 145010 12200 145066 13000 4 mprj_adr_o_user[27]
port 823 nsew
rlabel metal2 s 145378 12200 145434 13000 4 mprj_adr_o_user[28]
port 824 nsew
rlabel metal2 s 145746 12200 145802 13000 4 mprj_adr_o_user[29]
port 825 nsew
rlabel metal2 s 146114 12200 146170 13000 4 mprj_adr_o_user[2]
port 826 nsew
rlabel metal2 s 146482 12200 146538 13000 4 mprj_adr_o_user[30]
port 827 nsew
rlabel metal2 s 146850 12200 146906 13000 4 mprj_adr_o_user[31]
port 828 nsew
rlabel metal2 s 147218 12200 147274 13000 4 mprj_adr_o_user[3]
port 829 nsew
rlabel metal2 s 147586 12200 147642 13000 4 mprj_adr_o_user[4]
port 830 nsew
rlabel metal2 s 147954 12200 148010 13000 4 mprj_adr_o_user[5]
port 831 nsew
rlabel metal2 s 148322 12200 148378 13000 4 mprj_adr_o_user[6]
port 832 nsew
rlabel metal2 s 148690 12200 148746 13000 4 mprj_adr_o_user[7]
port 833 nsew
rlabel metal2 s 149058 12200 149114 13000 4 mprj_adr_o_user[8]
port 834 nsew
rlabel metal2 s 149426 12200 149482 13000 4 mprj_adr_o_user[9]
port 835 nsew
rlabel metal2 s 151082 0 151138 800 4 mprj_cyc_o_core
port 836 nsew
rlabel metal2 s 149794 12200 149850 13000 4 mprj_cyc_o_user
port 837 nsew
rlabel metal2 s 151450 0 151506 800 4 mprj_dat_o_core[0]
port 838 nsew
rlabel metal2 s 151818 0 151874 800 4 mprj_dat_o_core[10]
port 839 nsew
rlabel metal2 s 152186 0 152242 800 4 mprj_dat_o_core[11]
port 840 nsew
rlabel metal2 s 152554 0 152610 800 4 mprj_dat_o_core[12]
port 841 nsew
rlabel metal2 s 152922 0 152978 800 4 mprj_dat_o_core[13]
port 842 nsew
rlabel metal2 s 153290 0 153346 800 4 mprj_dat_o_core[14]
port 843 nsew
rlabel metal2 s 153658 0 153714 800 4 mprj_dat_o_core[15]
port 844 nsew
rlabel metal2 s 154026 0 154082 800 4 mprj_dat_o_core[16]
port 845 nsew
rlabel metal2 s 154394 0 154450 800 4 mprj_dat_o_core[17]
port 846 nsew
rlabel metal2 s 154762 0 154818 800 4 mprj_dat_o_core[18]
port 847 nsew
rlabel metal2 s 155130 0 155186 800 4 mprj_dat_o_core[19]
port 848 nsew
rlabel metal2 s 155498 0 155554 800 4 mprj_dat_o_core[1]
port 849 nsew
rlabel metal2 s 155866 0 155922 800 4 mprj_dat_o_core[20]
port 850 nsew
rlabel metal2 s 156234 0 156290 800 4 mprj_dat_o_core[21]
port 851 nsew
rlabel metal2 s 156602 0 156658 800 4 mprj_dat_o_core[22]
port 852 nsew
rlabel metal2 s 156970 0 157026 800 4 mprj_dat_o_core[23]
port 853 nsew
rlabel metal2 s 157338 0 157394 800 4 mprj_dat_o_core[24]
port 854 nsew
rlabel metal2 s 157706 0 157762 800 4 mprj_dat_o_core[25]
port 855 nsew
rlabel metal2 s 158074 0 158130 800 4 mprj_dat_o_core[26]
port 856 nsew
rlabel metal2 s 158442 0 158498 800 4 mprj_dat_o_core[27]
port 857 nsew
rlabel metal2 s 158810 0 158866 800 4 mprj_dat_o_core[28]
port 858 nsew
rlabel metal2 s 159178 0 159234 800 4 mprj_dat_o_core[29]
port 859 nsew
rlabel metal2 s 159546 0 159602 800 4 mprj_dat_o_core[2]
port 860 nsew
rlabel metal2 s 159914 0 159970 800 4 mprj_dat_o_core[30]
port 861 nsew
rlabel metal2 s 160282 0 160338 800 4 mprj_dat_o_core[31]
port 862 nsew
rlabel metal2 s 160650 0 160706 800 4 mprj_dat_o_core[3]
port 863 nsew
rlabel metal2 s 161018 0 161074 800 4 mprj_dat_o_core[4]
port 864 nsew
rlabel metal2 s 161386 0 161442 800 4 mprj_dat_o_core[5]
port 865 nsew
rlabel metal2 s 161754 0 161810 800 4 mprj_dat_o_core[6]
port 866 nsew
rlabel metal2 s 162122 0 162178 800 4 mprj_dat_o_core[7]
port 867 nsew
rlabel metal2 s 162490 0 162546 800 4 mprj_dat_o_core[8]
port 868 nsew
rlabel metal2 s 162858 0 162914 800 4 mprj_dat_o_core[9]
port 869 nsew
rlabel metal2 s 150162 12200 150218 13000 4 mprj_dat_o_user[0]
port 870 nsew
rlabel metal2 s 150530 12200 150586 13000 4 mprj_dat_o_user[10]
port 871 nsew
rlabel metal2 s 150898 12200 150954 13000 4 mprj_dat_o_user[11]
port 872 nsew
rlabel metal2 s 151266 12200 151322 13000 4 mprj_dat_o_user[12]
port 873 nsew
rlabel metal2 s 151634 12200 151690 13000 4 mprj_dat_o_user[13]
port 874 nsew
rlabel metal2 s 152002 12200 152058 13000 4 mprj_dat_o_user[14]
port 875 nsew
rlabel metal2 s 152370 12200 152426 13000 4 mprj_dat_o_user[15]
port 876 nsew
rlabel metal2 s 152738 12200 152794 13000 4 mprj_dat_o_user[16]
port 877 nsew
rlabel metal2 s 153106 12200 153162 13000 4 mprj_dat_o_user[17]
port 878 nsew
rlabel metal2 s 153474 12200 153530 13000 4 mprj_dat_o_user[18]
port 879 nsew
rlabel metal2 s 153842 12200 153898 13000 4 mprj_dat_o_user[19]
port 880 nsew
rlabel metal2 s 154210 12200 154266 13000 4 mprj_dat_o_user[1]
port 881 nsew
rlabel metal2 s 154578 12200 154634 13000 4 mprj_dat_o_user[20]
port 882 nsew
rlabel metal2 s 154946 12200 155002 13000 4 mprj_dat_o_user[21]
port 883 nsew
rlabel metal2 s 155314 12200 155370 13000 4 mprj_dat_o_user[22]
port 884 nsew
rlabel metal2 s 155682 12200 155738 13000 4 mprj_dat_o_user[23]
port 885 nsew
rlabel metal2 s 156050 12200 156106 13000 4 mprj_dat_o_user[24]
port 886 nsew
rlabel metal2 s 156418 12200 156474 13000 4 mprj_dat_o_user[25]
port 887 nsew
rlabel metal2 s 156786 12200 156842 13000 4 mprj_dat_o_user[26]
port 888 nsew
rlabel metal2 s 157154 12200 157210 13000 4 mprj_dat_o_user[27]
port 889 nsew
rlabel metal2 s 157522 12200 157578 13000 4 mprj_dat_o_user[28]
port 890 nsew
rlabel metal2 s 157890 12200 157946 13000 4 mprj_dat_o_user[29]
port 891 nsew
rlabel metal2 s 158258 12200 158314 13000 4 mprj_dat_o_user[2]
port 892 nsew
rlabel metal2 s 158626 12200 158682 13000 4 mprj_dat_o_user[30]
port 893 nsew
rlabel metal2 s 158994 12200 159050 13000 4 mprj_dat_o_user[31]
port 894 nsew
rlabel metal2 s 159362 12200 159418 13000 4 mprj_dat_o_user[3]
port 895 nsew
rlabel metal2 s 159730 12200 159786 13000 4 mprj_dat_o_user[4]
port 896 nsew
rlabel metal2 s 160098 12200 160154 13000 4 mprj_dat_o_user[5]
port 897 nsew
rlabel metal2 s 160466 12200 160522 13000 4 mprj_dat_o_user[6]
port 898 nsew
rlabel metal2 s 160834 12200 160890 13000 4 mprj_dat_o_user[7]
port 899 nsew
rlabel metal2 s 161202 12200 161258 13000 4 mprj_dat_o_user[8]
port 900 nsew
rlabel metal2 s 161570 12200 161626 13000 4 mprj_dat_o_user[9]
port 901 nsew
rlabel metal2 s 163226 0 163282 800 4 mprj_sel_o_core[0]
port 902 nsew
rlabel metal2 s 163594 0 163650 800 4 mprj_sel_o_core[1]
port 903 nsew
rlabel metal2 s 163962 0 164018 800 4 mprj_sel_o_core[2]
port 904 nsew
rlabel metal2 s 164330 0 164386 800 4 mprj_sel_o_core[3]
port 905 nsew
rlabel metal2 s 161938 12200 161994 13000 4 mprj_sel_o_user[0]
port 906 nsew
rlabel metal2 s 162306 12200 162362 13000 4 mprj_sel_o_user[1]
port 907 nsew
rlabel metal2 s 162674 12200 162730 13000 4 mprj_sel_o_user[2]
port 908 nsew
rlabel metal2 s 163042 12200 163098 13000 4 mprj_sel_o_user[3]
port 909 nsew
rlabel metal2 s 164698 0 164754 800 4 mprj_stb_o_core
port 910 nsew
rlabel metal2 s 163410 12200 163466 13000 4 mprj_stb_o_user
port 911 nsew
rlabel metal2 s 165066 0 165122 800 4 mprj_we_o_core
port 912 nsew
rlabel metal2 s 163778 12200 163834 13000 4 mprj_we_o_user
port 913 nsew
rlabel metal2 s 165434 0 165490 800 4 user1_vcc_powergood
port 914 nsew
rlabel metal2 s 165802 0 165858 800 4 user1_vdd_powergood
port 915 nsew
rlabel metal2 s 166170 0 166226 800 4 user2_vcc_powergood
port 916 nsew
rlabel metal2 s 166538 0 166594 800 4 user2_vdd_powergood
port 917 nsew
rlabel metal2 s 164146 12200 164202 13000 4 user_clock
port 918 nsew
rlabel metal2 s 164514 12200 164570 13000 4 user_clock2
port 919 nsew
rlabel metal2 s 164882 12200 164938 13000 4 user_reset
port 920 nsew
rlabel metal2 s 754 0 810 800 4 user_resetn
port 921 nsew
rlabel metal1 s 368 11376 169556 11472 4 VPWR
port 922 nsew
rlabel metal1 s 368 11920 169556 12016 4 VGND
port 923 nsew
<< properties >>
string FIXED_BBOX 0 0 169594 13025
string GDS_FILE /project/openlane/mgmt_protect/runs/mgmt_protect/results/magic/mgmt_protect.gds
string GDS_END 4538328
string GDS_START 130836
<< end >>
