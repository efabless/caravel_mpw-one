sky130_ef_io__vssio_hvc_clamped_pad.cdl