VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 598.760 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.860 597.600 2.140 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.640 597.600 159.920 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.280 597.600 175.560 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.920 597.600 191.200 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.020 597.600 207.300 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.660 597.600 222.940 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 238.300 597.600 238.580 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.400 597.600 254.680 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 270.040 597.600 270.320 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 285.680 597.600 285.960 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.780 597.600 302.060 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.500 597.600 17.780 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.420 597.600 317.700 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.060 597.600 333.340 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 348.700 597.600 348.980 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.800 597.600 365.080 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 380.440 597.600 380.720 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.080 597.600 396.360 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 412.180 597.600 412.460 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 427.820 597.600 428.100 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.460 597.600 443.740 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 459.560 597.600 459.840 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.140 597.600 33.420 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 475.200 597.600 475.480 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.840 597.600 491.120 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.940 597.600 507.220 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 522.580 597.600 522.860 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 538.220 597.600 538.500 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.320 597.600 554.600 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.960 597.600 570.240 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.600 597.600 585.880 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.780 597.600 49.060 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.880 597.600 65.160 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.520 597.600 80.800 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.160 597.600 96.440 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.260 597.600 112.540 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.900 597.600 128.180 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.540 597.600 143.820 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.920 597.600 7.200 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.700 597.600 164.980 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.340 597.600 180.620 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.440 597.600 196.720 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.080 597.600 212.360 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 227.720 597.600 228.000 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.820 597.600 244.100 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.460 597.600 259.740 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 275.100 597.600 275.380 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.200 597.600 291.480 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 306.840 597.600 307.120 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.560 597.600 22.840 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.480 597.600 322.760 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 338.580 597.600 338.860 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.220 597.600 354.500 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 369.860 597.600 370.140 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 385.960 597.600 386.240 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.600 597.600 401.880 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 417.240 597.600 417.520 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 432.880 597.600 433.160 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.980 597.600 449.260 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 464.620 597.600 464.900 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.660 597.600 38.940 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 480.260 597.600 480.540 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.360 597.600 496.640 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 512.000 597.600 512.280 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 527.640 597.600 527.920 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 543.740 597.600 544.020 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 559.380 597.600 559.660 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.020 597.600 575.300 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.120 597.600 591.400 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.300 597.600 54.580 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.940 597.600 70.220 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.040 597.600 86.320 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.680 597.600 101.960 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.320 597.600 117.600 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.960 597.600 133.240 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.060 597.600 149.340 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.980 597.600 12.260 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.220 597.600 170.500 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.860 597.600 186.140 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.500 597.600 201.780 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 217.140 597.600 217.420 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 233.240 597.600 233.520 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.880 597.600 249.160 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.520 597.600 264.800 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 280.620 597.600 280.900 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.260 597.600 296.540 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.900 597.600 312.180 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.080 597.600 28.360 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.000 597.600 328.280 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.640 597.600 343.920 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.280 597.600 359.560 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 375.380 597.600 375.660 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 391.020 597.600 391.300 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 406.660 597.600 406.940 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 422.760 597.600 423.040 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.400 597.600 438.680 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 454.040 597.600 454.320 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 470.140 597.600 470.420 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.720 597.600 44.000 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 485.780 597.600 486.060 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 501.420 597.600 501.700 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 517.060 597.600 517.340 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.160 597.600 533.440 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 548.800 597.600 549.080 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 564.440 597.600 564.720 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 580.540 597.600 580.820 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.180 597.600 596.460 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.360 597.600 59.640 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.460 597.600 75.740 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.100 597.600 91.380 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.740 597.600 107.020 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.840 597.600 123.120 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.480 597.600 138.760 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.120 597.600 154.400 600.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.740 0.000 130.020 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.820 0.000 497.100 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.500 0.000 500.780 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.180 0.000 504.460 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.860 0.000 508.140 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 511.540 0.000 511.820 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 515.220 0.000 515.500 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.900 0.000 519.180 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 522.580 0.000 522.860 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 526.260 0.000 526.540 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 529.940 0.000 530.220 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.080 0.000 166.360 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.620 0.000 533.900 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 537.300 0.000 537.580 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.980 0.000 541.260 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.660 0.000 544.940 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 548.340 0.000 548.620 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 552.020 0.000 552.300 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 555.700 0.000 555.980 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 559.380 0.000 559.660 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 563.060 0.000 563.340 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 566.740 0.000 567.020 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.760 0.000 170.040 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 570.420 0.000 570.700 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.100 0.000 574.380 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 577.780 0.000 578.060 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.460 0.000 581.740 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.140 0.000 585.420 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 588.820 0.000 589.100 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.500 0.000 592.780 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.180 0.000 596.460 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.440 0.000 173.720 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.120 0.000 177.400 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.800 0.000 181.080 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.480 0.000 184.760 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.160 0.000 188.440 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.840 0.000 192.120 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.520 0.000 195.800 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.200 0.000 199.480 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.420 0.000 133.700 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.880 0.000 203.160 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.560 0.000 206.840 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.240 0.000 210.520 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.920 0.000 214.200 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.600 0.000 217.880 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 221.280 0.000 221.560 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.960 0.000 225.240 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.640 0.000 228.920 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.320 0.000 232.600 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.000 0.000 236.280 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.100 0.000 137.380 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.680 0.000 239.960 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 243.360 0.000 243.640 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.040 0.000 247.320 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 250.720 0.000 251.000 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.400 0.000 254.680 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.080 0.000 258.360 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 261.760 0.000 262.040 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.440 0.000 265.720 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.120 0.000 269.400 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 272.800 0.000 273.080 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.780 0.000 141.060 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.480 0.000 276.760 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.160 0.000 280.440 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 283.840 0.000 284.120 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 287.520 0.000 287.800 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.200 0.000 291.480 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.880 0.000 295.160 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.560 0.000 298.840 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.240 0.000 302.520 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.920 0.000 306.200 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 309.600 0.000 309.880 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.460 0.000 144.740 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 313.280 0.000 313.560 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.960 0.000 317.240 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 320.640 0.000 320.920 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.320 0.000 324.600 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.000 0.000 328.280 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.680 0.000 331.960 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.360 0.000 335.640 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.040 0.000 339.320 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 342.720 0.000 343.000 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.400 0.000 346.680 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.140 0.000 148.420 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.080 0.000 350.360 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.760 0.000 354.040 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.440 0.000 357.720 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 361.120 0.000 361.400 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.800 0.000 365.080 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.480 0.000 368.760 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.160 0.000 372.440 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 375.380 0.000 375.660 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.060 0.000 379.340 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.740 0.000 383.020 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.360 0.000 151.640 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.420 0.000 386.700 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.100 0.000 390.380 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 393.780 0.000 394.060 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.460 0.000 397.740 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.140 0.000 401.420 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.820 0.000 405.100 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.500 0.000 408.780 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 412.180 0.000 412.460 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 415.860 0.000 416.140 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.540 0.000 419.820 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.040 0.000 155.320 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 423.220 0.000 423.500 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.900 0.000 427.180 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 430.580 0.000 430.860 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 434.260 0.000 434.540 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.940 0.000 438.220 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 441.620 0.000 441.900 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 445.300 0.000 445.580 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.980 0.000 449.260 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.660 0.000 452.940 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 456.340 0.000 456.620 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.720 0.000 159.000 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.020 0.000 460.300 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 463.700 0.000 463.980 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 467.380 0.000 467.660 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.060 0.000 471.340 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.740 0.000 475.020 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.420 0.000 478.700 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 482.100 0.000 482.380 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 485.780 0.000 486.060 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 489.460 0.000 489.740 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 493.140 0.000 493.420 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.400 0.000 162.680 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.660 0.000 130.940 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 498.200 0.000 498.480 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 501.880 0.000 502.160 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.560 0.000 505.840 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 509.240 0.000 509.520 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 512.920 0.000 513.200 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 516.600 0.000 516.880 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.280 0.000 520.560 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.960 0.000 524.240 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 527.180 0.000 527.460 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.860 0.000 531.140 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.460 0.000 167.740 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.540 0.000 534.820 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 538.220 0.000 538.500 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 541.900 0.000 542.180 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.580 0.000 545.860 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.260 0.000 549.540 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 552.940 0.000 553.220 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.620 0.000 556.900 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 560.300 0.000 560.580 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.980 0.000 564.260 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 567.660 0.000 567.940 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 171.140 0.000 171.420 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 571.340 0.000 571.620 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.020 0.000 575.300 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 578.700 0.000 578.980 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.380 0.000 582.660 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.060 0.000 586.340 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 589.740 0.000 590.020 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.420 0.000 593.700 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 597.100 0.000 597.380 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.820 0.000 175.100 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 178.500 0.000 178.780 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 182.180 0.000 182.460 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.860 0.000 186.140 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 189.540 0.000 189.820 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.220 0.000 193.500 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.900 0.000 197.180 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 200.580 0.000 200.860 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.340 0.000 134.620 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 204.260 0.000 204.540 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 207.940 0.000 208.220 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 211.620 0.000 211.900 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 215.300 0.000 215.580 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 218.980 0.000 219.260 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.660 0.000 222.940 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 226.340 0.000 226.620 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.020 0.000 230.300 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 233.700 0.000 233.980 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.380 0.000 237.660 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.020 0.000 138.300 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 241.060 0.000 241.340 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.740 0.000 245.020 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.420 0.000 248.700 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.100 0.000 252.380 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 255.780 0.000 256.060 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.460 0.000 259.740 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 263.140 0.000 263.420 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.820 0.000 267.100 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.500 0.000 270.780 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.180 0.000 274.460 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.700 0.000 141.980 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.860 0.000 278.140 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 281.540 0.000 281.820 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.220 0.000 285.500 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.900 0.000 289.180 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.580 0.000 292.860 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.260 0.000 296.540 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 299.940 0.000 300.220 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 303.160 0.000 303.440 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 306.840 0.000 307.120 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 310.520 0.000 310.800 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.380 0.000 145.660 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 314.200 0.000 314.480 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 317.880 0.000 318.160 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.560 0.000 321.840 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.240 0.000 325.520 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.920 0.000 329.200 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 332.600 0.000 332.880 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.280 0.000 336.560 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 339.960 0.000 340.240 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.640 0.000 343.920 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.320 0.000 347.600 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.060 0.000 149.340 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.000 0.000 351.280 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.680 0.000 354.960 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 358.360 0.000 358.640 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.040 0.000 362.320 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.720 0.000 366.000 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 369.400 0.000 369.680 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 373.080 0.000 373.360 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 376.760 0.000 377.040 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 380.440 0.000 380.720 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 384.120 0.000 384.400 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.740 0.000 153.020 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 387.800 0.000 388.080 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 391.480 0.000 391.760 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.160 0.000 395.440 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.840 0.000 399.120 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.520 0.000 402.800 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 406.200 0.000 406.480 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.880 0.000 410.160 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.560 0.000 413.840 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 417.240 0.000 417.520 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.920 0.000 421.200 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.420 0.000 156.700 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 424.600 0.000 424.880 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 428.280 0.000 428.560 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.960 0.000 432.240 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.640 0.000 435.920 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 439.320 0.000 439.600 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 443.000 0.000 443.280 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.680 0.000 446.960 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.360 0.000 450.640 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 454.040 0.000 454.320 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.720 0.000 458.000 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.100 0.000 160.380 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 461.400 0.000 461.680 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 465.080 0.000 465.360 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 468.760 0.000 469.040 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.440 0.000 472.720 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 476.120 0.000 476.400 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 479.800 0.000 480.080 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.480 0.000 483.760 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 487.160 0.000 487.440 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 490.840 0.000 491.120 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 494.520 0.000 494.800 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.780 0.000 164.060 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.040 0.000 132.320 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 499.120 0.000 499.400 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 502.800 0.000 503.080 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.480 0.000 506.760 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 510.160 0.000 510.440 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.840 0.000 514.120 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.520 0.000 517.800 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 521.200 0.000 521.480 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.880 0.000 525.160 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 528.560 0.000 528.840 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 532.240 0.000 532.520 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 168.840 0.000 169.120 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 535.920 0.000 536.200 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 539.600 0.000 539.880 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.280 0.000 543.560 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.960 0.000 547.240 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.640 0.000 550.920 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.320 0.000 554.600 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 558.000 0.000 558.280 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.680 0.000 561.960 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.360 0.000 565.640 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.040 0.000 569.320 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.520 0.000 172.800 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.720 0.000 573.000 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 576.400 0.000 576.680 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 580.080 0.000 580.360 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 583.760 0.000 584.040 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.440 0.000 587.720 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 591.120 0.000 591.400 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 594.800 0.000 595.080 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.480 0.000 598.760 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.200 0.000 176.480 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.880 0.000 180.160 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 183.560 0.000 183.840 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.240 0.000 187.520 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.920 0.000 191.200 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.600 0.000 194.880 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.280 0.000 198.560 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 201.960 0.000 202.240 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.720 0.000 136.000 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.640 0.000 205.920 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.320 0.000 209.600 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.000 0.000 213.280 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.680 0.000 216.960 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.360 0.000 220.640 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.040 0.000 224.320 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.260 0.000 227.540 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.940 0.000 231.220 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 234.620 0.000 234.900 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 238.300 0.000 238.580 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.400 0.000 139.680 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.980 0.000 242.260 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 245.660 0.000 245.940 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.340 0.000 249.620 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.020 0.000 253.300 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.700 0.000 256.980 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 260.380 0.000 260.660 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.060 0.000 264.340 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 267.740 0.000 268.020 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.420 0.000 271.700 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.100 0.000 275.380 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.080 0.000 143.360 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.780 0.000 279.060 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.460 0.000 282.740 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 286.140 0.000 286.420 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.820 0.000 290.100 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.500 0.000 293.780 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.180 0.000 297.460 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.860 0.000 301.140 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 304.540 0.000 304.820 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 308.220 0.000 308.500 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.900 0.000 312.180 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 146.760 0.000 147.040 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.580 0.000 315.860 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.260 0.000 319.540 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.940 0.000 323.220 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.620 0.000 326.900 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.300 0.000 330.580 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.980 0.000 334.260 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.660 0.000 337.940 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 341.340 0.000 341.620 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.020 0.000 345.300 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 348.700 0.000 348.980 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.440 0.000 150.720 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.380 0.000 352.660 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.060 0.000 356.340 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.740 0.000 360.020 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.420 0.000 363.700 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.100 0.000 367.380 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.780 0.000 371.060 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.460 0.000 374.740 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 378.140 0.000 378.420 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.820 0.000 382.100 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.500 0.000 385.780 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.120 0.000 154.400 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.180 0.000 389.460 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.860 0.000 393.140 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.540 0.000 396.820 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.220 0.000 400.500 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.900 0.000 404.180 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.580 0.000 407.860 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 411.260 0.000 411.540 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.940 0.000 415.220 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.620 0.000 418.900 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.300 0.000 422.580 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.800 0.000 158.080 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.980 0.000 426.260 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 429.660 0.000 429.940 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.340 0.000 433.620 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.020 0.000 437.300 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.700 0.000 440.980 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.380 0.000 444.660 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.060 0.000 448.340 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.280 0.000 451.560 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.960 0.000 455.240 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 458.640 0.000 458.920 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.480 0.000 161.760 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.320 0.000 462.600 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.000 0.000 466.280 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.680 0.000 469.960 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 473.360 0.000 473.640 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.040 0.000 477.320 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.720 0.000 481.000 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.400 0.000 484.680 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 488.080 0.000 488.360 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 491.760 0.000 492.040 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.440 0.000 495.720 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.160 0.000 165.440 2.400 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.940 0.000 1.220 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.320 0.000 2.600 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.920 0.000 7.200 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.780 0.000 49.060 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.460 0.000 52.740 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.140 0.000 56.420 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.820 0.000 60.100 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.500 0.000 63.780 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.180 0.000 67.460 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.860 0.000 71.140 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.540 0.000 74.820 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.220 0.000 78.500 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.900 0.000 82.180 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.980 0.000 12.260 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.580 0.000 85.860 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.260 0.000 89.540 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.940 0.000 93.220 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.620 0.000 96.900 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.300 0.000 100.580 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.980 0.000 104.260 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.660 0.000 107.940 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.340 0.000 111.620 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.020 0.000 115.300 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.700 0.000 118.980 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.040 0.000 17.320 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.380 0.000 122.660 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.060 0.000 126.340 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.640 0.000 21.920 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.700 0.000 26.980 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.380 0.000 30.660 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.060 0.000 34.340 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.740 0.000 38.020 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.420 0.000 41.700 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.100 0.000 45.380 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.240 0.000 3.520 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.300 0.000 8.580 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.160 0.000 50.440 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.840 0.000 54.120 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.520 0.000 57.800 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.200 0.000 61.480 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.880 0.000 65.160 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.560 0.000 68.840 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.240 0.000 72.520 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.460 0.000 75.740 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.140 0.000 79.420 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.820 0.000 83.100 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.360 0.000 13.640 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.500 0.000 86.780 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.180 0.000 90.460 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.860 0.000 94.140 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.540 0.000 97.820 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.220 0.000 101.500 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.900 0.000 105.180 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.580 0.000 108.860 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.260 0.000 112.540 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.940 0.000 116.220 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.620 0.000 119.900 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.960 0.000 18.240 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.300 0.000 123.580 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.980 0.000 127.260 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.020 0.000 23.300 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.080 0.000 28.360 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.760 0.000 32.040 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.440 0.000 35.720 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.120 0.000 39.400 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.800 0.000 43.080 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.480 0.000 46.760 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.680 0.000 9.960 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.080 0.000 51.360 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.760 0.000 55.040 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.440 0.000 58.720 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.120 0.000 62.400 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.800 0.000 66.080 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.480 0.000 69.760 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.160 0.000 73.440 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.840 0.000 77.120 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.520 0.000 80.800 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.200 0.000 84.480 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.280 0.000 14.560 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.880 0.000 88.160 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.560 0.000 91.840 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.240 0.000 95.520 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.920 0.000 99.200 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.600 0.000 102.880 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.280 0.000 106.560 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.960 0.000 110.240 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.640 0.000 113.920 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.320 0.000 117.600 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.000 0.000 121.280 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.340 0.000 19.620 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.680 0.000 124.960 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.360 0.000 128.640 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.400 0.000 24.680 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.000 0.000 29.280 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.680 0.000 32.960 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.360 0.000 36.640 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.040 0.000 40.320 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.720 0.000 44.000 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.400 0.000 47.680 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.600 0.000 10.880 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.660 0.000 15.940 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.720 0.000 21.000 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.320 0.000 25.600 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.620 0.000 4.900 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.000 0.000 6.280 2.400 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.510 10.640 22.110 587.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.310 10.640 98.910 587.760 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.990 6.545 593.790 587.605 ;
      LAYER met1 ;
        RECT 0.000 5.140 597.400 587.760 ;
      LAYER met2 ;
        RECT 0.030 597.320 1.580 597.600 ;
        RECT 2.420 597.320 6.640 597.600 ;
        RECT 7.480 597.320 11.700 597.600 ;
        RECT 12.540 597.320 17.220 597.600 ;
        RECT 18.060 597.320 22.280 597.600 ;
        RECT 23.120 597.320 27.800 597.600 ;
        RECT 28.640 597.320 32.860 597.600 ;
        RECT 33.700 597.320 38.380 597.600 ;
        RECT 39.220 597.320 43.440 597.600 ;
        RECT 44.280 597.320 48.500 597.600 ;
        RECT 49.340 597.320 54.020 597.600 ;
        RECT 54.860 597.320 59.080 597.600 ;
        RECT 59.920 597.320 64.600 597.600 ;
        RECT 65.440 597.320 69.660 597.600 ;
        RECT 70.500 597.320 75.180 597.600 ;
        RECT 76.020 597.320 80.240 597.600 ;
        RECT 81.080 597.320 85.760 597.600 ;
        RECT 86.600 597.320 90.820 597.600 ;
        RECT 91.660 597.320 95.880 597.600 ;
        RECT 96.720 597.320 101.400 597.600 ;
        RECT 102.240 597.320 106.460 597.600 ;
        RECT 107.300 597.320 111.980 597.600 ;
        RECT 112.820 597.320 117.040 597.600 ;
        RECT 117.880 597.320 122.560 597.600 ;
        RECT 123.400 597.320 127.620 597.600 ;
        RECT 128.460 597.320 132.680 597.600 ;
        RECT 133.520 597.320 138.200 597.600 ;
        RECT 139.040 597.320 143.260 597.600 ;
        RECT 144.100 597.320 148.780 597.600 ;
        RECT 149.620 597.320 153.840 597.600 ;
        RECT 154.680 597.320 159.360 597.600 ;
        RECT 160.200 597.320 164.420 597.600 ;
        RECT 165.260 597.320 169.940 597.600 ;
        RECT 170.780 597.320 175.000 597.600 ;
        RECT 175.840 597.320 180.060 597.600 ;
        RECT 180.900 597.320 185.580 597.600 ;
        RECT 186.420 597.320 190.640 597.600 ;
        RECT 191.480 597.320 196.160 597.600 ;
        RECT 197.000 597.320 201.220 597.600 ;
        RECT 202.060 597.320 206.740 597.600 ;
        RECT 207.580 597.320 211.800 597.600 ;
        RECT 212.640 597.320 216.860 597.600 ;
        RECT 217.700 597.320 222.380 597.600 ;
        RECT 223.220 597.320 227.440 597.600 ;
        RECT 228.280 597.320 232.960 597.600 ;
        RECT 233.800 597.320 238.020 597.600 ;
        RECT 238.860 597.320 243.540 597.600 ;
        RECT 244.380 597.320 248.600 597.600 ;
        RECT 249.440 597.320 254.120 597.600 ;
        RECT 254.960 597.320 259.180 597.600 ;
        RECT 260.020 597.320 264.240 597.600 ;
        RECT 265.080 597.320 269.760 597.600 ;
        RECT 270.600 597.320 274.820 597.600 ;
        RECT 275.660 597.320 280.340 597.600 ;
        RECT 281.180 597.320 285.400 597.600 ;
        RECT 286.240 597.320 290.920 597.600 ;
        RECT 291.760 597.320 295.980 597.600 ;
        RECT 296.820 597.320 301.500 597.600 ;
        RECT 302.340 597.320 306.560 597.600 ;
        RECT 307.400 597.320 311.620 597.600 ;
        RECT 312.460 597.320 317.140 597.600 ;
        RECT 317.980 597.320 322.200 597.600 ;
        RECT 323.040 597.320 327.720 597.600 ;
        RECT 328.560 597.320 332.780 597.600 ;
        RECT 333.620 597.320 338.300 597.600 ;
        RECT 339.140 597.320 343.360 597.600 ;
        RECT 344.200 597.320 348.420 597.600 ;
        RECT 349.260 597.320 353.940 597.600 ;
        RECT 354.780 597.320 359.000 597.600 ;
        RECT 359.840 597.320 364.520 597.600 ;
        RECT 365.360 597.320 369.580 597.600 ;
        RECT 370.420 597.320 375.100 597.600 ;
        RECT 375.940 597.320 380.160 597.600 ;
        RECT 381.000 597.320 385.680 597.600 ;
        RECT 386.520 597.320 390.740 597.600 ;
        RECT 391.580 597.320 395.800 597.600 ;
        RECT 396.640 597.320 401.320 597.600 ;
        RECT 402.160 597.320 406.380 597.600 ;
        RECT 407.220 597.320 411.900 597.600 ;
        RECT 412.740 597.320 416.960 597.600 ;
        RECT 417.800 597.320 422.480 597.600 ;
        RECT 423.320 597.320 427.540 597.600 ;
        RECT 428.380 597.320 432.600 597.600 ;
        RECT 433.440 597.320 438.120 597.600 ;
        RECT 438.960 597.320 443.180 597.600 ;
        RECT 444.020 597.320 448.700 597.600 ;
        RECT 449.540 597.320 453.760 597.600 ;
        RECT 454.600 597.320 459.280 597.600 ;
        RECT 460.120 597.320 464.340 597.600 ;
        RECT 465.180 597.320 469.860 597.600 ;
        RECT 470.700 597.320 474.920 597.600 ;
        RECT 475.760 597.320 479.980 597.600 ;
        RECT 480.820 597.320 485.500 597.600 ;
        RECT 486.340 597.320 490.560 597.600 ;
        RECT 491.400 597.320 496.080 597.600 ;
        RECT 496.920 597.320 501.140 597.600 ;
        RECT 501.980 597.320 506.660 597.600 ;
        RECT 507.500 597.320 511.720 597.600 ;
        RECT 512.560 597.320 516.780 597.600 ;
        RECT 517.620 597.320 522.300 597.600 ;
        RECT 523.140 597.320 527.360 597.600 ;
        RECT 528.200 597.320 532.880 597.600 ;
        RECT 533.720 597.320 537.940 597.600 ;
        RECT 538.780 597.320 543.460 597.600 ;
        RECT 544.300 597.320 548.520 597.600 ;
        RECT 549.360 597.320 554.040 597.600 ;
        RECT 554.880 597.320 559.100 597.600 ;
        RECT 559.940 597.320 564.160 597.600 ;
        RECT 565.000 597.320 569.680 597.600 ;
        RECT 570.520 597.320 574.740 597.600 ;
        RECT 575.580 597.320 580.260 597.600 ;
        RECT 581.100 597.320 585.320 597.600 ;
        RECT 586.160 597.320 590.840 597.600 ;
        RECT 591.680 597.320 595.900 597.600 ;
        RECT 596.740 597.320 597.370 597.600 ;
        RECT 0.030 2.680 597.370 597.320 ;
        RECT 0.580 2.400 0.660 2.680 ;
        RECT 1.500 2.400 2.040 2.680 ;
        RECT 2.880 2.400 2.960 2.680 ;
        RECT 3.800 2.400 4.340 2.680 ;
        RECT 5.180 2.400 5.720 2.680 ;
        RECT 6.560 2.400 6.640 2.680 ;
        RECT 7.480 2.400 8.020 2.680 ;
        RECT 8.860 2.400 9.400 2.680 ;
        RECT 10.240 2.400 10.320 2.680 ;
        RECT 11.160 2.400 11.700 2.680 ;
        RECT 12.540 2.400 13.080 2.680 ;
        RECT 13.920 2.400 14.000 2.680 ;
        RECT 14.840 2.400 15.380 2.680 ;
        RECT 16.220 2.400 16.760 2.680 ;
        RECT 17.600 2.400 17.680 2.680 ;
        RECT 18.520 2.400 19.060 2.680 ;
        RECT 19.900 2.400 20.440 2.680 ;
        RECT 21.280 2.400 21.360 2.680 ;
        RECT 22.200 2.400 22.740 2.680 ;
        RECT 23.580 2.400 24.120 2.680 ;
        RECT 24.960 2.400 25.040 2.680 ;
        RECT 25.880 2.400 26.420 2.680 ;
        RECT 27.260 2.400 27.800 2.680 ;
        RECT 28.640 2.400 28.720 2.680 ;
        RECT 29.560 2.400 30.100 2.680 ;
        RECT 30.940 2.400 31.480 2.680 ;
        RECT 32.320 2.400 32.400 2.680 ;
        RECT 33.240 2.400 33.780 2.680 ;
        RECT 34.620 2.400 35.160 2.680 ;
        RECT 36.000 2.400 36.080 2.680 ;
        RECT 36.920 2.400 37.460 2.680 ;
        RECT 38.300 2.400 38.840 2.680 ;
        RECT 39.680 2.400 39.760 2.680 ;
        RECT 40.600 2.400 41.140 2.680 ;
        RECT 41.980 2.400 42.520 2.680 ;
        RECT 43.360 2.400 43.440 2.680 ;
        RECT 44.280 2.400 44.820 2.680 ;
        RECT 45.660 2.400 46.200 2.680 ;
        RECT 47.040 2.400 47.120 2.680 ;
        RECT 47.960 2.400 48.500 2.680 ;
        RECT 49.340 2.400 49.880 2.680 ;
        RECT 50.720 2.400 50.800 2.680 ;
        RECT 51.640 2.400 52.180 2.680 ;
        RECT 53.020 2.400 53.560 2.680 ;
        RECT 54.400 2.400 54.480 2.680 ;
        RECT 55.320 2.400 55.860 2.680 ;
        RECT 56.700 2.400 57.240 2.680 ;
        RECT 58.080 2.400 58.160 2.680 ;
        RECT 59.000 2.400 59.540 2.680 ;
        RECT 60.380 2.400 60.920 2.680 ;
        RECT 61.760 2.400 61.840 2.680 ;
        RECT 62.680 2.400 63.220 2.680 ;
        RECT 64.060 2.400 64.600 2.680 ;
        RECT 65.440 2.400 65.520 2.680 ;
        RECT 66.360 2.400 66.900 2.680 ;
        RECT 67.740 2.400 68.280 2.680 ;
        RECT 69.120 2.400 69.200 2.680 ;
        RECT 70.040 2.400 70.580 2.680 ;
        RECT 71.420 2.400 71.960 2.680 ;
        RECT 72.800 2.400 72.880 2.680 ;
        RECT 73.720 2.400 74.260 2.680 ;
        RECT 75.100 2.400 75.180 2.680 ;
        RECT 76.020 2.400 76.560 2.680 ;
        RECT 77.400 2.400 77.940 2.680 ;
        RECT 78.780 2.400 78.860 2.680 ;
        RECT 79.700 2.400 80.240 2.680 ;
        RECT 81.080 2.400 81.620 2.680 ;
        RECT 82.460 2.400 82.540 2.680 ;
        RECT 83.380 2.400 83.920 2.680 ;
        RECT 84.760 2.400 85.300 2.680 ;
        RECT 86.140 2.400 86.220 2.680 ;
        RECT 87.060 2.400 87.600 2.680 ;
        RECT 88.440 2.400 88.980 2.680 ;
        RECT 89.820 2.400 89.900 2.680 ;
        RECT 90.740 2.400 91.280 2.680 ;
        RECT 92.120 2.400 92.660 2.680 ;
        RECT 93.500 2.400 93.580 2.680 ;
        RECT 94.420 2.400 94.960 2.680 ;
        RECT 95.800 2.400 96.340 2.680 ;
        RECT 97.180 2.400 97.260 2.680 ;
        RECT 98.100 2.400 98.640 2.680 ;
        RECT 99.480 2.400 100.020 2.680 ;
        RECT 100.860 2.400 100.940 2.680 ;
        RECT 101.780 2.400 102.320 2.680 ;
        RECT 103.160 2.400 103.700 2.680 ;
        RECT 104.540 2.400 104.620 2.680 ;
        RECT 105.460 2.400 106.000 2.680 ;
        RECT 106.840 2.400 107.380 2.680 ;
        RECT 108.220 2.400 108.300 2.680 ;
        RECT 109.140 2.400 109.680 2.680 ;
        RECT 110.520 2.400 111.060 2.680 ;
        RECT 111.900 2.400 111.980 2.680 ;
        RECT 112.820 2.400 113.360 2.680 ;
        RECT 114.200 2.400 114.740 2.680 ;
        RECT 115.580 2.400 115.660 2.680 ;
        RECT 116.500 2.400 117.040 2.680 ;
        RECT 117.880 2.400 118.420 2.680 ;
        RECT 119.260 2.400 119.340 2.680 ;
        RECT 120.180 2.400 120.720 2.680 ;
        RECT 121.560 2.400 122.100 2.680 ;
        RECT 122.940 2.400 123.020 2.680 ;
        RECT 123.860 2.400 124.400 2.680 ;
        RECT 125.240 2.400 125.780 2.680 ;
        RECT 126.620 2.400 126.700 2.680 ;
        RECT 127.540 2.400 128.080 2.680 ;
        RECT 128.920 2.400 129.460 2.680 ;
        RECT 130.300 2.400 130.380 2.680 ;
        RECT 131.220 2.400 131.760 2.680 ;
        RECT 132.600 2.400 133.140 2.680 ;
        RECT 133.980 2.400 134.060 2.680 ;
        RECT 134.900 2.400 135.440 2.680 ;
        RECT 136.280 2.400 136.820 2.680 ;
        RECT 137.660 2.400 137.740 2.680 ;
        RECT 138.580 2.400 139.120 2.680 ;
        RECT 139.960 2.400 140.500 2.680 ;
        RECT 141.340 2.400 141.420 2.680 ;
        RECT 142.260 2.400 142.800 2.680 ;
        RECT 143.640 2.400 144.180 2.680 ;
        RECT 145.020 2.400 145.100 2.680 ;
        RECT 145.940 2.400 146.480 2.680 ;
        RECT 147.320 2.400 147.860 2.680 ;
        RECT 148.700 2.400 148.780 2.680 ;
        RECT 149.620 2.400 150.160 2.680 ;
        RECT 151.000 2.400 151.080 2.680 ;
        RECT 151.920 2.400 152.460 2.680 ;
        RECT 153.300 2.400 153.840 2.680 ;
        RECT 154.680 2.400 154.760 2.680 ;
        RECT 155.600 2.400 156.140 2.680 ;
        RECT 156.980 2.400 157.520 2.680 ;
        RECT 158.360 2.400 158.440 2.680 ;
        RECT 159.280 2.400 159.820 2.680 ;
        RECT 160.660 2.400 161.200 2.680 ;
        RECT 162.040 2.400 162.120 2.680 ;
        RECT 162.960 2.400 163.500 2.680 ;
        RECT 164.340 2.400 164.880 2.680 ;
        RECT 165.720 2.400 165.800 2.680 ;
        RECT 166.640 2.400 167.180 2.680 ;
        RECT 168.020 2.400 168.560 2.680 ;
        RECT 169.400 2.400 169.480 2.680 ;
        RECT 170.320 2.400 170.860 2.680 ;
        RECT 171.700 2.400 172.240 2.680 ;
        RECT 173.080 2.400 173.160 2.680 ;
        RECT 174.000 2.400 174.540 2.680 ;
        RECT 175.380 2.400 175.920 2.680 ;
        RECT 176.760 2.400 176.840 2.680 ;
        RECT 177.680 2.400 178.220 2.680 ;
        RECT 179.060 2.400 179.600 2.680 ;
        RECT 180.440 2.400 180.520 2.680 ;
        RECT 181.360 2.400 181.900 2.680 ;
        RECT 182.740 2.400 183.280 2.680 ;
        RECT 184.120 2.400 184.200 2.680 ;
        RECT 185.040 2.400 185.580 2.680 ;
        RECT 186.420 2.400 186.960 2.680 ;
        RECT 187.800 2.400 187.880 2.680 ;
        RECT 188.720 2.400 189.260 2.680 ;
        RECT 190.100 2.400 190.640 2.680 ;
        RECT 191.480 2.400 191.560 2.680 ;
        RECT 192.400 2.400 192.940 2.680 ;
        RECT 193.780 2.400 194.320 2.680 ;
        RECT 195.160 2.400 195.240 2.680 ;
        RECT 196.080 2.400 196.620 2.680 ;
        RECT 197.460 2.400 198.000 2.680 ;
        RECT 198.840 2.400 198.920 2.680 ;
        RECT 199.760 2.400 200.300 2.680 ;
        RECT 201.140 2.400 201.680 2.680 ;
        RECT 202.520 2.400 202.600 2.680 ;
        RECT 203.440 2.400 203.980 2.680 ;
        RECT 204.820 2.400 205.360 2.680 ;
        RECT 206.200 2.400 206.280 2.680 ;
        RECT 207.120 2.400 207.660 2.680 ;
        RECT 208.500 2.400 209.040 2.680 ;
        RECT 209.880 2.400 209.960 2.680 ;
        RECT 210.800 2.400 211.340 2.680 ;
        RECT 212.180 2.400 212.720 2.680 ;
        RECT 213.560 2.400 213.640 2.680 ;
        RECT 214.480 2.400 215.020 2.680 ;
        RECT 215.860 2.400 216.400 2.680 ;
        RECT 217.240 2.400 217.320 2.680 ;
        RECT 218.160 2.400 218.700 2.680 ;
        RECT 219.540 2.400 220.080 2.680 ;
        RECT 220.920 2.400 221.000 2.680 ;
        RECT 221.840 2.400 222.380 2.680 ;
        RECT 223.220 2.400 223.760 2.680 ;
        RECT 224.600 2.400 224.680 2.680 ;
        RECT 225.520 2.400 226.060 2.680 ;
        RECT 226.900 2.400 226.980 2.680 ;
        RECT 227.820 2.400 228.360 2.680 ;
        RECT 229.200 2.400 229.740 2.680 ;
        RECT 230.580 2.400 230.660 2.680 ;
        RECT 231.500 2.400 232.040 2.680 ;
        RECT 232.880 2.400 233.420 2.680 ;
        RECT 234.260 2.400 234.340 2.680 ;
        RECT 235.180 2.400 235.720 2.680 ;
        RECT 236.560 2.400 237.100 2.680 ;
        RECT 237.940 2.400 238.020 2.680 ;
        RECT 238.860 2.400 239.400 2.680 ;
        RECT 240.240 2.400 240.780 2.680 ;
        RECT 241.620 2.400 241.700 2.680 ;
        RECT 242.540 2.400 243.080 2.680 ;
        RECT 243.920 2.400 244.460 2.680 ;
        RECT 245.300 2.400 245.380 2.680 ;
        RECT 246.220 2.400 246.760 2.680 ;
        RECT 247.600 2.400 248.140 2.680 ;
        RECT 248.980 2.400 249.060 2.680 ;
        RECT 249.900 2.400 250.440 2.680 ;
        RECT 251.280 2.400 251.820 2.680 ;
        RECT 252.660 2.400 252.740 2.680 ;
        RECT 253.580 2.400 254.120 2.680 ;
        RECT 254.960 2.400 255.500 2.680 ;
        RECT 256.340 2.400 256.420 2.680 ;
        RECT 257.260 2.400 257.800 2.680 ;
        RECT 258.640 2.400 259.180 2.680 ;
        RECT 260.020 2.400 260.100 2.680 ;
        RECT 260.940 2.400 261.480 2.680 ;
        RECT 262.320 2.400 262.860 2.680 ;
        RECT 263.700 2.400 263.780 2.680 ;
        RECT 264.620 2.400 265.160 2.680 ;
        RECT 266.000 2.400 266.540 2.680 ;
        RECT 267.380 2.400 267.460 2.680 ;
        RECT 268.300 2.400 268.840 2.680 ;
        RECT 269.680 2.400 270.220 2.680 ;
        RECT 271.060 2.400 271.140 2.680 ;
        RECT 271.980 2.400 272.520 2.680 ;
        RECT 273.360 2.400 273.900 2.680 ;
        RECT 274.740 2.400 274.820 2.680 ;
        RECT 275.660 2.400 276.200 2.680 ;
        RECT 277.040 2.400 277.580 2.680 ;
        RECT 278.420 2.400 278.500 2.680 ;
        RECT 279.340 2.400 279.880 2.680 ;
        RECT 280.720 2.400 281.260 2.680 ;
        RECT 282.100 2.400 282.180 2.680 ;
        RECT 283.020 2.400 283.560 2.680 ;
        RECT 284.400 2.400 284.940 2.680 ;
        RECT 285.780 2.400 285.860 2.680 ;
        RECT 286.700 2.400 287.240 2.680 ;
        RECT 288.080 2.400 288.620 2.680 ;
        RECT 289.460 2.400 289.540 2.680 ;
        RECT 290.380 2.400 290.920 2.680 ;
        RECT 291.760 2.400 292.300 2.680 ;
        RECT 293.140 2.400 293.220 2.680 ;
        RECT 294.060 2.400 294.600 2.680 ;
        RECT 295.440 2.400 295.980 2.680 ;
        RECT 296.820 2.400 296.900 2.680 ;
        RECT 297.740 2.400 298.280 2.680 ;
        RECT 299.120 2.400 299.660 2.680 ;
        RECT 300.500 2.400 300.580 2.680 ;
        RECT 301.420 2.400 301.960 2.680 ;
        RECT 302.800 2.400 302.880 2.680 ;
        RECT 303.720 2.400 304.260 2.680 ;
        RECT 305.100 2.400 305.640 2.680 ;
        RECT 306.480 2.400 306.560 2.680 ;
        RECT 307.400 2.400 307.940 2.680 ;
        RECT 308.780 2.400 309.320 2.680 ;
        RECT 310.160 2.400 310.240 2.680 ;
        RECT 311.080 2.400 311.620 2.680 ;
        RECT 312.460 2.400 313.000 2.680 ;
        RECT 313.840 2.400 313.920 2.680 ;
        RECT 314.760 2.400 315.300 2.680 ;
        RECT 316.140 2.400 316.680 2.680 ;
        RECT 317.520 2.400 317.600 2.680 ;
        RECT 318.440 2.400 318.980 2.680 ;
        RECT 319.820 2.400 320.360 2.680 ;
        RECT 321.200 2.400 321.280 2.680 ;
        RECT 322.120 2.400 322.660 2.680 ;
        RECT 323.500 2.400 324.040 2.680 ;
        RECT 324.880 2.400 324.960 2.680 ;
        RECT 325.800 2.400 326.340 2.680 ;
        RECT 327.180 2.400 327.720 2.680 ;
        RECT 328.560 2.400 328.640 2.680 ;
        RECT 329.480 2.400 330.020 2.680 ;
        RECT 330.860 2.400 331.400 2.680 ;
        RECT 332.240 2.400 332.320 2.680 ;
        RECT 333.160 2.400 333.700 2.680 ;
        RECT 334.540 2.400 335.080 2.680 ;
        RECT 335.920 2.400 336.000 2.680 ;
        RECT 336.840 2.400 337.380 2.680 ;
        RECT 338.220 2.400 338.760 2.680 ;
        RECT 339.600 2.400 339.680 2.680 ;
        RECT 340.520 2.400 341.060 2.680 ;
        RECT 341.900 2.400 342.440 2.680 ;
        RECT 343.280 2.400 343.360 2.680 ;
        RECT 344.200 2.400 344.740 2.680 ;
        RECT 345.580 2.400 346.120 2.680 ;
        RECT 346.960 2.400 347.040 2.680 ;
        RECT 347.880 2.400 348.420 2.680 ;
        RECT 349.260 2.400 349.800 2.680 ;
        RECT 350.640 2.400 350.720 2.680 ;
        RECT 351.560 2.400 352.100 2.680 ;
        RECT 352.940 2.400 353.480 2.680 ;
        RECT 354.320 2.400 354.400 2.680 ;
        RECT 355.240 2.400 355.780 2.680 ;
        RECT 356.620 2.400 357.160 2.680 ;
        RECT 358.000 2.400 358.080 2.680 ;
        RECT 358.920 2.400 359.460 2.680 ;
        RECT 360.300 2.400 360.840 2.680 ;
        RECT 361.680 2.400 361.760 2.680 ;
        RECT 362.600 2.400 363.140 2.680 ;
        RECT 363.980 2.400 364.520 2.680 ;
        RECT 365.360 2.400 365.440 2.680 ;
        RECT 366.280 2.400 366.820 2.680 ;
        RECT 367.660 2.400 368.200 2.680 ;
        RECT 369.040 2.400 369.120 2.680 ;
        RECT 369.960 2.400 370.500 2.680 ;
        RECT 371.340 2.400 371.880 2.680 ;
        RECT 372.720 2.400 372.800 2.680 ;
        RECT 373.640 2.400 374.180 2.680 ;
        RECT 375.020 2.400 375.100 2.680 ;
        RECT 375.940 2.400 376.480 2.680 ;
        RECT 377.320 2.400 377.860 2.680 ;
        RECT 378.700 2.400 378.780 2.680 ;
        RECT 379.620 2.400 380.160 2.680 ;
        RECT 381.000 2.400 381.540 2.680 ;
        RECT 382.380 2.400 382.460 2.680 ;
        RECT 383.300 2.400 383.840 2.680 ;
        RECT 384.680 2.400 385.220 2.680 ;
        RECT 386.060 2.400 386.140 2.680 ;
        RECT 386.980 2.400 387.520 2.680 ;
        RECT 388.360 2.400 388.900 2.680 ;
        RECT 389.740 2.400 389.820 2.680 ;
        RECT 390.660 2.400 391.200 2.680 ;
        RECT 392.040 2.400 392.580 2.680 ;
        RECT 393.420 2.400 393.500 2.680 ;
        RECT 394.340 2.400 394.880 2.680 ;
        RECT 395.720 2.400 396.260 2.680 ;
        RECT 397.100 2.400 397.180 2.680 ;
        RECT 398.020 2.400 398.560 2.680 ;
        RECT 399.400 2.400 399.940 2.680 ;
        RECT 400.780 2.400 400.860 2.680 ;
        RECT 401.700 2.400 402.240 2.680 ;
        RECT 403.080 2.400 403.620 2.680 ;
        RECT 404.460 2.400 404.540 2.680 ;
        RECT 405.380 2.400 405.920 2.680 ;
        RECT 406.760 2.400 407.300 2.680 ;
        RECT 408.140 2.400 408.220 2.680 ;
        RECT 409.060 2.400 409.600 2.680 ;
        RECT 410.440 2.400 410.980 2.680 ;
        RECT 411.820 2.400 411.900 2.680 ;
        RECT 412.740 2.400 413.280 2.680 ;
        RECT 414.120 2.400 414.660 2.680 ;
        RECT 415.500 2.400 415.580 2.680 ;
        RECT 416.420 2.400 416.960 2.680 ;
        RECT 417.800 2.400 418.340 2.680 ;
        RECT 419.180 2.400 419.260 2.680 ;
        RECT 420.100 2.400 420.640 2.680 ;
        RECT 421.480 2.400 422.020 2.680 ;
        RECT 422.860 2.400 422.940 2.680 ;
        RECT 423.780 2.400 424.320 2.680 ;
        RECT 425.160 2.400 425.700 2.680 ;
        RECT 426.540 2.400 426.620 2.680 ;
        RECT 427.460 2.400 428.000 2.680 ;
        RECT 428.840 2.400 429.380 2.680 ;
        RECT 430.220 2.400 430.300 2.680 ;
        RECT 431.140 2.400 431.680 2.680 ;
        RECT 432.520 2.400 433.060 2.680 ;
        RECT 433.900 2.400 433.980 2.680 ;
        RECT 434.820 2.400 435.360 2.680 ;
        RECT 436.200 2.400 436.740 2.680 ;
        RECT 437.580 2.400 437.660 2.680 ;
        RECT 438.500 2.400 439.040 2.680 ;
        RECT 439.880 2.400 440.420 2.680 ;
        RECT 441.260 2.400 441.340 2.680 ;
        RECT 442.180 2.400 442.720 2.680 ;
        RECT 443.560 2.400 444.100 2.680 ;
        RECT 444.940 2.400 445.020 2.680 ;
        RECT 445.860 2.400 446.400 2.680 ;
        RECT 447.240 2.400 447.780 2.680 ;
        RECT 448.620 2.400 448.700 2.680 ;
        RECT 449.540 2.400 450.080 2.680 ;
        RECT 450.920 2.400 451.000 2.680 ;
        RECT 451.840 2.400 452.380 2.680 ;
        RECT 453.220 2.400 453.760 2.680 ;
        RECT 454.600 2.400 454.680 2.680 ;
        RECT 455.520 2.400 456.060 2.680 ;
        RECT 456.900 2.400 457.440 2.680 ;
        RECT 458.280 2.400 458.360 2.680 ;
        RECT 459.200 2.400 459.740 2.680 ;
        RECT 460.580 2.400 461.120 2.680 ;
        RECT 461.960 2.400 462.040 2.680 ;
        RECT 462.880 2.400 463.420 2.680 ;
        RECT 464.260 2.400 464.800 2.680 ;
        RECT 465.640 2.400 465.720 2.680 ;
        RECT 466.560 2.400 467.100 2.680 ;
        RECT 467.940 2.400 468.480 2.680 ;
        RECT 469.320 2.400 469.400 2.680 ;
        RECT 470.240 2.400 470.780 2.680 ;
        RECT 471.620 2.400 472.160 2.680 ;
        RECT 473.000 2.400 473.080 2.680 ;
        RECT 473.920 2.400 474.460 2.680 ;
        RECT 475.300 2.400 475.840 2.680 ;
        RECT 476.680 2.400 476.760 2.680 ;
        RECT 477.600 2.400 478.140 2.680 ;
        RECT 478.980 2.400 479.520 2.680 ;
        RECT 480.360 2.400 480.440 2.680 ;
        RECT 481.280 2.400 481.820 2.680 ;
        RECT 482.660 2.400 483.200 2.680 ;
        RECT 484.040 2.400 484.120 2.680 ;
        RECT 484.960 2.400 485.500 2.680 ;
        RECT 486.340 2.400 486.880 2.680 ;
        RECT 487.720 2.400 487.800 2.680 ;
        RECT 488.640 2.400 489.180 2.680 ;
        RECT 490.020 2.400 490.560 2.680 ;
        RECT 491.400 2.400 491.480 2.680 ;
        RECT 492.320 2.400 492.860 2.680 ;
        RECT 493.700 2.400 494.240 2.680 ;
        RECT 495.080 2.400 495.160 2.680 ;
        RECT 496.000 2.400 496.540 2.680 ;
        RECT 497.380 2.400 497.920 2.680 ;
        RECT 498.760 2.400 498.840 2.680 ;
        RECT 499.680 2.400 500.220 2.680 ;
        RECT 501.060 2.400 501.600 2.680 ;
        RECT 502.440 2.400 502.520 2.680 ;
        RECT 503.360 2.400 503.900 2.680 ;
        RECT 504.740 2.400 505.280 2.680 ;
        RECT 506.120 2.400 506.200 2.680 ;
        RECT 507.040 2.400 507.580 2.680 ;
        RECT 508.420 2.400 508.960 2.680 ;
        RECT 509.800 2.400 509.880 2.680 ;
        RECT 510.720 2.400 511.260 2.680 ;
        RECT 512.100 2.400 512.640 2.680 ;
        RECT 513.480 2.400 513.560 2.680 ;
        RECT 514.400 2.400 514.940 2.680 ;
        RECT 515.780 2.400 516.320 2.680 ;
        RECT 517.160 2.400 517.240 2.680 ;
        RECT 518.080 2.400 518.620 2.680 ;
        RECT 519.460 2.400 520.000 2.680 ;
        RECT 520.840 2.400 520.920 2.680 ;
        RECT 521.760 2.400 522.300 2.680 ;
        RECT 523.140 2.400 523.680 2.680 ;
        RECT 524.520 2.400 524.600 2.680 ;
        RECT 525.440 2.400 525.980 2.680 ;
        RECT 526.820 2.400 526.900 2.680 ;
        RECT 527.740 2.400 528.280 2.680 ;
        RECT 529.120 2.400 529.660 2.680 ;
        RECT 530.500 2.400 530.580 2.680 ;
        RECT 531.420 2.400 531.960 2.680 ;
        RECT 532.800 2.400 533.340 2.680 ;
        RECT 534.180 2.400 534.260 2.680 ;
        RECT 535.100 2.400 535.640 2.680 ;
        RECT 536.480 2.400 537.020 2.680 ;
        RECT 537.860 2.400 537.940 2.680 ;
        RECT 538.780 2.400 539.320 2.680 ;
        RECT 540.160 2.400 540.700 2.680 ;
        RECT 541.540 2.400 541.620 2.680 ;
        RECT 542.460 2.400 543.000 2.680 ;
        RECT 543.840 2.400 544.380 2.680 ;
        RECT 545.220 2.400 545.300 2.680 ;
        RECT 546.140 2.400 546.680 2.680 ;
        RECT 547.520 2.400 548.060 2.680 ;
        RECT 548.900 2.400 548.980 2.680 ;
        RECT 549.820 2.400 550.360 2.680 ;
        RECT 551.200 2.400 551.740 2.680 ;
        RECT 552.580 2.400 552.660 2.680 ;
        RECT 553.500 2.400 554.040 2.680 ;
        RECT 554.880 2.400 555.420 2.680 ;
        RECT 556.260 2.400 556.340 2.680 ;
        RECT 557.180 2.400 557.720 2.680 ;
        RECT 558.560 2.400 559.100 2.680 ;
        RECT 559.940 2.400 560.020 2.680 ;
        RECT 560.860 2.400 561.400 2.680 ;
        RECT 562.240 2.400 562.780 2.680 ;
        RECT 563.620 2.400 563.700 2.680 ;
        RECT 564.540 2.400 565.080 2.680 ;
        RECT 565.920 2.400 566.460 2.680 ;
        RECT 567.300 2.400 567.380 2.680 ;
        RECT 568.220 2.400 568.760 2.680 ;
        RECT 569.600 2.400 570.140 2.680 ;
        RECT 570.980 2.400 571.060 2.680 ;
        RECT 571.900 2.400 572.440 2.680 ;
        RECT 573.280 2.400 573.820 2.680 ;
        RECT 574.660 2.400 574.740 2.680 ;
        RECT 575.580 2.400 576.120 2.680 ;
        RECT 576.960 2.400 577.500 2.680 ;
        RECT 578.340 2.400 578.420 2.680 ;
        RECT 579.260 2.400 579.800 2.680 ;
        RECT 580.640 2.400 581.180 2.680 ;
        RECT 582.020 2.400 582.100 2.680 ;
        RECT 582.940 2.400 583.480 2.680 ;
        RECT 584.320 2.400 584.860 2.680 ;
        RECT 585.700 2.400 585.780 2.680 ;
        RECT 586.620 2.400 587.160 2.680 ;
        RECT 588.000 2.400 588.540 2.680 ;
        RECT 589.380 2.400 589.460 2.680 ;
        RECT 590.300 2.400 590.840 2.680 ;
        RECT 591.680 2.400 592.220 2.680 ;
        RECT 593.060 2.400 593.140 2.680 ;
        RECT 593.980 2.400 594.520 2.680 ;
        RECT 595.360 2.400 595.900 2.680 ;
        RECT 596.740 2.400 596.820 2.680 ;
      LAYER met3 ;
        RECT 0.915 9.695 559.710 587.685 ;
      LAYER met4 ;
        RECT 134.085 9.695 559.710 587.760 ;
  END
END user_proj_example
END LIBRARY

