.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/top_gpiov2/sky130_fd_io__top_gpiov2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/amuxsplitv2_delay/sky130_fd_io__amuxsplitv2_delay.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/amuxsplitv2_switch_levelshifter/sky130_fd_io__amuxsplitv2_switch_levelshifter.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/amuxsplitv2_switch_s0/sky130_fd_io__amuxsplitv2_switch_s0.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/amuxsplitv2_switch/sky130_fd_io__amuxsplitv2_switch.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/amuxsplitv2_switch_sl/sky130_fd_io__amuxsplitv2_switch_sl.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/amx_inv1/sky130_fd_io__amx_inv1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_cclat_hvnand3/sky130_fd_io__com_cclat_hvnand3.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_cclat_hvnor3/sky130_fd_io__com_cclat_hvnor3.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_cclat_i2c_fix/sky130_fd_io__com_cclat_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_cclat_inv_in/sky130_fd_io__com_cclat_inv_in.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_cclat_inv_out/sky130_fd_io__com_cclat_inv_out.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_cclat/sky130_fd_io__com_cclat.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_ctl_ls/sky130_fd_io__com_ctl_ls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_inv_x1_dnw/sky130_fd_io__com_inv_x1_dnw.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_nand2_dnw/sky130_fd_io__com_nand2_dnw.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_nor2_dnw/sky130_fd_io__com_nor2_dnw.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pad/sky130_fd_io__com_pad.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pddrvr_unit_2_5/sky130_fd_io__com_pddrvr_unit_2_5.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pdpredrvr_pbias/sky130_fd_io__com_pdpredrvr_pbias.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pdpredrvr_strong_slow/sky130_fd_io__com_pdpredrvr_strong_slow.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pdpredrvr_weak/sky130_fd_io__com_pdpredrvr_weak.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pudrvr_strong_slow/sky130_fd_io__com_pudrvr_strong_slow.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pudrvr_weak/sky130_fd_io__com_pudrvr_weak.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pupredrvr_nbias/sky130_fd_io__com_pupredrvr_nbias.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pupredrvr_strong_slow/sky130_fd_io__com_pupredrvr_strong_slow.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_pupredrvr_weak/sky130_fd_io__com_pupredrvr_weak.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_res_strong_slow/sky130_fd_io__com_res_strong_slow.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_res_weak/sky130_fd_io__com_res_weak.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/com_xres_weak_pu/sky130_fd_io__com_xres_weak_pu.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/enh_nand2_1/sky130_fd_io__enh_nand2_1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/enh_nand2_1_sp/sky130_fd_io__enh_nand2_1_sp.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/enh_nor2_x1/sky130_fd_io__enh_nor2_x1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_buf_localesd/sky130_fd_io__gpio_buf_localesd.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ctlv2_i2c_fix/sky130_fd_io__gpio_ctlv2_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_dat_ls_i2c_fix/sky130_fd_io__gpio_dat_ls_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_dat_ls/sky130_fd_io__gpio_dat_ls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_amux_i2c_fix/sky130_fd_io__gpio_ovtv2_amux_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_amux_switch/sky130_fd_io__gpio_ovtv2_amux_switch.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_buf_localesd/sky130_fd_io__gpio_ovtv2_buf_localesd.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_ctl_hld_i2c_fix/sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_ctl_lsbank_i2c_fix/sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_bias/sky130_fd_io__gpio_ovtv2_hotswap_bias.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_ctl_i2c_fix/sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_i2c_fix_leak_fix/sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_latch/sky130_fd_io__gpio_ovtv2_hotswap_latch.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_nonoverlap_leak_fix/sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_pghs_i2c_fix/sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_pghspu/sky130_fd_io__gpio_ovtv2_hotswap_pghspu.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_pug_ovtfix/sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_pug/sky130_fd_io__gpio_ovtv2_hotswap_pug.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_vpb_bias/sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_hotswap_vpb_bias_unit/sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_ibuf_se/sky130_fd_io__gpio_ovtv2_ibuf_se.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_ictl_logic/sky130_fd_io__gpio_ovtv2_ictl_logic.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_in_buf/sky130_fd_io__gpio_ovtv2_in_buf.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_ipath_hvls/sky130_fd_io__gpio_ovtv2_ipath_hvls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_ipath_lvls/sky130_fd_io__gpio_ovtv2_ipath_lvls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_ipath/sky130_fd_io__gpio_ovtv2_ipath.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_obpredrvr_leak_fix/sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_obpredrvr_new_leak_fix/sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_obpredrvr_old/sky130_fd_io__gpio_ovtv2_obpredrvr_old.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_octl_dat_i2c_fix_leak_fix/sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_octl_i2c_fix/sky130_fd_io__gpio_ovtv2_octl_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_odrvr_i2c_fix_leak_fix/sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_odrvr_sub/sky130_fd_io__gpio_ovtv2_odrvr_sub.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_opath_datoe_i2c_fix/sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_opath_i2c_fix_leak_fix/sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pddrvr/sky130_fd_io__gpio_ovtv2_pddrvr.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pddrvr_unit/sky130_fd_io__gpio_ovtv2_pddrvr_unit.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pdpredrvr_pbias/sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pdpredrvr_strong_cmos/sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pdpredrvr_strong_leak_fix/sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pdpredrvr_strong_nr2/sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pdpredrvr_strong_nr3/sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_predrvr_switch/sky130_fd_io__gpio_ovtv2_predrvr_switch.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pudrvr_strong/sky130_fd_io__gpio_ovtv2_pudrvr_strong.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pudrvr_strong_slow/sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pudrvr_unit_2_5/sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pudrvr_weak/sky130_fd_io__gpio_ovtv2_pudrvr_weak.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pupredrvr_strong_nd2/sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pupredrvr_strong_nd3/sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_ovtv2_pupredrvr_strong/sky130_fd_io__gpio_ovtv2_pupredrvr_strong.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_pddrvr_strong/sky130_fd_io__gpio_pddrvr_strong.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_pddrvr_strong_slow/sky130_fd_io__gpio_pddrvr_strong_slow.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_pddrvr_weak/sky130_fd_io__gpio_pddrvr_weak.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_pudrvr_strong/sky130_fd_io__gpio_pudrvr_strong.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpio_pudrvr_unit_2_5/sky130_fd_io__gpio_pudrvr_unit_2_5.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ctl_inv_1/sky130_fd_io__gpiov2_amux_ctl_inv_1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ctl_logic_i2c_fix/sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ctl_logic/sky130_fd_io__gpiov2_amux_ctl_logic.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ctl_lshv2hv/sky130_fd_io__gpiov2_amux_ctl_lshv2hv.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ctl_ls_i2c_fix/sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ctl_ls/sky130_fd_io__gpiov2_amux_ctl_ls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_decoder/sky130_fd_io__gpiov2_amux_decoder.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_drvr_i2c_fix/sky130_fd_io__gpiov2_amux_drvr_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_drvr_lshv2hv/sky130_fd_io__gpiov2_amux_drvr_lshv2hv.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_drvr_ls_i2c_fix3/sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_drvr_ls_i2c_fix3_ver2/sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_drvr_ls/sky130_fd_io__gpiov2_amux_drvr_ls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_drvr/sky130_fd_io__gpiov2_amux_drvr.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ls_i2c_fix/sky130_fd_io__gpiov2_amux_ls_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ls_inv_x1/sky130_fd_io__gpiov2_amux_ls_inv_x1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_ls/sky130_fd_io__gpiov2_amux_ls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_nand4/sky130_fd_io__gpiov2_amux_nand4.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_nand5/sky130_fd_io__gpiov2_amux_nand5.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux/sky130_fd_io__gpiov2_amux.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amux_switch/sky130_fd_io__gpiov2_amux_switch.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amx_inv4/sky130_fd_io__gpiov2_amx_inv4.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amx_pdcsd_inv/sky130_fd_io__gpiov2_amx_pdcsd_inv.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amx_pucsd_buf/sky130_fd_io__gpiov2_amx_pucsd_buf.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_amx_pucsd_inv/sky130_fd_io__gpiov2_amx_pucsd_inv.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_ctl_hld/sky130_fd_io__gpiov2_ctl_hld.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_ctl_lsbank/sky130_fd_io__gpiov2_ctl_lsbank.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_ctl/sky130_fd_io__gpiov2_ctl.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_ibuf_se/sky130_fd_io__gpiov2_ibuf_se.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_ictl_logic/sky130_fd_io__gpiov2_ictl_logic.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_inbuf_lvinv_x1/sky130_fd_io__gpiov2_inbuf_lvinv_x1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_in_buf/sky130_fd_io__gpiov2_in_buf.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_ipath_hvls/sky130_fd_io__gpiov2_ipath_hvls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_ipath_lvls/sky130_fd_io__gpiov2_ipath_lvls.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_ipath/sky130_fd_io__gpiov2_ipath.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_obpredrvr/sky130_fd_io__gpiov2_obpredrvr.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_octl_dat/sky130_fd_io__gpiov2_octl_dat.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_octl_mux/sky130_fd_io__gpiov2_octl_mux.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_octl/sky130_fd_io__gpiov2_octl.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_odrvr/sky130_fd_io__gpiov2_odrvr.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_odrvr_sub/sky130_fd_io__gpiov2_odrvr_sub.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_opath_datoe/sky130_fd_io__gpiov2_opath_datoe.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_opath/sky130_fd_io__gpiov2_opath.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_pddrvr_strong/sky130_fd_io__gpiov2_pddrvr_strong.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_pdpredrvr_strong_nr2/sky130_fd_io__gpiov2_pdpredrvr_strong_nr2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_pdpredrvr_strong_nr3/sky130_fd_io__gpiov2_pdpredrvr_strong_nr3.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_pdpredrvr_strong/sky130_fd_io__gpiov2_pdpredrvr_strong.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_pupredrvr_strong_nd2/sky130_fd_io__gpiov2_pupredrvr_strong_nd2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_pupredrvr_strong/sky130_fd_io__gpiov2_pupredrvr_strong.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/gpiov2_vcchib_in_buf/sky130_fd_io__gpiov2_vcchib_in_buf.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/hvsbt_inv_x1/sky130_fd_io__hvsbt_inv_x1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/hvsbt_inv_x2/sky130_fd_io__hvsbt_inv_x2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/hvsbt_inv_x4/sky130_fd_io__hvsbt_inv_x4.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/hvsbt_inv_x8/sky130_fd_io__hvsbt_inv_x8.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/hvsbt_nand2/sky130_fd_io__hvsbt_nand2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/hvsbt_nor/sky130_fd_io__hvsbt_nor.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/hvsbt_xor/sky130_fd_io__hvsbt_xor.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/inv_1/sky130_fd_io__inv_1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/nand2_1/sky130_fd_io__nand2_1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/nand2_2_enhpath/sky130_fd_io__nand2_2_enhpath.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/nor2_1/sky130_fd_io__nor2_1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/nor2_4_enhpath/sky130_fd_io__nor2_4_enhpath.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/nor3_dnw/sky130_fd_io__nor3_dnw.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/res250only_small/sky130_fd_io__res250only_small.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/res75only_small/sky130_fd_io__res75only_small.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/signal_5_sym_hv_local_5term/sky130_fd_io__signal_5_sym_hv_local_5term.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hotswap_dly/sky130_fd_io__sio_hotswap_dly.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hotswap_hys/sky130_fd_io__sio_hotswap_hys.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hotswap_log_i2c_fix/sky130_fd_io__sio_hotswap_log_i2c_fix.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hotswap_pghspd/sky130_fd_io__sio_hotswap_pghspd.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hotswap_wpd/sky130_fd_io__sio_hotswap_wpd.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hvsbt_inv_x1/sky130_fd_io__sio_hvsbt_inv_x1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hvsbt_inv_x2/sky130_fd_io__sio_hvsbt_inv_x2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hvsbt_inv_x4/sky130_fd_io__sio_hvsbt_inv_x4.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hvsbt_nand2/sky130_fd_io__sio_hvsbt_nand2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_hvsbt_nor/sky130_fd_io__sio_hvsbt_nor.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_tk_em1o/sky130_fd_io__sio_tk_em1o.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_tk_em1s/sky130_fd_io__sio_tk_em1s.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/sio_tk_tie_r_out_esd/sky130_fd_io__sio_tk_tie_r_out_esd.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/tk_em1o/sky130_fd_io__tk_em1o.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/tk_em1s/sky130_fd_io__tk_em1s.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/tk_em2o/sky130_fd_io__tk_em2o.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/tk_em2s/sky130_fd_io__tk_em2s.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/tk_opti/sky130_fd_io__tk_opti.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/tk_opto/sky130_fd_io__tk_opto.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/tk_tie_r_out_esd/sky130_fd_io__tk_tie_r_out_esd.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/top_amuxsplitv2/sky130_fd_io__top_amuxsplitv2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/top_gpio_ovtv2/sky130_fd_io__top_gpio_ovtv2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/top_ground_hvc_wpad/sky130_fd_io__top_ground_hvc_wpad.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/top_hvclamp_wopadv2/sky130_fd_io__top_hvclamp_wopadv2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/top_power_hvc_wpadv2/sky130_fd_io__top_power_hvc_wpadv2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/top_vrefcapv2/sky130_fd_io__top_vrefcapv2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/top_xres4v2/sky130_fd_io__top_xres4v2.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xor2_1/sky130_fd_io__xor2_1.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres4v2_in_buf/sky130_fd_io__xres4v2_in_buf.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres_esd/sky130_fd_io__xres_esd.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres_inv_hys/sky130_fd_io__xres_inv_hys.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres_rcfilter_lpf_rcunit/sky130_fd_io__xres_rcfilter_lpf_rcunit.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres_rcfilter_lpf_res_sub/sky130_fd_io__xres_rcfilter_lpf_res_sub.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres_rcfilter_lpf/sky130_fd_io__xres_rcfilter_lpf.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres_tk_emlc/sky130_fd_io__xres_tk_emlc.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres_tk_emlo/sky130_fd_io__xres_tk_emlo.spice
.include ../../../../../../pdks/skywater-pdk-scratch/libraries/sky130_fd_io/v0.2.1/cells/xres_wpu/sky130_fd_io__xres_wpu.spice
