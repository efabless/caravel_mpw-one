* NGSPICE file created from mprj_logic_high.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[46] HI[47]
+ HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57] HI[58]
+ HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68] HI[69]
+ HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79] HI[7]
+ HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8] HI[90]
+ HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1 vssd1
Xinsts\[308\] vssd1 vssd1 vccd1 vccd1 HI[308] insts\[308\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[210\] vssd1 vssd1 vccd1 vccd1 HI[210] insts\[210\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[425\] vssd1 vssd1 vccd1 vccd1 HI[425] insts\[425\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[258\] vssd1 vssd1 vccd1 vccd1 HI[258] insts\[258\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[160\] vssd1 vssd1 vccd1 vccd1 HI[160] insts\[160\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[40\] vssd1 vssd1 vccd1 vccd1 HI[40] insts\[40\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[375\] vssd1 vssd1 vccd1 vccd1 HI[375] insts\[375\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[88\] vssd1 vssd1 vccd1 vccd1 HI[88] insts\[88\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[123\] vssd1 vssd1 vccd1 vccd1 HI[123] insts\[123\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[240\] vssd1 vssd1 vccd1 vccd1 HI[240] insts\[240\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[338\] vssd1 vssd1 vccd1 vccd1 HI[338] insts\[338\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[9\] vssd1 vssd1 vccd1 vccd1 HI[9] insts\[9\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[455\] vssd1 vssd1 vccd1 vccd1 HI[455] insts\[455\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[288\] vssd1 vssd1 vccd1 vccd1 HI[288] insts\[288\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[190\] vssd1 vssd1 vccd1 vccd1 HI[190] insts\[190\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[70\] vssd1 vssd1 vccd1 vccd1 HI[70] insts\[70\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[203\] vssd1 vssd1 vccd1 vccd1 HI[203] insts\[203\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[418\] vssd1 vssd1 vccd1 vccd1 HI[418] insts\[418\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[153\] vssd1 vssd1 vccd1 vccd1 HI[153] insts\[153\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[320\] vssd1 vssd1 vccd1 vccd1 HI[320] insts\[320\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[33\] vssd1 vssd1 vccd1 vccd1 HI[33] insts\[33\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[270\] vssd1 vssd1 vccd1 vccd1 HI[270] insts\[270\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[368\] vssd1 vssd1 vccd1 vccd1 HI[368] insts\[368\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[116\] vssd1 vssd1 vccd1 vccd1 HI[116] insts\[116\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[233\] vssd1 vssd1 vccd1 vccd1 HI[233] insts\[233\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[400\] vssd1 vssd1 vccd1 vccd1 HI[400] insts\[400\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[183\] vssd1 vssd1 vccd1 vccd1 HI[183] insts\[183\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[448\] vssd1 vssd1 vccd1 vccd1 HI[448] insts\[448\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[350\] vssd1 vssd1 vccd1 vccd1 HI[350] insts\[350\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[63\] vssd1 vssd1 vccd1 vccd1 HI[63] insts\[63\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[398\] vssd1 vssd1 vccd1 vccd1 HI[398] insts\[398\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[146\] vssd1 vssd1 vccd1 vccd1 HI[146] insts\[146\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[313\] vssd1 vssd1 vccd1 vccd1 HI[313] insts\[313\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[26\] vssd1 vssd1 vccd1 vccd1 HI[26] insts\[26\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[430\] vssd1 vssd1 vccd1 vccd1 HI[430] insts\[430\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[263\] vssd1 vssd1 vccd1 vccd1 HI[263] insts\[263\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[109\] vssd1 vssd1 vccd1 vccd1 HI[109] insts\[109\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[380\] vssd1 vssd1 vccd1 vccd1 HI[380] insts\[380\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[93\] vssd1 vssd1 vccd1 vccd1 HI[93] insts\[93\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[226\] vssd1 vssd1 vccd1 vccd1 HI[226] insts\[226\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[343\] vssd1 vssd1 vccd1 vccd1 HI[343] insts\[343\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[176\] vssd1 vssd1 vccd1 vccd1 HI[176] insts\[176\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[56\] vssd1 vssd1 vccd1 vccd1 HI[56] insts\[56\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[460\] vssd1 vssd1 vccd1 vccd1 HI[460] insts\[460\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[293\] vssd1 vssd1 vccd1 vccd1 HI[293] insts\[293\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[139\] vssd1 vssd1 vccd1 vccd1 HI[139] insts\[139\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[306\] vssd1 vssd1 vccd1 vccd1 HI[306] insts\[306\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[19\] vssd1 vssd1 vccd1 vccd1 HI[19] insts\[19\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[423\] vssd1 vssd1 vccd1 vccd1 HI[423] insts\[423\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[256\] vssd1 vssd1 vccd1 vccd1 HI[256] insts\[256\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[373\] vssd1 vssd1 vccd1 vccd1 HI[373] insts\[373\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[86\] vssd1 vssd1 vccd1 vccd1 HI[86] insts\[86\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[219\] vssd1 vssd1 vccd1 vccd1 HI[219] insts\[219\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[121\] vssd1 vssd1 vccd1 vccd1 HI[121] insts\[121\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[336\] vssd1 vssd1 vccd1 vccd1 HI[336] insts\[336\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[169\] vssd1 vssd1 vccd1 vccd1 HI[169] insts\[169\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[49\] vssd1 vssd1 vccd1 vccd1 HI[49] insts\[49\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[286\] vssd1 vssd1 vccd1 vccd1 HI[286] insts\[286\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[7\] vssd1 vssd1 vccd1 vccd1 HI[7] insts\[7\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[453\] vssd1 vssd1 vccd1 vccd1 HI[453] insts\[453\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[201\] vssd1 vssd1 vccd1 vccd1 HI[201] insts\[201\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[416\] vssd1 vssd1 vccd1 vccd1 HI[416] insts\[416\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[249\] vssd1 vssd1 vccd1 vccd1 HI[249] insts\[249\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[151\] vssd1 vssd1 vccd1 vccd1 HI[151] insts\[151\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[31\] vssd1 vssd1 vccd1 vccd1 HI[31] insts\[31\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[199\] vssd1 vssd1 vccd1 vccd1 HI[199] insts\[199\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[366\] vssd1 vssd1 vccd1 vccd1 HI[366] insts\[366\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[79\] vssd1 vssd1 vccd1 vccd1 HI[79] insts\[79\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[114\] vssd1 vssd1 vccd1 vccd1 HI[114] insts\[114\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[231\] vssd1 vssd1 vccd1 vccd1 HI[231] insts\[231\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[329\] vssd1 vssd1 vccd1 vccd1 HI[329] insts\[329\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[446\] vssd1 vssd1 vccd1 vccd1 HI[446] insts\[446\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[279\] vssd1 vssd1 vccd1 vccd1 HI[279] insts\[279\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[181\] vssd1 vssd1 vccd1 vccd1 HI[181] insts\[181\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[61\] vssd1 vssd1 vccd1 vccd1 HI[61] insts\[61\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[396\] vssd1 vssd1 vccd1 vccd1 HI[396] insts\[396\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[144\] vssd1 vssd1 vccd1 vccd1 HI[144] insts\[144\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[311\] vssd1 vssd1 vccd1 vccd1 HI[311] insts\[311\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[409\] vssd1 vssd1 vccd1 vccd1 HI[409] insts\[409\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[24\] vssd1 vssd1 vccd1 vccd1 HI[24] insts\[24\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[261\] vssd1 vssd1 vccd1 vccd1 HI[261] insts\[261\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[359\] vssd1 vssd1 vccd1 vccd1 HI[359] insts\[359\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[107\] vssd1 vssd1 vccd1 vccd1 HI[107] insts\[107\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[91\] vssd1 vssd1 vccd1 vccd1 HI[91] insts\[91\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[224\] vssd1 vssd1 vccd1 vccd1 HI[224] insts\[224\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[439\] vssd1 vssd1 vccd1 vccd1 HI[439] insts\[439\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[174\] vssd1 vssd1 vccd1 vccd1 HI[174] insts\[174\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[341\] vssd1 vssd1 vccd1 vccd1 HI[341] insts\[341\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[54\] vssd1 vssd1 vccd1 vccd1 HI[54] insts\[54\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[291\] vssd1 vssd1 vccd1 vccd1 HI[291] insts\[291\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[389\] vssd1 vssd1 vccd1 vccd1 HI[389] insts\[389\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[304\] vssd1 vssd1 vccd1 vccd1 HI[304] insts\[304\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[137\] vssd1 vssd1 vccd1 vccd1 HI[137] insts\[137\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[17\] vssd1 vssd1 vccd1 vccd1 HI[17] insts\[17\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[421\] vssd1 vssd1 vccd1 vccd1 HI[421] insts\[421\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[254\] vssd1 vssd1 vccd1 vccd1 HI[254] insts\[254\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[371\] vssd1 vssd1 vccd1 vccd1 HI[371] insts\[371\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[84\] vssd1 vssd1 vccd1 vccd1 HI[84] insts\[84\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[217\] vssd1 vssd1 vccd1 vccd1 HI[217] insts\[217\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[167\] vssd1 vssd1 vccd1 vccd1 HI[167] insts\[167\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[334\] vssd1 vssd1 vccd1 vccd1 HI[334] insts\[334\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[47\] vssd1 vssd1 vccd1 vccd1 HI[47] insts\[47\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[5\] vssd1 vssd1 vccd1 vccd1 HI[5] insts\[5\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[451\] vssd1 vssd1 vccd1 vccd1 HI[451] insts\[451\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[284\] vssd1 vssd1 vccd1 vccd1 HI[284] insts\[284\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[247\] vssd1 vssd1 vccd1 vccd1 HI[247] insts\[247\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[414\] vssd1 vssd1 vccd1 vccd1 HI[414] insts\[414\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[197\] vssd1 vssd1 vccd1 vccd1 HI[197] insts\[197\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[364\] vssd1 vssd1 vccd1 vccd1 HI[364] insts\[364\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[77\] vssd1 vssd1 vccd1 vccd1 HI[77] insts\[77\]/LO sky130_fd_sc_hd__conb_1
XPHY_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[112\] vssd1 vssd1 vccd1 vccd1 HI[112] insts\[112\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[327\] vssd1 vssd1 vccd1 vccd1 HI[327] insts\[327\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[444\] vssd1 vssd1 vccd1 vccd1 HI[444] insts\[444\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[277\] vssd1 vssd1 vccd1 vccd1 HI[277] insts\[277\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[394\] vssd1 vssd1 vccd1 vccd1 HI[394] insts\[394\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[407\] vssd1 vssd1 vccd1 vccd1 HI[407] insts\[407\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[142\] vssd1 vssd1 vccd1 vccd1 HI[142] insts\[142\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[22\] vssd1 vssd1 vccd1 vccd1 HI[22] insts\[22\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[357\] vssd1 vssd1 vccd1 vccd1 HI[357] insts\[357\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[105\] vssd1 vssd1 vccd1 vccd1 HI[105] insts\[105\]/LO sky130_fd_sc_hd__conb_1
XPHY_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[222\] vssd1 vssd1 vccd1 vccd1 HI[222] insts\[222\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[437\] vssd1 vssd1 vccd1 vccd1 HI[437] insts\[437\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[172\] vssd1 vssd1 vccd1 vccd1 HI[172] insts\[172\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[52\] vssd1 vssd1 vccd1 vccd1 HI[52] insts\[52\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[387\] vssd1 vssd1 vccd1 vccd1 HI[387] insts\[387\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[302\] vssd1 vssd1 vccd1 vccd1 HI[302] insts\[302\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[135\] vssd1 vssd1 vccd1 vccd1 HI[135] insts\[135\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[15\] vssd1 vssd1 vccd1 vccd1 HI[15] insts\[15\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[252\] vssd1 vssd1 vccd1 vccd1 HI[252] insts\[252\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[82\] vssd1 vssd1 vccd1 vccd1 HI[82] insts\[82\]/LO sky130_fd_sc_hd__conb_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[215\] vssd1 vssd1 vccd1 vccd1 HI[215] insts\[215\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[165\] vssd1 vssd1 vccd1 vccd1 HI[165] insts\[165\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[332\] vssd1 vssd1 vccd1 vccd1 HI[332] insts\[332\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[45\] vssd1 vssd1 vccd1 vccd1 HI[45] insts\[45\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[282\] vssd1 vssd1 vccd1 vccd1 HI[282] insts\[282\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[3\] vssd1 vssd1 vccd1 vccd1 HI[3] insts\[3\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[128\] vssd1 vssd1 vccd1 vccd1 HI[128] insts\[128\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[245\] vssd1 vssd1 vccd1 vccd1 HI[245] insts\[245\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[412\] vssd1 vssd1 vccd1 vccd1 HI[412] insts\[412\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[195\] vssd1 vssd1 vccd1 vccd1 HI[195] insts\[195\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[362\] vssd1 vssd1 vccd1 vccd1 HI[362] insts\[362\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[75\] vssd1 vssd1 vccd1 vccd1 HI[75] insts\[75\]/LO sky130_fd_sc_hd__conb_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[208\] vssd1 vssd1 vccd1 vccd1 HI[208] insts\[208\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[110\] vssd1 vssd1 vccd1 vccd1 HI[110] insts\[110\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[158\] vssd1 vssd1 vccd1 vccd1 HI[158] insts\[158\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[325\] vssd1 vssd1 vccd1 vccd1 HI[325] insts\[325\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[38\] vssd1 vssd1 vccd1 vccd1 HI[38] insts\[38\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[442\] vssd1 vssd1 vccd1 vccd1 HI[442] insts\[442\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[275\] vssd1 vssd1 vccd1 vccd1 HI[275] insts\[275\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[392\] vssd1 vssd1 vccd1 vccd1 HI[392] insts\[392\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[238\] vssd1 vssd1 vccd1 vccd1 HI[238] insts\[238\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[140\] vssd1 vssd1 vccd1 vccd1 HI[140] insts\[140\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[405\] vssd1 vssd1 vccd1 vccd1 HI[405] insts\[405\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[20\] vssd1 vssd1 vccd1 vccd1 HI[20] insts\[20\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[188\] vssd1 vssd1 vccd1 vccd1 HI[188] insts\[188\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[355\] vssd1 vssd1 vccd1 vccd1 HI[355] insts\[355\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[68\] vssd1 vssd1 vccd1 vccd1 HI[68] insts\[68\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[103\] vssd1 vssd1 vccd1 vccd1 HI[103] insts\[103\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[220\] vssd1 vssd1 vccd1 vccd1 HI[220] insts\[220\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[318\] vssd1 vssd1 vccd1 vccd1 HI[318] insts\[318\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[170\] vssd1 vssd1 vccd1 vccd1 HI[170] insts\[170\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[435\] vssd1 vssd1 vccd1 vccd1 HI[435] insts\[435\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[268\] vssd1 vssd1 vccd1 vccd1 HI[268] insts\[268\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[50\] vssd1 vssd1 vccd1 vccd1 HI[50] insts\[50\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[385\] vssd1 vssd1 vccd1 vccd1 HI[385] insts\[385\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[98\] vssd1 vssd1 vccd1 vccd1 HI[98] insts\[98\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[300\] vssd1 vssd1 vccd1 vccd1 HI[300] insts\[300\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[133\] vssd1 vssd1 vccd1 vccd1 HI[133] insts\[133\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[13\] vssd1 vssd1 vccd1 vccd1 HI[13] insts\[13\]/LO sky130_fd_sc_hd__conb_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[250\] vssd1 vssd1 vccd1 vccd1 HI[250] insts\[250\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[348\] vssd1 vssd1 vccd1 vccd1 HI[348] insts\[348\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[298\] vssd1 vssd1 vccd1 vccd1 HI[298] insts\[298\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[80\] vssd1 vssd1 vccd1 vccd1 HI[80] insts\[80\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[213\] vssd1 vssd1 vccd1 vccd1 HI[213] insts\[213\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[428\] vssd1 vssd1 vccd1 vccd1 HI[428] insts\[428\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[163\] vssd1 vssd1 vccd1 vccd1 HI[163] insts\[163\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[330\] vssd1 vssd1 vccd1 vccd1 HI[330] insts\[330\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[43\] vssd1 vssd1 vccd1 vccd1 HI[43] insts\[43\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[280\] vssd1 vssd1 vccd1 vccd1 HI[280] insts\[280\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[1\] vssd1 vssd1 vccd1 vccd1 HI[1] insts\[1\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[378\] vssd1 vssd1 vccd1 vccd1 HI[378] insts\[378\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[126\] vssd1 vssd1 vccd1 vccd1 HI[126] insts\[126\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[243\] vssd1 vssd1 vccd1 vccd1 HI[243] insts\[243\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[410\] vssd1 vssd1 vccd1 vccd1 HI[410] insts\[410\]/LO sky130_fd_sc_hd__conb_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[458\] vssd1 vssd1 vccd1 vccd1 HI[458] insts\[458\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[193\] vssd1 vssd1 vccd1 vccd1 HI[193] insts\[193\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[360\] vssd1 vssd1 vccd1 vccd1 HI[360] insts\[360\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[73\] vssd1 vssd1 vccd1 vccd1 HI[73] insts\[73\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[206\] vssd1 vssd1 vccd1 vccd1 HI[206] insts\[206\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[156\] vssd1 vssd1 vccd1 vccd1 HI[156] insts\[156\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[323\] vssd1 vssd1 vccd1 vccd1 HI[323] insts\[323\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[36\] vssd1 vssd1 vccd1 vccd1 HI[36] insts\[36\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[273\] vssd1 vssd1 vccd1 vccd1 HI[273] insts\[273\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[440\] vssd1 vssd1 vccd1 vccd1 HI[440] insts\[440\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[119\] vssd1 vssd1 vccd1 vccd1 HI[119] insts\[119\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[390\] vssd1 vssd1 vccd1 vccd1 HI[390] insts\[390\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[236\] vssd1 vssd1 vccd1 vccd1 HI[236] insts\[236\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[403\] vssd1 vssd1 vccd1 vccd1 HI[403] insts\[403\]/LO sky130_fd_sc_hd__conb_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[353\] vssd1 vssd1 vccd1 vccd1 HI[353] insts\[353\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[186\] vssd1 vssd1 vccd1 vccd1 HI[186] insts\[186\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[66\] vssd1 vssd1 vccd1 vccd1 HI[66] insts\[66\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[101\] vssd1 vssd1 vccd1 vccd1 HI[101] insts\[101\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[316\] vssd1 vssd1 vccd1 vccd1 HI[316] insts\[316\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[149\] vssd1 vssd1 vccd1 vccd1 HI[149] insts\[149\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[29\] vssd1 vssd1 vccd1 vccd1 HI[29] insts\[29\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[433\] vssd1 vssd1 vccd1 vccd1 HI[433] insts\[433\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[266\] vssd1 vssd1 vccd1 vccd1 HI[266] insts\[266\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[383\] vssd1 vssd1 vccd1 vccd1 HI[383] insts\[383\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[96\] vssd1 vssd1 vccd1 vccd1 HI[96] insts\[96\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[229\] vssd1 vssd1 vccd1 vccd1 HI[229] insts\[229\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[131\] vssd1 vssd1 vccd1 vccd1 HI[131] insts\[131\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[11\] vssd1 vssd1 vccd1 vccd1 HI[11] insts\[11\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[179\] vssd1 vssd1 vccd1 vccd1 HI[179] insts\[179\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[346\] vssd1 vssd1 vccd1 vccd1 HI[346] insts\[346\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[59\] vssd1 vssd1 vccd1 vccd1 HI[59] insts\[59\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[296\] vssd1 vssd1 vccd1 vccd1 HI[296] insts\[296\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[211\] vssd1 vssd1 vccd1 vccd1 HI[211] insts\[211\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[309\] vssd1 vssd1 vccd1 vccd1 HI[309] insts\[309\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[426\] vssd1 vssd1 vccd1 vccd1 HI[426] insts\[426\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[259\] vssd1 vssd1 vccd1 vccd1 HI[259] insts\[259\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[161\] vssd1 vssd1 vccd1 vccd1 HI[161] insts\[161\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[41\] vssd1 vssd1 vccd1 vccd1 HI[41] insts\[41\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[376\] vssd1 vssd1 vccd1 vccd1 HI[376] insts\[376\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[89\] vssd1 vssd1 vccd1 vccd1 HI[89] insts\[89\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[124\] vssd1 vssd1 vccd1 vccd1 HI[124] insts\[124\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[241\] vssd1 vssd1 vccd1 vccd1 HI[241] insts\[241\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[339\] vssd1 vssd1 vccd1 vccd1 HI[339] insts\[339\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[456\] vssd1 vssd1 vccd1 vccd1 HI[456] insts\[456\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[289\] vssd1 vssd1 vccd1 vccd1 HI[289] insts\[289\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[191\] vssd1 vssd1 vccd1 vccd1 HI[191] insts\[191\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[71\] vssd1 vssd1 vccd1 vccd1 HI[71] insts\[71\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[204\] vssd1 vssd1 vccd1 vccd1 HI[204] insts\[204\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[419\] vssd1 vssd1 vccd1 vccd1 HI[419] insts\[419\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[154\] vssd1 vssd1 vccd1 vccd1 HI[154] insts\[154\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[321\] vssd1 vssd1 vccd1 vccd1 HI[321] insts\[321\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[34\] vssd1 vssd1 vccd1 vccd1 HI[34] insts\[34\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[271\] vssd1 vssd1 vccd1 vccd1 HI[271] insts\[271\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[369\] vssd1 vssd1 vccd1 vccd1 HI[369] insts\[369\]/LO sky130_fd_sc_hd__conb_1
XPHY_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[117\] vssd1 vssd1 vccd1 vccd1 HI[117] insts\[117\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[234\] vssd1 vssd1 vccd1 vccd1 HI[234] insts\[234\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[401\] vssd1 vssd1 vccd1 vccd1 HI[401] insts\[401\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[449\] vssd1 vssd1 vccd1 vccd1 HI[449] insts\[449\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[184\] vssd1 vssd1 vccd1 vccd1 HI[184] insts\[184\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[351\] vssd1 vssd1 vccd1 vccd1 HI[351] insts\[351\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[64\] vssd1 vssd1 vccd1 vccd1 HI[64] insts\[64\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[399\] vssd1 vssd1 vccd1 vccd1 HI[399] insts\[399\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[314\] vssd1 vssd1 vccd1 vccd1 HI[314] insts\[314\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[147\] vssd1 vssd1 vccd1 vccd1 HI[147] insts\[147\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[27\] vssd1 vssd1 vccd1 vccd1 HI[27] insts\[27\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[431\] vssd1 vssd1 vccd1 vccd1 HI[431] insts\[431\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[264\] vssd1 vssd1 vccd1 vccd1 HI[264] insts\[264\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[381\] vssd1 vssd1 vccd1 vccd1 HI[381] insts\[381\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[94\] vssd1 vssd1 vccd1 vccd1 HI[94] insts\[94\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[227\] vssd1 vssd1 vccd1 vccd1 HI[227] insts\[227\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[177\] vssd1 vssd1 vccd1 vccd1 HI[177] insts\[177\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[344\] vssd1 vssd1 vccd1 vccd1 HI[344] insts\[344\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[57\] vssd1 vssd1 vccd1 vccd1 HI[57] insts\[57\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[461\] vssd1 vssd1 vccd1 vccd1 HI[461] insts\[461\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[294\] vssd1 vssd1 vccd1 vccd1 HI[294] insts\[294\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[307\] vssd1 vssd1 vccd1 vccd1 HI[307] insts\[307\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[424\] vssd1 vssd1 vccd1 vccd1 HI[424] insts\[424\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[257\] vssd1 vssd1 vccd1 vccd1 HI[257] insts\[257\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[374\] vssd1 vssd1 vccd1 vccd1 HI[374] insts\[374\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[87\] vssd1 vssd1 vccd1 vccd1 HI[87] insts\[87\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[122\] vssd1 vssd1 vccd1 vccd1 HI[122] insts\[122\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[337\] vssd1 vssd1 vccd1 vccd1 HI[337] insts\[337\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[8\] vssd1 vssd1 vccd1 vccd1 HI[8] insts\[8\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[454\] vssd1 vssd1 vccd1 vccd1 HI[454] insts\[454\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[287\] vssd1 vssd1 vccd1 vccd1 HI[287] insts\[287\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[202\] vssd1 vssd1 vccd1 vccd1 HI[202] insts\[202\]/LO sky130_fd_sc_hd__conb_1
XPHY_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[417\] vssd1 vssd1 vccd1 vccd1 HI[417] insts\[417\]/LO sky130_fd_sc_hd__conb_1
XPHY_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[152\] vssd1 vssd1 vccd1 vccd1 HI[152] insts\[152\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[32\] vssd1 vssd1 vccd1 vccd1 HI[32] insts\[32\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[367\] vssd1 vssd1 vccd1 vccd1 HI[367] insts\[367\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[115\] vssd1 vssd1 vccd1 vccd1 HI[115] insts\[115\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[232\] vssd1 vssd1 vccd1 vccd1 HI[232] insts\[232\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[447\] vssd1 vssd1 vccd1 vccd1 HI[447] insts\[447\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[182\] vssd1 vssd1 vccd1 vccd1 HI[182] insts\[182\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[62\] vssd1 vssd1 vccd1 vccd1 HI[62] insts\[62\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[397\] vssd1 vssd1 vccd1 vccd1 HI[397] insts\[397\]/LO sky130_fd_sc_hd__conb_1
XPHY_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[145\] vssd1 vssd1 vccd1 vccd1 HI[145] insts\[145\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[312\] vssd1 vssd1 vccd1 vccd1 HI[312] insts\[312\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[25\] vssd1 vssd1 vccd1 vccd1 HI[25] insts\[25\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[262\] vssd1 vssd1 vccd1 vccd1 HI[262] insts\[262\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[108\] vssd1 vssd1 vccd1 vccd1 HI[108] insts\[108\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[92\] vssd1 vssd1 vccd1 vccd1 HI[92] insts\[92\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[225\] vssd1 vssd1 vccd1 vccd1 HI[225] insts\[225\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[175\] vssd1 vssd1 vccd1 vccd1 HI[175] insts\[175\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[342\] vssd1 vssd1 vccd1 vccd1 HI[342] insts\[342\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[55\] vssd1 vssd1 vccd1 vccd1 HI[55] insts\[55\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[292\] vssd1 vssd1 vccd1 vccd1 HI[292] insts\[292\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[305\] vssd1 vssd1 vccd1 vccd1 HI[305] insts\[305\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[138\] vssd1 vssd1 vccd1 vccd1 HI[138] insts\[138\]/LO sky130_fd_sc_hd__conb_1
XPHY_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_51 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[18\] vssd1 vssd1 vccd1 vccd1 HI[18] insts\[18\]/LO sky130_fd_sc_hd__conb_1
XPHY_40 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[422\] vssd1 vssd1 vccd1 vccd1 HI[422] insts\[422\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[255\] vssd1 vssd1 vccd1 vccd1 HI[255] insts\[255\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[372\] vssd1 vssd1 vccd1 vccd1 HI[372] insts\[372\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[85\] vssd1 vssd1 vccd1 vccd1 HI[85] insts\[85\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[218\] vssd1 vssd1 vccd1 vccd1 HI[218] insts\[218\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[120\] vssd1 vssd1 vccd1 vccd1 HI[120] insts\[120\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[168\] vssd1 vssd1 vccd1 vccd1 HI[168] insts\[168\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[335\] vssd1 vssd1 vccd1 vccd1 HI[335] insts\[335\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[48\] vssd1 vssd1 vccd1 vccd1 HI[48] insts\[48\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[6\] vssd1 vssd1 vccd1 vccd1 HI[6] insts\[6\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[452\] vssd1 vssd1 vccd1 vccd1 HI[452] insts\[452\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[285\] vssd1 vssd1 vccd1 vccd1 HI[285] insts\[285\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[200\] vssd1 vssd1 vccd1 vccd1 HI[200] insts\[200\]/LO sky130_fd_sc_hd__conb_1
XPHY_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_52 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[415\] vssd1 vssd1 vccd1 vccd1 HI[415] insts\[415\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[248\] vssd1 vssd1 vccd1 vccd1 HI[248] insts\[248\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[150\] vssd1 vssd1 vccd1 vccd1 HI[150] insts\[150\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[30\] vssd1 vssd1 vccd1 vccd1 HI[30] insts\[30\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[198\] vssd1 vssd1 vccd1 vccd1 HI[198] insts\[198\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[365\] vssd1 vssd1 vccd1 vccd1 HI[365] insts\[365\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[78\] vssd1 vssd1 vccd1 vccd1 HI[78] insts\[78\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[113\] vssd1 vssd1 vccd1 vccd1 HI[113] insts\[113\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[230\] vssd1 vssd1 vccd1 vccd1 HI[230] insts\[230\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[328\] vssd1 vssd1 vccd1 vccd1 HI[328] insts\[328\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[445\] vssd1 vssd1 vccd1 vccd1 HI[445] insts\[445\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[278\] vssd1 vssd1 vccd1 vccd1 HI[278] insts\[278\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[180\] vssd1 vssd1 vccd1 vccd1 HI[180] insts\[180\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[60\] vssd1 vssd1 vccd1 vccd1 HI[60] insts\[60\]/LO sky130_fd_sc_hd__conb_1
XPHY_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[395\] vssd1 vssd1 vccd1 vccd1 HI[395] insts\[395\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[310\] vssd1 vssd1 vccd1 vccd1 HI[310] insts\[310\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[143\] vssd1 vssd1 vccd1 vccd1 HI[143] insts\[143\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[408\] vssd1 vssd1 vccd1 vccd1 HI[408] insts\[408\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[23\] vssd1 vssd1 vccd1 vccd1 HI[23] insts\[23\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[260\] vssd1 vssd1 vccd1 vccd1 HI[260] insts\[260\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[358\] vssd1 vssd1 vccd1 vccd1 HI[358] insts\[358\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[106\] vssd1 vssd1 vccd1 vccd1 HI[106] insts\[106\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[90\] vssd1 vssd1 vccd1 vccd1 HI[90] insts\[90\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[223\] vssd1 vssd1 vccd1 vccd1 HI[223] insts\[223\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[438\] vssd1 vssd1 vccd1 vccd1 HI[438] insts\[438\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[173\] vssd1 vssd1 vccd1 vccd1 HI[173] insts\[173\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[340\] vssd1 vssd1 vccd1 vccd1 HI[340] insts\[340\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[53\] vssd1 vssd1 vccd1 vccd1 HI[53] insts\[53\]/LO sky130_fd_sc_hd__conb_1
XPHY_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[290\] vssd1 vssd1 vccd1 vccd1 HI[290] insts\[290\]/LO sky130_fd_sc_hd__conb_1
XPHY_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[388\] vssd1 vssd1 vccd1 vccd1 HI[388] insts\[388\]/LO sky130_fd_sc_hd__conb_1
XPHY_32 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[303\] vssd1 vssd1 vccd1 vccd1 HI[303] insts\[303\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[136\] vssd1 vssd1 vccd1 vccd1 HI[136] insts\[136\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[16\] vssd1 vssd1 vccd1 vccd1 HI[16] insts\[16\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[420\] vssd1 vssd1 vccd1 vccd1 HI[420] insts\[420\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[253\] vssd1 vssd1 vccd1 vccd1 HI[253] insts\[253\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[370\] vssd1 vssd1 vccd1 vccd1 HI[370] insts\[370\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[83\] vssd1 vssd1 vccd1 vccd1 HI[83] insts\[83\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[216\] vssd1 vssd1 vccd1 vccd1 HI[216] insts\[216\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[166\] vssd1 vssd1 vccd1 vccd1 HI[166] insts\[166\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[333\] vssd1 vssd1 vccd1 vccd1 HI[333] insts\[333\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[46\] vssd1 vssd1 vccd1 vccd1 HI[46] insts\[46\]/LO sky130_fd_sc_hd__conb_1
XPHY_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[450\] vssd1 vssd1 vccd1 vccd1 HI[450] insts\[450\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[283\] vssd1 vssd1 vccd1 vccd1 HI[283] insts\[283\]/LO sky130_fd_sc_hd__conb_1
XPHY_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[4\] vssd1 vssd1 vccd1 vccd1 HI[4] insts\[4\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[129\] vssd1 vssd1 vccd1 vccd1 HI[129] insts\[129\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[413\] vssd1 vssd1 vccd1 vccd1 HI[413] insts\[413\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[246\] vssd1 vssd1 vccd1 vccd1 HI[246] insts\[246\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[196\] vssd1 vssd1 vccd1 vccd1 HI[196] insts\[196\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[363\] vssd1 vssd1 vccd1 vccd1 HI[363] insts\[363\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[76\] vssd1 vssd1 vccd1 vccd1 HI[76] insts\[76\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[209\] vssd1 vssd1 vccd1 vccd1 HI[209] insts\[209\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[111\] vssd1 vssd1 vccd1 vccd1 HI[111] insts\[111\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[159\] vssd1 vssd1 vccd1 vccd1 HI[159] insts\[159\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[326\] vssd1 vssd1 vccd1 vccd1 HI[326] insts\[326\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[39\] vssd1 vssd1 vccd1 vccd1 HI[39] insts\[39\]/LO sky130_fd_sc_hd__conb_1
XPHY_12 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[443\] vssd1 vssd1 vccd1 vccd1 HI[443] insts\[443\]/LO sky130_fd_sc_hd__conb_1
XPHY_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[276\] vssd1 vssd1 vccd1 vccd1 HI[276] insts\[276\]/LO sky130_fd_sc_hd__conb_1
XPHY_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_23 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[393\] vssd1 vssd1 vccd1 vccd1 HI[393] insts\[393\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[239\] vssd1 vssd1 vccd1 vccd1 HI[239] insts\[239\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[141\] vssd1 vssd1 vccd1 vccd1 HI[141] insts\[141\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[406\] vssd1 vssd1 vccd1 vccd1 HI[406] insts\[406\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[21\] vssd1 vssd1 vccd1 vccd1 HI[21] insts\[21\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[189\] vssd1 vssd1 vccd1 vccd1 HI[189] insts\[189\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[356\] vssd1 vssd1 vccd1 vccd1 HI[356] insts\[356\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[69\] vssd1 vssd1 vccd1 vccd1 HI[69] insts\[69\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[104\] vssd1 vssd1 vccd1 vccd1 HI[104] insts\[104\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[221\] vssd1 vssd1 vccd1 vccd1 HI[221] insts\[221\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[319\] vssd1 vssd1 vccd1 vccd1 HI[319] insts\[319\]/LO sky130_fd_sc_hd__conb_1
XPHY_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[436\] vssd1 vssd1 vccd1 vccd1 HI[436] insts\[436\]/LO sky130_fd_sc_hd__conb_1
XPHY_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[269\] vssd1 vssd1 vccd1 vccd1 HI[269] insts\[269\]/LO sky130_fd_sc_hd__conb_1
XPHY_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[171\] vssd1 vssd1 vccd1 vccd1 HI[171] insts\[171\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[51\] vssd1 vssd1 vccd1 vccd1 HI[51] insts\[51\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[386\] vssd1 vssd1 vccd1 vccd1 HI[386] insts\[386\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[99\] vssd1 vssd1 vccd1 vccd1 HI[99] insts\[99\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[301\] vssd1 vssd1 vccd1 vccd1 HI[301] insts\[301\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[134\] vssd1 vssd1 vccd1 vccd1 HI[134] insts\[134\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[14\] vssd1 vssd1 vccd1 vccd1 HI[14] insts\[14\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[251\] vssd1 vssd1 vccd1 vccd1 HI[251] insts\[251\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[349\] vssd1 vssd1 vccd1 vccd1 HI[349] insts\[349\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[299\] vssd1 vssd1 vccd1 vccd1 HI[299] insts\[299\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[81\] vssd1 vssd1 vccd1 vccd1 HI[81] insts\[81\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[214\] vssd1 vssd1 vccd1 vccd1 HI[214] insts\[214\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[429\] vssd1 vssd1 vccd1 vccd1 HI[429] insts\[429\]/LO sky130_fd_sc_hd__conb_1
XPHY_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[164\] vssd1 vssd1 vccd1 vccd1 HI[164] insts\[164\]/LO sky130_fd_sc_hd__conb_1
XPHY_25 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[331\] vssd1 vssd1 vccd1 vccd1 HI[331] insts\[331\]/LO sky130_fd_sc_hd__conb_1
XPHY_47 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[44\] vssd1 vssd1 vccd1 vccd1 HI[44] insts\[44\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[2\] vssd1 vssd1 vccd1 vccd1 HI[2] insts\[2\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[281\] vssd1 vssd1 vccd1 vccd1 HI[281] insts\[281\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[379\] vssd1 vssd1 vccd1 vccd1 HI[379] insts\[379\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[127\] vssd1 vssd1 vccd1 vccd1 HI[127] insts\[127\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[244\] vssd1 vssd1 vccd1 vccd1 HI[244] insts\[244\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[411\] vssd1 vssd1 vccd1 vccd1 HI[411] insts\[411\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[459\] vssd1 vssd1 vccd1 vccd1 HI[459] insts\[459\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[194\] vssd1 vssd1 vccd1 vccd1 HI[194] insts\[194\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[361\] vssd1 vssd1 vccd1 vccd1 HI[361] insts\[361\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[74\] vssd1 vssd1 vccd1 vccd1 HI[74] insts\[74\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[207\] vssd1 vssd1 vccd1 vccd1 HI[207] insts\[207\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[157\] vssd1 vssd1 vccd1 vccd1 HI[157] insts\[157\]/LO sky130_fd_sc_hd__conb_1
XPHY_15 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[324\] vssd1 vssd1 vccd1 vccd1 HI[324] insts\[324\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[37\] vssd1 vssd1 vccd1 vccd1 HI[37] insts\[37\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[441\] vssd1 vssd1 vccd1 vccd1 HI[441] insts\[441\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[274\] vssd1 vssd1 vccd1 vccd1 HI[274] insts\[274\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[391\] vssd1 vssd1 vccd1 vccd1 HI[391] insts\[391\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[237\] vssd1 vssd1 vccd1 vccd1 HI[237] insts\[237\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[404\] vssd1 vssd1 vccd1 vccd1 HI[404] insts\[404\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[354\] vssd1 vssd1 vccd1 vccd1 HI[354] insts\[354\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[187\] vssd1 vssd1 vccd1 vccd1 HI[187] insts\[187\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[67\] vssd1 vssd1 vccd1 vccd1 HI[67] insts\[67\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[102\] vssd1 vssd1 vccd1 vccd1 HI[102] insts\[102\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_38 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[317\] vssd1 vssd1 vccd1 vccd1 HI[317] insts\[317\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[434\] vssd1 vssd1 vccd1 vccd1 HI[434] insts\[434\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[267\] vssd1 vssd1 vccd1 vccd1 HI[267] insts\[267\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[384\] vssd1 vssd1 vccd1 vccd1 HI[384] insts\[384\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[97\] vssd1 vssd1 vccd1 vccd1 HI[97] insts\[97\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[132\] vssd1 vssd1 vccd1 vccd1 HI[132] insts\[132\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[12\] vssd1 vssd1 vccd1 vccd1 HI[12] insts\[12\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[347\] vssd1 vssd1 vccd1 vccd1 HI[347] insts\[347\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[297\] vssd1 vssd1 vccd1 vccd1 HI[297] insts\[297\]/LO sky130_fd_sc_hd__conb_1
XPHY_17 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[212\] vssd1 vssd1 vccd1 vccd1 HI[212] insts\[212\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[162\] vssd1 vssd1 vccd1 vccd1 HI[162] insts\[162\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[427\] vssd1 vssd1 vccd1 vccd1 HI[427] insts\[427\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[42\] vssd1 vssd1 vccd1 vccd1 HI[42] insts\[42\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[377\] vssd1 vssd1 vccd1 vccd1 HI[377] insts\[377\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[0\] vssd1 vssd1 vccd1 vccd1 HI[0] insts\[0\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[125\] vssd1 vssd1 vccd1 vccd1 HI[125] insts\[125\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[242\] vssd1 vssd1 vccd1 vccd1 HI[242] insts\[242\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[457\] vssd1 vssd1 vccd1 vccd1 HI[457] insts\[457\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[192\] vssd1 vssd1 vccd1 vccd1 HI[192] insts\[192\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[72\] vssd1 vssd1 vccd1 vccd1 HI[72] insts\[72\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[205\] vssd1 vssd1 vccd1 vccd1 HI[205] insts\[205\]/LO sky130_fd_sc_hd__conb_1
XPHY_18 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_29 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinsts\[155\] vssd1 vssd1 vccd1 vccd1 HI[155] insts\[155\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[322\] vssd1 vssd1 vccd1 vccd1 HI[322] insts\[322\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[35\] vssd1 vssd1 vccd1 vccd1 HI[35] insts\[35\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[272\] vssd1 vssd1 vccd1 vccd1 HI[272] insts\[272\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[118\] vssd1 vssd1 vccd1 vccd1 HI[118] insts\[118\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[235\] vssd1 vssd1 vccd1 vccd1 HI[235] insts\[235\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[402\] vssd1 vssd1 vccd1 vccd1 HI[402] insts\[402\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[185\] vssd1 vssd1 vccd1 vccd1 HI[185] insts\[185\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[352\] vssd1 vssd1 vccd1 vccd1 HI[352] insts\[352\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[65\] vssd1 vssd1 vccd1 vccd1 HI[65] insts\[65\]/LO sky130_fd_sc_hd__conb_1
XPHY_19 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinsts\[100\] vssd1 vssd1 vccd1 vccd1 HI[100] insts\[100\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[148\] vssd1 vssd1 vccd1 vccd1 HI[148] insts\[148\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[315\] vssd1 vssd1 vccd1 vccd1 HI[315] insts\[315\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[28\] vssd1 vssd1 vccd1 vccd1 HI[28] insts\[28\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[265\] vssd1 vssd1 vccd1 vccd1 HI[265] insts\[265\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[432\] vssd1 vssd1 vccd1 vccd1 HI[432] insts\[432\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[382\] vssd1 vssd1 vccd1 vccd1 HI[382] insts\[382\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[95\] vssd1 vssd1 vccd1 vccd1 HI[95] insts\[95\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[228\] vssd1 vssd1 vccd1 vccd1 HI[228] insts\[228\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[130\] vssd1 vssd1 vccd1 vccd1 HI[130] insts\[130\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[10\] vssd1 vssd1 vccd1 vccd1 HI[10] insts\[10\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[178\] vssd1 vssd1 vccd1 vccd1 HI[178] insts\[178\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[345\] vssd1 vssd1 vccd1 vccd1 HI[345] insts\[345\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinsts\[58\] vssd1 vssd1 vccd1 vccd1 HI[58] insts\[58\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[295\] vssd1 vssd1 vccd1 vccd1 HI[295] insts\[295\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
.ends

