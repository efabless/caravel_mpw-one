VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sram_1rw1r_32_256_8_sky130
  CLASS BLOCK ;
  FOREIGN sram_1rw1r_32_256_8_sky130 ;
  ORIGIN 0.000 0.000 ;
  SIZE 386.480 BY 456.235 ;
  SYMMETRY X Y R90 ;
  PIN din0[0]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 63.210000 0.000000 63.510000 4.600000 ;
    END
  END din0[0]

  PIN din0[1]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 69.050000 0.000000 69.350000 4.600000 ;
    END
  END din0[1]

  PIN din0[2]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 74.890000 0.000000 75.190000 4.600000 ;
    END
  END din0[2]

  PIN din0[3]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 80.730000 0.000000 81.030000 4.600000 ;
    END
  END din0[3]

  PIN din0[4]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 86.570000 0.000000 86.870000 4.600000 ;
    END
  END din0[4]

  PIN din0[5]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 92.410000 0.000000 92.710000 4.600000 ;
    END
  END din0[5]

  PIN din0[6]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 98.250000 0.000000 98.550000 4.600000 ;
    END
  END din0[6]

  PIN din0[7]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 104.090000 0.000000 104.390000 4.600000 ;
    END
  END din0[7]

  PIN din0[8]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 109.930000 0.000000 110.230000 4.600000 ;
    END
  END din0[8]

  PIN din0[9]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 115.770000 0.000000 116.070000 4.600000 ;
    END
  END din0[9]

  PIN din0[10]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 121.610000 0.000000 121.910000 4.600000 ;
    END
  END din0[10]

  PIN din0[11]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 127.450000 0.000000 127.750000 4.600000 ;
    END
  END din0[11]

  PIN din0[12]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 133.290000 0.000000 133.590000 4.600000 ;
    END
  END din0[12]

  PIN din0[13]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 139.130000 0.000000 139.430000 4.600000 ;
    END
  END din0[13]

  PIN din0[14]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 144.970000 0.000000 145.270000 4.600000 ;
    END
  END din0[14]

  PIN din0[15]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 150.810000 0.000000 151.110000 4.600000 ;
    END
  END din0[15]

  PIN din0[16]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 156.650000 0.000000 156.950000 4.600000 ;
    END
  END din0[16]

  PIN din0[17]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 162.490000 0.000000 162.790000 4.600000 ;
    END
  END din0[17]

  PIN din0[18]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 168.330000 0.000000 168.630000 4.600000 ;
    END
  END din0[18]

  PIN din0[19]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 174.170000 0.000000 174.470000 4.600000 ;
    END
  END din0[19]

  PIN din0[20]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 180.010000 0.000000 180.310000 4.600000 ;
    END
  END din0[20]

  PIN din0[21]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 185.850000 0.000000 186.150000 4.600000 ;
    END
  END din0[21]

  PIN din0[22]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 191.690000 0.000000 191.990000 4.600000 ;
    END
  END din0[22]

  PIN din0[23]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 197.530000 0.000000 197.830000 4.600000 ;
    END
  END din0[23]

  PIN din0[24]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 203.370000 0.000000 203.670000 4.600000 ;
    END
  END din0[24]

  PIN din0[25]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 209.210000 0.000000 209.510000 4.600000 ;
    END
  END din0[25]

  PIN din0[26]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 215.050000 0.000000 215.350000 4.600000 ;
    END
  END din0[26]

  PIN din0[27]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 220.890000 0.000000 221.190000 4.600000 ;
    END
  END din0[27]

  PIN din0[28]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 226.730000 0.000000 227.030000 4.600000 ;
    END
  END din0[28]

  PIN din0[29]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 232.570000 0.000000 232.870000 4.600000 ;
    END
  END din0[29]

  PIN din0[30]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 238.410000 0.000000 238.710000 4.600000 ;
    END
  END din0[30]

  PIN din0[31]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 244.250000 0.000000 244.550000 4.600000 ;
    END
  END din0[31]

  PIN addr0[0]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 34.010000 0.000000 34.310000 4.600000 ;
    END
  END addr0[0]

  PIN addr0[1]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 390.365000 4.600000 390.665000 ;
    END
  END addr0[1]

  PIN addr0[2]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 398.865000 4.600000 399.165000 ;
    END
  END addr0[2]

  PIN addr0[3]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 404.505000 4.600000 404.805000 ;
    END
  END addr0[3]

  PIN addr0[4]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 413.005000 4.600000 413.305000 ;
    END
  END addr0[4]

  PIN addr0[5]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 418.645000 4.600000 418.945000 ;
    END
  END addr0[5]

  PIN addr0[6]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 427.145000 4.600000 427.445000 ;
    END
  END addr0[6]

  PIN addr0[7]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 432.785000 4.600000 433.085000 ;
    END
  END addr0[7]

  PIN addr1[0]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 342.890000 452.035000 343.190000 456.235000 ;
    END
  END addr1[0]

  PIN addr1[1]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 382.180000 146.910000 386.480000 147.210000 ;
    END
  END addr1[1]

  PIN addr1[2]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 382.180000 138.410000 386.480000 138.710000 ;
    END
  END addr1[2]

  PIN addr1[3]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 382.180000 132.770000 386.480000 133.070000 ;
    END
  END addr1[3]

  PIN addr1[4]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 382.180000 124.270000 386.480000 124.570000 ;
    END
  END addr1[4]

  PIN addr1[5]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 382.180000 118.630000 386.480000 118.930000 ;
    END
  END addr1[5]

  PIN addr1[6]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 382.180000 110.130000 386.480000 110.430000 ;
    END
  END addr1[6]

  PIN addr1[7]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 382.180000 104.490000 386.480000 104.790000 ;
    END
  END addr1[7]

  PIN csb0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.625000 4.600000 92.925000 ;
    END
  END csb0

  PIN csb1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 382.180000 448.265000 386.480000 448.565000 ;
    END
  END csb1

  PIN web0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.125000 4.600000 101.425000 ;
    END
  END web0

  PIN clk0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER met4 ;
        RECT 19.015000 0.000000 19.315000 4.600000 ;
    END
  END clk0

  PIN clk1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER met4 ;
        RECT 367.865000 452.035000 368.165000 456.235000 ;
    END
  END clk1

  PIN wmask0[0]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 39.850000 0.000000 40.150000 4.600000 ;
    END
  END wmask0[0]

  PIN wmask0[1]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 45.690000 0.000000 45.990000 4.600000 ;
    END
  END wmask0[1]

  PIN wmask0[2]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 51.530000 0.000000 51.830000 4.600000 ;
    END
  END wmask0[2]

  PIN wmask0[3]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met4 ;
        RECT 57.370000 0.000000 57.670000 4.600000 ;
    END
  END wmask0[3]

  PIN dout0[0]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 63.830000 0.000000 64.130000 4.600000 ;
    END
  END dout0[0]

  PIN dout0[1]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 69.670000 0.000000 69.970000 4.600000 ;
    END
  END dout0[1]

  PIN dout0[2]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 75.510000 0.000000 75.810000 4.600000 ;
    END
  END dout0[2]

  PIN dout0[3]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 81.350000 0.000000 81.650000 4.600000 ;
    END
  END dout0[3]

  PIN dout0[4]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 87.190000 0.000000 87.490000 4.600000 ;
    END
  END dout0[4]

  PIN dout0[5]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 93.030000 0.000000 93.330000 4.600000 ;
    END
  END dout0[5]

  PIN dout0[6]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 98.870000 0.000000 99.170000 4.600000 ;
    END
  END dout0[6]

  PIN dout0[7]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 104.710000 0.000000 105.010000 4.600000 ;
    END
  END dout0[7]

  PIN dout0[8]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 110.550000 0.000000 110.850000 4.600000 ;
    END
  END dout0[8]

  PIN dout0[9]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 116.390000 0.000000 116.690000 4.600000 ;
    END
  END dout0[9]

  PIN dout0[10]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 122.230000 0.000000 122.530000 4.600000 ;
    END
  END dout0[10]

  PIN dout0[11]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 128.070000 0.000000 128.370000 4.600000 ;
    END
  END dout0[11]

  PIN dout0[12]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 133.910000 0.000000 134.210000 4.600000 ;
    END
  END dout0[12]

  PIN dout0[13]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 139.750000 0.000000 140.050000 4.600000 ;
    END
  END dout0[13]

  PIN dout0[14]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 145.590000 0.000000 145.890000 4.600000 ;
    END
  END dout0[14]

  PIN dout0[15]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 151.430000 0.000000 151.730000 4.600000 ;
    END
  END dout0[15]

  PIN dout0[16]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 157.270000 0.000000 157.570000 4.600000 ;
    END
  END dout0[16]

  PIN dout0[17]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 163.110000 0.000000 163.410000 4.600000 ;
    END
  END dout0[17]

  PIN dout0[18]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 168.950000 0.000000 169.250000 4.600000 ;
    END
  END dout0[18]

  PIN dout0[19]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 174.790000 0.000000 175.090000 4.600000 ;
    END
  END dout0[19]

  PIN dout0[20]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 180.630000 0.000000 180.930000 4.600000 ;
    END
  END dout0[20]

  PIN dout0[21]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 186.470000 0.000000 186.770000 4.600000 ;
    END
  END dout0[21]

  PIN dout0[22]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 192.310000 0.000000 192.610000 4.600000 ;
    END
  END dout0[22]

  PIN dout0[23]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 198.150000 0.000000 198.450000 4.600000 ;
    END
  END dout0[23]

  PIN dout0[24]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 203.990000 0.000000 204.290000 4.600000 ;
    END
  END dout0[24]

  PIN dout0[25]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 209.830000 0.000000 210.130000 4.600000 ;
    END
  END dout0[25]

  PIN dout0[26]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 215.670000 0.000000 215.970000 4.600000 ;
    END
  END dout0[26]

  PIN dout0[27]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 221.510000 0.000000 221.810000 4.600000 ;
    END
  END dout0[27]

  PIN dout0[28]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 227.350000 0.000000 227.650000 4.600000 ;
    END
  END dout0[28]

  PIN dout0[29]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 233.190000 0.000000 233.490000 4.600000 ;
    END
  END dout0[29]

  PIN dout0[30]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 239.030000 0.000000 239.330000 4.600000 ;
    END
  END dout0[30]

  PIN dout0[31]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 244.870000 0.000000 245.170000 4.600000 ;
    END
  END dout0[31]

  PIN dout1[0]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 94.025000 452.035000 94.325000 456.235000 ;
    END
  END dout1[0]

  PIN dout1[1]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 100.265000 452.035000 100.565000 456.235000 ;
    END
  END dout1[1]

  PIN dout1[2]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 106.505000 452.035000 106.805000 456.235000 ;
    END
  END dout1[2]

  PIN dout1[3]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 112.745000 452.035000 113.045000 456.235000 ;
    END
  END dout1[3]

  PIN dout1[4]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 118.985000 452.035000 119.285000 456.235000 ;
    END
  END dout1[4]

  PIN dout1[5]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 125.225000 452.035000 125.525000 456.235000 ;
    END
  END dout1[5]

  PIN dout1[6]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 131.465000 452.035000 131.765000 456.235000 ;
    END
  END dout1[6]

  PIN dout1[7]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 137.705000 452.035000 138.005000 456.235000 ;
    END
  END dout1[7]

  PIN dout1[8]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 143.945000 452.035000 144.245000 456.235000 ;
    END
  END dout1[8]

  PIN dout1[9]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 150.185000 452.035000 150.485000 456.235000 ;
    END
  END dout1[9]

  PIN dout1[10]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 156.425000 452.035000 156.725000 456.235000 ;
    END
  END dout1[10]

  PIN dout1[11]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 162.665000 452.035000 162.965000 456.235000 ;
    END
  END dout1[11]

  PIN dout1[12]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 168.905000 452.035000 169.205000 456.235000 ;
    END
  END dout1[12]

  PIN dout1[13]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 175.145000 452.035000 175.445000 456.235000 ;
    END
  END dout1[13]

  PIN dout1[14]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 181.385000 452.035000 181.685000 456.235000 ;
    END
  END dout1[14]

  PIN dout1[15]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 187.625000 452.035000 187.925000 456.235000 ;
    END
  END dout1[15]

  PIN dout1[16]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 193.865000 452.035000 194.165000 456.235000 ;
    END
  END dout1[16]

  PIN dout1[17]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 200.105000 452.035000 200.405000 456.235000 ;
    END
  END dout1[17]

  PIN dout1[18]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 206.345000 452.035000 206.645000 456.235000 ;
    END
  END dout1[18]

  PIN dout1[19]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 212.585000 452.035000 212.885000 456.235000 ;
    END
  END dout1[19]

  PIN dout1[20]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 218.825000 452.035000 219.125000 456.235000 ;
    END
  END dout1[20]

  PIN dout1[21]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 225.065000 452.035000 225.365000 456.235000 ;
    END
  END dout1[21]

  PIN dout1[22]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 231.305000 452.035000 231.605000 456.235000 ;
    END
  END dout1[22]

  PIN dout1[23]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 237.545000 452.035000 237.845000 456.235000 ;
    END
  END dout1[23]

  PIN dout1[24]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 243.785000 452.035000 244.085000 456.235000 ;
    END
  END dout1[24]

  PIN dout1[25]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 250.025000 452.035000 250.325000 456.235000 ;
    END
  END dout1[25]

  PIN dout1[26]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 256.265000 452.035000 256.565000 456.235000 ;
    END
  END dout1[26]

  PIN dout1[27]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 262.505000 452.035000 262.805000 456.235000 ;
    END
  END dout1[27]

  PIN dout1[28]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 268.745000 452.035000 269.045000 456.235000 ;
    END
  END dout1[28]

  PIN dout1[29]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 274.985000 452.035000 275.285000 456.235000 ;
    END
  END dout1[29]

  PIN dout1[30]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 281.225000 452.035000 281.525000 456.235000 ;
    END
  END dout1[30]

  PIN dout1[31]
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.553900 ;
    PORT
      LAYER met4 ;
        RECT 287.465000 452.035000 287.765000 456.235000 ;
    END
  END dout1[31]

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 381.040 443.600 384.050 444.660 ;
      LAYER via3 ;
        RECT 382.500 443.620 384.020 444.630 ;
      LAYER met4 ;
        RECT 382.470 3.670 384.070 444.680 ;
    END
  END vdd

  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 359.280 451.080 361.020 452.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.040 450.400 386.300 452.140 ;
      LAYER via3 ;
        RECT 384.720 450.440 386.240 452.050 ;
      LAYER met4 ;
        RECT 384.690 4.060 386.310 452.140 ;
    END
  END gnd

  OBS
     LAYER li1 ;
       RECT 5.000 5.000 381.780 451.535 ;
     LAYER met1 ;
       RECT 5.000 5.000 381.780 451.535 ;
     LAYER met2 ;
       RECT 5.000 5.000 381.780 451.535 ;
     LAYER met3 ;
       RECT 5.000 5.000 381.780 451.535 ;
     LAYER met4 ;
       RECT 5.000 5.000 381.780 451.535 ;
  END
END sram_1rw1r_32_256_8_sky130
END LIBRARY

