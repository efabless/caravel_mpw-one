magic
tech sky130A
magscale 1 2
timestamp 1619659917
<< error_s >>
rect 78120 1031109 91280 1031322
rect 78120 1018304 78290 1031109
rect 78440 1030789 90960 1031002
rect 78440 1018624 78610 1030789
rect 90778 1018624 90960 1030789
rect 78440 1018512 90960 1018624
rect 91098 1018304 91280 1031109
rect 78120 1018192 91280 1018304
rect 129520 1031109 142680 1031322
rect 129520 1018304 129690 1031109
rect 129840 1030789 142360 1031002
rect 129840 1018624 130010 1030789
rect 142178 1018624 142360 1030789
rect 129840 1018512 142360 1018624
rect 142498 1018304 142680 1031109
rect 129520 1018192 142680 1018304
rect 180920 1031109 194080 1031322
rect 232320 1031245 245480 1031322
rect 283920 1031245 297080 1031322
rect 385720 1031245 398880 1031322
rect 180920 1018304 181090 1031109
rect 181240 1030789 193760 1031002
rect 181240 1018624 181410 1030789
rect 193578 1018624 193760 1030789
rect 181240 1018512 193760 1018624
rect 193898 1018304 194080 1031109
rect 474720 1031109 487880 1031322
rect 232640 1030925 245160 1031002
rect 284240 1030925 296760 1031002
rect 386040 1030925 398560 1031002
rect 180920 1018192 194080 1018304
rect 474720 1018304 474890 1031109
rect 475040 1030789 487560 1031002
rect 475040 1018624 475210 1030789
rect 487378 1018624 487560 1030789
rect 475040 1018512 487560 1018624
rect 487698 1018304 487880 1031109
rect 474720 1018192 487880 1018304
rect 526120 1031109 539280 1031322
rect 526120 1018304 526290 1031109
rect 526440 1030789 538960 1031002
rect 526440 1018624 526610 1030789
rect 538778 1018624 538960 1030789
rect 526440 1018512 538960 1018624
rect 539098 1018304 539280 1031109
rect 526120 1018192 539280 1018304
rect 627920 1031109 641080 1031322
rect 627920 1018304 628090 1031109
rect 628240 1030789 640760 1031002
rect 628240 1018624 628410 1030789
rect 640578 1018624 640760 1030789
rect 628240 1018512 640760 1018624
rect 640898 1018304 641080 1031109
rect 627920 1018192 641080 1018304
rect 6278 969098 19408 969280
rect 6278 956290 6491 969098
rect 6598 968778 19088 968960
rect 6598 956610 6811 968778
rect 18976 956610 19088 968778
rect 6598 956440 19088 956610
rect 19296 956290 19408 969098
rect 6278 956120 19408 956290
rect 698192 965510 711322 965680
rect 698192 952702 698304 965510
rect 698512 965190 711002 965360
rect 698512 953022 698624 965190
rect 710789 953022 711002 965190
rect 698512 952840 711002 953022
rect 711109 952702 711322 965510
rect 698192 952520 711322 952702
rect 141667 39934 141813 40000
rect 145091 39934 145143 40000
rect 145464 39289 145492 39299
rect 145436 39285 145492 39289
rect 145436 39271 145489 39285
rect 144523 39241 144579 39269
rect 144623 39261 144653 39269
rect 144523 39233 144551 39241
rect 144571 39233 144579 39241
rect 144597 39241 144653 39261
rect 145436 39261 145442 39271
rect 145436 39247 145461 39261
rect 145464 39247 145489 39271
rect 145436 39243 145464 39247
rect 145502 39242 145558 39247
rect 144523 39215 144571 39233
rect 144597 39215 144625 39241
rect 144523 39213 144625 39215
rect 145433 39219 145558 39242
rect 145433 39214 145489 39219
rect 144551 39205 144599 39213
rect 144543 39187 144599 39205
rect 145461 39191 145525 39214
rect 145530 39191 145558 39219
rect 144543 39159 144571 39187
rect 145461 39186 145489 39191
rect 145497 39163 145530 39178
rect 145497 39150 145553 39163
rect 145525 39122 145553 39150
rect 145571 39150 145627 39178
rect 145571 39135 145591 39150
rect 145599 39135 145627 39150
rect 145591 39122 145627 39135
rect 145573 39084 145591 39085
rect 141748 39020 141804 39048
rect 141847 39039 143068 39077
rect 143128 39039 144423 39077
rect 145601 39056 145619 39085
rect 141748 39011 141776 39020
rect 141784 39011 141804 39020
rect 141822 39020 141878 39039
rect 141748 38992 141784 39011
rect 141822 38992 141850 39020
rect 141682 38954 141738 38982
rect 141776 38969 141812 38982
rect 141684 38934 141712 38954
rect 141736 38934 141738 38954
rect 141684 38928 141738 38934
rect 141756 38954 141812 38969
rect 141684 38926 141736 38928
rect 141756 38926 141784 38954
rect 143002 38377 143122 38433
rect 143355 38420 143448 38433
rect 143328 38377 143448 38420
rect 142946 38373 143448 38377
rect 142946 38317 143079 38373
rect 143272 38317 143392 38373
rect 142946 38300 143006 38317
rect 143019 38313 143332 38317
rect 143019 38300 143066 38313
rect 142946 38257 143019 38300
rect 143272 38257 143332 38313
rect 145505 38178 145561 38188
rect 145601 38178 145635 38188
rect 143006 38120 143019 38161
rect 145505 38148 145567 38178
rect 145579 38160 145635 38178
rect 145579 38148 145607 38160
rect 145465 38136 145607 38148
rect 145465 38132 145533 38136
rect 145539 38132 145607 38136
rect 145465 38120 145521 38132
rect 145539 38120 145595 38132
rect 142959 38101 143006 38120
rect 143019 38101 143066 38120
rect 145465 38108 145493 38120
rect 145501 38108 145521 38120
rect 145533 38108 145567 38120
rect 143006 38060 143019 38101
rect 145465 38092 145501 38108
rect 145539 38092 145567 38108
rect 145493 38080 145529 38082
rect 145473 38054 145529 38080
rect 141813 37971 141933 38031
rect 145473 38026 145501 38054
rect 141813 37911 141820 37971
rect 141873 37911 141933 37971
rect 141656 37805 141684 37811
rect 141736 37795 141748 37811
rect 141684 37783 141748 37795
rect 141692 37767 141748 37783
rect 141684 37755 141720 37767
rect 141692 37739 141720 37755
rect 141594 36821 141629 36832
rect 141573 36804 141629 36821
rect 141573 36776 141601 36804
rect 145902 36801 146022 36861
rect 145902 36771 145934 36801
rect 145962 36771 146022 36801
rect 145902 36743 146112 36771
rect 145874 36711 146112 36743
rect 145874 36683 145994 36711
rect 145934 36651 146026 36683
rect 146052 36651 146112 36711
rect 145934 36623 145994 36651
rect 146142 36621 146202 36651
rect 146082 36536 146141 36591
rect 146142 36536 146201 36591
rect 146082 36531 146201 36536
rect 145418 34371 145470 34398
rect 145418 34343 145470 34370
rect 145318 33775 145374 33782
rect 145318 33737 145375 33775
rect 145273 33733 145403 33737
rect 145273 33710 145346 33733
rect 145347 33710 145403 33733
rect 145273 33709 145403 33710
rect 145296 33704 145376 33709
rect 145296 33682 145375 33704
rect 145296 33681 145348 33682
rect 145964 33624 146084 33684
rect 146141 33669 146230 33684
rect 145964 33609 146024 33624
rect 146027 33609 146084 33624
rect 146110 33624 146230 33669
rect 145964 33564 146027 33609
rect 146110 33564 146170 33624
rect 145821 33481 145941 33541
rect 146024 33519 146087 33541
rect 145821 33459 145881 33481
rect 145910 33459 145941 33481
rect 145967 33481 146087 33519
rect 145821 33424 145910 33459
rect 145967 33424 146027 33481
rect 145704 33421 146027 33424
rect 145704 33364 145824 33421
rect 145881 33399 145970 33421
rect 145721 33351 145781 33364
rect 145806 33351 145824 33364
rect 143145 33321 145824 33351
rect 145850 33364 145970 33399
rect 143145 33320 145837 33321
rect 145850 33320 145910 33364
rect 143145 33304 145910 33320
rect 143145 33260 145866 33304
rect 143145 33231 145806 33260
rect 143145 33175 145721 33231
rect 145746 33200 145806 33231
rect 132948 30016 133162 30063
rect 132948 29956 133162 30003
rect 133762 26500 133822 26510
rect 133422 26480 133822 26500
rect 133422 26450 133799 26480
rect 133422 26440 133542 26450
rect 133482 26390 133739 26440
rect 133762 26390 133799 26450
rect 133482 26380 133542 26390
rect 133889 26300 134009 26353
rect 133739 26293 134009 26300
rect 133739 26270 133942 26293
rect 133949 26270 134009 26293
rect 133739 26243 134009 26270
rect 133679 26233 134009 26243
rect 133679 26210 134002 26233
rect 133679 26183 133799 26210
rect 133739 26180 133929 26183
rect 133949 26180 133989 26210
rect 133739 26150 133949 26180
rect 133739 26123 133799 26150
rect 134122 26120 134182 26150
rect 133929 26090 134122 26120
rect 133929 26053 134122 26060
rect 133869 26000 134122 26053
rect 133869 25993 133989 26000
rect 133929 25940 134122 25993
rect 133929 25933 133989 25940
rect 134392 25860 134452 25880
rect 134062 25850 134452 25860
rect 134062 25820 134424 25850
rect 134062 25800 134182 25820
rect 134122 25760 134364 25800
rect 134392 25760 134424 25820
rect 134122 25740 134182 25760
rect 134304 25584 134368 25618
rect 134304 25558 134424 25584
rect 134364 25520 134424 25558
rect 134402 25498 134424 25520
rect 147800 21003 147920 25993
<< metal1 >>
rect 673454 875168 673460 875220
rect 673512 875208 673518 875220
rect 675386 875208 675392 875220
rect 673512 875180 675392 875208
rect 673512 875168 673518 875180
rect 675386 875168 675392 875180
rect 675444 875168 675450 875220
rect 673546 874488 673552 874540
rect 673604 874528 673610 874540
rect 675386 874528 675392 874540
rect 673604 874500 675392 874528
rect 673604 874488 673610 874500
rect 675386 874488 675392 874500
rect 675444 874488 675450 874540
rect 673730 870136 673736 870188
rect 673788 870176 673794 870188
rect 675386 870176 675392 870188
rect 673788 870148 675392 870176
rect 673788 870136 673794 870148
rect 675386 870136 675392 870148
rect 675444 870136 675450 870188
rect 673638 864424 673644 864476
rect 673696 864464 673702 864476
rect 675386 864464 675392 864476
rect 673696 864436 675392 864464
rect 673696 864424 673702 864436
rect 675386 864424 675392 864436
rect 675444 864424 675450 864476
rect 673730 863200 673736 863252
rect 673788 863240 673794 863252
rect 675386 863240 675392 863252
rect 673788 863212 675392 863240
rect 673788 863200 673794 863212
rect 675386 863200 675392 863212
rect 675444 863200 675450 863252
rect 675294 818320 675300 818372
rect 675352 818360 675358 818372
rect 677502 818360 677508 818372
rect 675352 818332 677508 818360
rect 675352 818320 675358 818332
rect 677502 818320 677508 818332
rect 677560 818320 677566 818372
rect 41782 799552 41788 799604
rect 41840 799592 41846 799604
rect 42334 799592 42340 799604
rect 41840 799564 42340 799592
rect 41840 799552 41846 799564
rect 42334 799552 42340 799564
rect 42392 799552 42398 799604
rect 41782 797716 41788 797768
rect 41840 797756 41846 797768
rect 42702 797756 42708 797768
rect 41840 797728 42708 797756
rect 41840 797716 41846 797728
rect 42702 797716 42708 797728
rect 42760 797716 42766 797768
rect 41782 792548 41788 792600
rect 41840 792588 41846 792600
rect 42334 792588 42340 792600
rect 41840 792560 42340 792588
rect 41840 792548 41846 792560
rect 42334 792548 42340 792560
rect 42392 792548 42398 792600
rect 41782 787244 41788 787296
rect 41840 787284 41846 787296
rect 42610 787284 42616 787296
rect 41840 787256 42616 787284
rect 41840 787244 41846 787256
rect 42610 787244 42616 787256
rect 42668 787244 42674 787296
rect 41782 786632 41788 786684
rect 41840 786672 41846 786684
rect 42518 786672 42524 786684
rect 41840 786644 42524 786672
rect 41840 786632 41846 786644
rect 42518 786632 42524 786644
rect 42576 786632 42582 786684
rect 673454 786564 673460 786616
rect 673512 786604 673518 786616
rect 674006 786604 674012 786616
rect 673512 786576 674012 786604
rect 673512 786564 673518 786576
rect 674006 786564 674012 786576
rect 674064 786604 674070 786616
rect 675386 786604 675392 786616
rect 674064 786576 675392 786604
rect 674064 786564 674070 786576
rect 675386 786564 675392 786576
rect 675444 786564 675450 786616
rect 673546 786360 673552 786412
rect 673604 786400 673610 786412
rect 675386 786400 675392 786412
rect 673604 786372 675392 786400
rect 673604 786360 673610 786372
rect 675386 786360 675392 786372
rect 675444 786360 675450 786412
rect 675294 781600 675300 781652
rect 675352 781600 675358 781652
rect 675312 781448 675340 781600
rect 675294 781396 675300 781448
rect 675352 781396 675358 781448
rect 673454 774868 673460 774920
rect 673512 774908 673518 774920
rect 673638 774908 673644 774920
rect 673512 774880 673644 774908
rect 673512 774868 673518 774880
rect 673638 774868 673644 774880
rect 673696 774908 673702 774920
rect 675386 774908 675392 774920
rect 673696 774880 675392 774908
rect 673696 774868 673702 774880
rect 675386 774868 675392 774880
rect 675444 774868 675450 774920
rect 675202 773984 675208 774036
rect 675260 774024 675266 774036
rect 675386 774024 675392 774036
rect 675260 773996 675392 774024
rect 675260 773984 675266 773996
rect 675386 773984 675392 773996
rect 675444 773984 675450 774036
rect 673730 772760 673736 772812
rect 673788 772800 673794 772812
rect 674006 772800 674012 772812
rect 673788 772772 674012 772800
rect 673788 772760 673794 772772
rect 674006 772760 674012 772772
rect 674064 772760 674070 772812
rect 42426 767320 42432 767372
rect 42484 767360 42490 767372
rect 42702 767360 42708 767372
rect 42484 767332 42708 767360
rect 42484 767320 42490 767332
rect 42702 767320 42708 767332
rect 42760 767320 42766 767372
rect 42518 758956 42524 759008
rect 42576 758996 42582 759008
rect 42794 758996 42800 759008
rect 42576 758968 42800 758996
rect 42576 758956 42582 758968
rect 42794 758956 42800 758968
rect 42852 758956 42858 759008
rect 41782 756372 41788 756424
rect 41840 756412 41846 756424
rect 42334 756412 42340 756424
rect 41840 756384 42340 756412
rect 41840 756372 41846 756384
rect 42334 756372 42340 756384
rect 42392 756372 42398 756424
rect 41782 754468 41788 754520
rect 41840 754508 41846 754520
rect 42426 754508 42432 754520
rect 41840 754480 42432 754508
rect 41840 754468 41846 754480
rect 42426 754468 42432 754480
rect 42484 754468 42490 754520
rect 673730 753516 673736 753568
rect 673788 753556 673794 753568
rect 673914 753556 673920 753568
rect 673788 753528 673920 753556
rect 673788 753516 673794 753528
rect 673914 753516 673920 753528
rect 673972 753516 673978 753568
rect 42518 753448 42524 753500
rect 42576 753488 42582 753500
rect 42794 753488 42800 753500
rect 42576 753460 42800 753488
rect 42576 753448 42582 753460
rect 42794 753448 42800 753460
rect 42852 753448 42858 753500
rect 41782 749368 41788 749420
rect 41840 749408 41846 749420
rect 42334 749408 42340 749420
rect 41840 749380 42340 749408
rect 41840 749368 41846 749380
rect 42334 749368 42340 749380
rect 42392 749368 42398 749420
rect 41782 744132 41788 744184
rect 41840 744172 41846 744184
rect 42334 744172 42340 744184
rect 41840 744144 42340 744172
rect 41840 744132 41846 744144
rect 42334 744132 42340 744144
rect 42392 744172 42398 744184
rect 42610 744172 42616 744184
rect 42392 744144 42616 744172
rect 42392 744132 42398 744144
rect 42610 744132 42616 744144
rect 42668 744132 42674 744184
rect 41782 743996 41788 744048
rect 41840 744036 41846 744048
rect 42518 744036 42524 744048
rect 41840 744008 42524 744036
rect 41840 743996 41846 744008
rect 42518 743996 42524 744008
rect 42576 744036 42582 744048
rect 42978 744036 42984 744048
rect 42576 744008 42984 744036
rect 42576 743996 42582 744008
rect 42978 743996 42984 744008
rect 43036 743996 43042 744048
rect 673638 741956 673644 742008
rect 673696 741996 673702 742008
rect 673914 741996 673920 742008
rect 673696 741968 673920 741996
rect 673696 741956 673702 741968
rect 673914 741956 673920 741968
rect 673972 741996 673978 742008
rect 673972 741968 675432 741996
rect 673972 741956 673978 741968
rect 675404 741940 675432 741968
rect 675386 741888 675392 741940
rect 675444 741888 675450 741940
rect 673546 740664 673552 740716
rect 673604 740704 673610 740716
rect 675386 740704 675392 740716
rect 673604 740676 675392 740704
rect 673604 740664 673610 740676
rect 675386 740664 675392 740676
rect 675444 740664 675450 740716
rect 673638 739780 673644 739832
rect 673696 739780 673702 739832
rect 673656 739696 673684 739780
rect 673638 739644 673644 739696
rect 673696 739644 673702 739696
rect 42334 739576 42340 739628
rect 42392 739616 42398 739628
rect 42610 739616 42616 739628
rect 42392 739588 42616 739616
rect 42392 739576 42398 739588
rect 42610 739576 42616 739588
rect 42668 739576 42674 739628
rect 42518 734136 42524 734188
rect 42576 734176 42582 734188
rect 42978 734176 42984 734188
rect 42576 734148 42984 734176
rect 42576 734136 42582 734148
rect 42978 734136 42984 734148
rect 43036 734136 43042 734188
rect 673454 730124 673460 730176
rect 673512 730164 673518 730176
rect 675386 730164 675392 730176
rect 673512 730136 675392 730164
rect 673512 730124 673518 730136
rect 675386 730124 675392 730136
rect 675444 730124 675450 730176
rect 42518 720332 42524 720384
rect 42576 720372 42582 720384
rect 42886 720372 42892 720384
rect 42576 720344 42892 720372
rect 42576 720332 42582 720344
rect 42886 720332 42892 720344
rect 42944 720332 42950 720384
rect 41782 713124 41788 713176
rect 41840 713164 41846 713176
rect 42334 713164 42340 713176
rect 41840 713136 42340 713164
rect 41840 713124 41846 713136
rect 42334 713124 42340 713136
rect 42392 713124 42398 713176
rect 41782 711288 41788 711340
rect 41840 711328 41846 711340
rect 42426 711328 42432 711340
rect 41840 711300 42432 711328
rect 41840 711288 41846 711300
rect 42426 711288 42432 711300
rect 42484 711328 42490 711340
rect 42702 711328 42708 711340
rect 42484 711300 42708 711328
rect 42484 711288 42490 711300
rect 42702 711288 42708 711300
rect 42760 711288 42766 711340
rect 41782 706188 41788 706240
rect 41840 706228 41846 706240
rect 42334 706228 42340 706240
rect 41840 706200 42340 706228
rect 41840 706188 41846 706200
rect 42334 706188 42340 706200
rect 42392 706188 42398 706240
rect 673638 701020 673644 701072
rect 673696 701060 673702 701072
rect 673822 701060 673828 701072
rect 673696 701032 673828 701060
rect 673696 701020 673702 701032
rect 673822 701020 673828 701032
rect 673880 701020 673886 701072
rect 41782 700952 41788 701004
rect 41840 700992 41846 701004
rect 42610 700992 42616 701004
rect 41840 700964 42616 700992
rect 41840 700952 41846 700964
rect 42610 700952 42616 700964
rect 42668 700952 42674 701004
rect 41782 700816 41788 700868
rect 41840 700856 41846 700868
rect 42886 700856 42892 700868
rect 41840 700828 42892 700856
rect 41840 700816 41846 700828
rect 42886 700816 42892 700828
rect 42944 700816 42950 700868
rect 675386 695920 675392 695972
rect 675444 695920 675450 695972
rect 673638 695852 673644 695904
rect 673696 695892 673702 695904
rect 675404 695892 675432 695920
rect 673696 695864 675432 695892
rect 673696 695852 673702 695864
rect 42426 695512 42432 695564
rect 42484 695552 42490 695564
rect 42886 695552 42892 695564
rect 42484 695524 42892 695552
rect 42484 695512 42490 695524
rect 42886 695512 42892 695524
rect 42944 695512 42950 695564
rect 673546 695308 673552 695360
rect 673604 695348 673610 695360
rect 675386 695348 675392 695360
rect 673604 695320 675392 695348
rect 673604 695308 673610 695320
rect 675386 695308 675392 695320
rect 675444 695308 675450 695360
rect 673454 685176 673460 685228
rect 673512 685216 673518 685228
rect 675386 685216 675392 685228
rect 673512 685188 675392 685216
rect 673512 685176 673518 685188
rect 675386 685176 675392 685188
rect 675444 685176 675450 685228
rect 42426 681640 42432 681692
rect 42484 681640 42490 681692
rect 42444 681612 42472 681640
rect 42794 681612 42800 681624
rect 42444 681584 42800 681612
rect 42794 681572 42800 681584
rect 42852 681572 42858 681624
rect 42610 678512 42616 678564
rect 42668 678552 42674 678564
rect 42978 678552 42984 678564
rect 42668 678524 42984 678552
rect 42668 678512 42674 678524
rect 42978 678512 42984 678524
rect 43036 678512 43042 678564
rect 42426 676132 42432 676184
rect 42484 676172 42490 676184
rect 42978 676172 42984 676184
rect 42484 676144 42984 676172
rect 42484 676132 42490 676144
rect 42978 676132 42984 676144
rect 43036 676132 43042 676184
rect 41782 669944 41788 669996
rect 41840 669984 41846 669996
rect 42334 669984 42340 669996
rect 41840 669956 42340 669984
rect 41840 669944 41846 669956
rect 42334 669944 42340 669956
rect 42392 669944 42398 669996
rect 41782 669060 41788 669112
rect 41840 669100 41846 669112
rect 42518 669100 42524 669112
rect 41840 669072 42524 669100
rect 41840 669060 41846 669072
rect 42518 669060 42524 669072
rect 42576 669060 42582 669112
rect 41782 663008 41788 663060
rect 41840 663048 41846 663060
rect 42334 663048 42340 663060
rect 41840 663020 42340 663048
rect 41840 663008 41846 663020
rect 42334 663008 42340 663020
rect 42392 663008 42398 663060
rect 41782 658656 41788 658708
rect 41840 658696 41846 658708
rect 42426 658696 42432 658708
rect 41840 658668 42432 658696
rect 41840 658656 41846 658668
rect 42426 658656 42432 658668
rect 42484 658696 42490 658708
rect 42702 658696 42708 658708
rect 42484 658668 42708 658696
rect 42484 658656 42490 658668
rect 42702 658656 42708 658668
rect 42760 658656 42766 658708
rect 41782 658044 41788 658096
rect 41840 658084 41846 658096
rect 42794 658084 42800 658096
rect 41840 658056 42800 658084
rect 41840 658044 41846 658056
rect 42794 658044 42800 658056
rect 42852 658044 42858 658096
rect 673638 651720 673644 651772
rect 673696 651760 673702 651772
rect 675386 651760 675392 651772
rect 673696 651732 675392 651760
rect 673696 651720 673702 651732
rect 675386 651720 675392 651732
rect 675444 651720 675450 651772
rect 42426 651380 42432 651432
rect 42484 651420 42490 651432
rect 42794 651420 42800 651432
rect 42484 651392 42800 651420
rect 42484 651380 42490 651392
rect 42794 651380 42800 651392
rect 42852 651380 42858 651432
rect 673546 651108 673552 651160
rect 673604 651148 673610 651160
rect 675386 651148 675392 651160
rect 673604 651120 675392 651148
rect 673604 651108 673610 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 675202 646008 675208 646060
rect 675260 646008 675266 646060
rect 675220 645776 675248 646008
rect 675294 645776 675300 645788
rect 675220 645748 675300 645776
rect 675294 645736 675300 645748
rect 675352 645736 675358 645788
rect 673454 639684 673460 639736
rect 673512 639724 673518 639736
rect 673914 639724 673920 639736
rect 673512 639696 673920 639724
rect 673512 639684 673518 639696
rect 673914 639684 673920 639696
rect 673972 639724 673978 639736
rect 675386 639724 675392 639736
rect 673972 639696 675392 639724
rect 673972 639684 673978 639696
rect 675386 639684 675392 639696
rect 675444 639684 675450 639736
rect 675202 638800 675208 638852
rect 675260 638840 675266 638852
rect 675386 638840 675392 638852
rect 675260 638812 675392 638840
rect 675260 638800 675266 638812
rect 675386 638800 675392 638812
rect 675444 638800 675450 638852
rect 42518 632000 42524 632052
rect 42576 632000 42582 632052
rect 42702 632000 42708 632052
rect 42760 632040 42766 632052
rect 42978 632040 42984 632052
rect 42760 632012 42984 632040
rect 42760 632000 42766 632012
rect 42978 632000 42984 632012
rect 43036 632000 43042 632052
rect 42536 631904 42564 632000
rect 42794 631904 42800 631916
rect 42536 631876 42800 631904
rect 42794 631864 42800 631876
rect 42852 631864 42858 631916
rect 41782 626764 41788 626816
rect 41840 626804 41846 626816
rect 42334 626804 42340 626816
rect 41840 626776 42340 626804
rect 41840 626764 41846 626776
rect 42334 626764 42340 626776
rect 42392 626764 42398 626816
rect 41782 624928 41788 624980
rect 41840 624968 41846 624980
rect 42794 624968 42800 624980
rect 41840 624940 42800 624968
rect 41840 624928 41846 624940
rect 42794 624928 42800 624940
rect 42852 624928 42858 624980
rect 41782 619760 41788 619812
rect 41840 619800 41846 619812
rect 42334 619800 42340 619812
rect 41840 619772 42340 619800
rect 41840 619760 41846 619772
rect 42334 619760 42340 619772
rect 42392 619760 42398 619812
rect 41782 615476 41788 615528
rect 41840 615516 41846 615528
rect 42978 615516 42984 615528
rect 41840 615488 42984 615516
rect 41840 615476 41846 615488
rect 42978 615476 42984 615488
rect 43036 615476 43042 615528
rect 41782 614796 41788 614848
rect 41840 614836 41846 614848
rect 42518 614836 42524 614848
rect 41840 614808 42524 614836
rect 41840 614796 41846 614808
rect 42518 614796 42524 614808
rect 42576 614796 42582 614848
rect 42794 612824 42800 612876
rect 42852 612824 42858 612876
rect 42610 612756 42616 612808
rect 42668 612796 42674 612808
rect 42812 612796 42840 612824
rect 42668 612768 42840 612796
rect 42668 612756 42674 612768
rect 42610 612620 42616 612672
rect 42668 612660 42674 612672
rect 42794 612660 42800 612672
rect 42668 612632 42800 612660
rect 42668 612620 42674 612632
rect 42794 612620 42800 612632
rect 42852 612620 42858 612672
rect 673638 606704 673644 606756
rect 673696 606744 673702 606756
rect 675386 606744 675392 606756
rect 673696 606716 675392 606744
rect 673696 606704 673702 606716
rect 675386 606704 675392 606716
rect 675444 606704 675450 606756
rect 673546 606160 673552 606212
rect 673604 606200 673610 606212
rect 675018 606200 675024 606212
rect 673604 606172 675024 606200
rect 673604 606160 673610 606172
rect 675018 606160 675024 606172
rect 675076 606200 675082 606212
rect 675386 606200 675392 606212
rect 675076 606172 675392 606200
rect 675076 606160 675082 606172
rect 675386 606160 675392 606172
rect 675444 606160 675450 606212
rect 675202 600788 675208 600840
rect 675260 600828 675266 600840
rect 675386 600828 675392 600840
rect 675260 600800 675392 600828
rect 675260 600788 675266 600800
rect 675386 600788 675392 600800
rect 675444 600788 675450 600840
rect 673638 594872 673644 594924
rect 673696 594912 673702 594924
rect 673914 594912 673920 594924
rect 673696 594884 673920 594912
rect 673696 594872 673702 594884
rect 673914 594872 673920 594884
rect 673972 594912 673978 594924
rect 675386 594912 675392 594924
rect 673972 594884 675392 594912
rect 673972 594872 673978 594884
rect 675386 594872 675392 594884
rect 675444 594872 675450 594924
rect 673730 594736 673736 594788
rect 673788 594776 673794 594788
rect 675018 594776 675024 594788
rect 673788 594748 675024 594776
rect 673788 594736 673794 594748
rect 675018 594736 675024 594748
rect 675076 594736 675082 594788
rect 675294 593376 675300 593428
rect 675352 593376 675358 593428
rect 675312 593224 675340 593376
rect 675294 593172 675300 593224
rect 675352 593172 675358 593224
rect 673546 585148 673552 585200
rect 673604 585188 673610 585200
rect 673822 585188 673828 585200
rect 673604 585160 673828 585188
rect 673604 585148 673610 585160
rect 673822 585148 673828 585160
rect 673880 585148 673886 585200
rect 41782 583516 41788 583568
rect 41840 583556 41846 583568
rect 42334 583556 42340 583568
rect 41840 583528 42340 583556
rect 41840 583516 41846 583528
rect 42334 583516 42340 583528
rect 42392 583516 42398 583568
rect 41782 582632 41788 582684
rect 41840 582672 41846 582684
rect 42794 582672 42800 582684
rect 41840 582644 42800 582672
rect 41840 582632 41846 582644
rect 42794 582632 42800 582644
rect 42852 582632 42858 582684
rect 41782 576580 41788 576632
rect 41840 576620 41846 576632
rect 42334 576620 42340 576632
rect 41840 576592 42340 576620
rect 41840 576580 41846 576592
rect 42334 576580 42340 576592
rect 42392 576580 42398 576632
rect 673730 575424 673736 575476
rect 673788 575464 673794 575476
rect 674374 575464 674380 575476
rect 673788 575436 674380 575464
rect 673788 575424 673794 575436
rect 674374 575424 674380 575436
rect 674432 575424 674438 575476
rect 42334 574064 42340 574116
rect 42392 574104 42398 574116
rect 42794 574104 42800 574116
rect 42392 574076 42800 574104
rect 42392 574064 42398 574076
rect 42794 574064 42800 574076
rect 42852 574064 42858 574116
rect 41782 571208 41788 571260
rect 41840 571248 41846 571260
rect 42794 571248 42800 571260
rect 41840 571220 42800 571248
rect 41840 571208 41846 571220
rect 42794 571208 42800 571220
rect 42852 571208 42858 571260
rect 41782 570664 41788 570716
rect 41840 570704 41846 570716
rect 42518 570704 42524 570716
rect 41840 570676 42524 570704
rect 41840 570664 41846 570676
rect 42518 570664 42524 570676
rect 42576 570704 42582 570716
rect 42702 570704 42708 570716
rect 42576 570676 42708 570704
rect 42576 570664 42582 570676
rect 42702 570664 42708 570676
rect 42760 570664 42766 570716
rect 673546 560532 673552 560584
rect 673604 560572 673610 560584
rect 673822 560572 673828 560584
rect 673604 560544 673828 560572
rect 673604 560532 673610 560544
rect 673822 560532 673828 560544
rect 673880 560572 673886 560584
rect 675386 560572 675392 560584
rect 673880 560544 675392 560572
rect 673880 560532 673886 560544
rect 675386 560532 675392 560544
rect 675444 560532 675450 560584
rect 674006 559920 674012 559972
rect 674064 559960 674070 559972
rect 674374 559960 674380 559972
rect 674064 559932 674380 559960
rect 674064 559920 674070 559932
rect 674374 559920 674380 559932
rect 674432 559960 674438 559972
rect 675386 559960 675392 559972
rect 674432 559932 675392 559960
rect 674432 559920 674438 559932
rect 675386 559920 675392 559932
rect 675444 559920 675450 559972
rect 42610 554752 42616 554804
rect 42668 554792 42674 554804
rect 42794 554792 42800 554804
rect 42668 554764 42800 554792
rect 42668 554752 42674 554764
rect 42794 554752 42800 554764
rect 42852 554752 42858 554804
rect 673638 550468 673644 550520
rect 673696 550508 673702 550520
rect 675386 550508 675392 550520
rect 673696 550480 675392 550508
rect 673696 550468 673702 550480
rect 675386 550468 675392 550480
rect 675444 550468 675450 550520
rect 673546 546388 673552 546440
rect 673604 546388 673610 546440
rect 673564 546360 673592 546388
rect 673822 546360 673828 546372
rect 673564 546332 673828 546360
rect 673822 546320 673828 546332
rect 673880 546320 673886 546372
rect 41782 540336 41788 540388
rect 41840 540376 41846 540388
rect 42334 540376 42340 540388
rect 41840 540348 42340 540376
rect 41840 540336 41846 540348
rect 42334 540336 42340 540348
rect 42392 540336 42398 540388
rect 41782 539452 41788 539504
rect 41840 539492 41846 539504
rect 42518 539492 42524 539504
rect 41840 539464 42524 539492
rect 41840 539452 41846 539464
rect 42518 539452 42524 539464
rect 42576 539452 42582 539504
rect 41782 533400 41788 533452
rect 41840 533440 41846 533452
rect 42334 533440 42340 533452
rect 41840 533412 42340 533440
rect 41840 533400 41846 533412
rect 42334 533400 42340 533412
rect 42392 533400 42398 533452
rect 41782 528028 41788 528080
rect 41840 528068 41846 528080
rect 42610 528068 42616 528080
rect 41840 528040 42616 528068
rect 41840 528028 41846 528040
rect 42610 528028 42616 528040
rect 42668 528028 42674 528080
rect 41782 527484 41788 527536
rect 41840 527524 41846 527536
rect 42426 527524 42432 527536
rect 41840 527496 42432 527524
rect 41840 527484 41846 527496
rect 42426 527484 42432 527496
rect 42484 527524 42490 527536
rect 42702 527524 42708 527536
rect 42484 527496 42708 527524
rect 42484 527484 42490 527496
rect 42702 527484 42708 527496
rect 42760 527484 42766 527536
rect 675294 513748 675300 513800
rect 675352 513788 675358 513800
rect 677686 513788 677692 513800
rect 675352 513760 677692 513788
rect 675352 513748 675358 513760
rect 677686 513748 677692 513760
rect 677744 513748 677750 513800
rect 673730 502324 673736 502376
rect 673788 502364 673794 502376
rect 673914 502364 673920 502376
rect 673788 502336 673920 502364
rect 673788 502324 673794 502336
rect 673914 502324 673920 502336
rect 673972 502324 673978 502376
rect 673546 498176 673552 498228
rect 673604 498216 673610 498228
rect 673822 498216 673828 498228
rect 673604 498188 673828 498216
rect 673604 498176 673610 498188
rect 673822 498176 673828 498188
rect 673880 498176 673886 498228
rect 673822 469316 673828 469328
rect 673748 469288 673828 469316
rect 673748 469192 673776 469288
rect 673822 469276 673828 469288
rect 673880 469276 673886 469328
rect 673730 469140 673736 469192
rect 673788 469140 673794 469192
rect 673730 463632 673736 463684
rect 673788 463672 673794 463684
rect 674006 463672 674012 463684
rect 673788 463644 674012 463672
rect 673788 463632 673794 463644
rect 674006 463632 674012 463644
rect 674064 463632 674070 463684
rect 673546 449556 673552 449608
rect 673604 449596 673610 449608
rect 673822 449596 673828 449608
rect 673604 449568 673828 449596
rect 673604 449556 673610 449568
rect 673822 449556 673828 449568
rect 673880 449556 673886 449608
rect 42610 444320 42616 444372
rect 42668 444360 42674 444372
rect 42794 444360 42800 444372
rect 42668 444332 42800 444360
rect 42668 444320 42674 444332
rect 42794 444320 42800 444332
rect 42852 444320 42858 444372
rect 673730 444320 673736 444372
rect 673788 444360 673794 444372
rect 674006 444360 674012 444372
rect 673788 444332 674012 444360
rect 673788 444320 673794 444332
rect 674006 444320 674012 444332
rect 674064 444320 674070 444372
rect 42702 441532 42708 441584
rect 42760 441572 42766 441584
rect 42794 441572 42800 441584
rect 42760 441544 42800 441572
rect 42760 441532 42766 441544
rect 42794 441532 42800 441544
rect 42852 441532 42858 441584
rect 42610 422288 42616 422340
rect 42668 422328 42674 422340
rect 42702 422328 42708 422340
rect 42668 422300 42708 422328
rect 42668 422288 42674 422300
rect 42702 422288 42708 422300
rect 42760 422288 42766 422340
rect 673638 420724 673644 420776
rect 673696 420764 673702 420776
rect 673822 420764 673828 420776
rect 673696 420736 673828 420764
rect 673696 420724 673702 420736
rect 673822 420724 673828 420736
rect 673880 420724 673886 420776
rect 41782 412768 41788 412820
rect 41840 412808 41846 412820
rect 42334 412808 42340 412820
rect 41840 412780 42340 412808
rect 41840 412768 41846 412780
rect 42334 412768 42340 412780
rect 42392 412768 42398 412820
rect 41782 411204 41788 411256
rect 41840 411244 41846 411256
rect 42518 411244 42524 411256
rect 41840 411216 42524 411244
rect 41840 411204 41846 411216
rect 42518 411204 42524 411216
rect 42576 411204 42582 411256
rect 41782 405764 41788 405816
rect 41840 405804 41846 405816
rect 42334 405804 42340 405816
rect 41840 405776 42340 405804
rect 41840 405764 41846 405776
rect 42334 405764 42340 405776
rect 42392 405764 42398 405816
rect 42610 405696 42616 405748
rect 42668 405736 42674 405748
rect 42886 405736 42892 405748
rect 42668 405708 42892 405736
rect 42668 405696 42674 405708
rect 42886 405696 42892 405708
rect 42944 405696 42950 405748
rect 673822 401548 673828 401600
rect 673880 401588 673886 401600
rect 675294 401588 675300 401600
rect 673880 401560 675300 401588
rect 673880 401548 673886 401560
rect 675294 401548 675300 401560
rect 675352 401548 675358 401600
rect 41782 401344 41788 401396
rect 41840 401384 41846 401396
rect 42886 401384 42892 401396
rect 41840 401356 42892 401384
rect 41840 401344 41846 401356
rect 42886 401344 42892 401356
rect 42944 401344 42950 401396
rect 41782 400800 41788 400852
rect 41840 400840 41846 400852
rect 42426 400840 42432 400852
rect 41840 400812 42432 400840
rect 41840 400800 41846 400812
rect 42426 400800 42432 400812
rect 42484 400800 42490 400852
rect 42610 386316 42616 386368
rect 42668 386356 42674 386368
rect 42886 386356 42892 386368
rect 42668 386328 42892 386356
rect 42668 386316 42674 386328
rect 42886 386316 42892 386328
rect 42944 386316 42950 386368
rect 673730 384276 673736 384328
rect 673788 384316 673794 384328
rect 675386 384316 675392 384328
rect 673788 384288 675392 384316
rect 673788 384276 673794 384288
rect 675386 384276 675392 384288
rect 675444 384276 675450 384328
rect 673638 383188 673644 383240
rect 673696 383228 673702 383240
rect 675294 383228 675300 383240
rect 673696 383200 675300 383228
rect 673696 383188 673702 383200
rect 675294 383188 675300 383200
rect 675352 383188 675358 383240
rect 673546 380876 673552 380928
rect 673604 380916 673610 380928
rect 673730 380916 673736 380928
rect 673604 380888 673736 380916
rect 673604 380876 673610 380888
rect 673730 380876 673736 380888
rect 673788 380876 673794 380928
rect 42794 372580 42800 372632
rect 42852 372620 42858 372632
rect 42978 372620 42984 372632
rect 42852 372592 42984 372620
rect 42852 372580 42858 372592
rect 42978 372580 42984 372592
rect 43036 372580 43042 372632
rect 673730 372308 673736 372360
rect 673788 372348 673794 372360
rect 675386 372348 675392 372360
rect 673788 372320 675392 372348
rect 673788 372308 673794 372320
rect 675386 372308 675392 372320
rect 675444 372308 675450 372360
rect 41782 369520 41788 369572
rect 41840 369560 41846 369572
rect 42334 369560 42340 369572
rect 41840 369532 42340 369560
rect 41840 369520 41846 369532
rect 42334 369520 42340 369532
rect 42392 369520 42398 369572
rect 41782 368636 41788 368688
rect 41840 368676 41846 368688
rect 42886 368676 42892 368688
rect 41840 368648 42892 368676
rect 41840 368636 41846 368648
rect 42886 368636 42892 368648
rect 42944 368636 42950 368688
rect 42518 367820 42524 367872
rect 42576 367860 42582 367872
rect 42794 367860 42800 367872
rect 42576 367832 42800 367860
rect 42576 367820 42582 367832
rect 42794 367820 42800 367832
rect 42852 367820 42858 367872
rect 41782 362584 41788 362636
rect 41840 362624 41846 362636
rect 42334 362624 42340 362636
rect 41840 362596 42340 362624
rect 41840 362584 41846 362596
rect 42334 362584 42340 362596
rect 42392 362584 42398 362636
rect 41782 358232 41788 358284
rect 41840 358272 41846 358284
rect 42518 358272 42524 358284
rect 41840 358244 42524 358272
rect 41840 358232 41846 358244
rect 42518 358232 42524 358244
rect 42576 358232 42582 358284
rect 41782 357620 41788 357672
rect 41840 357660 41846 357672
rect 42426 357660 42432 357672
rect 41840 357632 42432 357660
rect 41840 357620 41846 357632
rect 42426 357620 42432 357632
rect 42484 357660 42490 357672
rect 42610 357660 42616 357672
rect 42484 357632 42616 357660
rect 42484 357620 42490 357632
rect 42610 357620 42616 357632
rect 42668 357620 42674 357672
rect 673546 338104 673552 338156
rect 673604 338144 673610 338156
rect 675386 338144 675392 338156
rect 673604 338116 675392 338144
rect 673604 338104 673610 338116
rect 675386 338104 675392 338116
rect 675444 338104 675450 338156
rect 673638 337492 673644 337544
rect 673696 337532 673702 337544
rect 675386 337532 675392 337544
rect 673696 337504 675392 337532
rect 673696 337492 673702 337504
rect 675386 337492 675392 337504
rect 675444 337492 675450 337544
rect 673730 328040 673736 328092
rect 673788 328080 673794 328092
rect 675386 328080 675392 328092
rect 673788 328052 675392 328080
rect 673788 328040 673794 328052
rect 675386 328040 675392 328052
rect 675444 328040 675450 328092
rect 41782 326340 41788 326392
rect 41840 326380 41846 326392
rect 42334 326380 42340 326392
rect 41840 326352 42340 326380
rect 41840 326340 41846 326352
rect 42334 326340 42340 326352
rect 42392 326340 42398 326392
rect 41782 325456 41788 325508
rect 41840 325496 41846 325508
rect 42426 325496 42432 325508
rect 41840 325468 42432 325496
rect 41840 325456 41846 325468
rect 42426 325456 42432 325468
rect 42484 325496 42490 325508
rect 42702 325496 42708 325508
rect 42484 325468 42708 325496
rect 42484 325456 42490 325468
rect 42702 325456 42708 325468
rect 42760 325456 42766 325508
rect 42426 322872 42432 322924
rect 42484 322912 42490 322924
rect 42484 322884 42748 322912
rect 42484 322872 42490 322884
rect 42720 322856 42748 322884
rect 42610 322804 42616 322856
rect 42668 322804 42674 322856
rect 42702 322804 42708 322856
rect 42760 322804 42766 322856
rect 42628 322776 42656 322804
rect 42886 322776 42892 322788
rect 42628 322748 42892 322776
rect 42886 322736 42892 322748
rect 42944 322736 42950 322788
rect 41782 319404 41788 319456
rect 41840 319444 41846 319456
rect 42334 319444 42340 319456
rect 41840 319416 42340 319444
rect 41840 319404 41846 319416
rect 42334 319404 42340 319416
rect 42392 319404 42398 319456
rect 42334 314168 42340 314220
rect 42392 314208 42398 314220
rect 42702 314208 42708 314220
rect 42392 314180 42708 314208
rect 42392 314168 42398 314180
rect 42702 314168 42708 314180
rect 42760 314168 42766 314220
rect 41782 314032 41788 314084
rect 41840 314072 41846 314084
rect 42518 314072 42524 314084
rect 41840 314044 42524 314072
rect 41840 314032 41846 314044
rect 42518 314032 42524 314044
rect 42576 314072 42582 314084
rect 42702 314072 42708 314084
rect 42576 314044 42708 314072
rect 42576 314032 42582 314044
rect 42702 314032 42708 314044
rect 42760 314032 42766 314084
rect 41782 313488 41788 313540
rect 41840 313488 41846 313540
rect 41800 313460 41828 313488
rect 42794 313460 42800 313472
rect 41800 313432 42800 313460
rect 42794 313420 42800 313432
rect 42852 313420 42858 313472
rect 673546 303560 673552 303612
rect 673604 303600 673610 303612
rect 675294 303600 675300 303612
rect 673604 303572 675300 303600
rect 673604 303560 673610 303572
rect 675294 303560 675300 303572
rect 675352 303560 675358 303612
rect 673638 293564 673644 293616
rect 673696 293604 673702 293616
rect 673914 293604 673920 293616
rect 673696 293576 673920 293604
rect 673696 293564 673702 293576
rect 673914 293564 673920 293576
rect 673972 293604 673978 293616
rect 675386 293604 675392 293616
rect 673972 293576 675392 293604
rect 673972 293564 673978 293576
rect 675386 293564 675392 293576
rect 675444 293564 675450 293616
rect 673638 293428 673644 293480
rect 673696 293468 673702 293480
rect 675294 293468 675300 293480
rect 673696 293440 675300 293468
rect 673696 293428 673702 293440
rect 675294 293428 675300 293440
rect 675352 293428 675358 293480
rect 41782 283160 41788 283212
rect 41840 283200 41846 283212
rect 42334 283200 42340 283212
rect 41840 283172 42340 283200
rect 41840 283160 41846 283172
rect 42334 283160 42340 283172
rect 42392 283160 42398 283212
rect 41782 282276 41788 282328
rect 41840 282316 41846 282328
rect 42518 282316 42524 282328
rect 41840 282288 42524 282316
rect 41840 282276 41846 282288
rect 42518 282276 42524 282288
rect 42576 282276 42582 282328
rect 673730 282072 673736 282124
rect 673788 282112 673794 282124
rect 675386 282112 675392 282124
rect 673788 282084 675392 282112
rect 673788 282072 673794 282084
rect 675386 282072 675392 282084
rect 675444 282072 675450 282124
rect 41782 276156 41788 276208
rect 41840 276196 41846 276208
rect 42334 276196 42340 276208
rect 41840 276168 42340 276196
rect 41840 276156 41846 276168
rect 42334 276156 42340 276168
rect 42392 276156 42398 276208
rect 41782 271872 41788 271924
rect 41840 271912 41846 271924
rect 42702 271912 42708 271924
rect 41840 271884 42708 271912
rect 41840 271872 41846 271884
rect 42702 271872 42708 271884
rect 42760 271872 42766 271924
rect 41782 271192 41788 271244
rect 41840 271232 41846 271244
rect 42518 271232 42524 271244
rect 41840 271204 42524 271232
rect 41840 271192 41846 271204
rect 42518 271192 42524 271204
rect 42576 271232 42582 271244
rect 42794 271232 42800 271244
rect 42576 271204 42800 271232
rect 42576 271192 42582 271204
rect 42794 271192 42800 271204
rect 42852 271192 42858 271244
rect 673454 264936 673460 264988
rect 673512 264976 673518 264988
rect 673638 264976 673644 264988
rect 673512 264948 673644 264976
rect 673512 264936 673518 264948
rect 673638 264936 673644 264948
rect 673696 264936 673702 264988
rect 673454 248684 673460 248736
rect 673512 248724 673518 248736
rect 675294 248724 675300 248736
rect 673512 248696 675300 248724
rect 673512 248684 673518 248696
rect 675294 248684 675300 248696
rect 675352 248684 675358 248736
rect 673638 247460 673644 247512
rect 673696 247500 673702 247512
rect 673914 247500 673920 247512
rect 673696 247472 673920 247500
rect 673696 247460 673702 247472
rect 673914 247460 673920 247472
rect 673972 247500 673978 247512
rect 675386 247500 675392 247512
rect 673972 247472 675392 247500
rect 673972 247460 673978 247472
rect 675386 247460 675392 247472
rect 675444 247460 675450 247512
rect 42334 245556 42340 245608
rect 42392 245596 42398 245608
rect 42886 245596 42892 245608
rect 42392 245568 42892 245596
rect 42392 245556 42398 245568
rect 42886 245556 42892 245568
rect 42944 245556 42950 245608
rect 42518 245488 42524 245540
rect 42576 245528 42582 245540
rect 42794 245528 42800 245540
rect 42576 245500 42800 245528
rect 42576 245488 42582 245500
rect 42794 245488 42800 245500
rect 42852 245488 42858 245540
rect 673822 243788 673828 243840
rect 673880 243828 673886 243840
rect 675294 243828 675300 243840
rect 673880 243800 675300 243828
rect 673880 243788 673886 243800
rect 675294 243788 675300 243800
rect 675352 243788 675358 243840
rect 41782 239912 41788 239964
rect 41840 239952 41846 239964
rect 42334 239952 42340 239964
rect 41840 239924 42340 239952
rect 41840 239912 41846 239924
rect 42334 239912 42340 239924
rect 42392 239912 42398 239964
rect 41782 238076 41788 238128
rect 41840 238116 41846 238128
rect 42610 238116 42616 238128
rect 41840 238088 42616 238116
rect 41840 238076 41846 238088
rect 42610 238076 42616 238088
rect 42668 238116 42674 238128
rect 42886 238116 42892 238128
rect 42668 238088 42892 238116
rect 42668 238076 42674 238088
rect 42886 238076 42892 238088
rect 42944 238076 42950 238128
rect 673914 237668 673920 237720
rect 673972 237708 673978 237720
rect 675386 237708 675392 237720
rect 673972 237680 675392 237708
rect 673972 237668 673978 237680
rect 675386 237668 675392 237680
rect 675444 237668 675450 237720
rect 673914 237328 673920 237380
rect 673972 237368 673978 237380
rect 674098 237368 674104 237380
rect 673972 237340 674104 237368
rect 673972 237328 673978 237340
rect 674098 237328 674104 237340
rect 674156 237328 674162 237380
rect 41782 232976 41788 233028
rect 41840 233016 41846 233028
rect 42334 233016 42340 233028
rect 41840 232988 42340 233016
rect 41840 232976 41846 232988
rect 42334 232976 42340 232988
rect 42392 232976 42398 233028
rect 42334 232840 42340 232892
rect 42392 232880 42398 232892
rect 42610 232880 42616 232892
rect 42392 232852 42616 232880
rect 42392 232840 42398 232852
rect 42610 232840 42616 232852
rect 42668 232840 42674 232892
rect 674098 231752 674104 231804
rect 674156 231792 674162 231804
rect 674282 231792 674288 231804
rect 674156 231764 674288 231792
rect 674156 231752 674162 231764
rect 674282 231752 674288 231764
rect 674340 231752 674346 231804
rect 41782 228624 41788 228676
rect 41840 228664 41846 228676
rect 42702 228664 42708 228676
rect 41840 228636 42708 228664
rect 41840 228624 41846 228636
rect 42702 228624 42708 228636
rect 42760 228624 42766 228676
rect 41782 228012 41788 228064
rect 41840 228052 41846 228064
rect 42610 228052 42616 228064
rect 41840 228024 42616 228052
rect 41840 228012 41846 228024
rect 42610 228012 42616 228024
rect 42668 228052 42674 228064
rect 42794 228052 42800 228064
rect 42668 228024 42800 228052
rect 42668 228012 42674 228024
rect 42794 228012 42800 228024
rect 42852 228012 42858 228064
rect 673822 218084 673828 218136
rect 673880 218084 673886 218136
rect 673840 218000 673868 218084
rect 673822 217948 673828 218000
rect 673880 217948 673886 218000
rect 673730 212508 673736 212560
rect 673788 212548 673794 212560
rect 673822 212548 673828 212560
rect 673788 212520 673828 212548
rect 673788 212508 673794 212520
rect 673822 212508 673828 212520
rect 673880 212508 673886 212560
rect 674006 212508 674012 212560
rect 674064 212548 674070 212560
rect 674282 212548 674288 212560
rect 674064 212520 674288 212548
rect 674064 212508 674070 212520
rect 674282 212508 674288 212520
rect 674340 212508 674346 212560
rect 42334 208360 42340 208412
rect 42392 208400 42398 208412
rect 42886 208400 42892 208412
rect 42392 208372 42892 208400
rect 42392 208360 42398 208372
rect 42886 208360 42892 208372
rect 42944 208360 42950 208412
rect 673730 203872 673736 203924
rect 673788 203912 673794 203924
rect 675386 203912 675392 203924
rect 673788 203884 675392 203912
rect 673788 203872 673794 203884
rect 675386 203872 675392 203884
rect 675444 203872 675450 203924
rect 673638 203328 673644 203380
rect 673696 203368 673702 203380
rect 675386 203368 675392 203380
rect 673696 203340 675392 203368
rect 673696 203328 673702 203340
rect 675386 203328 675392 203340
rect 675444 203328 675450 203380
rect 674006 198704 674012 198756
rect 674064 198744 674070 198756
rect 675202 198744 675208 198756
rect 674064 198716 675208 198744
rect 674064 198704 674070 198716
rect 675202 198704 675208 198716
rect 675260 198704 675266 198756
rect 41782 196732 41788 196784
rect 41840 196772 41846 196784
rect 42334 196772 42340 196784
rect 41840 196744 42340 196772
rect 41840 196732 41846 196744
rect 42334 196732 42340 196744
rect 42392 196732 42398 196784
rect 41782 194896 41788 194948
rect 41840 194936 41846 194948
rect 42426 194936 42432 194948
rect 41840 194908 42432 194936
rect 41840 194896 41846 194908
rect 42426 194896 42432 194908
rect 42484 194936 42490 194948
rect 42886 194936 42892 194948
rect 42484 194908 42892 194936
rect 42484 194896 42490 194908
rect 42886 194896 42892 194908
rect 42944 194896 42950 194948
rect 674742 192108 674748 192160
rect 674800 192148 674806 192160
rect 675202 192148 675208 192160
rect 674800 192120 675208 192148
rect 674800 192108 674806 192120
rect 675202 192108 675208 192120
rect 675260 192148 675266 192160
rect 675386 192148 675392 192160
rect 675260 192120 675392 192148
rect 675260 192108 675266 192120
rect 675386 192108 675392 192120
rect 675444 192108 675450 192160
rect 41782 189796 41788 189848
rect 41840 189836 41846 189848
rect 42334 189836 42340 189848
rect 41840 189808 42340 189836
rect 41840 189796 41846 189808
rect 42334 189796 42340 189808
rect 42392 189796 42398 189848
rect 41782 185444 41788 185496
rect 41840 185484 41846 185496
rect 42334 185484 42340 185496
rect 41840 185456 42340 185484
rect 41840 185444 41846 185456
rect 42334 185444 42340 185456
rect 42392 185484 42398 185496
rect 42702 185484 42708 185496
rect 42392 185456 42708 185484
rect 42392 185444 42398 185456
rect 42702 185444 42708 185456
rect 42760 185444 42766 185496
rect 42426 185308 42432 185360
rect 42484 185348 42490 185360
rect 42702 185348 42708 185360
rect 42484 185320 42708 185348
rect 42484 185308 42490 185320
rect 42702 185308 42708 185320
rect 42760 185308 42766 185360
rect 41782 184832 41788 184884
rect 41840 184872 41846 184884
rect 42426 184872 42432 184884
rect 41840 184844 42432 184872
rect 41840 184832 41846 184844
rect 42426 184832 42432 184844
rect 42484 184872 42490 184884
rect 42610 184872 42616 184884
rect 42484 184844 42616 184872
rect 42484 184832 42490 184844
rect 42610 184832 42616 184844
rect 42668 184832 42674 184884
rect 673822 173884 673828 173936
rect 673880 173924 673886 173936
rect 674742 173924 674748 173936
rect 673880 173896 674748 173924
rect 673880 173884 673886 173896
rect 674742 173884 674748 173896
rect 674800 173884 674806 173936
rect 673546 158312 673552 158364
rect 673604 158352 673610 158364
rect 675386 158352 675392 158364
rect 673604 158324 675392 158352
rect 673604 158312 673610 158324
rect 675386 158312 675392 158324
rect 675444 158312 675450 158364
rect 673454 157292 673460 157344
rect 673512 157332 673518 157344
rect 675386 157332 675392 157344
rect 673512 157304 675392 157332
rect 673512 157292 673518 157304
rect 675386 157292 675392 157304
rect 675444 157292 675450 157344
rect 42518 149064 42524 149116
rect 42576 149104 42582 149116
rect 42702 149104 42708 149116
rect 42576 149076 42708 149104
rect 42576 149064 42582 149076
rect 42702 149064 42708 149076
rect 42760 149064 42766 149116
rect 673638 147092 673644 147144
rect 673696 147132 673702 147144
rect 675018 147132 675024 147144
rect 673696 147104 675024 147132
rect 673696 147092 673702 147104
rect 675018 147092 675024 147104
rect 675076 147132 675082 147144
rect 675386 147132 675392 147144
rect 675076 147104 675392 147132
rect 675076 147092 675082 147104
rect 675386 147092 675392 147104
rect 675444 147092 675450 147144
rect 674006 140632 674012 140684
rect 674064 140672 674070 140684
rect 675018 140672 675024 140684
rect 674064 140644 675024 140672
rect 674064 140632 674070 140644
rect 675018 140632 675024 140644
rect 675076 140632 675082 140684
rect 42242 121456 42248 121508
rect 42300 121496 42306 121508
rect 44726 121496 44732 121508
rect 42300 121468 44732 121496
rect 42300 121456 42306 121468
rect 44726 121456 44732 121468
rect 44784 121456 44790 121508
rect 673822 115948 673828 116000
rect 673880 115988 673886 116000
rect 674006 115988 674012 116000
rect 673880 115960 674012 115988
rect 673880 115948 673886 115960
rect 674006 115948 674012 115960
rect 674064 115948 674070 116000
rect 42978 115880 42984 115932
rect 43036 115920 43042 115932
rect 44726 115920 44732 115932
rect 43036 115892 44732 115920
rect 43036 115880 43042 115892
rect 44726 115880 44732 115892
rect 44784 115880 44790 115932
rect 673822 115812 673828 115864
rect 673880 115852 673886 115864
rect 675018 115852 675024 115864
rect 673880 115824 675024 115852
rect 673880 115812 673886 115824
rect 675018 115812 675024 115824
rect 675076 115812 675082 115864
rect 673546 112752 673552 112804
rect 673604 112792 673610 112804
rect 675386 112792 675392 112804
rect 673604 112764 675392 112792
rect 673604 112752 673610 112764
rect 675386 112752 675392 112764
rect 675444 112752 675450 112804
rect 673454 112072 673460 112124
rect 673512 112112 673518 112124
rect 675386 112112 675392 112124
rect 673512 112084 675392 112112
rect 673512 112072 673518 112084
rect 675386 112072 675392 112084
rect 675444 112072 675450 112124
rect 42518 110440 42524 110492
rect 42576 110480 42582 110492
rect 42702 110480 42708 110492
rect 42576 110452 42708 110480
rect 42576 110440 42582 110452
rect 42702 110440 42708 110452
rect 42760 110440 42766 110492
rect 673638 102280 673644 102332
rect 673696 102320 673702 102332
rect 675018 102320 675024 102332
rect 673696 102292 675024 102320
rect 673696 102280 673702 102292
rect 675018 102280 675024 102292
rect 675076 102320 675082 102332
rect 675386 102320 675392 102332
rect 675076 102292 675392 102320
rect 675076 102280 675082 102292
rect 675386 102280 675392 102292
rect 675444 102280 675450 102332
rect 44634 82832 44640 82884
rect 44692 82832 44698 82884
rect 44652 82804 44680 82832
rect 44818 82804 44824 82816
rect 44652 82776 44824 82804
rect 44818 82764 44824 82776
rect 44876 82764 44882 82816
rect 42334 45704 42340 45756
rect 42392 45744 42398 45756
rect 140958 45744 140964 45756
rect 42392 45716 140964 45744
rect 42392 45704 42398 45716
rect 140958 45704 140964 45716
rect 141016 45704 141022 45756
rect 42426 45636 42432 45688
rect 42484 45676 42490 45688
rect 143626 45676 143632 45688
rect 42484 45648 143632 45676
rect 42484 45636 42490 45648
rect 143626 45636 143632 45648
rect 143684 45636 143690 45688
rect 42702 45568 42708 45620
rect 42760 45608 42766 45620
rect 143534 45608 143540 45620
rect 42760 45580 143540 45608
rect 42760 45568 42766 45580
rect 143534 45568 143540 45580
rect 143592 45568 143598 45620
rect 527450 45568 527456 45620
rect 527508 45608 527514 45620
rect 673546 45608 673552 45620
rect 527508 45580 673552 45608
rect 527508 45568 527514 45580
rect 673546 45568 673552 45580
rect 673604 45568 673610 45620
rect 44910 45500 44916 45552
rect 44968 45540 44974 45552
rect 195974 45540 195980 45552
rect 44968 45512 195980 45540
rect 44968 45500 44974 45512
rect 195974 45500 195980 45512
rect 196032 45500 196038 45552
rect 516318 45500 516324 45552
rect 516376 45540 516382 45552
rect 673638 45540 673644 45552
rect 516376 45512 673644 45540
rect 516376 45500 516382 45512
rect 673638 45500 673644 45512
rect 673696 45500 673702 45552
rect 405642 44752 405648 44804
rect 405700 44792 405706 44804
rect 411254 44792 411260 44804
rect 405700 44764 411260 44792
rect 405700 44752 405706 44764
rect 411254 44752 411260 44764
rect 411312 44752 411318 44804
rect 359366 44724 359372 44736
rect 342272 44696 359372 44724
rect 195974 44412 195980 44464
rect 196032 44452 196038 44464
rect 304534 44452 304540 44464
rect 196032 44424 304540 44452
rect 196032 44412 196038 44424
rect 304534 44412 304540 44424
rect 304592 44452 304598 44464
rect 342272 44452 342300 44696
rect 359366 44684 359372 44696
rect 359424 44684 359430 44736
rect 406746 44684 406752 44736
rect 406804 44724 406810 44736
rect 406804 44696 411300 44724
rect 406804 44684 406810 44696
rect 411272 44588 411300 44696
rect 425054 44684 425060 44736
rect 425112 44724 425118 44736
rect 444190 44724 444196 44736
rect 425112 44696 444196 44724
rect 425112 44684 425118 44696
rect 444190 44684 444196 44696
rect 444248 44684 444254 44736
rect 483014 44656 483020 44668
rect 473280 44628 483020 44656
rect 425054 44588 425060 44600
rect 411272 44560 425060 44588
rect 425054 44548 425060 44560
rect 425112 44548 425118 44600
rect 461486 44588 461492 44600
rect 449820 44560 461492 44588
rect 354398 44480 354404 44532
rect 354456 44520 354462 44532
rect 360562 44520 360568 44532
rect 354456 44492 360568 44520
rect 354456 44480 354462 44492
rect 360562 44480 360568 44492
rect 360620 44480 360626 44532
rect 360654 44480 360660 44532
rect 360712 44520 360718 44532
rect 386414 44520 386420 44532
rect 360712 44492 386420 44520
rect 360712 44480 360718 44492
rect 386414 44480 386420 44492
rect 386472 44480 386478 44532
rect 399662 44480 399668 44532
rect 399720 44520 399726 44532
rect 406746 44520 406752 44532
rect 399720 44492 406752 44520
rect 399720 44480 399726 44492
rect 406746 44480 406752 44492
rect 406804 44480 406810 44532
rect 411254 44480 411260 44532
rect 411312 44520 411318 44532
rect 411312 44492 414244 44520
rect 411312 44480 411318 44492
rect 414216 44464 414244 44492
rect 444282 44480 444288 44532
rect 444340 44520 444346 44532
rect 449820 44520 449848 44560
rect 461486 44548 461492 44560
rect 461544 44588 461550 44600
rect 469122 44588 469128 44600
rect 461544 44560 469128 44588
rect 461544 44548 461550 44560
rect 469122 44548 469128 44560
rect 469180 44548 469186 44600
rect 469214 44548 469220 44600
rect 469272 44588 469278 44600
rect 473280 44588 473308 44628
rect 483014 44616 483020 44628
rect 483072 44616 483078 44668
rect 469272 44560 473308 44588
rect 502260 44560 502380 44588
rect 469272 44548 469278 44560
rect 502260 44532 502288 44560
rect 444340 44492 449848 44520
rect 444340 44480 444346 44492
rect 502242 44480 502248 44532
rect 502300 44480 502306 44532
rect 502352 44520 502380 44560
rect 516318 44520 516324 44532
rect 502352 44492 516324 44520
rect 516318 44480 516324 44492
rect 516376 44480 516382 44532
rect 304592 44424 342300 44452
rect 304592 44412 304598 44424
rect 414198 44412 414204 44464
rect 414256 44452 414262 44464
rect 419810 44452 419816 44464
rect 414256 44424 419816 44452
rect 414256 44412 414262 44424
rect 419810 44412 419816 44424
rect 419868 44412 419874 44464
rect 143626 44344 143632 44396
rect 143684 44384 143690 44396
rect 145098 44384 145104 44396
rect 143684 44356 145104 44384
rect 143684 44344 143690 44356
rect 145098 44344 145104 44356
rect 145156 44384 145162 44396
rect 195330 44384 195336 44396
rect 145156 44356 195336 44384
rect 145156 44344 145162 44356
rect 195330 44344 195336 44356
rect 195388 44384 195394 44396
rect 199654 44384 199660 44396
rect 195388 44356 199660 44384
rect 195388 44344 195394 44356
rect 199654 44344 199660 44356
rect 199712 44344 199718 44396
rect 200850 44344 200856 44396
rect 200908 44384 200914 44396
rect 241330 44384 241336 44396
rect 200908 44356 241336 44384
rect 200908 44344 200914 44356
rect 241330 44344 241336 44356
rect 241388 44384 241394 44396
rect 251082 44384 251088 44396
rect 241388 44356 251088 44384
rect 241388 44344 241394 44356
rect 251082 44344 251088 44356
rect 251140 44344 251146 44396
rect 306374 44344 306380 44396
rect 306432 44384 306438 44396
rect 309410 44384 309416 44396
rect 306432 44356 309416 44384
rect 306432 44344 306438 44356
rect 309410 44344 309416 44356
rect 309468 44384 309474 44396
rect 352558 44384 352564 44396
rect 309468 44356 352564 44384
rect 309468 44344 309474 44356
rect 352558 44344 352564 44356
rect 352616 44384 352622 44396
rect 355410 44384 355416 44396
rect 352616 44356 355416 44384
rect 352616 44344 352622 44356
rect 355410 44344 355416 44356
rect 355468 44344 355474 44396
rect 359366 44344 359372 44396
rect 359424 44384 359430 44396
rect 360654 44384 360660 44396
rect 359424 44356 360660 44384
rect 359424 44344 359430 44356
rect 360654 44344 360660 44356
rect 360712 44344 360718 44396
rect 364242 44344 364248 44396
rect 364300 44384 364306 44396
rect 407390 44384 407396 44396
rect 364300 44356 407396 44384
rect 364300 44344 364306 44356
rect 407390 44344 407396 44356
rect 407448 44384 407454 44396
rect 410426 44384 410432 44396
rect 407448 44356 410432 44384
rect 407448 44344 407454 44356
rect 410426 44344 410432 44356
rect 410484 44344 410490 44396
rect 419074 44344 419080 44396
rect 419132 44384 419138 44396
rect 462130 44384 462136 44396
rect 419132 44356 462136 44384
rect 419132 44344 419138 44356
rect 462130 44344 462136 44356
rect 462188 44384 462194 44396
rect 465166 44384 465172 44396
rect 462188 44356 465172 44384
rect 462188 44344 462194 44356
rect 465166 44344 465172 44356
rect 465224 44344 465230 44396
rect 473814 44344 473820 44396
rect 473872 44384 473878 44396
rect 516962 44384 516968 44396
rect 473872 44356 516968 44384
rect 473872 44344 473878 44356
rect 516962 44344 516968 44356
rect 517020 44384 517026 44396
rect 519998 44384 520004 44396
rect 517020 44356 520004 44384
rect 517020 44344 517026 44356
rect 519998 44344 520004 44356
rect 520056 44344 520062 44396
rect 188522 44276 188528 44328
rect 188580 44316 188586 44328
rect 192846 44316 192852 44328
rect 188580 44288 192852 44316
rect 188580 44276 188586 44288
rect 192846 44276 192852 44288
rect 192904 44316 192910 44328
rect 201494 44316 201500 44328
rect 192904 44288 201500 44316
rect 192904 44276 192910 44288
rect 201494 44276 201500 44288
rect 201552 44316 201558 44328
rect 297082 44316 297088 44328
rect 201552 44288 297088 44316
rect 201552 44276 201558 44288
rect 297082 44276 297088 44288
rect 297140 44316 297146 44328
rect 299566 44316 299572 44328
rect 297140 44288 299572 44316
rect 297140 44276 297146 44288
rect 299566 44276 299572 44288
rect 299624 44316 299630 44328
rect 305730 44316 305736 44328
rect 299624 44288 305736 44316
rect 299624 44276 299630 44288
rect 305730 44276 305736 44288
rect 305788 44316 305794 44328
rect 351914 44316 351920 44328
rect 305788 44288 351920 44316
rect 305788 44276 305794 44288
rect 351914 44276 351920 44288
rect 351972 44316 351978 44328
rect 354398 44316 354404 44328
rect 351972 44288 354404 44316
rect 351972 44276 351978 44288
rect 354398 44276 354404 44288
rect 354456 44276 354462 44328
rect 358722 44316 358728 44328
rect 355520 44288 358728 44316
rect 186682 44208 186688 44260
rect 186740 44248 186746 44260
rect 194686 44248 194692 44260
rect 186740 44220 194692 44248
rect 186740 44208 186746 44220
rect 194686 44208 194692 44220
rect 194744 44208 194750 44260
rect 199654 44208 199660 44260
rect 199712 44248 199718 44260
rect 303890 44248 303896 44260
rect 199712 44220 303896 44248
rect 199712 44208 199718 44220
rect 303890 44208 303896 44220
rect 303948 44248 303954 44260
rect 308214 44248 308220 44260
rect 303948 44220 308220 44248
rect 303948 44208 303954 44220
rect 308214 44208 308220 44220
rect 308272 44248 308278 44260
rect 355520 44248 355548 44288
rect 358722 44276 358728 44288
rect 358780 44276 358786 44328
rect 360562 44276 360568 44328
rect 360620 44316 360626 44328
rect 399662 44316 399668 44328
rect 360620 44288 399668 44316
rect 360620 44276 360626 44288
rect 399662 44276 399668 44288
rect 399720 44276 399726 44328
rect 413554 44316 413560 44328
rect 399772 44288 413560 44316
rect 308272 44220 355548 44248
rect 308272 44208 308278 44220
rect 355594 44208 355600 44260
rect 355652 44248 355658 44260
rect 359918 44248 359924 44260
rect 355652 44220 359924 44248
rect 355652 44208 355658 44220
rect 359918 44208 359924 44220
rect 359976 44208 359982 44260
rect 363046 44208 363052 44260
rect 363104 44248 363110 44260
rect 399772 44248 399800 44288
rect 413554 44276 413560 44288
rect 413612 44316 413618 44328
rect 417878 44316 417884 44328
rect 413612 44288 417884 44316
rect 413612 44276 413618 44288
rect 417878 44276 417884 44288
rect 417936 44316 417942 44328
rect 468294 44316 468300 44328
rect 417936 44288 468300 44316
rect 417936 44276 417942 44288
rect 468294 44276 468300 44288
rect 468352 44316 468358 44328
rect 472618 44316 472624 44328
rect 468352 44288 472624 44316
rect 468352 44276 468358 44288
rect 472618 44276 472624 44288
rect 472676 44316 472682 44328
rect 523126 44316 523132 44328
rect 472676 44288 523132 44316
rect 472676 44276 472682 44288
rect 523126 44276 523132 44288
rect 523184 44276 523190 44328
rect 363104 44220 399800 44248
rect 363104 44208 363110 44220
rect 411070 44208 411076 44260
rect 411128 44248 411134 44260
rect 419718 44248 419724 44260
rect 411128 44220 419724 44248
rect 411128 44208 411134 44220
rect 419718 44208 419724 44220
rect 419776 44208 419782 44260
rect 419810 44208 419816 44260
rect 419868 44248 419874 44260
rect 468938 44248 468944 44260
rect 419868 44220 468944 44248
rect 419868 44208 419874 44220
rect 468938 44208 468944 44220
rect 468996 44248 469002 44260
rect 523770 44248 523776 44260
rect 468996 44220 523776 44248
rect 468996 44208 469002 44220
rect 523770 44208 523776 44220
rect 523828 44208 523834 44260
rect 295242 44140 295248 44192
rect 295300 44180 295306 44192
rect 303246 44180 303252 44192
rect 295300 44152 303252 44180
rect 295300 44140 295306 44152
rect 303246 44140 303252 44152
rect 303304 44140 303310 44192
rect 350074 44140 350080 44192
rect 350132 44180 350138 44192
rect 358078 44180 358084 44192
rect 350132 44152 358084 44180
rect 350132 44140 350138 44152
rect 358078 44140 358084 44152
rect 358136 44140 358142 44192
rect 358722 44140 358728 44192
rect 358780 44180 358786 44192
rect 363064 44180 363092 44208
rect 358780 44152 363092 44180
rect 358780 44140 358786 44152
rect 404906 44140 404912 44192
rect 404964 44180 404970 44192
rect 412910 44180 412916 44192
rect 404964 44152 412916 44180
rect 404964 44140 404970 44152
rect 412910 44140 412916 44152
rect 412968 44140 412974 44192
rect 459646 44140 459652 44192
rect 459704 44180 459710 44192
rect 467650 44180 467656 44192
rect 459704 44152 467656 44180
rect 459704 44140 459710 44152
rect 467650 44140 467656 44152
rect 467708 44140 467714 44192
rect 514478 44140 514484 44192
rect 514536 44180 514542 44192
rect 522482 44180 522488 44192
rect 514536 44152 522488 44180
rect 514536 44140 514542 44152
rect 522482 44140 522488 44152
rect 522540 44140 522546 44192
rect 523126 44140 523132 44192
rect 523184 44180 523190 44192
rect 527450 44180 527456 44192
rect 523184 44152 527456 44180
rect 523184 44140 523190 44152
rect 527450 44140 527456 44152
rect 527508 44140 527514 44192
rect 576762 42712 576768 42764
rect 576820 42752 576826 42764
rect 673454 42752 673460 42764
rect 576820 42724 673460 42752
rect 576820 42712 576826 42724
rect 673454 42712 673460 42724
rect 673512 42712 673518 42764
rect 251082 42032 251088 42084
rect 251140 42072 251146 42084
rect 255222 42072 255228 42084
rect 251140 42044 255228 42072
rect 251140 42032 251146 42044
rect 255222 42032 255228 42044
rect 255280 42032 255286 42084
rect 146294 41964 146300 42016
rect 146352 42004 146358 42016
rect 569126 42004 569132 42016
rect 146352 41976 569132 42004
rect 146352 41964 146358 41976
rect 569126 41964 569132 41976
rect 569184 42004 569190 42016
rect 576762 42004 576768 42016
rect 569184 41976 576768 42004
rect 569184 41964 569190 41976
rect 576762 41964 576768 41976
rect 576820 41964 576826 42016
rect 187694 41896 187700 41948
rect 187752 41936 187758 41948
rect 188430 41936 188436 41948
rect 187752 41908 188436 41936
rect 187752 41896 187758 41908
rect 188430 41896 188436 41908
rect 188488 41896 188494 41948
rect 198918 41896 198924 41948
rect 198976 41936 198982 41948
rect 307478 41936 307484 41948
rect 198976 41908 307484 41936
rect 198976 41896 198982 41908
rect 198458 41828 198464 41880
rect 198516 41868 198522 41880
rect 200114 41868 200120 41880
rect 198516 41840 200120 41868
rect 198516 41828 198522 41840
rect 200114 41828 200120 41840
rect 200172 41828 200178 41880
rect 255222 41828 255228 41880
rect 255280 41868 255286 41880
rect 297634 41868 297640 41880
rect 255280 41840 297640 41868
rect 255280 41828 255286 41840
rect 297634 41828 297640 41840
rect 297692 41868 297698 41880
rect 300670 41868 300676 41880
rect 297692 41840 300676 41868
rect 297692 41828 297698 41840
rect 300670 41828 300676 41840
rect 300728 41828 300734 41880
rect 149606 41760 149612 41812
rect 149664 41800 149670 41812
rect 187694 41800 187700 41812
rect 149664 41772 187700 41800
rect 149664 41760 149670 41772
rect 187694 41760 187700 41772
rect 187752 41760 187758 41812
rect 189258 41760 189264 41812
rect 189316 41800 189322 41812
rect 191098 41800 191104 41812
rect 189316 41772 191104 41800
rect 189316 41760 189322 41772
rect 191098 41760 191104 41772
rect 191156 41800 191162 41812
rect 192294 41800 192300 41812
rect 191156 41772 192300 41800
rect 191156 41760 191162 41772
rect 192294 41760 192300 41772
rect 192352 41800 192358 41812
rect 193582 41800 193588 41812
rect 192352 41772 193588 41800
rect 192352 41760 192358 41772
rect 193582 41760 193588 41772
rect 193640 41800 193646 41812
rect 196434 41800 196440 41812
rect 193640 41772 196440 41800
rect 193640 41760 193646 41772
rect 196434 41760 196440 41772
rect 196492 41760 196498 41812
rect 198826 41800 198832 41812
rect 198752 41772 198832 41800
rect 168282 41732 168288 41744
rect 160020 41704 168288 41732
rect 160020 41664 160048 41704
rect 168282 41692 168288 41704
rect 168340 41692 168346 41744
rect 154500 41636 160048 41664
rect 93762 41556 93768 41608
rect 93820 41596 93826 41608
rect 93820 41568 102180 41596
rect 93820 41556 93826 41568
rect 102152 41528 102180 41568
rect 121546 41556 121552 41608
rect 121604 41596 121610 41608
rect 121604 41568 135300 41596
rect 121604 41556 121610 41568
rect 121270 41528 121276 41540
rect 102152 41500 121276 41528
rect 121270 41488 121276 41500
rect 121328 41488 121334 41540
rect 135272 41528 135300 41568
rect 140866 41556 140872 41608
rect 140924 41596 140930 41608
rect 154500 41596 154528 41636
rect 140924 41568 154528 41596
rect 140924 41556 140930 41568
rect 140682 41528 140688 41540
rect 135272 41500 140688 41528
rect 140682 41488 140688 41500
rect 140740 41488 140746 41540
rect 168282 41488 168288 41540
rect 168340 41528 168346 41540
rect 198752 41528 198780 41772
rect 198826 41760 198832 41772
rect 198884 41760 198890 41812
rect 302234 41760 302240 41812
rect 302292 41800 302298 41812
rect 304994 41800 305000 41812
rect 302292 41772 305000 41800
rect 302292 41760 302298 41772
rect 304994 41760 305000 41772
rect 305052 41800 305058 41812
rect 306282 41800 306288 41812
rect 305052 41772 306288 41800
rect 305052 41760 305058 41772
rect 306282 41760 306288 41772
rect 306340 41760 306346 41812
rect 307404 41732 307432 41908
rect 307478 41896 307484 41908
rect 307536 41896 307542 41948
rect 362494 41896 362500 41948
rect 362552 41936 362558 41948
rect 367094 41936 367100 41948
rect 362552 41908 367100 41936
rect 362552 41896 362558 41908
rect 367094 41896 367100 41908
rect 367152 41896 367158 41948
rect 360010 41828 360016 41880
rect 360068 41868 360074 41880
rect 361114 41868 361120 41880
rect 360068 41840 361120 41868
rect 360068 41828 360074 41840
rect 361114 41828 361120 41840
rect 361172 41868 361178 41880
rect 363506 41868 363512 41880
rect 361172 41840 363512 41868
rect 361172 41828 361178 41840
rect 363506 41828 363512 41840
rect 363564 41828 363570 41880
rect 410518 41828 410524 41880
rect 410576 41868 410582 41880
rect 411806 41868 411812 41880
rect 410576 41840 411812 41868
rect 410576 41828 410582 41840
rect 411806 41828 411812 41840
rect 411864 41868 411870 41880
rect 414842 41868 414848 41880
rect 411864 41840 414848 41868
rect 411864 41828 411870 41840
rect 414842 41828 414848 41840
rect 414900 41868 414906 41880
rect 416130 41868 416136 41880
rect 414900 41840 416136 41868
rect 414900 41828 414906 41840
rect 416130 41828 416136 41840
rect 416188 41868 416194 41880
rect 418522 41868 418528 41880
rect 416188 41840 418528 41868
rect 416188 41828 416194 41840
rect 418522 41828 418528 41840
rect 418580 41828 418586 41880
rect 464154 41828 464160 41880
rect 464212 41868 464218 41880
rect 467190 41868 467196 41880
rect 464212 41840 467196 41868
rect 464212 41828 464218 41840
rect 467190 41828 467196 41840
rect 467248 41868 467254 41880
rect 470042 41868 470048 41880
rect 467248 41840 470048 41868
rect 467248 41828 467254 41840
rect 470042 41828 470048 41840
rect 470100 41828 470106 41880
rect 470962 41868 470968 41880
rect 470152 41840 470968 41868
rect 409322 41760 409328 41812
rect 409380 41800 409386 41812
rect 412358 41800 412364 41812
rect 409380 41772 412364 41800
rect 409380 41760 409386 41772
rect 412358 41760 412364 41772
rect 412416 41800 412422 41812
rect 415210 41800 415216 41812
rect 412416 41772 415216 41800
rect 412416 41760 412422 41772
rect 415210 41760 415216 41772
rect 415268 41760 415274 41812
rect 417050 41760 417056 41812
rect 417108 41800 417114 41812
rect 417108 41772 417280 41800
rect 417108 41760 417114 41772
rect 307404 41704 309180 41732
rect 309152 41664 309180 41704
rect 314562 41664 314568 41676
rect 309152 41636 314568 41664
rect 314562 41624 314568 41636
rect 314620 41624 314626 41676
rect 314654 41624 314660 41676
rect 314712 41664 314718 41676
rect 314712 41636 328408 41664
rect 314712 41624 314718 41636
rect 328380 41596 328408 41636
rect 386322 41624 386328 41676
rect 386380 41664 386386 41676
rect 417252 41664 417280 41772
rect 465350 41760 465356 41812
rect 465408 41800 465414 41812
rect 466362 41800 466368 41812
rect 465408 41772 466368 41800
rect 465408 41760 465414 41772
rect 466362 41760 466368 41772
rect 466420 41800 466426 41812
rect 469674 41800 469680 41812
rect 466420 41772 469680 41800
rect 466420 41760 466426 41772
rect 469674 41760 469680 41772
rect 469732 41800 469738 41812
rect 470152 41800 470180 41840
rect 470962 41828 470968 41840
rect 471020 41868 471026 41880
rect 473078 41868 473084 41880
rect 471020 41840 473084 41868
rect 471020 41828 471026 41840
rect 473078 41828 473084 41840
rect 473136 41828 473142 41880
rect 520090 41828 520096 41880
rect 520148 41868 520154 41880
rect 521194 41868 521200 41880
rect 520148 41840 521200 41868
rect 520148 41828 520154 41840
rect 521194 41828 521200 41840
rect 521252 41868 521258 41880
rect 524230 41868 524236 41880
rect 521252 41840 524236 41868
rect 521252 41828 521258 41840
rect 524230 41828 524236 41840
rect 524288 41868 524294 41880
rect 525518 41868 525524 41880
rect 524288 41840 525524 41868
rect 524288 41828 524294 41840
rect 525518 41828 525524 41840
rect 525576 41868 525582 41880
rect 527910 41868 527916 41880
rect 525576 41840 527916 41868
rect 525576 41828 525582 41840
rect 527910 41828 527916 41840
rect 527968 41828 527974 41880
rect 469732 41772 470180 41800
rect 469732 41760 469738 41772
rect 471882 41760 471888 41812
rect 471940 41800 471946 41812
rect 471940 41772 472112 41800
rect 471940 41760 471946 41772
rect 472084 41664 472112 41772
rect 526714 41760 526720 41812
rect 526772 41760 526778 41812
rect 386380 41636 391888 41664
rect 386380 41624 386386 41636
rect 349614 41596 349620 41608
rect 328380 41568 333928 41596
rect 168340 41500 198780 41528
rect 333900 41528 333928 41568
rect 333992 41568 349620 41596
rect 333992 41528 334020 41568
rect 349614 41556 349620 41568
rect 349672 41556 349678 41608
rect 333900 41500 334020 41528
rect 168340 41488 168346 41500
rect 391860 41460 391888 41636
rect 417252 41636 430528 41664
rect 417252 41460 417280 41636
rect 430500 41528 430528 41636
rect 472084 41636 488488 41664
rect 472084 41528 472112 41636
rect 488460 41596 488488 41636
rect 488460 41568 502380 41596
rect 430500 41500 472112 41528
rect 502352 41528 502380 41568
rect 507854 41556 507860 41608
rect 507912 41596 507918 41608
rect 507912 41568 521608 41596
rect 507912 41556 507918 41568
rect 507762 41528 507768 41540
rect 502352 41500 507768 41528
rect 507762 41488 507768 41500
rect 507820 41488 507826 41540
rect 521580 41528 521608 41568
rect 526732 41528 526760 41760
rect 521580 41500 526760 41528
rect 391860 41432 417280 41460
rect 144638 40740 144644 40792
rect 144696 40780 144702 40792
rect 146294 40780 146300 40792
rect 144696 40752 146300 40780
rect 144696 40740 144702 40752
rect 146294 40740 146300 40752
rect 146352 40740 146358 40792
rect 135162 40196 135168 40248
rect 135220 40236 135226 40248
rect 143534 40236 143540 40248
rect 135220 40208 143540 40236
rect 135220 40196 135226 40208
rect 143534 40196 143540 40208
rect 143592 40196 143598 40248
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143074 40100 143080 40112
rect 141048 40072 143080 40100
rect 141048 40060 141054 40072
rect 142586 39950 142614 40072
rect 143074 40060 143080 40072
rect 143132 40100 143138 40112
rect 144638 40100 144644 40112
rect 143132 40072 144644 40100
rect 143132 40060 143138 40072
rect 144638 40060 144644 40072
rect 144696 40060 144702 40112
rect 145091 39934 145143 40000
<< via1 >>
rect 673460 875168 673512 875220
rect 675392 875168 675444 875220
rect 673552 874488 673604 874540
rect 675392 874488 675444 874540
rect 673736 870136 673788 870188
rect 675392 870136 675444 870188
rect 673644 864424 673696 864476
rect 675392 864424 675444 864476
rect 673736 863200 673788 863252
rect 675392 863200 675444 863252
rect 675300 818320 675352 818372
rect 677508 818320 677560 818372
rect 41788 799552 41840 799604
rect 42340 799552 42392 799604
rect 41788 797716 41840 797768
rect 42708 797716 42760 797768
rect 41788 792548 41840 792600
rect 42340 792548 42392 792600
rect 41788 787244 41840 787296
rect 42616 787244 42668 787296
rect 41788 786632 41840 786684
rect 42524 786632 42576 786684
rect 673460 786564 673512 786616
rect 674012 786564 674064 786616
rect 675392 786564 675444 786616
rect 673552 786360 673604 786412
rect 675392 786360 675444 786412
rect 675300 781600 675352 781652
rect 675300 781396 675352 781448
rect 673460 774868 673512 774920
rect 673644 774868 673696 774920
rect 675392 774868 675444 774920
rect 675208 773984 675260 774036
rect 675392 773984 675444 774036
rect 673736 772760 673788 772812
rect 674012 772760 674064 772812
rect 42432 767320 42484 767372
rect 42708 767320 42760 767372
rect 42524 758956 42576 759008
rect 42800 758956 42852 759008
rect 41788 756372 41840 756424
rect 42340 756372 42392 756424
rect 41788 754468 41840 754520
rect 42432 754468 42484 754520
rect 673736 753516 673788 753568
rect 673920 753516 673972 753568
rect 42524 753448 42576 753500
rect 42800 753448 42852 753500
rect 41788 749368 41840 749420
rect 42340 749368 42392 749420
rect 41788 744132 41840 744184
rect 42340 744132 42392 744184
rect 42616 744132 42668 744184
rect 41788 743996 41840 744048
rect 42524 743996 42576 744048
rect 42984 743996 43036 744048
rect 673644 741956 673696 742008
rect 673920 741956 673972 742008
rect 675392 741888 675444 741940
rect 673552 740664 673604 740716
rect 675392 740664 675444 740716
rect 673644 739780 673696 739832
rect 673644 739644 673696 739696
rect 42340 739576 42392 739628
rect 42616 739576 42668 739628
rect 42524 734136 42576 734188
rect 42984 734136 43036 734188
rect 673460 730124 673512 730176
rect 675392 730124 675444 730176
rect 42524 720332 42576 720384
rect 42892 720332 42944 720384
rect 41788 713124 41840 713176
rect 42340 713124 42392 713176
rect 41788 711288 41840 711340
rect 42432 711288 42484 711340
rect 42708 711288 42760 711340
rect 41788 706188 41840 706240
rect 42340 706188 42392 706240
rect 673644 701020 673696 701072
rect 673828 701020 673880 701072
rect 41788 700952 41840 701004
rect 42616 700952 42668 701004
rect 41788 700816 41840 700868
rect 42892 700816 42944 700868
rect 675392 695920 675444 695972
rect 673644 695852 673696 695904
rect 42432 695512 42484 695564
rect 42892 695512 42944 695564
rect 673552 695308 673604 695360
rect 675392 695308 675444 695360
rect 673460 685176 673512 685228
rect 675392 685176 675444 685228
rect 42432 681640 42484 681692
rect 42800 681572 42852 681624
rect 42616 678512 42668 678564
rect 42984 678512 43036 678564
rect 42432 676132 42484 676184
rect 42984 676132 43036 676184
rect 41788 669944 41840 669996
rect 42340 669944 42392 669996
rect 41788 669060 41840 669112
rect 42524 669060 42576 669112
rect 41788 663008 41840 663060
rect 42340 663008 42392 663060
rect 41788 658656 41840 658708
rect 42432 658656 42484 658708
rect 42708 658656 42760 658708
rect 41788 658044 41840 658096
rect 42800 658044 42852 658096
rect 673644 651720 673696 651772
rect 675392 651720 675444 651772
rect 42432 651380 42484 651432
rect 42800 651380 42852 651432
rect 673552 651108 673604 651160
rect 675392 651108 675444 651160
rect 675208 646008 675260 646060
rect 675300 645736 675352 645788
rect 673460 639684 673512 639736
rect 673920 639684 673972 639736
rect 675392 639684 675444 639736
rect 675208 638800 675260 638852
rect 675392 638800 675444 638852
rect 42524 632000 42576 632052
rect 42708 632000 42760 632052
rect 42984 632000 43036 632052
rect 42800 631864 42852 631916
rect 41788 626764 41840 626816
rect 42340 626764 42392 626816
rect 41788 624928 41840 624980
rect 42800 624928 42852 624980
rect 41788 619760 41840 619812
rect 42340 619760 42392 619812
rect 41788 615476 41840 615528
rect 42984 615476 43036 615528
rect 41788 614796 41840 614848
rect 42524 614796 42576 614848
rect 42800 612824 42852 612876
rect 42616 612756 42668 612808
rect 42616 612620 42668 612672
rect 42800 612620 42852 612672
rect 673644 606704 673696 606756
rect 675392 606704 675444 606756
rect 673552 606160 673604 606212
rect 675024 606160 675076 606212
rect 675392 606160 675444 606212
rect 675208 600788 675260 600840
rect 675392 600788 675444 600840
rect 673644 594872 673696 594924
rect 673920 594872 673972 594924
rect 675392 594872 675444 594924
rect 673736 594736 673788 594788
rect 675024 594736 675076 594788
rect 675300 593376 675352 593428
rect 675300 593172 675352 593224
rect 673552 585148 673604 585200
rect 673828 585148 673880 585200
rect 41788 583516 41840 583568
rect 42340 583516 42392 583568
rect 41788 582632 41840 582684
rect 42800 582632 42852 582684
rect 41788 576580 41840 576632
rect 42340 576580 42392 576632
rect 673736 575424 673788 575476
rect 674380 575424 674432 575476
rect 42340 574064 42392 574116
rect 42800 574064 42852 574116
rect 41788 571208 41840 571260
rect 42800 571208 42852 571260
rect 41788 570664 41840 570716
rect 42524 570664 42576 570716
rect 42708 570664 42760 570716
rect 673552 560532 673604 560584
rect 673828 560532 673880 560584
rect 675392 560532 675444 560584
rect 674012 559920 674064 559972
rect 674380 559920 674432 559972
rect 675392 559920 675444 559972
rect 42616 554752 42668 554804
rect 42800 554752 42852 554804
rect 673644 550468 673696 550520
rect 675392 550468 675444 550520
rect 673552 546388 673604 546440
rect 673828 546320 673880 546372
rect 41788 540336 41840 540388
rect 42340 540336 42392 540388
rect 41788 539452 41840 539504
rect 42524 539452 42576 539504
rect 41788 533400 41840 533452
rect 42340 533400 42392 533452
rect 41788 528028 41840 528080
rect 42616 528028 42668 528080
rect 41788 527484 41840 527536
rect 42432 527484 42484 527536
rect 42708 527484 42760 527536
rect 675300 513748 675352 513800
rect 677692 513748 677744 513800
rect 673736 502324 673788 502376
rect 673920 502324 673972 502376
rect 673552 498176 673604 498228
rect 673828 498176 673880 498228
rect 673828 469276 673880 469328
rect 673736 469140 673788 469192
rect 673736 463632 673788 463684
rect 674012 463632 674064 463684
rect 673552 449556 673604 449608
rect 673828 449556 673880 449608
rect 42616 444320 42668 444372
rect 42800 444320 42852 444372
rect 673736 444320 673788 444372
rect 674012 444320 674064 444372
rect 42708 441532 42760 441584
rect 42800 441532 42852 441584
rect 42616 422288 42668 422340
rect 42708 422288 42760 422340
rect 673644 420724 673696 420776
rect 673828 420724 673880 420776
rect 41788 412768 41840 412820
rect 42340 412768 42392 412820
rect 41788 411204 41840 411256
rect 42524 411204 42576 411256
rect 41788 405764 41840 405816
rect 42340 405764 42392 405816
rect 42616 405696 42668 405748
rect 42892 405696 42944 405748
rect 673828 401548 673880 401600
rect 675300 401548 675352 401600
rect 41788 401344 41840 401396
rect 42892 401344 42944 401396
rect 41788 400800 41840 400852
rect 42432 400800 42484 400852
rect 42616 386316 42668 386368
rect 42892 386316 42944 386368
rect 673736 384276 673788 384328
rect 675392 384276 675444 384328
rect 673644 383188 673696 383240
rect 675300 383188 675352 383240
rect 673552 380876 673604 380928
rect 673736 380876 673788 380928
rect 42800 372580 42852 372632
rect 42984 372580 43036 372632
rect 673736 372308 673788 372360
rect 675392 372308 675444 372360
rect 41788 369520 41840 369572
rect 42340 369520 42392 369572
rect 41788 368636 41840 368688
rect 42892 368636 42944 368688
rect 42524 367820 42576 367872
rect 42800 367820 42852 367872
rect 41788 362584 41840 362636
rect 42340 362584 42392 362636
rect 41788 358232 41840 358284
rect 42524 358232 42576 358284
rect 41788 357620 41840 357672
rect 42432 357620 42484 357672
rect 42616 357620 42668 357672
rect 673552 338104 673604 338156
rect 675392 338104 675444 338156
rect 673644 337492 673696 337544
rect 675392 337492 675444 337544
rect 673736 328040 673788 328092
rect 675392 328040 675444 328092
rect 41788 326340 41840 326392
rect 42340 326340 42392 326392
rect 41788 325456 41840 325508
rect 42432 325456 42484 325508
rect 42708 325456 42760 325508
rect 42432 322872 42484 322924
rect 42616 322804 42668 322856
rect 42708 322804 42760 322856
rect 42892 322736 42944 322788
rect 41788 319404 41840 319456
rect 42340 319404 42392 319456
rect 42340 314168 42392 314220
rect 42708 314168 42760 314220
rect 41788 314032 41840 314084
rect 42524 314032 42576 314084
rect 42708 314032 42760 314084
rect 41788 313488 41840 313540
rect 42800 313420 42852 313472
rect 673552 303560 673604 303612
rect 675300 303560 675352 303612
rect 673644 293564 673696 293616
rect 673920 293564 673972 293616
rect 675392 293564 675444 293616
rect 673644 293428 673696 293480
rect 675300 293428 675352 293480
rect 41788 283160 41840 283212
rect 42340 283160 42392 283212
rect 41788 282276 41840 282328
rect 42524 282276 42576 282328
rect 673736 282072 673788 282124
rect 675392 282072 675444 282124
rect 41788 276156 41840 276208
rect 42340 276156 42392 276208
rect 41788 271872 41840 271924
rect 42708 271872 42760 271924
rect 41788 271192 41840 271244
rect 42524 271192 42576 271244
rect 42800 271192 42852 271244
rect 673460 264936 673512 264988
rect 673644 264936 673696 264988
rect 673460 248684 673512 248736
rect 675300 248684 675352 248736
rect 673644 247460 673696 247512
rect 673920 247460 673972 247512
rect 675392 247460 675444 247512
rect 42340 245556 42392 245608
rect 42892 245556 42944 245608
rect 42524 245488 42576 245540
rect 42800 245488 42852 245540
rect 673828 243788 673880 243840
rect 675300 243788 675352 243840
rect 41788 239912 41840 239964
rect 42340 239912 42392 239964
rect 41788 238076 41840 238128
rect 42616 238076 42668 238128
rect 42892 238076 42944 238128
rect 673920 237668 673972 237720
rect 675392 237668 675444 237720
rect 673920 237328 673972 237380
rect 674104 237328 674156 237380
rect 41788 232976 41840 233028
rect 42340 232976 42392 233028
rect 42340 232840 42392 232892
rect 42616 232840 42668 232892
rect 674104 231752 674156 231804
rect 674288 231752 674340 231804
rect 41788 228624 41840 228676
rect 42708 228624 42760 228676
rect 41788 228012 41840 228064
rect 42616 228012 42668 228064
rect 42800 228012 42852 228064
rect 673828 218084 673880 218136
rect 673828 217948 673880 218000
rect 673736 212508 673788 212560
rect 673828 212508 673880 212560
rect 674012 212508 674064 212560
rect 674288 212508 674340 212560
rect 42340 208360 42392 208412
rect 42892 208360 42944 208412
rect 673736 203872 673788 203924
rect 675392 203872 675444 203924
rect 673644 203328 673696 203380
rect 675392 203328 675444 203380
rect 674012 198704 674064 198756
rect 675208 198704 675260 198756
rect 41788 196732 41840 196784
rect 42340 196732 42392 196784
rect 41788 194896 41840 194948
rect 42432 194896 42484 194948
rect 42892 194896 42944 194948
rect 674748 192108 674800 192160
rect 675208 192108 675260 192160
rect 675392 192108 675444 192160
rect 41788 189796 41840 189848
rect 42340 189796 42392 189848
rect 41788 185444 41840 185496
rect 42340 185444 42392 185496
rect 42708 185444 42760 185496
rect 42432 185308 42484 185360
rect 42708 185308 42760 185360
rect 41788 184832 41840 184884
rect 42432 184832 42484 184884
rect 42616 184832 42668 184884
rect 673828 173884 673880 173936
rect 674748 173884 674800 173936
rect 673552 158312 673604 158364
rect 675392 158312 675444 158364
rect 673460 157292 673512 157344
rect 675392 157292 675444 157344
rect 42524 149064 42576 149116
rect 42708 149064 42760 149116
rect 673644 147092 673696 147144
rect 675024 147092 675076 147144
rect 675392 147092 675444 147144
rect 674012 140632 674064 140684
rect 675024 140632 675076 140684
rect 42248 121456 42300 121508
rect 44732 121456 44784 121508
rect 673828 115948 673880 116000
rect 674012 115948 674064 116000
rect 42984 115880 43036 115932
rect 44732 115880 44784 115932
rect 673828 115812 673880 115864
rect 675024 115812 675076 115864
rect 673552 112752 673604 112804
rect 675392 112752 675444 112804
rect 673460 112072 673512 112124
rect 675392 112072 675444 112124
rect 42524 110440 42576 110492
rect 42708 110440 42760 110492
rect 673644 102280 673696 102332
rect 675024 102280 675076 102332
rect 675392 102280 675444 102332
rect 44640 82832 44692 82884
rect 44824 82764 44876 82816
rect 42340 45704 42392 45756
rect 140964 45704 141016 45756
rect 42432 45636 42484 45688
rect 143632 45636 143684 45688
rect 42708 45568 42760 45620
rect 143540 45568 143592 45620
rect 527456 45568 527508 45620
rect 673552 45568 673604 45620
rect 44916 45500 44968 45552
rect 195980 45500 196032 45552
rect 516324 45500 516376 45552
rect 673644 45500 673696 45552
rect 405648 44752 405700 44804
rect 411260 44752 411312 44804
rect 195980 44412 196032 44464
rect 304540 44412 304592 44464
rect 359372 44684 359424 44736
rect 406752 44684 406804 44736
rect 425060 44684 425112 44736
rect 444196 44684 444248 44736
rect 425060 44548 425112 44600
rect 354404 44480 354456 44532
rect 360568 44480 360620 44532
rect 360660 44480 360712 44532
rect 386420 44480 386472 44532
rect 399668 44480 399720 44532
rect 406752 44480 406804 44532
rect 411260 44480 411312 44532
rect 444288 44480 444340 44532
rect 461492 44548 461544 44600
rect 469128 44548 469180 44600
rect 469220 44548 469272 44600
rect 483020 44616 483072 44668
rect 502248 44480 502300 44532
rect 516324 44480 516376 44532
rect 414204 44412 414256 44464
rect 419816 44412 419868 44464
rect 143632 44344 143684 44396
rect 145104 44344 145156 44396
rect 195336 44344 195388 44396
rect 199660 44344 199712 44396
rect 200856 44344 200908 44396
rect 241336 44344 241388 44396
rect 251088 44344 251140 44396
rect 306380 44344 306432 44396
rect 309416 44344 309468 44396
rect 352564 44344 352616 44396
rect 355416 44344 355468 44396
rect 359372 44344 359424 44396
rect 360660 44344 360712 44396
rect 364248 44344 364300 44396
rect 407396 44344 407448 44396
rect 410432 44344 410484 44396
rect 419080 44344 419132 44396
rect 462136 44344 462188 44396
rect 465172 44344 465224 44396
rect 473820 44344 473872 44396
rect 516968 44344 517020 44396
rect 520004 44344 520056 44396
rect 188528 44276 188580 44328
rect 192852 44276 192904 44328
rect 201500 44276 201552 44328
rect 297088 44276 297140 44328
rect 299572 44276 299624 44328
rect 305736 44276 305788 44328
rect 351920 44276 351972 44328
rect 354404 44276 354456 44328
rect 186688 44208 186740 44260
rect 194692 44208 194744 44260
rect 199660 44208 199712 44260
rect 303896 44208 303948 44260
rect 308220 44208 308272 44260
rect 358728 44276 358780 44328
rect 360568 44276 360620 44328
rect 399668 44276 399720 44328
rect 355600 44208 355652 44260
rect 359924 44208 359976 44260
rect 363052 44208 363104 44260
rect 413560 44276 413612 44328
rect 417884 44276 417936 44328
rect 468300 44276 468352 44328
rect 472624 44276 472676 44328
rect 523132 44276 523184 44328
rect 411076 44208 411128 44260
rect 419724 44208 419776 44260
rect 419816 44208 419868 44260
rect 468944 44208 468996 44260
rect 523776 44208 523828 44260
rect 295248 44140 295300 44192
rect 303252 44140 303304 44192
rect 350080 44140 350132 44192
rect 358084 44140 358136 44192
rect 358728 44140 358780 44192
rect 404912 44140 404964 44192
rect 412916 44140 412968 44192
rect 459652 44140 459704 44192
rect 467656 44140 467708 44192
rect 514484 44140 514536 44192
rect 522488 44140 522540 44192
rect 523132 44140 523184 44192
rect 527456 44140 527508 44192
rect 576768 42712 576820 42764
rect 673460 42712 673512 42764
rect 251088 42032 251140 42084
rect 255228 42032 255280 42084
rect 146300 41964 146352 42016
rect 569132 41964 569184 42016
rect 576768 41964 576820 42016
rect 187700 41896 187752 41948
rect 188436 41896 188488 41948
rect 198924 41896 198976 41948
rect 198464 41828 198516 41880
rect 200120 41828 200172 41880
rect 255228 41828 255280 41880
rect 297640 41828 297692 41880
rect 300676 41828 300728 41880
rect 149612 41760 149664 41812
rect 187700 41760 187752 41812
rect 189264 41760 189316 41812
rect 191104 41760 191156 41812
rect 192300 41760 192352 41812
rect 193588 41760 193640 41812
rect 196440 41760 196492 41812
rect 168288 41692 168340 41744
rect 93768 41556 93820 41608
rect 121552 41556 121604 41608
rect 121276 41488 121328 41540
rect 140872 41556 140924 41608
rect 140688 41488 140740 41540
rect 168288 41488 168340 41540
rect 198832 41760 198884 41812
rect 302240 41760 302292 41812
rect 305000 41760 305052 41812
rect 306288 41760 306340 41812
rect 307484 41896 307536 41948
rect 362500 41896 362552 41948
rect 367100 41896 367152 41948
rect 360016 41828 360068 41880
rect 361120 41828 361172 41880
rect 363512 41828 363564 41880
rect 410524 41828 410576 41880
rect 411812 41828 411864 41880
rect 414848 41828 414900 41880
rect 416136 41828 416188 41880
rect 418528 41828 418580 41880
rect 464160 41828 464212 41880
rect 467196 41828 467248 41880
rect 470048 41828 470100 41880
rect 409328 41760 409380 41812
rect 412364 41760 412416 41812
rect 415216 41760 415268 41812
rect 417056 41760 417108 41812
rect 314568 41624 314620 41676
rect 314660 41624 314712 41676
rect 386328 41624 386380 41676
rect 465356 41760 465408 41812
rect 466368 41760 466420 41812
rect 469680 41760 469732 41812
rect 470968 41828 471020 41880
rect 473084 41828 473136 41880
rect 520096 41828 520148 41880
rect 521200 41828 521252 41880
rect 524236 41828 524288 41880
rect 525524 41828 525576 41880
rect 527916 41828 527968 41880
rect 471888 41760 471940 41812
rect 526720 41760 526772 41812
rect 349620 41556 349672 41608
rect 507860 41556 507912 41608
rect 507768 41488 507820 41540
rect 144644 40740 144696 40792
rect 146300 40740 146352 40792
rect 135168 40196 135220 40248
rect 143540 40196 143592 40248
rect 140996 40060 141048 40112
rect 143080 40060 143132 40112
rect 144644 40060 144696 40112
<< metal2 >>
rect 342164 997474 342224 997483
rect 342164 997405 342224 997414
rect 342180 997192 342208 997405
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 673472 875226 673500 875276
rect 675404 875226 675432 875683
rect 673460 875220 673512 875226
rect 673460 875162 673512 875168
rect 675392 875220 675444 875226
rect 675392 875162 675444 875168
rect 42246 870088 42302 870097
rect 42246 870023 42302 870032
rect 41722 800075 41828 800103
rect 41800 799610 41828 800075
rect 41788 799604 41840 799610
rect 41788 799546 41840 799552
rect 41713 799417 42193 799473
rect 41722 798238 41828 798266
rect 41800 797774 41828 798238
rect 41788 797768 41840 797774
rect 41788 797710 41840 797716
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41788 792600 41840 792606
rect 41788 792542 41840 792548
rect 41800 792099 41828 792542
rect 41722 792071 41828 792099
rect 41713 791413 42193 791469
rect 41713 790769 42193 790825
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 41800 787302 41828 787752
rect 41788 787296 41840 787302
rect 41788 787238 41840 787244
rect 41800 786690 41828 787122
rect 41788 786684 41840 786690
rect 41788 786626 41840 786632
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 41722 756894 41828 756922
rect 41800 756430 41828 756894
rect 41788 756424 41840 756430
rect 41788 756366 41840 756372
rect 41713 756217 42193 756273
rect 41722 755035 41828 755063
rect 41800 754526 41828 755035
rect 41788 754520 41840 754526
rect 41788 754462 41840 754468
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41788 749420 41840 749426
rect 41788 749362 41840 749368
rect 41800 748898 41828 749362
rect 41722 748870 41828 748898
rect 41713 748213 42193 748269
rect 41713 747569 42193 747625
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41722 744547 41828 744575
rect 41800 744190 41828 744547
rect 41788 744184 41840 744190
rect 41788 744126 41840 744132
rect 41788 744048 41840 744054
rect 41788 743990 41840 743996
rect 41800 743931 41828 743990
rect 41722 743903 41828 743931
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 41722 713675 41828 713703
rect 41800 713182 41828 713675
rect 41788 713176 41840 713182
rect 41788 713118 41840 713124
rect 41713 713017 42193 713073
rect 41722 711835 41828 711863
rect 41800 711346 41828 711835
rect 41788 711340 41840 711346
rect 41788 711282 41840 711288
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41788 706240 41840 706246
rect 41788 706182 41840 706188
rect 41800 705699 41828 706182
rect 41722 705671 41828 705699
rect 41713 705013 42193 705069
rect 41713 704369 42193 704425
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41722 701347 41828 701375
rect 41800 701010 41828 701347
rect 41788 701004 41840 701010
rect 41788 700946 41840 700952
rect 41788 700868 41840 700874
rect 41788 700810 41840 700816
rect 41800 700712 41828 700810
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41722 670475 41828 670503
rect 41800 670002 41828 670475
rect 41788 669996 41840 670002
rect 41788 669938 41840 669944
rect 41713 669817 42193 669873
rect 41788 669112 41840 669118
rect 41788 669054 41840 669060
rect 41800 668658 41828 669054
rect 41722 668630 41828 668658
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 41788 663060 41840 663066
rect 41788 663002 41840 663008
rect 41800 662499 41828 663002
rect 41722 662471 41828 662499
rect 41713 661813 42193 661869
rect 41713 661169 42193 661225
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41788 658708 41840 658714
rect 41788 658650 41840 658656
rect 41800 658186 41828 658650
rect 41722 658158 41828 658186
rect 41788 658096 41840 658102
rect 41788 658038 41840 658044
rect 41800 657522 41828 658038
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 41722 627286 41828 627314
rect 41800 626822 41828 627286
rect 41788 626816 41840 626822
rect 41788 626758 41840 626764
rect 41713 626617 42193 626673
rect 41722 625435 41828 625463
rect 41800 624986 41828 625435
rect 41788 624980 41840 624986
rect 41788 624922 41840 624928
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 41788 619812 41840 619818
rect 41788 619754 41840 619760
rect 41800 619290 41828 619754
rect 41722 619262 41828 619290
rect 41713 618613 42193 618669
rect 41713 617969 42193 618025
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41788 615528 41840 615534
rect 41788 615470 41840 615476
rect 41800 614975 41828 615470
rect 41722 614947 41828 614975
rect 41788 614848 41840 614854
rect 41788 614790 41840 614796
rect 41800 614331 41828 614790
rect 41722 614303 41828 614331
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 41722 584075 41828 584103
rect 41800 583574 41828 584075
rect 41788 583568 41840 583574
rect 41788 583510 41840 583516
rect 41713 583417 42193 583473
rect 41788 582684 41840 582690
rect 41788 582626 41840 582632
rect 41800 582263 41828 582626
rect 41722 582235 41828 582263
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41788 576632 41840 576638
rect 41788 576574 41840 576580
rect 41800 576099 41828 576574
rect 41722 576071 41828 576099
rect 41713 575413 42193 575469
rect 41713 574769 42193 574825
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41722 571747 41828 571775
rect 41800 571266 41828 571747
rect 41788 571260 41840 571266
rect 41788 571202 41840 571208
rect 41800 570722 41828 571108
rect 41788 570716 41840 570722
rect 41788 570658 41840 570664
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41722 540875 41828 540903
rect 41800 540394 41828 540875
rect 41788 540388 41840 540394
rect 41788 540330 41840 540336
rect 41713 540217 42193 540273
rect 41788 539504 41840 539510
rect 41788 539446 41840 539452
rect 41800 539050 41828 539446
rect 41722 539022 41828 539050
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41788 533452 41840 533458
rect 41788 533394 41840 533400
rect 41800 532899 41828 533394
rect 41722 532871 41828 532899
rect 41713 532213 42193 532269
rect 41713 531569 42193 531625
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41722 528550 41828 528578
rect 41800 528086 41828 528550
rect 41788 528080 41840 528086
rect 41788 528022 41840 528028
rect 41722 527903 41828 527931
rect 41800 527542 41828 527903
rect 41788 527536 41840 527542
rect 41788 527478 41840 527484
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41722 413275 41828 413303
rect 41800 412826 41828 413275
rect 41788 412820 41840 412826
rect 41788 412762 41840 412768
rect 41713 412617 42193 412673
rect 41800 411262 41828 411432
rect 41788 411256 41840 411262
rect 41788 411198 41840 411204
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 41788 405816 41840 405822
rect 41788 405758 41840 405764
rect 41800 405299 41828 405758
rect 41722 405271 41828 405299
rect 41713 404613 42193 404669
rect 41713 403969 42193 404025
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41788 401396 41840 401402
rect 41788 401338 41840 401344
rect 41800 400975 41828 401338
rect 41722 400947 41828 400975
rect 41788 400852 41840 400858
rect 41788 400794 41840 400800
rect 41800 400330 41828 400794
rect 41722 400302 41828 400330
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41722 370075 41828 370103
rect 41800 369578 41828 370075
rect 41788 369572 41840 369578
rect 41788 369514 41840 369520
rect 41713 369417 42193 369473
rect 41788 368688 41840 368694
rect 41788 368630 41840 368636
rect 41800 368263 41828 368630
rect 41722 368235 41828 368263
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41788 362636 41840 362642
rect 41788 362578 41840 362584
rect 41800 362076 41828 362578
rect 41713 361413 42193 361469
rect 41713 360769 42193 360825
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41788 358284 41840 358290
rect 41788 358226 41840 358232
rect 41800 357762 41828 358226
rect 41722 357734 41828 357762
rect 41788 357672 41840 357678
rect 41788 357614 41840 357620
rect 41800 357131 41828 357614
rect 41722 357103 41828 357131
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 41722 326862 41828 326890
rect 41800 326398 41828 326862
rect 41788 326392 41840 326398
rect 41788 326334 41840 326340
rect 41713 326217 42193 326273
rect 41788 325508 41840 325514
rect 41788 325450 41840 325456
rect 41800 325063 41828 325450
rect 41722 325035 41828 325063
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41788 319456 41840 319462
rect 41788 319398 41840 319404
rect 41800 318899 41828 319398
rect 41722 318871 41828 318899
rect 41713 318213 42193 318269
rect 41713 317569 42193 317625
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41722 314547 41828 314575
rect 41800 314090 41828 314547
rect 41788 314084 41840 314090
rect 41788 314026 41840 314032
rect 41722 313903 41828 313931
rect 41800 313546 41828 313903
rect 41788 313540 41840 313546
rect 41788 313482 41840 313488
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 41722 283675 41828 283703
rect 41800 283218 41828 283675
rect 41788 283212 41840 283218
rect 41788 283154 41840 283160
rect 41713 283017 42193 283073
rect 41788 282328 41840 282334
rect 41788 282270 41840 282276
rect 41800 281874 41828 282270
rect 41722 281846 41828 281874
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41788 276208 41840 276214
rect 41788 276150 41840 276156
rect 41800 275699 41828 276150
rect 41722 275671 41828 275699
rect 41713 275013 42193 275069
rect 41713 274369 42193 274425
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41788 271924 41840 271930
rect 41788 271866 41840 271872
rect 41800 271356 41828 271866
rect 41788 271244 41840 271250
rect 41788 271186 41840 271192
rect 41800 270722 41828 271186
rect 41722 270694 41828 270722
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 41722 240502 41828 240530
rect 41800 239970 41828 240502
rect 41788 239964 41840 239970
rect 41788 239906 41840 239912
rect 41713 239817 42193 239873
rect 41722 238635 41828 238663
rect 41800 238134 41828 238635
rect 41788 238128 41840 238134
rect 41788 238070 41840 238076
rect 41713 237977 42193 238033
rect 41713 237333 42193 237389
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 41788 233028 41840 233034
rect 41788 232970 41840 232976
rect 41800 232506 41828 232970
rect 41722 232478 41828 232506
rect 41713 231813 42193 231869
rect 41713 231169 42193 231225
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41788 228676 41840 228682
rect 41788 228618 41840 228624
rect 41800 228166 41828 228618
rect 41788 228064 41840 228070
rect 41788 228006 41840 228012
rect 41800 227531 41828 228006
rect 41722 227503 41828 227531
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41800 196790 41828 197300
rect 41788 196784 41840 196790
rect 41788 196726 41840 196732
rect 41713 196617 42193 196673
rect 41722 195435 41828 195463
rect 41800 194954 41828 195435
rect 41788 194948 41840 194954
rect 41788 194890 41840 194896
rect 41713 194777 42193 194833
rect 41713 194133 42193 194189
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41788 189848 41840 189854
rect 41788 189790 41840 189796
rect 41800 189299 41828 189790
rect 41722 189271 41828 189299
rect 41713 188613 42193 188669
rect 41713 187969 42193 188025
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41788 185496 41840 185502
rect 41788 185438 41840 185444
rect 41800 184975 41828 185438
rect 41722 184947 41828 184975
rect 41788 184884 41840 184890
rect 41788 184826 41840 184832
rect 41800 184331 41828 184826
rect 41722 184303 41828 184331
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 42260 121514 42288 870023
rect 42340 799604 42392 799610
rect 42340 799546 42392 799552
rect 42352 792606 42380 799546
rect 42708 797768 42760 797774
rect 42708 797710 42760 797716
rect 42340 792600 42392 792606
rect 42340 792542 42392 792548
rect 42616 787296 42668 787302
rect 42616 787238 42668 787244
rect 42524 786684 42576 786690
rect 42524 786626 42576 786632
rect 42432 767372 42484 767378
rect 42432 767314 42484 767320
rect 42340 756424 42392 756430
rect 42340 756366 42392 756372
rect 42352 749426 42380 756366
rect 42444 754526 42472 767314
rect 42536 759014 42564 786626
rect 42524 759008 42576 759014
rect 42524 758950 42576 758956
rect 42432 754520 42484 754526
rect 42432 754462 42484 754468
rect 42340 749420 42392 749426
rect 42340 749362 42392 749368
rect 42340 744184 42392 744190
rect 42340 744126 42392 744132
rect 42352 739634 42380 744126
rect 42340 739628 42392 739634
rect 42340 739570 42392 739576
rect 42340 713176 42392 713182
rect 42340 713118 42392 713124
rect 42352 706246 42380 713118
rect 42444 711346 42472 754462
rect 42524 753500 42576 753506
rect 42524 753442 42576 753448
rect 42536 744054 42564 753442
rect 42628 744190 42656 787238
rect 42720 767378 42748 797710
rect 673472 786622 673500 875162
rect 673564 874546 673592 874568
rect 675404 874546 675432 875039
rect 673552 874540 673604 874546
rect 673552 874482 673604 874488
rect 675392 874540 675444 874546
rect 675392 874482 675444 874488
rect 673460 786616 673512 786622
rect 673460 786558 673512 786564
rect 673564 786418 673592 874482
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871975 675887 872031
rect 675407 871331 675887 871387
rect 675404 870194 675432 870740
rect 673736 870188 673788 870194
rect 673736 870130 673788 870136
rect 675392 870188 675444 870194
rect 675392 870130 675444 870136
rect 673656 864482 673684 864518
rect 673644 864476 673696 864482
rect 673644 864418 673696 864424
rect 673552 786412 673604 786418
rect 673552 786354 673604 786360
rect 673460 774920 673512 774926
rect 673460 774862 673512 774868
rect 42708 767372 42760 767378
rect 42708 767314 42760 767320
rect 42800 759008 42852 759014
rect 42800 758950 42852 758956
rect 42812 753506 42840 758950
rect 42800 753500 42852 753506
rect 42800 753442 42852 753448
rect 42616 744184 42668 744190
rect 42616 744126 42668 744132
rect 42524 744048 42576 744054
rect 42524 743990 42576 743996
rect 42984 744048 43036 744054
rect 42984 743990 43036 743996
rect 42616 739628 42668 739634
rect 42616 739570 42668 739576
rect 42524 734188 42576 734194
rect 42524 734130 42576 734136
rect 42536 720390 42564 734130
rect 42524 720384 42576 720390
rect 42524 720326 42576 720332
rect 42432 711340 42484 711346
rect 42432 711282 42484 711288
rect 42340 706240 42392 706246
rect 42340 706182 42392 706188
rect 42628 701010 42656 739570
rect 42996 734194 43024 743990
rect 42984 734188 43036 734194
rect 42984 734130 43036 734136
rect 673472 730182 673500 774862
rect 673564 740722 673592 786354
rect 673656 774926 673684 864418
rect 673748 863258 673776 870130
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675404 864482 675432 864551
rect 675392 864476 675444 864482
rect 675392 864418 675444 864424
rect 675407 863327 675887 863383
rect 673736 863252 673788 863258
rect 673736 863194 673788 863200
rect 675392 863252 675444 863258
rect 675392 863194 675444 863200
rect 675404 862716 675432 863194
rect 677506 818408 677562 818417
rect 675300 818372 675352 818378
rect 677506 818343 677508 818352
rect 675300 818314 675352 818320
rect 677560 818343 677562 818352
rect 677508 818314 677560 818320
rect 674012 786616 674064 786622
rect 674012 786558 674064 786564
rect 673644 774920 673696 774926
rect 673644 774862 673696 774868
rect 674024 772818 674052 786558
rect 675312 781658 675340 818314
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675392 786616 675444 786622
rect 675392 786558 675444 786564
rect 675404 786483 675432 786558
rect 675392 786412 675444 786418
rect 675392 786354 675444 786360
rect 675404 785839 675432 786354
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782775 675887 782831
rect 675407 782131 675887 782187
rect 675300 781652 675352 781658
rect 675300 781594 675352 781600
rect 675220 781510 675418 781538
rect 675220 774042 675248 781510
rect 675300 781448 675352 781454
rect 675300 781390 675352 781396
rect 675208 774036 675260 774042
rect 675208 773978 675260 773984
rect 673736 772812 673788 772818
rect 673736 772754 673788 772760
rect 674012 772812 674064 772818
rect 674012 772754 674064 772760
rect 673748 753574 673776 772754
rect 673736 753568 673788 753574
rect 673736 753510 673788 753516
rect 673920 753568 673972 753574
rect 673920 753510 673972 753516
rect 673932 742014 673960 753510
rect 673644 742008 673696 742014
rect 673644 741950 673696 741956
rect 673920 742008 673972 742014
rect 673920 741950 673972 741956
rect 673552 740716 673604 740722
rect 673552 740658 673604 740664
rect 673460 730176 673512 730182
rect 673460 730118 673512 730124
rect 42892 720384 42944 720390
rect 42892 720326 42944 720332
rect 42708 711340 42760 711346
rect 42708 711282 42760 711288
rect 42616 701004 42668 701010
rect 42616 700946 42668 700952
rect 42432 695564 42484 695570
rect 42432 695506 42484 695512
rect 42444 681698 42472 695506
rect 42432 681692 42484 681698
rect 42432 681634 42484 681640
rect 42628 678570 42656 700946
rect 42616 678564 42668 678570
rect 42616 678506 42668 678512
rect 42720 678450 42748 711282
rect 42904 700874 42932 720326
rect 42892 700868 42944 700874
rect 42892 700810 42944 700816
rect 42904 695570 42932 700810
rect 42892 695564 42944 695570
rect 42892 695506 42944 695512
rect 673472 685234 673500 730118
rect 673564 695366 673592 740658
rect 673656 739838 673684 741950
rect 673644 739832 673696 739838
rect 673644 739774 673696 739780
rect 673644 739696 673696 739702
rect 673644 739638 673696 739644
rect 673656 720338 673684 739638
rect 675312 736658 675340 781390
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675404 774926 675432 775351
rect 675392 774920 675444 774926
rect 675392 774862 675444 774868
rect 675407 774127 675887 774183
rect 675392 774036 675444 774042
rect 675392 773978 675444 773984
rect 675404 773500 675432 773978
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 675392 741940 675444 741946
rect 675392 741882 675444 741888
rect 675404 741483 675432 741882
rect 675404 740722 675432 740860
rect 675392 740716 675444 740722
rect 675392 740658 675444 740664
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737775 675887 737831
rect 675407 737131 675887 737187
rect 675220 736630 675340 736658
rect 675220 728362 675248 736630
rect 675312 736494 675418 736522
rect 675312 729042 675340 736494
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675404 730182 675432 730351
rect 675392 730176 675444 730182
rect 675392 730118 675444 730124
rect 675407 729127 675887 729183
rect 675312 729014 675432 729042
rect 675404 728484 675432 729014
rect 675220 728334 675340 728362
rect 673656 720310 673868 720338
rect 673840 701078 673868 720310
rect 673644 701072 673696 701078
rect 673644 701014 673696 701020
rect 673828 701072 673880 701078
rect 673828 701014 673880 701020
rect 673656 695910 673684 701014
rect 673644 695904 673696 695910
rect 673644 695846 673696 695852
rect 673552 695360 673604 695366
rect 673552 695302 673604 695308
rect 673460 685228 673512 685234
rect 673460 685170 673512 685176
rect 42800 681624 42852 681630
rect 42800 681566 42852 681572
rect 42628 678422 42748 678450
rect 42432 676184 42484 676190
rect 42432 676126 42484 676132
rect 42340 669996 42392 670002
rect 42340 669938 42392 669944
rect 42352 663066 42380 669938
rect 42340 663060 42392 663066
rect 42340 663002 42392 663008
rect 42444 658714 42472 676126
rect 42628 672194 42656 678422
rect 42536 672166 42656 672194
rect 42536 669118 42564 672166
rect 42524 669112 42576 669118
rect 42524 669054 42576 669060
rect 42432 658708 42484 658714
rect 42432 658650 42484 658656
rect 42432 651432 42484 651438
rect 42432 651374 42484 651380
rect 42444 631938 42472 651374
rect 42536 632058 42564 669054
rect 42708 658708 42760 658714
rect 42708 658650 42760 658656
rect 42720 632058 42748 658650
rect 42812 658102 42840 681566
rect 42984 678564 43036 678570
rect 42984 678506 43036 678512
rect 42996 676190 43024 678506
rect 42984 676184 43036 676190
rect 42984 676126 43036 676132
rect 42800 658096 42852 658102
rect 42800 658038 42852 658044
rect 42812 651438 42840 658038
rect 42800 651432 42852 651438
rect 42800 651374 42852 651380
rect 673472 639742 673500 685170
rect 673564 651166 673592 695302
rect 673656 651778 673684 695846
rect 675312 691642 675340 728334
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675404 695978 675432 696483
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675404 695366 675432 695844
rect 675392 695360 675444 695366
rect 675392 695302 675444 695308
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692775 675887 692831
rect 675407 692131 675887 692187
rect 675220 691614 675340 691642
rect 675220 683346 675248 691614
rect 675418 691478 675524 691506
rect 675496 690962 675524 691478
rect 675312 690934 675524 690962
rect 675312 683525 675340 690934
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675404 685234 675432 685372
rect 675392 685228 675444 685234
rect 675392 685170 675444 685176
rect 675407 684127 675887 684183
rect 675312 683497 675418 683525
rect 675220 683318 675340 683346
rect 673644 651772 673696 651778
rect 673644 651714 673696 651720
rect 673552 651160 673604 651166
rect 673552 651102 673604 651108
rect 673460 639736 673512 639742
rect 673460 639678 673512 639684
rect 42524 632052 42576 632058
rect 42524 631994 42576 632000
rect 42708 632052 42760 632058
rect 42708 631994 42760 632000
rect 42984 632052 43036 632058
rect 42984 631994 43036 632000
rect 42444 631910 42564 631938
rect 42340 626816 42392 626822
rect 42340 626758 42392 626764
rect 42352 619818 42380 626758
rect 42340 619812 42392 619818
rect 42340 619754 42392 619760
rect 42536 614854 42564 631910
rect 42800 631916 42852 631922
rect 42800 631858 42852 631864
rect 42812 624986 42840 631858
rect 42800 624980 42852 624986
rect 42800 624922 42852 624928
rect 42524 614848 42576 614854
rect 42524 614790 42576 614796
rect 42340 583568 42392 583574
rect 42340 583510 42392 583516
rect 42352 576638 42380 583510
rect 42340 576632 42392 576638
rect 42340 576574 42392 576580
rect 42340 574116 42392 574122
rect 42340 574058 42392 574064
rect 42352 540546 42380 574058
rect 42536 570722 42564 614790
rect 42812 612882 42840 624922
rect 42996 615534 43024 631994
rect 42984 615528 43036 615534
rect 42984 615470 43036 615476
rect 42800 612876 42852 612882
rect 42800 612818 42852 612824
rect 42616 612808 42668 612814
rect 42996 612762 43024 615470
rect 42616 612750 42668 612756
rect 42628 612678 42656 612750
rect 42720 612734 43024 612762
rect 42616 612672 42668 612678
rect 42616 612614 42668 612620
rect 42720 571282 42748 612734
rect 42800 612672 42852 612678
rect 42800 612614 42852 612620
rect 42812 582690 42840 612614
rect 673564 606218 673592 651102
rect 673656 606762 673684 651714
rect 675312 646898 675340 683318
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675392 651772 675444 651778
rect 675392 651714 675444 651720
rect 675404 651283 675432 651714
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 675404 650639 675432 651102
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 647575 675887 647631
rect 675407 646931 675887 646987
rect 675220 646870 675340 646898
rect 675220 646066 675248 646870
rect 675208 646060 675260 646066
rect 675208 646002 675260 646008
rect 675404 645946 675432 646340
rect 675220 645918 675432 645946
rect 673920 639736 673972 639742
rect 673920 639678 673972 639684
rect 673644 606756 673696 606762
rect 673644 606698 673696 606704
rect 673552 606212 673604 606218
rect 673552 606154 673604 606160
rect 673656 595082 673684 606698
rect 673564 595054 673684 595082
rect 673564 585206 673592 595054
rect 673932 594930 673960 639678
rect 675220 638858 675248 645918
rect 675300 645788 675352 645794
rect 675300 645730 675352 645736
rect 675208 638852 675260 638858
rect 675208 638794 675260 638800
rect 675024 606212 675076 606218
rect 675024 606154 675076 606160
rect 673644 594924 673696 594930
rect 673644 594866 673696 594872
rect 673920 594924 673972 594930
rect 673920 594866 673972 594872
rect 673552 585200 673604 585206
rect 673552 585142 673604 585148
rect 42800 582684 42852 582690
rect 42800 582626 42852 582632
rect 42812 574122 42840 582626
rect 42800 574116 42852 574122
rect 42800 574058 42852 574064
rect 42720 571266 42840 571282
rect 42720 571260 42852 571266
rect 42720 571254 42800 571260
rect 42800 571202 42852 571208
rect 42524 570716 42576 570722
rect 42524 570658 42576 570664
rect 42708 570716 42760 570722
rect 42708 570658 42760 570664
rect 42616 554804 42668 554810
rect 42616 554746 42668 554752
rect 42352 540518 42564 540546
rect 42340 540388 42392 540394
rect 42340 540330 42392 540336
rect 42352 533458 42380 540330
rect 42536 539510 42564 540518
rect 42524 539504 42576 539510
rect 42524 539446 42576 539452
rect 42340 533452 42392 533458
rect 42340 533394 42392 533400
rect 42432 527536 42484 527542
rect 42432 527478 42484 527484
rect 42340 412820 42392 412826
rect 42340 412762 42392 412768
rect 42352 405822 42380 412762
rect 42340 405816 42392 405822
rect 42340 405758 42392 405764
rect 42444 400858 42472 527478
rect 42536 411262 42564 539446
rect 42628 528086 42656 554746
rect 42616 528080 42668 528086
rect 42616 528022 42668 528028
rect 42628 444378 42656 528022
rect 42720 527542 42748 570658
rect 42812 554810 42840 571202
rect 673552 560584 673604 560590
rect 673552 560526 673604 560532
rect 42800 554804 42852 554810
rect 42800 554746 42852 554752
rect 673564 546446 673592 560526
rect 673656 550526 673684 594866
rect 675036 594794 675064 606154
rect 675208 600840 675260 600846
rect 675208 600782 675260 600788
rect 673736 594788 673788 594794
rect 673736 594730 673788 594736
rect 675024 594788 675076 594794
rect 675024 594730 675076 594736
rect 673748 575482 673776 594730
rect 675220 593314 675248 600782
rect 675312 593434 675340 645730
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675404 639742 675432 640151
rect 675392 639736 675444 639742
rect 675392 639678 675444 639684
rect 675407 638927 675887 638983
rect 675392 638852 675444 638858
rect 675392 638794 675444 638800
rect 675404 638316 675432 638794
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675392 606756 675444 606762
rect 675392 606698 675444 606704
rect 675404 606283 675432 606698
rect 675392 606212 675444 606218
rect 675392 606154 675444 606160
rect 675404 605639 675432 606154
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 602575 675887 602631
rect 675407 601931 675887 601987
rect 675404 600846 675432 601324
rect 675392 600840 675444 600846
rect 675392 600782 675444 600788
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675404 594930 675432 595151
rect 675392 594924 675444 594930
rect 675392 594866 675444 594872
rect 675407 593927 675887 593983
rect 675300 593428 675352 593434
rect 675300 593370 675352 593376
rect 675220 593286 675418 593314
rect 675300 593224 675352 593230
rect 675300 593166 675352 593172
rect 673828 585200 673880 585206
rect 673828 585142 673880 585148
rect 673736 575476 673788 575482
rect 673736 575418 673788 575424
rect 673840 560590 673868 585142
rect 674380 575476 674432 575482
rect 674380 575418 674432 575424
rect 673828 560584 673880 560590
rect 673828 560526 673880 560532
rect 674392 559978 674420 575418
rect 674012 559972 674064 559978
rect 674012 559914 674064 559920
rect 674380 559972 674432 559978
rect 674380 559914 674432 559920
rect 673644 550520 673696 550526
rect 673644 550462 673696 550468
rect 673552 546440 673604 546446
rect 673552 546382 673604 546388
rect 673828 546372 673880 546378
rect 673828 546314 673880 546320
rect 42708 527536 42760 527542
rect 42708 527478 42760 527484
rect 673734 521656 673790 521665
rect 673734 521591 673790 521600
rect 673748 502382 673776 521591
rect 673736 502376 673788 502382
rect 673736 502318 673788 502324
rect 673840 498234 673868 546314
rect 674024 521665 674052 559914
rect 675312 556186 675340 593166
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675404 560590 675432 561068
rect 675392 560584 675444 560590
rect 675392 560526 675444 560532
rect 675404 559978 675432 560439
rect 675392 559972 675444 559978
rect 675392 559914 675444 559920
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 557375 675887 557431
rect 675407 556731 675887 556787
rect 675220 556158 675340 556186
rect 675220 548298 675248 556158
rect 675312 556101 675418 556129
rect 675312 548570 675340 556101
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675392 550520 675444 550526
rect 675392 550462 675444 550468
rect 675404 549951 675432 550462
rect 675407 548727 675887 548783
rect 675312 548542 675432 548570
rect 675220 548270 675340 548298
rect 674010 521656 674066 521665
rect 674010 521591 674066 521600
rect 675312 513806 675340 548270
rect 675404 548111 675432 548542
rect 675300 513800 675352 513806
rect 677692 513800 677744 513806
rect 675300 513742 675352 513748
rect 677690 513768 677692 513777
rect 677744 513768 677746 513777
rect 677690 513703 677746 513712
rect 673920 502376 673972 502382
rect 673920 502318 673972 502324
rect 673552 498228 673604 498234
rect 673552 498170 673604 498176
rect 673828 498228 673880 498234
rect 673828 498170 673880 498176
rect 673564 449614 673592 498170
rect 673932 488458 673960 502318
rect 673840 488430 673960 488458
rect 673840 469334 673868 488430
rect 673828 469328 673880 469334
rect 673828 469270 673880 469276
rect 673736 469192 673788 469198
rect 673736 469134 673788 469140
rect 673748 463690 673776 469134
rect 673736 463684 673788 463690
rect 673736 463626 673788 463632
rect 674012 463684 674064 463690
rect 674012 463626 674064 463632
rect 673552 449608 673604 449614
rect 673552 449550 673604 449556
rect 673828 449608 673880 449614
rect 673828 449550 673880 449556
rect 42616 444372 42668 444378
rect 42616 444314 42668 444320
rect 42800 444372 42852 444378
rect 42800 444314 42852 444320
rect 673736 444372 673788 444378
rect 673736 444314 673788 444320
rect 42812 441590 42840 444314
rect 42708 441584 42760 441590
rect 42708 441526 42760 441532
rect 42800 441584 42852 441590
rect 42800 441526 42852 441532
rect 42720 422346 42748 441526
rect 42616 422340 42668 422346
rect 42616 422282 42668 422288
rect 42708 422340 42760 422346
rect 42708 422282 42760 422288
rect 42524 411256 42576 411262
rect 42524 411198 42576 411204
rect 42432 400852 42484 400858
rect 42432 400794 42484 400800
rect 42340 369572 42392 369578
rect 42340 369514 42392 369520
rect 42352 362642 42380 369514
rect 42340 362636 42392 362642
rect 42340 362578 42392 362584
rect 42444 357678 42472 400794
rect 42536 391898 42564 411198
rect 42628 405754 42656 422282
rect 673748 421002 673776 444314
rect 673656 420974 673776 421002
rect 673656 420782 673684 420974
rect 673840 420866 673868 449550
rect 674024 444378 674052 463626
rect 674012 444372 674064 444378
rect 674012 444314 674064 444320
rect 673748 420838 673868 420866
rect 673644 420776 673696 420782
rect 673644 420718 673696 420724
rect 42616 405748 42668 405754
rect 42616 405690 42668 405696
rect 42892 405748 42944 405754
rect 42892 405690 42944 405696
rect 42904 401402 42932 405690
rect 42892 401396 42944 401402
rect 42892 401338 42944 401344
rect 42904 401282 42932 401338
rect 42904 401254 43024 401282
rect 42536 391870 42656 391898
rect 42628 386374 42656 391870
rect 42616 386368 42668 386374
rect 42616 386310 42668 386316
rect 42892 386368 42944 386374
rect 42892 386310 42944 386316
rect 42800 372632 42852 372638
rect 42800 372574 42852 372580
rect 42812 367878 42840 372574
rect 42904 368694 42932 386310
rect 42996 372638 43024 401254
rect 673748 384334 673776 420838
rect 673828 420776 673880 420782
rect 673828 420718 673880 420724
rect 673840 401606 673868 420718
rect 673828 401600 673880 401606
rect 673828 401542 673880 401548
rect 675300 401600 675352 401606
rect 675300 401542 675352 401548
rect 673736 384328 673788 384334
rect 673736 384270 673788 384276
rect 673644 383240 673696 383246
rect 673644 383182 673696 383188
rect 673552 380928 673604 380934
rect 673552 380870 673604 380876
rect 42984 372632 43036 372638
rect 42984 372574 43036 372580
rect 42892 368688 42944 368694
rect 42892 368630 42944 368636
rect 42524 367872 42576 367878
rect 42524 367814 42576 367820
rect 42800 367872 42852 367878
rect 42800 367814 42852 367820
rect 42536 358290 42564 367814
rect 42904 367724 42932 368630
rect 42812 367696 42932 367724
rect 42524 358284 42576 358290
rect 42524 358226 42576 358232
rect 42432 357672 42484 357678
rect 42432 357614 42484 357620
rect 42340 326392 42392 326398
rect 42340 326334 42392 326340
rect 42352 319462 42380 326334
rect 42432 325508 42484 325514
rect 42432 325450 42484 325456
rect 42444 322930 42472 325450
rect 42432 322924 42484 322930
rect 42432 322866 42484 322872
rect 42340 319456 42392 319462
rect 42340 319398 42392 319404
rect 42340 314220 42392 314226
rect 42340 314162 42392 314168
rect 42352 283703 42380 314162
rect 42536 314090 42564 358226
rect 42616 357672 42668 357678
rect 42616 357614 42668 357620
rect 42628 322862 42656 357614
rect 42812 342258 42840 367696
rect 42720 342230 42840 342258
rect 42720 325514 42748 342230
rect 673564 338162 673592 380870
rect 673552 338156 673604 338162
rect 673552 338098 673604 338104
rect 42708 325508 42760 325514
rect 42708 325450 42760 325456
rect 42616 322856 42668 322862
rect 42616 322798 42668 322804
rect 42708 322856 42760 322862
rect 42708 322798 42760 322804
rect 42720 314226 42748 322798
rect 42892 322788 42944 322794
rect 42892 322730 42944 322736
rect 42708 314220 42760 314226
rect 42708 314162 42760 314168
rect 42524 314084 42576 314090
rect 42524 314026 42576 314032
rect 42708 314084 42760 314090
rect 42708 314026 42760 314032
rect 42352 283675 42564 283703
rect 42340 283212 42392 283218
rect 42340 283154 42392 283160
rect 42352 276214 42380 283154
rect 42536 282334 42564 283675
rect 42524 282328 42576 282334
rect 42524 282270 42576 282276
rect 42340 276208 42392 276214
rect 42340 276150 42392 276156
rect 42536 276026 42564 282270
rect 42352 275998 42564 276026
rect 42352 245614 42380 275998
rect 42720 271930 42748 314026
rect 42800 313472 42852 313478
rect 42904 313426 42932 322730
rect 42852 313420 42932 313426
rect 42800 313414 42932 313420
rect 42812 313398 42932 313414
rect 42708 271924 42760 271930
rect 42708 271866 42760 271872
rect 42524 271244 42576 271250
rect 42524 271186 42576 271192
rect 42340 245608 42392 245614
rect 42340 245550 42392 245556
rect 42536 245546 42564 271186
rect 42524 245540 42576 245546
rect 42524 245482 42576 245488
rect 42340 239964 42392 239970
rect 42340 239906 42392 239912
rect 42352 233034 42380 239906
rect 42616 238128 42668 238134
rect 42616 238070 42668 238076
rect 42340 233028 42392 233034
rect 42340 232970 42392 232976
rect 42628 232898 42656 238070
rect 42340 232892 42392 232898
rect 42340 232834 42392 232840
rect 42616 232892 42668 232898
rect 42616 232834 42668 232840
rect 42352 208418 42380 232834
rect 42720 228682 42748 271866
rect 42812 271250 42840 313398
rect 673564 303618 673592 338098
rect 673656 337550 673684 383182
rect 673748 380934 673776 384270
rect 675312 383253 675340 401542
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675392 384328 675444 384334
rect 675392 384270 675444 384276
rect 675404 383860 675432 384270
rect 675312 383246 675418 383253
rect 675300 383240 675418 383246
rect 675352 383225 675418 383240
rect 675300 383182 675352 383188
rect 675312 383142 675340 383182
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 673736 380928 673788 380934
rect 673736 380870 673788 380876
rect 675407 380727 675887 380783
rect 675407 380175 675887 380231
rect 675407 379531 675887 379587
rect 675312 378901 675418 378929
rect 673736 372360 673788 372366
rect 673736 372302 673788 372308
rect 673644 337544 673696 337550
rect 673644 337486 673696 337492
rect 673552 303612 673604 303618
rect 673552 303554 673604 303560
rect 673656 293622 673684 337486
rect 673748 328098 673776 372302
rect 675312 370925 675340 378901
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675404 372366 675432 372751
rect 675392 372360 675444 372366
rect 675392 372302 675444 372308
rect 675407 371527 675887 371583
rect 675312 370897 675418 370925
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675404 338162 675432 338708
rect 675392 338156 675444 338162
rect 675392 338098 675444 338104
rect 675404 337550 675432 338028
rect 675392 337544 675444 337550
rect 675392 337486 675444 337492
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334975 675887 335031
rect 675407 334331 675887 334387
rect 675312 333701 675418 333729
rect 673736 328092 673788 328098
rect 673736 328034 673788 328040
rect 673644 293616 673696 293622
rect 673644 293558 673696 293564
rect 673644 293480 673696 293486
rect 673644 293422 673696 293428
rect 42800 271244 42852 271250
rect 42800 271186 42852 271192
rect 673656 264994 673684 293422
rect 673748 282130 673776 328034
rect 675312 325725 675340 333701
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675392 328092 675444 328098
rect 675392 328034 675444 328040
rect 675404 327556 675432 328034
rect 675407 326327 675887 326383
rect 675312 325697 675418 325725
rect 675300 303612 675352 303618
rect 675300 303554 675352 303560
rect 675312 293706 675340 303554
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675312 293678 675418 293706
rect 673920 293616 673972 293622
rect 673920 293558 673972 293564
rect 673736 282124 673788 282130
rect 673736 282066 673788 282072
rect 673460 264988 673512 264994
rect 673460 264930 673512 264936
rect 673644 264988 673696 264994
rect 673644 264930 673696 264936
rect 673472 248742 673500 264930
rect 673460 248736 673512 248742
rect 673460 248678 673512 248684
rect 673644 247512 673696 247518
rect 673644 247454 673696 247460
rect 42892 245608 42944 245614
rect 42892 245550 42944 245556
rect 42800 245540 42852 245546
rect 42800 245482 42852 245488
rect 42708 228676 42760 228682
rect 42708 228618 42760 228624
rect 42616 228064 42668 228070
rect 42616 228006 42668 228012
rect 42340 208412 42392 208418
rect 42340 208354 42392 208360
rect 42340 196784 42392 196790
rect 42340 196726 42392 196732
rect 42352 189854 42380 196726
rect 42432 194948 42484 194954
rect 42432 194890 42484 194896
rect 42340 189848 42392 189854
rect 42340 189790 42392 189796
rect 42340 185496 42392 185502
rect 42340 185438 42392 185444
rect 42248 121508 42300 121514
rect 42248 121450 42300 121456
rect 41418 80608 41474 80617
rect 41418 80543 41474 80552
rect 41432 78305 41460 80543
rect 41418 78296 41474 78305
rect 41418 78231 41474 78240
rect 42352 45762 42380 185438
rect 42444 185366 42472 194890
rect 42432 185360 42484 185366
rect 42432 185302 42484 185308
rect 42628 184890 42656 228006
rect 42720 185502 42748 228618
rect 42812 228070 42840 245482
rect 42904 238134 42932 245550
rect 42892 238128 42944 238134
rect 42892 238070 42944 238076
rect 42800 228064 42852 228070
rect 42800 228006 42852 228012
rect 42892 208412 42944 208418
rect 42892 208354 42944 208360
rect 42904 194954 42932 208354
rect 673656 203386 673684 247454
rect 673748 244066 673776 282066
rect 673932 247518 673960 293558
rect 675312 293486 675340 293678
rect 675392 293616 675444 293622
rect 675392 293558 675444 293564
rect 675300 293480 675352 293486
rect 675300 293422 675352 293428
rect 675404 293012 675432 293558
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289975 675887 290031
rect 675407 289331 675887 289387
rect 675312 288701 675418 288729
rect 675312 280725 675340 288701
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675404 282130 675432 282540
rect 675392 282124 675444 282130
rect 675392 282066 675444 282072
rect 675407 281327 675887 281383
rect 675312 280697 675418 280725
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675312 248742 675340 248773
rect 675300 248736 675352 248742
rect 675352 248684 675418 248690
rect 675300 248678 675418 248684
rect 675312 248662 675418 248678
rect 673920 247512 673972 247518
rect 673920 247454 673972 247460
rect 673748 244038 673960 244066
rect 673828 243840 673880 243846
rect 673828 243782 673880 243788
rect 673840 218142 673868 243782
rect 673932 237726 673960 244038
rect 675312 243846 675340 248662
rect 675404 247518 675432 248039
rect 675392 247512 675444 247518
rect 675392 247454 675444 247460
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244975 675887 245031
rect 675407 244331 675887 244387
rect 675300 243840 675352 243846
rect 675300 243782 675352 243788
rect 675312 243701 675418 243729
rect 673920 237720 673972 237726
rect 673920 237662 673972 237668
rect 673932 237386 673960 237662
rect 673920 237380 673972 237386
rect 673920 237322 673972 237328
rect 674104 237380 674156 237386
rect 674104 237322 674156 237328
rect 674116 231810 674144 237322
rect 675312 235725 675340 243701
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675392 237720 675444 237726
rect 675392 237662 675444 237668
rect 675404 237524 675432 237662
rect 675407 236327 675887 236383
rect 675312 235697 675418 235725
rect 674104 231804 674156 231810
rect 674104 231746 674156 231752
rect 674288 231804 674340 231810
rect 674288 231746 674340 231752
rect 673828 218136 673880 218142
rect 673828 218078 673880 218084
rect 673828 218000 673880 218006
rect 673828 217942 673880 217948
rect 673840 212566 673868 217942
rect 674300 212566 674328 231746
rect 673736 212560 673788 212566
rect 673736 212502 673788 212508
rect 673828 212560 673880 212566
rect 673828 212502 673880 212508
rect 674012 212560 674064 212566
rect 674012 212502 674064 212508
rect 674288 212560 674340 212566
rect 674288 212502 674340 212508
rect 673748 203930 673776 212502
rect 673736 203924 673788 203930
rect 673736 203866 673788 203872
rect 673644 203380 673696 203386
rect 673644 203322 673696 203328
rect 673656 203266 673684 203322
rect 673472 203238 673684 203266
rect 42892 194948 42944 194954
rect 42892 194890 42944 194896
rect 42708 185496 42760 185502
rect 42708 185438 42760 185444
rect 42708 185360 42760 185366
rect 42708 185302 42760 185308
rect 42432 184884 42484 184890
rect 42432 184826 42484 184832
rect 42616 184884 42668 184890
rect 42616 184826 42668 184832
rect 42340 45756 42392 45762
rect 42340 45698 42392 45704
rect 42444 45694 42472 184826
rect 42720 149122 42748 185302
rect 673472 157350 673500 203238
rect 673748 203130 673776 203866
rect 673564 203102 673776 203130
rect 673564 158370 673592 203102
rect 674024 198762 674052 212502
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675392 203924 675444 203930
rect 675392 203866 675444 203872
rect 675404 203483 675432 203866
rect 675392 203380 675444 203386
rect 675392 203322 675444 203328
rect 675404 202844 675432 203322
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199775 675887 199831
rect 675407 199131 675887 199187
rect 674012 198756 674064 198762
rect 674012 198698 674064 198704
rect 675208 198756 675260 198762
rect 675208 198698 675260 198704
rect 675220 192166 675248 198698
rect 675312 198614 675432 198642
rect 674748 192160 674800 192166
rect 674748 192102 674800 192108
rect 675208 192160 675260 192166
rect 675208 192102 675260 192108
rect 674760 173942 674788 192102
rect 675312 190525 675340 198614
rect 675404 198492 675432 198614
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675404 192166 675432 192372
rect 675392 192160 675444 192166
rect 675392 192102 675444 192108
rect 675407 191127 675887 191183
rect 675312 190497 675418 190525
rect 673828 173936 673880 173942
rect 673828 173878 673880 173884
rect 674748 173936 674800 173942
rect 674748 173878 674800 173884
rect 673552 158364 673604 158370
rect 673552 158306 673604 158312
rect 673460 157344 673512 157350
rect 673460 157286 673512 157292
rect 42524 149116 42576 149122
rect 42524 149058 42576 149064
rect 42708 149116 42760 149122
rect 42708 149058 42760 149064
rect 42536 129690 42564 149058
rect 42536 129662 42748 129690
rect 42720 110498 42748 129662
rect 44732 121508 44784 121514
rect 44732 121450 44784 121456
rect 44744 115938 44772 121450
rect 42984 115932 43036 115938
rect 42984 115874 43036 115880
rect 44732 115932 44784 115938
rect 44732 115874 44784 115880
rect 42524 110492 42576 110498
rect 42524 110434 42576 110440
rect 42708 110492 42760 110498
rect 42708 110434 42760 110440
rect 42536 91066 42564 110434
rect 42996 110401 43024 115874
rect 673472 112130 673500 157286
rect 673564 112810 673592 158306
rect 673840 154601 673868 173878
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675404 158370 675432 158508
rect 675392 158364 675444 158370
rect 675392 158306 675444 158312
rect 675404 157350 675432 157828
rect 675392 157344 675444 157350
rect 675392 157286 675444 157292
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154775 675887 154831
rect 673642 154592 673698 154601
rect 673642 154527 673698 154536
rect 673826 154592 673882 154601
rect 673826 154527 673882 154536
rect 673656 147150 673684 154527
rect 675407 154131 675887 154187
rect 675312 153501 675418 153529
rect 673644 147144 673696 147150
rect 673644 147086 673696 147092
rect 675024 147144 675076 147150
rect 675024 147086 675076 147092
rect 675036 140690 675064 147086
rect 675312 145525 675340 153501
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675404 147150 675432 147356
rect 675392 147144 675444 147150
rect 675392 147086 675444 147092
rect 675407 146127 675887 146183
rect 675312 145497 675418 145525
rect 674012 140684 674064 140690
rect 674012 140626 674064 140632
rect 675024 140684 675076 140690
rect 675024 140626 675076 140632
rect 674024 116006 674052 140626
rect 673828 116000 673880 116006
rect 673828 115942 673880 115948
rect 674012 116000 674064 116006
rect 674012 115942 674064 115948
rect 673840 115870 673868 115942
rect 673828 115864 673880 115870
rect 673828 115806 673880 115812
rect 675024 115864 675076 115870
rect 675024 115806 675076 115812
rect 673552 112804 673604 112810
rect 673552 112746 673604 112752
rect 673460 112124 673512 112130
rect 673460 112066 673512 112072
rect 42982 110392 43038 110401
rect 42982 110327 43038 110336
rect 42996 96665 43024 110327
rect 42982 96656 43038 96665
rect 42982 96591 43038 96600
rect 44638 96656 44694 96665
rect 44638 96591 44694 96600
rect 42536 91038 42748 91066
rect 42720 80617 42748 91038
rect 44652 82890 44680 96591
rect 44640 82884 44692 82890
rect 44640 82826 44692 82832
rect 44824 82816 44876 82822
rect 44824 82758 44876 82764
rect 44836 82634 44864 82758
rect 44836 82606 44956 82634
rect 42706 80608 42762 80617
rect 42706 80543 42762 80552
rect 42432 45688 42484 45694
rect 42432 45630 42484 45636
rect 42720 45626 42748 80543
rect 42708 45620 42760 45626
rect 42708 45562 42760 45568
rect 44928 45558 44956 82606
rect 140964 45756 141016 45762
rect 140964 45698 141016 45704
rect 44916 45552 44968 45558
rect 44916 45494 44968 45500
rect 93768 41608 93820 41614
rect 121552 41608 121604 41614
rect 93768 41550 93820 41556
rect 121288 41556 121552 41562
rect 140872 41608 140924 41614
rect 121288 41550 121604 41556
rect 140700 41556 140872 41562
rect 140700 41550 140924 41556
rect 93780 40225 93808 41550
rect 121288 41546 121592 41550
rect 140700 41546 140912 41550
rect 121276 41540 121592 41546
rect 121328 41534 121592 41540
rect 140688 41540 140912 41546
rect 121276 41482 121328 41488
rect 140740 41534 140912 41540
rect 140688 41482 140740 41488
rect 135168 40248 135220 40254
rect 93766 40216 93822 40225
rect 93766 40151 93822 40160
rect 135166 40216 135168 40225
rect 135220 40216 135222 40225
rect 140976 40202 141004 45698
rect 143632 45688 143684 45694
rect 143632 45630 143684 45636
rect 143540 45620 143592 45626
rect 143540 45562 143592 45568
rect 143552 40497 143580 45562
rect 143644 44402 143672 45630
rect 527456 45620 527508 45626
rect 527456 45562 527508 45568
rect 195980 45552 196032 45558
rect 195980 45494 196032 45500
rect 516324 45552 516376 45558
rect 516324 45494 516376 45500
rect 195992 44470 196020 45494
rect 405648 44804 405700 44810
rect 405648 44746 405700 44752
rect 411260 44804 411312 44810
rect 411260 44746 411312 44752
rect 359372 44736 359424 44742
rect 359372 44678 359424 44684
rect 354404 44532 354456 44538
rect 354404 44474 354456 44480
rect 195980 44464 196032 44470
rect 195980 44406 196032 44412
rect 304540 44464 304592 44470
rect 304540 44406 304592 44412
rect 143632 44396 143684 44402
rect 143632 44338 143684 44344
rect 145104 44396 145156 44402
rect 145104 44338 145156 44344
rect 195336 44396 195388 44402
rect 195336 44338 195388 44344
rect 144644 40792 144696 40798
rect 144644 40734 144696 40740
rect 143538 40488 143594 40497
rect 143538 40423 143594 40432
rect 143540 40248 143592 40254
rect 143078 40216 143134 40225
rect 140976 40174 141036 40202
rect 135166 40151 135222 40160
rect 141008 40118 141036 40174
rect 143078 40151 143134 40160
rect 143538 40216 143540 40225
rect 143592 40216 143594 40225
rect 143538 40151 143594 40160
rect 143092 40118 143120 40151
rect 144656 40118 144684 40734
rect 145116 40202 145144 44338
rect 188528 44328 188580 44334
rect 188528 44270 188580 44276
rect 192852 44328 192904 44334
rect 192852 44270 192904 44276
rect 186688 44260 186740 44266
rect 186688 44202 186740 44208
rect 146300 42016 146352 42022
rect 146300 41958 146352 41964
rect 146312 40798 146340 41958
rect 186700 41820 186728 44202
rect 149612 41812 149664 41818
rect 149612 41754 149664 41760
rect 146300 40792 146352 40798
rect 146300 40734 146352 40740
rect 149624 40361 149652 41754
rect 168288 41744 168340 41750
rect 187327 41713 187383 42193
rect 188540 41970 188568 44270
rect 188448 41954 188568 41970
rect 187700 41948 187752 41954
rect 187700 41890 187752 41896
rect 188436 41948 188568 41954
rect 188488 41942 188568 41948
rect 188436 41890 188488 41896
rect 187712 41818 187740 41890
rect 188540 41820 188568 41942
rect 189198 41818 189304 41834
rect 191038 41818 191144 41834
rect 192234 41818 192340 41834
rect 192864 41820 192892 44270
rect 194692 44260 194744 44266
rect 194692 44202 194744 44208
rect 193522 41818 193628 41834
rect 187700 41812 187752 41818
rect 189198 41812 189316 41818
rect 189198 41806 189264 41812
rect 187700 41754 187752 41760
rect 191038 41812 191156 41818
rect 191038 41806 191104 41812
rect 189264 41754 189316 41760
rect 192234 41812 192352 41818
rect 192234 41806 192300 41812
rect 191104 41754 191156 41760
rect 193522 41812 193640 41818
rect 193522 41806 193588 41812
rect 192300 41754 192352 41760
rect 193588 41754 193640 41760
rect 194043 41713 194099 42193
rect 194704 41820 194732 44202
rect 195348 41820 195376 44338
rect 195992 41820 196020 44406
rect 199660 44396 199712 44402
rect 199660 44338 199712 44344
rect 200856 44396 200908 44402
rect 200856 44338 200908 44344
rect 241336 44396 241388 44402
rect 241336 44338 241388 44344
rect 251088 44396 251140 44402
rect 251088 44338 251140 44344
rect 199672 44266 199700 44338
rect 199660 44260 199712 44266
rect 199660 44202 199712 44208
rect 198924 41948 198976 41954
rect 198924 41890 198976 41896
rect 198464 41880 198516 41886
rect 196452 41828 198464 41834
rect 198936 41834 198964 41890
rect 196452 41822 198516 41828
rect 196452 41818 198504 41822
rect 198844 41818 199042 41834
rect 199672 41820 199700 44202
rect 200120 41880 200172 41886
rect 200868 41834 200896 44338
rect 201500 44328 201552 44334
rect 201500 44270 201552 44276
rect 200172 41828 200896 41834
rect 200120 41822 200896 41828
rect 200132 41820 200896 41822
rect 201512 41820 201540 44270
rect 196440 41812 198504 41818
rect 196492 41806 198504 41812
rect 198832 41812 199042 41818
rect 196440 41754 196492 41760
rect 198884 41806 199042 41812
rect 200132 41806 200882 41820
rect 198832 41754 198884 41760
rect 168288 41686 168340 41692
rect 168300 41546 168328 41686
rect 168288 41540 168340 41546
rect 168288 41482 168340 41488
rect 241348 40510 241376 44338
rect 251100 42090 251128 44338
rect 297088 44328 297140 44334
rect 297088 44270 297140 44276
rect 299572 44328 299624 44334
rect 299572 44270 299624 44276
rect 295248 44192 295300 44198
rect 295248 44134 295300 44140
rect 251088 42084 251140 42090
rect 251088 42026 251140 42032
rect 255228 42084 255280 42090
rect 255228 42026 255280 42032
rect 255240 41886 255268 42026
rect 255228 41880 255280 41886
rect 255228 41822 255280 41828
rect 295260 41834 295288 44134
rect 297100 41834 297128 44270
rect 297640 41880 297692 41886
rect 295260 41806 295311 41834
rect 297100 41806 297151 41834
rect 299584 41834 299612 44270
rect 303896 44260 303948 44266
rect 303896 44202 303948 44208
rect 303252 44192 303304 44198
rect 303252 44134 303304 44140
rect 300676 41880 300728 41886
rect 297692 41828 297795 41834
rect 297640 41822 297795 41828
rect 297652 41806 297795 41822
rect 299584 41806 299635 41834
rect 300728 41828 302280 41834
rect 300676 41822 302280 41828
rect 300688 41818 302280 41822
rect 300688 41812 302292 41818
rect 300688 41806 302240 41812
rect 302240 41754 302292 41760
rect 302643 41713 302699 42193
rect 303264 41834 303292 44134
rect 303908 41834 303936 44202
rect 304552 41834 304580 44406
rect 306380 44396 306432 44402
rect 306380 44338 306432 44344
rect 309416 44396 309468 44402
rect 309416 44338 309468 44344
rect 352564 44396 352616 44402
rect 352564 44338 352616 44344
rect 305736 44328 305788 44334
rect 305736 44270 305788 44276
rect 305748 41834 305776 44270
rect 306392 41834 306420 44338
rect 308220 44260 308272 44266
rect 308220 44202 308272 44208
rect 303264 41806 303315 41834
rect 303908 41806 303959 41834
rect 304552 41806 304603 41834
rect 305012 41818 305155 41834
rect 305000 41812 305155 41818
rect 305052 41806 305155 41812
rect 305748 41806 305799 41834
rect 306300 41818 306443 41834
rect 306288 41812 306443 41818
rect 305000 41754 305052 41760
rect 306340 41806 306443 41812
rect 306288 41754 306340 41760
rect 306967 41713 307023 42193
rect 307484 41948 307536 41954
rect 307484 41890 307536 41896
rect 307496 41834 307524 41890
rect 308232 41834 308260 44202
rect 309428 41834 309456 44338
rect 351920 44328 351972 44334
rect 351920 44270 351972 44276
rect 350080 44192 350132 44198
rect 350080 44134 350132 44140
rect 307496 41806 307639 41834
rect 308232 41806 308283 41834
rect 308835 41806 309479 41834
rect 310095 41713 310151 42193
rect 349618 41848 349674 41857
rect 350092 41820 350120 44134
rect 351932 41820 351960 44270
rect 352576 41820 352604 44338
rect 354416 44334 354444 44474
rect 359384 44402 359412 44678
rect 405660 44577 405688 44746
rect 406752 44736 406804 44742
rect 406752 44678 406804 44684
rect 386418 44568 386474 44577
rect 360568 44532 360620 44538
rect 360568 44474 360620 44480
rect 360660 44532 360712 44538
rect 405646 44568 405702 44577
rect 386418 44503 386420 44512
rect 360660 44474 360712 44480
rect 386472 44503 386474 44512
rect 399668 44532 399720 44538
rect 386420 44474 386472 44480
rect 406764 44538 406792 44678
rect 411272 44538 411300 44746
rect 425060 44736 425112 44742
rect 425060 44678 425112 44684
rect 444196 44736 444248 44742
rect 444196 44678 444248 44684
rect 483018 44704 483074 44713
rect 425072 44606 425100 44678
rect 425060 44600 425112 44606
rect 425060 44542 425112 44548
rect 405646 44503 405702 44512
rect 406752 44532 406804 44538
rect 399668 44474 399720 44480
rect 406752 44474 406804 44480
rect 411260 44532 411312 44538
rect 411260 44474 411312 44480
rect 355416 44396 355468 44402
rect 355416 44338 355468 44344
rect 359372 44396 359424 44402
rect 359372 44338 359424 44344
rect 354404 44328 354456 44334
rect 354404 44270 354456 44276
rect 355428 44282 355456 44338
rect 358728 44328 358780 44334
rect 354416 41820 354444 44270
rect 355428 44266 355640 44282
rect 358728 44270 358780 44276
rect 355428 44260 355652 44266
rect 355428 44254 355600 44260
rect 355600 44202 355652 44208
rect 355612 41834 355640 44202
rect 358740 44198 358768 44270
rect 358084 44192 358136 44198
rect 358084 44134 358136 44140
rect 358728 44192 358780 44198
rect 358728 44134 358780 44140
rect 355612 41820 356914 41834
rect 355626 41806 356914 41820
rect 349618 41783 349674 41792
rect 314580 41682 314700 41698
rect 314568 41676 314712 41682
rect 314620 41670 314660 41676
rect 314568 41618 314620 41624
rect 314660 41618 314712 41624
rect 349632 41614 349660 41783
rect 357443 41713 357499 42193
rect 358096 41820 358124 44134
rect 358740 41820 358768 44134
rect 359384 41820 359412 44338
rect 360580 44334 360608 44474
rect 360672 44402 360700 44474
rect 360660 44396 360712 44402
rect 360660 44338 360712 44344
rect 364248 44396 364300 44402
rect 364248 44338 364300 44344
rect 360568 44328 360620 44334
rect 360568 44270 360620 44276
rect 359924 44260 359976 44266
rect 359924 44202 359976 44208
rect 359936 41834 359964 44202
rect 360016 41880 360068 41886
rect 359936 41828 360016 41834
rect 359936 41822 360068 41828
rect 359936 41820 360056 41822
rect 360580 41820 360608 44270
rect 363052 44260 363104 44266
rect 363052 44202 363104 44208
rect 361120 41880 361172 41886
rect 361172 41828 361238 41834
rect 361120 41822 361238 41828
rect 359950 41806 360056 41820
rect 361132 41806 361238 41822
rect 361767 41713 361823 42193
rect 362500 41948 362552 41954
rect 362420 41908 362500 41936
rect 362420 41857 362448 41908
rect 362500 41890 362552 41896
rect 362406 41848 362462 41857
rect 363064 41820 363092 44202
rect 363512 41880 363564 41886
rect 364260 41834 364288 44338
rect 399680 44334 399708 44474
rect 399668 44328 399720 44334
rect 399668 44270 399720 44276
rect 404912 44192 404964 44198
rect 404912 44134 404964 44140
rect 363564 41828 364288 41834
rect 363512 41822 364288 41828
rect 363524 41820 364288 41822
rect 363524 41806 364274 41820
rect 362406 41783 362462 41792
rect 364895 41713 364951 42193
rect 367098 41984 367154 41993
rect 367098 41919 367100 41928
rect 367152 41919 367154 41928
rect 386142 41984 386198 41993
rect 386142 41919 386198 41928
rect 367100 41890 367152 41896
rect 349620 41608 349672 41614
rect 349620 41550 349672 41556
rect 386156 41562 386184 41919
rect 404924 41820 404952 44134
rect 405527 41713 405583 42193
rect 406764 41820 406792 44474
rect 414204 44464 414256 44470
rect 414204 44406 414256 44412
rect 419816 44464 419868 44470
rect 419816 44406 419868 44412
rect 444208 44418 444236 44678
rect 483018 44639 483020 44648
rect 483072 44639 483074 44648
rect 502062 44704 502118 44713
rect 502062 44639 502118 44648
rect 483020 44610 483072 44616
rect 461492 44600 461544 44606
rect 461492 44542 461544 44548
rect 469128 44600 469180 44606
rect 469220 44600 469272 44606
rect 469180 44548 469220 44554
rect 469128 44542 469272 44548
rect 444288 44532 444340 44538
rect 444288 44474 444340 44480
rect 444300 44418 444328 44474
rect 407396 44396 407448 44402
rect 407396 44338 407448 44344
rect 410432 44396 410484 44402
rect 410432 44338 410484 44344
rect 407408 41820 407436 44338
rect 410444 41834 410472 44338
rect 413560 44328 413612 44334
rect 413560 44270 413612 44276
rect 411076 44260 411128 44266
rect 411076 44202 411128 44208
rect 410524 41880 410576 41886
rect 409262 41818 409368 41834
rect 410444 41828 410524 41834
rect 410444 41822 410576 41828
rect 410444 41820 410564 41822
rect 411088 41820 411116 44202
rect 412916 44192 412968 44198
rect 412916 44134 412968 44140
rect 411812 41880 411864 41886
rect 411746 41828 411812 41834
rect 411746 41822 411864 41828
rect 412243 41834 412299 42193
rect 409262 41812 409380 41818
rect 409262 41806 409328 41812
rect 410458 41806 410564 41820
rect 411746 41806 411852 41822
rect 412243 41818 412404 41834
rect 412928 41820 412956 44134
rect 413572 41820 413600 44270
rect 414216 41820 414244 44406
rect 419080 44396 419132 44402
rect 419080 44338 419132 44344
rect 417884 44328 417936 44334
rect 417884 44270 417936 44276
rect 414848 41880 414900 41886
rect 414782 41828 414848 41834
rect 416136 41880 416188 41886
rect 414782 41822 414900 41828
rect 412243 41812 412416 41818
rect 412243 41806 412364 41812
rect 409328 41754 409380 41760
rect 412243 41713 412299 41806
rect 414782 41806 414888 41822
rect 415228 41818 415426 41834
rect 415216 41812 415426 41818
rect 412364 41754 412416 41760
rect 415268 41806 415426 41812
rect 416070 41828 416136 41834
rect 416070 41822 416188 41828
rect 416070 41806 416176 41822
rect 415216 41754 415268 41760
rect 416567 41713 416623 42193
rect 417068 41818 417266 41834
rect 417896 41820 417924 44270
rect 418540 41886 418568 41917
rect 418528 41880 418580 41886
rect 418462 41828 418528 41834
rect 419092 41834 419120 44338
rect 419828 44266 419856 44406
rect 444208 44390 444328 44418
rect 419724 44260 419776 44266
rect 419724 44202 419776 44208
rect 419816 44260 419868 44266
rect 419816 44202 419868 44208
rect 419736 42193 419764 44202
rect 459652 44192 459704 44198
rect 459652 44134 459704 44140
rect 418580 41828 419120 41834
rect 418462 41820 419120 41828
rect 419695 41820 419764 42193
rect 459664 41834 459692 44134
rect 417056 41812 417266 41818
rect 417108 41806 417266 41812
rect 418462 41806 419106 41820
rect 417056 41754 417108 41760
rect 419695 41713 419751 41820
rect 459664 41806 459711 41834
rect 460327 41713 460383 42193
rect 461504 41834 461532 44542
rect 469140 44526 469260 44542
rect 502076 44418 502104 44639
rect 516336 44538 516364 45494
rect 502248 44532 502300 44538
rect 502248 44474 502300 44480
rect 516324 44532 516376 44538
rect 516324 44474 516376 44480
rect 502260 44418 502288 44474
rect 462136 44396 462188 44402
rect 462136 44338 462188 44344
rect 465172 44396 465224 44402
rect 465172 44338 465224 44344
rect 473820 44396 473872 44402
rect 502076 44390 502288 44418
rect 473820 44338 473872 44344
rect 462148 41834 462176 44338
rect 464160 41880 464212 41886
rect 461504 41806 461551 41834
rect 462148 41806 462195 41834
rect 464035 41828 464160 41834
rect 464035 41822 464212 41828
rect 465184 41834 465212 44338
rect 468300 44328 468352 44334
rect 465814 44296 465870 44305
rect 468300 44270 468352 44276
rect 472624 44328 472676 44334
rect 472624 44270 472676 44276
rect 465814 44231 465870 44240
rect 465828 41834 465856 44231
rect 467656 44192 467708 44198
rect 467656 44134 467708 44140
rect 467043 41834 467099 42193
rect 467196 41880 467248 41886
rect 464035 41806 464200 41822
rect 465184 41818 465396 41834
rect 465184 41812 465408 41818
rect 465184 41806 465356 41812
rect 465828 41806 465875 41834
rect 466380 41818 466519 41834
rect 466368 41812 466519 41818
rect 465356 41754 465408 41760
rect 466420 41806 466519 41812
rect 467043 41828 467196 41834
rect 467043 41822 467248 41828
rect 467668 41834 467696 44134
rect 468312 41834 468340 44270
rect 468944 44260 468996 44266
rect 468944 44202 468996 44208
rect 468956 41834 468984 44202
rect 470048 41880 470100 41886
rect 467043 41806 467236 41822
rect 467668 41806 467715 41834
rect 468312 41806 468359 41834
rect 468956 41806 469003 41834
rect 469555 41818 469720 41834
rect 470968 41880 471020 41886
rect 470100 41828 470199 41834
rect 470048 41822 470199 41828
rect 469555 41812 469732 41818
rect 469555 41806 469680 41812
rect 466368 41754 466420 41760
rect 467043 41713 467099 41806
rect 470060 41806 470199 41822
rect 470843 41828 470968 41834
rect 470843 41822 471020 41828
rect 470843 41806 471008 41822
rect 469680 41754 469732 41760
rect 471367 41713 471423 42193
rect 472636 41834 472664 44270
rect 473084 41880 473136 41886
rect 471900 41818 472039 41834
rect 471888 41812 472039 41818
rect 471940 41806 472039 41812
rect 472636 41806 472683 41834
rect 473832 41834 473860 44338
rect 474462 44296 474518 44305
rect 474462 44231 474518 44240
rect 474476 42193 474504 44231
rect 514484 44192 514536 44198
rect 514484 44134 514536 44140
rect 473136 41828 473879 41834
rect 473084 41822 473879 41828
rect 473096 41806 473879 41822
rect 474476 41806 474551 42193
rect 514496 41820 514524 44134
rect 471888 41754 471940 41760
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 516336 41820 516364 44474
rect 516968 44396 517020 44402
rect 516968 44338 517020 44344
rect 520004 44396 520056 44402
rect 520004 44338 520056 44344
rect 516980 41820 517008 44338
rect 518806 44296 518862 44305
rect 518806 44231 518862 44240
rect 518820 41820 518848 44231
rect 520016 41834 520044 44338
rect 523132 44328 523184 44334
rect 523132 44270 523184 44276
rect 524970 44296 525026 44305
rect 523144 44198 523172 44270
rect 523776 44260 523828 44266
rect 524970 44231 525026 44240
rect 523776 44202 523828 44208
rect 522488 44192 522540 44198
rect 522488 44134 522540 44140
rect 523132 44192 523184 44198
rect 523132 44134 523184 44140
rect 520096 41880 520148 41886
rect 520016 41828 520096 41834
rect 520016 41822 520148 41828
rect 520016 41820 520136 41822
rect 520030 41806 520136 41820
rect 520647 41713 520703 42193
rect 521200 41880 521252 41886
rect 521252 41828 521318 41834
rect 521200 41822 521318 41828
rect 521212 41806 521318 41822
rect 521843 41713 521899 42193
rect 522500 41820 522528 44134
rect 523144 41820 523172 44134
rect 523788 41820 523816 44202
rect 524984 42193 525012 44231
rect 527468 44198 527496 45562
rect 527456 44192 527508 44198
rect 527456 44134 527508 44140
rect 524236 41880 524288 41886
rect 524288 41828 524354 41834
rect 524236 41822 524354 41828
rect 524248 41806 524354 41822
rect 524971 41713 525027 42193
rect 525524 41880 525576 41886
rect 525576 41828 525642 41834
rect 525524 41822 525642 41828
rect 525536 41806 525642 41822
rect 526167 41713 526223 42193
rect 526732 41818 526838 41834
rect 527468 41820 527496 44134
rect 673472 42770 673500 112066
rect 673564 45626 673592 112746
rect 675036 102338 675064 115806
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675404 112810 675432 113283
rect 675392 112804 675444 112810
rect 675392 112746 675444 112752
rect 675404 112130 675432 112639
rect 675392 112124 675444 112130
rect 675392 112066 675444 112072
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 109575 675887 109631
rect 675407 108931 675887 108987
rect 675312 108310 675418 108338
rect 673644 102332 673696 102338
rect 673644 102274 673696 102280
rect 675024 102332 675076 102338
rect 675024 102274 675076 102280
rect 673552 45620 673604 45626
rect 673552 45562 673604 45568
rect 673656 45558 673684 102274
rect 675312 100314 675340 108310
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675392 102332 675444 102338
rect 675392 102274 675444 102280
rect 675404 102151 675432 102274
rect 675407 100927 675887 100983
rect 675312 100286 675418 100314
rect 673644 45552 673696 45558
rect 673644 45494 673696 45500
rect 576768 42764 576820 42770
rect 576768 42706 576820 42712
rect 673460 42764 673512 42770
rect 673460 42706 673512 42712
rect 527916 41880 527968 41886
rect 527968 41828 528678 41834
rect 527916 41822 528678 41828
rect 526720 41812 526838 41818
rect 526772 41806 526838 41812
rect 527928 41806 528678 41822
rect 526720 41754 526772 41760
rect 529295 41713 529351 42193
rect 576780 42022 576808 42706
rect 569132 42016 569184 42022
rect 569132 41958 569184 41964
rect 576768 42016 576820 42022
rect 576768 41958 576820 41964
rect 386328 41676 386380 41682
rect 386328 41618 386380 41624
rect 386340 41562 386368 41618
rect 507860 41608 507912 41614
rect 386156 41534 386368 41562
rect 507780 41556 507860 41562
rect 507780 41550 507912 41556
rect 507780 41546 507900 41550
rect 507768 41540 507900 41546
rect 507820 41534 507900 41540
rect 507768 41482 507820 41488
rect 240748 40482 241376 40510
rect 240748 40384 240776 40482
rect 149610 40352 149666 40361
rect 149610 40287 149666 40296
rect 145103 40174 145144 40202
rect 240560 40228 240950 40384
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143080 40112 143132 40118
rect 143080 40054 143132 40060
rect 144644 40112 144696 40118
rect 144644 40054 144696 40060
rect 141008 39984 141036 40054
rect 141667 39934 141813 40000
rect 143092 39916 143120 40054
rect 144656 39916 144684 40054
rect 145103 40000 145131 40174
rect 240560 40168 240732 40228
rect 240792 40168 240950 40228
rect 569144 40225 569172 41958
rect 240560 40008 240950 40168
rect 569130 40216 569186 40225
rect 569130 40151 569186 40160
rect 145091 39706 145143 40000
<< via2 >>
rect 342164 997414 342224 997474
rect 42246 870032 42302 870088
rect 677506 818372 677562 818408
rect 677506 818352 677508 818372
rect 677508 818352 677560 818372
rect 677560 818352 677562 818372
rect 673734 521600 673790 521656
rect 674010 521600 674066 521656
rect 677690 513748 677692 513768
rect 677692 513748 677744 513768
rect 677744 513748 677746 513768
rect 677690 513712 677746 513748
rect 41418 80552 41474 80608
rect 41418 78240 41474 78296
rect 673642 154536 673698 154592
rect 673826 154536 673882 154592
rect 42982 110336 43038 110392
rect 42982 96600 43038 96656
rect 44638 96600 44694 96656
rect 42706 80552 42762 80608
rect 93766 40160 93822 40216
rect 135166 40196 135168 40216
rect 135168 40196 135220 40216
rect 135220 40196 135222 40216
rect 135166 40160 135222 40196
rect 143538 40432 143594 40488
rect 143078 40160 143134 40216
rect 143538 40196 143540 40216
rect 143540 40196 143592 40216
rect 143592 40196 143594 40216
rect 143538 40160 143594 40196
rect 349618 41792 349674 41848
rect 386418 44532 386474 44568
rect 386418 44512 386420 44532
rect 386420 44512 386472 44532
rect 386472 44512 386474 44532
rect 405646 44512 405702 44568
rect 362406 41792 362462 41848
rect 367098 41948 367154 41984
rect 367098 41928 367100 41948
rect 367100 41928 367152 41948
rect 367152 41928 367154 41948
rect 386142 41928 386198 41984
rect 483018 44668 483074 44704
rect 483018 44648 483020 44668
rect 483020 44648 483072 44668
rect 483072 44648 483074 44668
rect 502062 44648 502118 44704
rect 465814 44240 465870 44296
rect 474462 44240 474518 44296
rect 518806 44240 518862 44296
rect 524970 44240 525026 44296
rect 149610 40296 149666 40352
rect 240732 40168 240792 40228
rect 569130 40160 569186 40216
<< metal3 >>
rect 333499 997600 338279 1002770
rect 343478 997600 348258 1002770
rect 575699 997600 580479 1004102
rect 585678 997600 590458 1004952
rect 342159 997478 342229 997479
rect 343590 997478 343650 997600
rect 342159 997474 343650 997478
rect 342159 997414 342164 997474
rect 342224 997418 343650 997474
rect 342224 997414 342229 997418
rect 342159 997409 342229 997414
rect 38220 922151 39600 926939
rect 678000 917700 679380 922500
rect 38220 912100 39600 916900
rect 678000 907660 679380 912448
rect 42241 870090 42307 870093
rect 39622 870088 42307 870090
rect 39622 870032 42246 870088
rect 42302 870032 42307 870088
rect 39622 870030 42307 870032
rect 39622 869924 39682 870030
rect 42241 870027 42307 870030
rect 32648 837678 40000 842458
rect 33497 827699 39999 832479
rect 677600 828521 680592 833301
rect 677600 818542 680592 823322
rect 677501 818410 677567 818413
rect 677734 818410 677794 818542
rect 677501 818408 677794 818410
rect 677501 818352 677506 818408
rect 677562 818352 677794 818408
rect 677501 818350 677794 818352
rect 677501 818347 677567 818350
rect 673729 521658 673795 521661
rect 674005 521658 674071 521661
rect 673729 521656 674071 521658
rect 673729 521600 673734 521656
rect 673790 521600 674010 521656
rect 674066 521600 674071 521656
rect 673729 521598 674071 521600
rect 673729 521595 673795 521598
rect 674005 521595 674071 521598
rect 677734 513773 677794 514012
rect 677685 513768 677794 513773
rect 677685 513712 677690 513768
rect 677746 513712 677794 513768
rect 677685 513710 677794 513712
rect 677685 513707 677751 513710
rect 37008 493078 40000 497858
rect 37008 483099 40000 487879
rect 678000 469900 685920 474700
rect 678000 459860 685920 464648
rect 31680 450951 39600 455739
rect 31680 440900 39600 445700
rect 673637 154594 673703 154597
rect 673821 154594 673887 154597
rect 673637 154592 673887 154594
rect 673637 154536 673642 154592
rect 673698 154536 673826 154592
rect 673882 154536 673887 154592
rect 673637 154534 673887 154536
rect 673637 154531 673703 154534
rect 673821 154531 673887 154534
rect 36040 120278 40000 125058
rect 36040 110394 40000 115079
rect 42977 110394 43043 110397
rect 36040 110392 43043 110394
rect 36040 110336 42982 110392
rect 43038 110336 43043 110392
rect 36040 110334 43043 110336
rect 36040 110299 40000 110334
rect 42977 110331 43043 110334
rect 42977 96658 43043 96661
rect 44633 96658 44699 96661
rect 42977 96656 44699 96658
rect 42977 96600 42982 96656
rect 43038 96600 44638 96656
rect 44694 96600 44699 96656
rect 42977 96598 44699 96600
rect 42977 96595 43043 96598
rect 44633 96595 44699 96598
rect 38220 78298 39600 82939
rect 41413 80610 41479 80613
rect 42701 80610 42767 80613
rect 41413 80608 42767 80610
rect 41413 80552 41418 80608
rect 41474 80552 42706 80608
rect 42762 80552 42767 80608
rect 41413 80550 42767 80552
rect 41413 80547 41479 80550
rect 42701 80547 42767 80550
rect 41413 78298 41479 78301
rect 38220 78296 41479 78298
rect 38220 78240 41418 78296
rect 41474 78240 41479 78296
rect 38220 78238 41479 78240
rect 38220 78151 39600 78238
rect 41413 78235 41479 78238
rect 38220 68100 39600 72900
rect 483013 44706 483079 44709
rect 502057 44706 502123 44709
rect 483013 44704 502123 44706
rect 483013 44648 483018 44704
rect 483074 44648 502062 44704
rect 502118 44648 502123 44704
rect 483013 44646 502123 44648
rect 483013 44643 483079 44646
rect 502057 44643 502123 44646
rect 386413 44570 386479 44573
rect 405641 44570 405707 44573
rect 386413 44568 405707 44570
rect 386413 44512 386418 44568
rect 386474 44512 405646 44568
rect 405702 44512 405707 44568
rect 386413 44510 405707 44512
rect 386413 44507 386479 44510
rect 405641 44507 405707 44510
rect 465809 44298 465875 44301
rect 474457 44298 474523 44301
rect 465809 44296 474523 44298
rect 465809 44240 465814 44296
rect 465870 44240 474462 44296
rect 474518 44240 474523 44296
rect 465809 44238 474523 44240
rect 465809 44235 465875 44238
rect 474457 44235 474523 44238
rect 518801 44298 518867 44301
rect 524965 44298 525031 44301
rect 518801 44296 525031 44298
rect 518801 44240 518806 44296
rect 518862 44240 524970 44296
rect 525026 44240 525031 44296
rect 518801 44238 525031 44240
rect 518801 44235 518867 44238
rect 524965 44235 525031 44238
rect 367093 41986 367159 41989
rect 386137 41986 386203 41989
rect 367093 41984 386203 41986
rect 367093 41928 367098 41984
rect 367154 41928 386142 41984
rect 386198 41928 386203 41984
rect 367093 41926 386203 41928
rect 367093 41923 367159 41926
rect 386137 41923 386203 41926
rect 349613 41850 349679 41853
rect 362401 41850 362467 41853
rect 349613 41848 362467 41850
rect 349613 41792 349618 41848
rect 349674 41792 362406 41848
rect 362462 41792 362467 41848
rect 349613 41790 362467 41792
rect 349613 41787 349679 41790
rect 362401 41787 362467 41790
rect 143533 40490 143599 40493
rect 143533 40488 145850 40490
rect 143533 40432 143538 40488
rect 143594 40432 145850 40488
rect 143533 40430 145850 40432
rect 143533 40427 143599 40430
rect 145790 40354 145850 40430
rect 149605 40354 149671 40357
rect 145790 40352 149671 40354
rect 145790 40296 149610 40352
rect 149666 40296 149671 40352
rect 145790 40294 149671 40296
rect 93761 40218 93827 40221
rect 135161 40218 135227 40221
rect 91142 40216 93827 40218
rect 91142 40160 93766 40216
rect 93822 40160 93827 40216
rect 91142 40158 93827 40160
rect 78942 32648 83722 40000
rect 91142 39999 91202 40158
rect 93761 40155 93827 40158
rect 133094 40216 135227 40218
rect 133094 40160 135166 40216
rect 135222 40160 135227 40216
rect 133094 40158 135227 40160
rect 88921 33497 93701 39999
rect 133094 39984 133154 40158
rect 135161 40155 135227 40158
rect 143073 40218 143139 40221
rect 143533 40218 143599 40221
rect 143073 40216 143458 40218
rect 143073 40160 143078 40216
rect 143134 40160 143458 40216
rect 143073 40158 143458 40160
rect 143073 40155 143139 40158
rect 141667 38178 141813 40000
rect 143398 39984 143458 40158
rect 143533 40216 144010 40218
rect 143533 40160 143538 40216
rect 143594 40160 144010 40216
rect 143533 40158 144010 40160
rect 143533 40155 143599 40158
rect 143950 39984 144010 40158
rect 145838 40014 145898 40294
rect 149605 40291 149671 40294
rect 145820 39954 145898 40014
rect 239730 40210 240114 40378
rect 239730 40146 239894 40210
rect 239958 40146 240114 40210
rect 239730 39990 240114 40146
rect 240560 40233 240950 40384
rect 240560 40163 240727 40233
rect 240797 40163 240950 40233
rect 240560 40008 240950 40163
rect 569125 40218 569191 40221
rect 569125 40216 569234 40218
rect 569125 40160 569130 40216
rect 569186 40160 569234 40216
rect 569125 40155 569234 40160
rect 569174 40000 569234 40155
rect 239896 39870 239956 39990
rect 239896 39810 241346 39870
rect 241286 39600 241346 39810
rect 241260 31680 246048 39600
rect 251300 31680 256100 39600
rect 569142 34830 573922 40000
rect 579121 34830 583901 40000
rect 622942 37008 627722 40000
rect 632921 37008 637701 40000
<< via3 >>
rect 239894 40146 239958 40210
rect 240727 40228 240797 40233
rect 240727 40168 240732 40228
rect 240732 40168 240792 40228
rect 240792 40168 240797 40228
rect 240727 40163 240797 40168
<< metal4 >>
rect 333400 1032757 333654 1037599
rect 348146 1032757 348400 1037599
rect 575600 1008881 575854 1008947
rect 590346 1008881 590600 1008947
rect 575600 1007929 575854 1008165
rect 590346 1007929 590600 1008165
rect 575600 1007147 575854 1007213
rect 590346 1007147 590600 1007213
rect 575600 1004947 575854 1005637
rect 590346 1004947 590600 1005637
rect 333400 1002767 333654 1003697
rect 348146 1002767 348400 1003697
rect 37293 926746 38223 927000
rect 679377 922346 680307 922600
rect 37293 912000 38223 912254
rect 679377 907600 680307 907854
rect 28653 842346 28719 842600
rect 29435 842346 29671 842600
rect 30387 842346 30453 842600
rect 31963 842346 32653 842600
rect 680587 833207 681277 833399
rect 28653 827600 28719 827854
rect 29435 827600 29671 827854
rect 30387 827600 30453 827854
rect 31963 827600 32653 827854
rect 680587 818400 681277 818592
rect 36323 497807 37013 497999
rect 36323 483000 37013 483192
rect 685917 474546 686847 474800
rect 685917 459800 686847 460054
rect 30753 455546 31683 455800
rect 30753 440800 31683 441054
rect 21000 124946 25992 125200
rect 35113 124946 36043 125200
rect 21000 110200 25992 110454
rect 35113 110200 36043 110454
rect 37293 82746 38223 83000
rect 37293 68000 38223 68254
rect 239730 40338 240114 40378
rect 239730 40018 239766 40338
rect 240086 40018 240114 40338
rect 239730 39990 240114 40018
rect 622800 36323 622992 37013
rect 637607 36323 637799 37013
rect 78800 31963 79054 32653
rect 93546 31963 93800 32653
rect 241200 30753 241454 31683
rect 255946 30753 256200 31683
rect 78800 30387 79054 30453
rect 93546 30387 93800 30453
rect 78800 29435 79054 29671
rect 93546 29435 93800 29671
rect 78800 28653 79054 28719
rect 93546 28653 93800 28719
<< via4 >>
rect 239766 40210 240086 40338
rect 239766 40146 239894 40210
rect 239894 40146 239958 40210
rect 239958 40146 240086 40210
rect 239766 40018 240086 40146
rect 240602 40233 240922 40358
rect 240602 40163 240727 40233
rect 240727 40163 240797 40233
rect 240797 40163 240922 40233
rect 240602 40038 240922 40163
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 575600 1007147 575854 1008947
rect 590346 1007147 590600 1008947
rect 575600 1004968 575854 1005616
rect 590346 1004968 590600 1005616
rect 333400 1002787 333654 1003677
rect 348146 1002787 348400 1003677
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 37313 926746 38203 927000
rect 6167 914054 19620 924934
rect 679397 922346 680287 922600
rect 37313 912000 38203 912254
rect 697980 909666 711433 920546
rect 679397 907600 680287 907854
rect 698512 863640 711002 876160
rect 28653 842346 30453 842600
rect 31983 842346 32631 842600
rect 6811 829010 18976 841178
rect 680607 833207 681257 833399
rect 28653 827600 30453 827854
rect 31983 827600 32631 827854
rect 698624 819822 710789 831990
rect 680607 818400 681257 818592
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 36343 497807 36993 497999
rect 6811 484410 18976 496578
rect 36343 483000 36993 483192
rect 685937 474546 686827 474800
rect 697980 461866 711433 472746
rect 685937 459800 686827 460054
rect 30773 455546 31663 455800
rect 6167 442854 19620 453734
rect 30773 440800 31663 441054
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 21003 124946 25993 125200
rect 35133 124946 36023 125200
rect 6811 111610 18976 123778
rect 21003 110200 25993 110454
rect 35133 110200 36023 110454
rect 698512 101240 711002 113760
rect 37313 82746 38203 83000
rect 6167 70054 19620 80934
rect 37313 68000 38203 68254
rect 240578 40380 240946 40382
rect 240206 40378 240946 40380
rect 239730 40358 240946 40378
rect 239730 40338 240602 40358
rect 239730 40018 239766 40338
rect 240086 40038 240602 40338
rect 240922 40038 240946 40358
rect 240086 40018 240946 40038
rect 239730 40014 240946 40018
rect 239730 40006 240866 40014
rect 239730 39990 240114 40006
rect 622800 36343 622992 36993
rect 637607 36343 637799 36993
rect 78800 31983 79054 32631
rect 93546 31983 93800 32631
rect 241200 30773 241454 31663
rect 255946 30773 256200 31663
rect 78800 28653 79054 30453
rect 93546 28653 93800 30453
rect 80222 6811 92390 18976
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use sky130_ef_io__com_bus_slice_20um  FILLER_177 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1619552202
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1619552202
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3
timestamp 1619552202
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_178 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_181
timestamp 1619552202
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_179 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_188
timestamp 1619552202
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1619552202
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1619552202
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1619552202
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_189
timestamp 1619552202
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1619552202
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_192
timestamp 1619552202
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_190
timestamp 1619552202
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_194
timestamp 1619552202
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_195
timestamp 1619552202
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_196
timestamp 1619552202
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1619552202
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_198
timestamp 1619552202
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1619552202
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1619552202
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1619552202
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1619552202
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1619552202
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1619552202
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_205
timestamp 1619552202
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_206
timestamp 1619552202
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1619552202
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_209
timestamp 1619552202
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_207
timestamp 1619552202
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 147600 0 -1 40000
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_211
timestamp 1619552202
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1619552202
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_212
timestamp 1619552202
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_214
timestamp 1619552202
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_215
timestamp 1619552202
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_213
timestamp 1619552202
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1619552202
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1619552202
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1619552202
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_222
timestamp 1619552202
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1619552202
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1619552202
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_223
timestamp 1619552202
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1619552202
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_226
timestamp 1619552202
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_224
timestamp 1619552202
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 202400 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_228
timestamp 1619552202
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1619552202
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_229
timestamp 1619552202
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_231
timestamp 1619552202
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_232
timestamp 1619552202
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_230
timestamp 1619552202
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1619552202
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1619552202
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1619552202
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1619552202
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1619552202
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_239
timestamp 1619552202
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_240
timestamp 1619552202
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1619552202
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_243
timestamp 1619552202
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_241
timestamp 1619552202
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 256200 0 -1 39593
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_245
timestamp 1619552202
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1619552202
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1619552202
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_246
timestamp 1619552202
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_248
timestamp 1619552202
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_249
timestamp 1619552202
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_247
timestamp 1619552202
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1619552202
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1619552202
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1619552202
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1619552202
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_256
timestamp 1619552202
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_257
timestamp 1619552202
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1619552202
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_260
timestamp 1619552202
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_258
timestamp 1619552202
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1619552202
transform -1 0 311000 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_262
timestamp 1619552202
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_263
timestamp 1619552202
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1619552202
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1619552202
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_266
timestamp 1619552202
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_264
timestamp 1619552202
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1619552202
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1619552202
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1619552202
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1619552202
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_273
timestamp 1619552202
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1619552202
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_274
timestamp 1619552202
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1619552202
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_277
timestamp 1619552202
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_275
timestamp 1619552202
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1619552202
transform -1 0 365800 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_279
timestamp 1619552202
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1619552202
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1619552202
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_280
timestamp 1619552202
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_282
timestamp 1619552202
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_283
timestamp 1619552202
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_281
timestamp 1619552202
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1619552202
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1619552202
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1619552202
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1619552202
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_290
timestamp 1619552202
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_291
timestamp 1619552202
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1619552202
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_294
timestamp 1619552202
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_292
timestamp 1619552202
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1619552202
transform -1 0 420600 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_296
timestamp 1619552202
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1619552202
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1619552202
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1619552202
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_297
timestamp 1619552202
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_299
timestamp 1619552202
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_300
timestamp 1619552202
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_298
timestamp 1619552202
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_307
timestamp 1619552202
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1619552202
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1619552202
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1619552202
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_308
timestamp 1619552202
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1619552202
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_311
timestamp 1619552202
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_309
timestamp 1619552202
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1619552202
transform -1 0 475400 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_313
timestamp 1619552202
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_314
timestamp 1619552202
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1619552202
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1619552202
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_317
timestamp 1619552202
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_315
timestamp 1619552202
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1619552202
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1619552202
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1619552202
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1619552202
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1619552202
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_324
timestamp 1619552202
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_325
timestamp 1619552202
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1619552202
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_328
timestamp 1619552202
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_326
timestamp 1619552202
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1619552202
transform -1 0 530200 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_330
timestamp 1619552202
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1619552202
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_331
timestamp 1619552202
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1619552202
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_334
timestamp 1619552202
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_332
timestamp 1619552202
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1619552202
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1619552202
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_341
timestamp 1619552202
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1619552202
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1619552202
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1619552202
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_342
timestamp 1619552202
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1619552202
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_345
timestamp 1619552202
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_343
timestamp 1619552202
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_347
timestamp 1619552202
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_348
timestamp 1619552202
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_349
timestamp 1619552202
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1619552202
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1619552202
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1619552202
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1619552202
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_350
timestamp 1619552202
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_351
timestamp 1619552202
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_358
timestamp 1619552202
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1619552202
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1619552202
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_359
timestamp 1619552202
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1619552202
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_362
timestamp 1619552202
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_360
timestamp 1619552202
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_364
timestamp 1619552202
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_365
timestamp 1619552202
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_367
timestamp 1619552202
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_366
timestamp 1619552202
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1619552202
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_368
timestamp 1619552202
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1619552202
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1619552202
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1619552202
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1619552202
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1619552202
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1619552202
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_376
timestamp 1619552202
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1619552202
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1619552202
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_1um  FILLER_378
timestamp 1619552202
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_379
timestamp 1619552202
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_380
timestamp 1619552202
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_377
timestamp 1619552202
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1619552202
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_383
timestamp 1619552202
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1619552202
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1619552202
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1619552202
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_387
timestamp 1619552202
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_389
timestamp 1619552202
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_388
timestamp 1619552202
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform 0 -1 39593 1 0 68000
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1619552202
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1619552202
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1619552202
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1619552202
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1619552202
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1619552202
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1619552202
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_619
timestamp 1619552202
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1619552198
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1619552198
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1619552202
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1619552202
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1619552202
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1619552202
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1619552202
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1619552202
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1619552202
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1619552202
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1619552202
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_397
timestamp 1619552202
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_399
timestamp 1619552202
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_398
timestamp 1619552202
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1619552202
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1619552202
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1619552202
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1619552202
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1619552202
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1619552202
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1619552202
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_629
timestamp 1619552202
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1619552202
transform 0 1 675407 -1 0 116000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1619552202
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1619552202
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1619552202
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1619552202
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1619552202
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_407
timestamp 1619552202
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1619552202
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_409
timestamp 1619552202
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_408
timestamp 1619552202
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_2
timestamp 1619552198
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1619552198
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1619552202
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1619552202
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1619552202
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1619552202
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1619552202
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1619552202
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1619552202
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1619552202
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1619552202
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_639
timestamp 1619552202
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_638
timestamp 1619552202
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1619552202
transform 0 1 675407 -1 0 161200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1619552202
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_417
timestamp 1619552202
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_418
timestamp 1619552202
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_420
timestamp 1619552202
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_419
timestamp 1619552202
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[18\]
timestamp 1619552202
transform 0 -1 42193 1 0 181600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1619552202
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1619552202
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1619552202
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1619552202
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1619552202
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1619552202
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1619552202
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1619552202
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1619552202
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1619552202
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1619552202
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_648
timestamp 1619552202
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1619552202
transform 0 1 675407 -1 0 206200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1619552202
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1619552202
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_428
timestamp 1619552202
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_430
timestamp 1619552202
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_429
timestamp 1619552202
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[17\]
timestamp 1619552202
transform 0 -1 42193 1 0 224800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1619552202
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1619552202
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1619552202
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1619552202
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1619552202
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1619552202
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1619552202
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1619552202
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1619552202
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_660
timestamp 1619552202
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_658
timestamp 1619552202
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_657
timestamp 1619552202
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1619552202
transform 0 1 675407 -1 0 251400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1619552202
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1619552202
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1619552202
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1619552202
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1619552202
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_438
timestamp 1619552202
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_440
timestamp 1619552202
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_439
timestamp 1619552202
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[16\]
timestamp 1619552202
transform 0 -1 42193 1 0 268000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1619552202
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1619552202
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1619552202
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1619552202
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1619552202
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1619552202
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_667
timestamp 1619552202
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1619552202
transform 0 1 675407 -1 0 296400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1619552202
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1619552202
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1619552202
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_448
timestamp 1619552202
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_450
timestamp 1619552202
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_449
timestamp 1619552202
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[15\]
timestamp 1619552202
transform 0 -1 42193 1 0 311200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1619552202
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1619552202
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1619552202
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_669
timestamp 1619552202
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_670
timestamp 1619552202
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1619552202
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1619552202
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1619552202
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1619552202
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1619552202
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_676
timestamp 1619552202
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1619552202
transform 0 1 675407 -1 0 341400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1619552202
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1619552202
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1619552202
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_458
timestamp 1619552202
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_459
timestamp 1619552202
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_460
timestamp 1619552202
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[14\]
timestamp 1619552202
transform 0 -1 42193 1 0 354400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1619552202
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1619552202
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1619552202
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1619552202
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1619552202
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1619552202
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1619552202
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1619552202
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1619552202
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1619552202
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_685
timestamp 1619552202
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_686
timestamp 1619552202
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1619552202
transform 0 1 675407 -1 0 386600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1619552202
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1619552202
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1619552202
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_468
timestamp 1619552202
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_470
timestamp 1619552202
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_469
timestamp 1619552202
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[13\]
timestamp 1619552202
transform 0 -1 42193 1 0 397600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1619552202
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1619552202
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1619552202
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1619552202
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1619552202
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1619552202
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1619552202
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1619552202
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1619552202
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1619552202
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_695
timestamp 1619552202
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1619552202
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1619552202
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1619552202
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1619552202
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_478
timestamp 1619552202
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1619552202
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_480
timestamp 1619552202
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_479
timestamp 1619552202
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__vssd_lvc_clamped2_pad  user2_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform 0 -1 39593 1 0 440800
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1619552202
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1619552202
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_697
timestamp 1619552202
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1619552202
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1619552202
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1619552202
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1619552202
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1619552202
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1619552202
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_705
timestamp 1619552202
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_704
timestamp 1619552202
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__vssd_lvc_clamped2_pad  user1_vssd_lvclmap_pad
timestamp 1619552202
transform 0 1 678007 -1 0 474800
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1619552202
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1619552202
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1619552202
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_488
timestamp 1619552202
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_490
timestamp 1619552202
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_489
timestamp 1619552202
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1619552202
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_492
timestamp 1619552202
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1619552202
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1619552202
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1619552202
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_708
timestamp 1619552202
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1619552202
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1619552202
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1619552202
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1619552202
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1619552202
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_714
timestamp 1619552202
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1619552202
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1619552202
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1619552202
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1619552202
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_502
timestamp 1619552202
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_503
timestamp 1619552202
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_498
timestamp 1619552202
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_500
timestamp 1619552202
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_499
timestamp 1619552202
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1619552202
transform 0 -1 42193 1 0 525200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1619552202
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1619552202
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1619552202
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1619552202
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1619552202
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1619552202
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1619552202
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_723
timestamp 1619552202
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1619552202
transform 0 1 675407 -1 0 563800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1619552202
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1619552202
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1619552202
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1619552202
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_508
timestamp 1619552202
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_510
timestamp 1619552202
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_509
timestamp 1619552202
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1619552202
transform 0 -1 42193 1 0 568400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1619552202
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_513
timestamp 1619552202
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1619552202
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1619552202
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1619552202
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1619552202
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1619552202
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1619552202
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1619552202
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_514
timestamp 1619552202
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1619552202
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1619552202
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1619552202
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_518
timestamp 1619552202
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_520
timestamp 1619552202
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_519
timestamp 1619552202
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1619552202
transform 0 -1 42193 1 0 611600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1619552202
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1619552202
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1619552202
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1619552202
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1619552202
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1619552202
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1619552202
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1619552202
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_733
timestamp 1619552202
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_732
timestamp 1619552202
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1619552202
transform 0 1 675407 -1 0 609000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_524
timestamp 1619552202
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1619552202
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1619552202
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1619552202
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_528
timestamp 1619552202
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_530
timestamp 1619552202
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_529
timestamp 1619552202
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1619552202
transform 0 -1 42193 1 0 654800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1619552202
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1619552202
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1619552202
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1619552202
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1619552202
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1619552202
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1619552202
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1619552202
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1619552202
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_742
timestamp 1619552202
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1619552202
transform 0 1 675407 -1 0 654000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1619552202
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1619552202
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1619552202
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1619552202
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1619552202
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_538
timestamp 1619552202
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_540
timestamp 1619552202
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_539
timestamp 1619552202
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1619552202
transform 0 -1 42193 1 0 698000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1619552202
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1619552202
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1619552202
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1619552202
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1619552202
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1619552202
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_752
timestamp 1619552202
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_751
timestamp 1619552202
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1619552202
transform 0 1 675407 -1 0 699200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1619552202
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1619552202
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1619552202
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1619552202
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1619552202
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_548
timestamp 1619552202
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_550
timestamp 1619552202
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_549
timestamp 1619552202
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1619552202
transform 0 -1 42193 1 0 741200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1619552202
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1619552202
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1619552202
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1619552202
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_764
timestamp 1619552202
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1619552202
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1619552202
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_761
timestamp 1619552202
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1619552202
transform 0 1 675407 -1 0 744200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1619552202
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1619552202
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1619552202
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1619552202
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1619552202
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_558
timestamp 1619552202
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_560
timestamp 1619552202
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_559
timestamp 1619552202
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1619552202
transform 0 -1 42193 1 0 784400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1619552202
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1619552202
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1619552202
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1619552202
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1619552202
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1619552202
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1619552202
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1619552202
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_770
timestamp 1619552202
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1619552202
transform 0 1 675407 -1 0 789200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1619552202
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1619552202
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1619552202
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1619552202
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1619552202
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_568
timestamp 1619552202
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_570
timestamp 1619552202
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_569
timestamp 1619552202
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1619552202
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1619552202
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1619552202
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1619552202
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_778
timestamp 1619552202
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1619552202
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1619552202
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1619552202
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_780
timestamp 1619552202
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_779
timestamp 1619552202
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1619552202
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1619552202
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1619552202
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1619552202
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1619552202
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1619552202
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_578
timestamp 1619552202
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_580
timestamp 1619552202
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_579
timestamp 1619552202
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1619552202
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1619552202
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1619552202
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1619552202
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1619552202
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_788
timestamp 1619552202
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_791
timestamp 1619552202
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_792
timestamp 1619552202
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_789
timestamp 1619552202
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1619552202
transform 0 1 675407 -1 0 878400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1619552202
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1619552202
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1619552202
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1619552202
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1619552202
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_588
timestamp 1619552202
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_590
timestamp 1619552202
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_589
timestamp 1619552202
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__vccd_lvc_clamped2_pad  user2_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform 0 -1 39593 1 0 912000
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_592
timestamp 1619552202
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_793
timestamp 1619552202
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1619552202
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1619552202
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1619552202
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1619552202
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_799
timestamp 1619552202
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_798
timestamp 1619552202
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__vccd_lvc_clamped2_pad  user1_vccd_lvclamp_pad
timestamp 1619552202
transform 0 1 678007 -1 0 922600
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_801
timestamp 1619552202
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_802
timestamp 1619552202
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1619552202
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1619552202
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1619552202
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1619552202
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[5\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform 0 -1 40000 1 0 955200
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1619552202
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_598
timestamp 1619552202
transform 0 -1 39593 1 0 951000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_600
timestamp 1619552202
transform 0 -1 39593 1 0 954000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_10
timestamp 1619552202
transform 0 -1 39593 1 0 954200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_599
timestamp 1619552202
transform 0 -1 39593 1 0 953000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_602
timestamp 1619552202
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[0\]
timestamp 1619552202
transform 0 1 677600 -1 0 966600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_803
timestamp 1619552202
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1619552202
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1619552202
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1619552202
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1619552202
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_810
timestamp 1619552202
transform 0 1 678007 -1 0 971600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_11
timestamp 1619552202
transform 0 1 678007 -1 0 967600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_808
timestamp 1619552202
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1619552202
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1619552202
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1619552202
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1619552202
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1619552202
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_608
timestamp 1619552202
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_610
timestamp 1619552202
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_611
timestamp 1619552202
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_609
timestamp 1619552202
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1619552202
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1619552202
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1619552202
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1619552202
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1619552202
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1619552202
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1619552202
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1619552202
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1619552202
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13
timestamp 1619552202
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1619552202
transform 1 0 75800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1619552202
transform 1 0 76000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_9
timestamp 1619552202
transform 1 0 76200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_14
timestamp 1619552202
transform 1 0 74800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[4\]
timestamp 1619552202
transform 1 0 77200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1619552202
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1619552202
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1619552202
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1619552202
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1619552202
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1619552202
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1619552202
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1619552202
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_26
timestamp 1619552202
transform 1 0 124200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_27
timestamp 1619552202
transform 1 0 126200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1619552202
transform 1 0 127200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1619552202
transform 1 0 127400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_8
timestamp 1619552202
transform 1 0 127600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[3\]
timestamp 1619552202
transform 1 0 128600 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1619552202
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1619552202
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1619552202
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1619552202
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1619552202
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1619552202
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1619552202
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1619552202
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_39
timestamp 1619552202
transform 1 0 175600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1619552202
transform 1 0 178600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1619552202
transform 1 0 178800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_7
timestamp 1619552202
transform 1 0 179000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_40
timestamp 1619552202
transform 1 0 177600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[2\]
timestamp 1619552202
transform 1 0 180000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1619552202
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1619552202
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1619552202
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1619552202
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1619552202
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1619552202
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1619552202
transform 1 0 219000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1619552202
transform 1 0 223000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_52
timestamp 1619552202
transform 1 0 227000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1619552202
transform 1 0 230000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1619552202
transform 1 0 230200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_6
timestamp 1619552202
transform 1 0 230400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1619552202
transform 1 0 229000 0 1 998007
box 0 0 1000 39593
use sky130_fd_io__top_power_hvc_wpadv2  user2_analog_pad\[1\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1619552202
transform 1 0 231400 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1619552202
transform 1 0 246400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1619552202
transform 1 0 250400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1619552202
transform 1 0 254400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1619552202
transform 1 0 258400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1619552202
transform 1 0 262400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1619552202
transform 1 0 266400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1619552202
transform 1 0 270400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1619552202
transform 1 0 274400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1619552202
transform 1 0 278400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1619552202
transform 1 0 281400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1619552202
transform 1 0 281600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1619552202
transform 1 0 281800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_5
timestamp 1619552202
transform 1 0 282000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1619552202
transform 1 0 280400 0 1 998007
box 0 0 1000 39593
use sky130_fd_io__top_power_hvc_wpadv2  user2_analog_pad\[0\]
timestamp 1619552202
transform 1 0 283000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1619552202
transform 1 0 298000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1619552202
transform 1 0 302000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1619552202
transform 1 0 306000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1619552202
transform 1 0 310000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1619552202
transform 1 0 314000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1619552202
transform 1 0 318000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1619552202
transform 1 0 322000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1619552202
transform 1 0 326000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_79
timestamp 1619552202
transform 1 0 330000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1619552202
transform 1 0 333000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1619552202
transform 1 0 333200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_80
timestamp 1619552202
transform 1 0 332000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\]
timestamp 1619552202
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_0
timestamp 1619552202
transform 1 0 348400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1619552202
transform 1 0 352400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_0
timestamp 1619552198
transform 1 0 351400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1619552198
transform 1 0 350400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1619552202
transform 1 0 356400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1619552202
transform 1 0 360400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1619552202
transform 1 0 364400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1619552202
transform 1 0 368400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1619552202
transform 1 0 372400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1619552202
transform 1 0 376400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_92
timestamp 1619552202
transform 1 0 380400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_94
timestamp 1619552202
transform 1 0 383400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1619552202
transform 1 0 383600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_4
timestamp 1619552202
transform 1 0 383800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_93
timestamp 1619552202
transform 1 0 382400 0 1 998007
box 0 0 1000 39593
use sky130_fd_io__top_power_hvc_wpadv2  user1_analog_pad\[4\]
timestamp 1619552202
transform 1 0 384800 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_97
timestamp 1619552202
transform 1 0 399800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1619552202
transform 1 0 403800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1619552202
transform 1 0 407800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1619552202
transform 1 0 411800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1619552202
transform 1 0 415800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1619552202
transform 1 0 419800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1619552202
transform 1 0 423800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1619552202
transform 1 0 427800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_0
timestamp 1619552202
transform 1 0 431800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1619552202
transform 1 0 437200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_0
timestamp 1619552202
transform 1 0 436800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_1
timestamp 1619552202
transform 1 0 437000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_0
timestamp 1619552202
transform 1 0 435800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1619552202
transform 1 0 441200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1619552202
transform 1 0 445200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1619552202
transform 1 0 449200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1619552202
transform 1 0 453200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1619552202
transform 1 0 457200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1619552202
transform 1 0 461200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1619552202
transform 1 0 465200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_119
timestamp 1619552202
transform 1 0 469200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_121
timestamp 1619552202
transform 1 0 472200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_122
timestamp 1619552202
transform 1 0 472400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_123
timestamp 1619552202
transform 1 0 472600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_3
timestamp 1619552202
transform 1 0 472800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_120
timestamp 1619552202
transform 1 0 471200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[3\]
timestamp 1619552202
transform 1 0 473800 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1619552202
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_126
timestamp 1619552202
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_127
timestamp 1619552202
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1619552202
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1619552202
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1619552202
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1619552202
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1619552202
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_133
timestamp 1619552202
transform 1 0 520800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_135
timestamp 1619552202
transform 1 0 523800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_136
timestamp 1619552202
transform 1 0 524000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_2
timestamp 1619552202
transform 1 0 524200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_134
timestamp 1619552202
transform 1 0 522800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[2\]
timestamp 1619552202
transform 1 0 525200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1619552202
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_139
timestamp 1619552202
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1619552202
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1619552202
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1619552202
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_143
timestamp 1619552202
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1619552202
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1619552202
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_146
timestamp 1619552202
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_148
timestamp 1619552202
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_149
timestamp 1619552202
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_147
timestamp 1619552202
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1619552202
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1619552202
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_152
timestamp 1619552202
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_153
timestamp 1619552202
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_154
timestamp 1619552202
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_155
timestamp 1619552202
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_156
timestamp 1619552202
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1619552202
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1619552202
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_159
timestamp 1619552202
transform 1 0 622600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_161
timestamp 1619552202
transform 1 0 625600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_162
timestamp 1619552202
transform 1 0 625800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_1
timestamp 1619552202
transform 1 0 626000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_160
timestamp 1619552202
transform 1 0 624600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[1\]
timestamp 1619552202
transform 1 0 627000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1619552202
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1619552202
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_166
timestamp 1619552202
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_167
timestamp 1619552202
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_168
timestamp 1619552202
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_169
timestamp 1619552202
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_170
timestamp 1619552202
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_171
timestamp 1619552202
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_172
timestamp 1619552202
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_811
timestamp 1619552202
transform 0 1 678007 -1 0 975600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_812
timestamp 1619552202
transform 0 1 678007 -1 0 979600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_813
timestamp 1619552202
transform 0 1 678007 -1 0 983600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_814
timestamp 1619552202
transform 0 1 678007 -1 0 987600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_815
timestamp 1619552202
transform 0 1 678007 -1 0 991600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_816
timestamp 1619552202
transform 0 1 678007 -1 0 995600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_818
timestamp 1619552202
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_817
timestamp 1619552202
transform 0 1 678007 -1 0 996600
box 0 0 1000 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1619552202
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_1um  FILLER_174
timestamp 1619552202
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_175
timestamp 1619552202
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_176
timestamp 1619552202
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_173
timestamp 1619552202
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 1 nsew signal tristate
rlabel metal2 s 194043 41713 194099 42193 6 por
port 2 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 3 nsew signal tristate
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 4 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 5 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 6 nsew signal input
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 7 nsew signal tristate
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 8 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 9 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 10 nsew signal input
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 11 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 12 nsew signal tristate
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 13 nsew signal input
rlabel metal2 s 412243 41713 412299 42193 6 flash_io0_ieb_core
port 14 nsew signal input
rlabel metal2 s 419695 41713 419751 42193 6 flash_io0_oeb_core
port 15 nsew signal input
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 16 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 17 nsew signal tristate
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 18 nsew signal input
rlabel metal2 s 467043 41713 467099 42193 6 flash_io1_ieb_core
port 19 nsew signal input
rlabel metal2 s 474495 41713 474551 42193 6 flash_io1_oeb_core
port 20 nsew signal input
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 21 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 22 nsew signal tristate
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 23 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 24 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 25 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 26 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 27 nsew signal input
rlabel metal4 s 37293 68000 38223 68254 6 vccd
port 28 nsew signal bidirectional
rlabel metal4 s 37293 82746 38223 83000 6 vccd
port 29 nsew signal bidirectional
rlabel metal5 s 37313 68000 38203 68254 6 vccd
port 30 nsew signal bidirectional
rlabel metal5 s 37313 82746 38203 83000 6 vccd
port 31 nsew signal bidirectional
rlabel metal3 s 38220 68100 39600 72900 6 vccd
port 32 nsew signal bidirectional
rlabel metal3 s 38220 78151 39600 82939 6 vccd
port 33 nsew signal bidirectional
rlabel metal4 s 637607 36323 637799 37013 6 vdda
port 35 nsew signal bidirectional
rlabel metal4 s 622800 36323 622992 37013 6 vdda
port 36 nsew signal bidirectional
rlabel metal5 s 637607 36343 637799 36993 6 vdda
port 37 nsew signal bidirectional
rlabel metal5 s 622800 36343 622992 36993 6 vdda
port 38 nsew signal bidirectional
rlabel metal3 s 632921 37008 637701 40000 6 vdda
port 39 nsew signal bidirectional
rlabel metal3 s 622942 37008 627722 40000 6 vdda
port 40 nsew signal bidirectional
rlabel metal4 s 21000 110200 25992 110454 6 vddio
port 42 nsew signal bidirectional
rlabel metal4 s 35113 110200 36043 110454 6 vddio
port 43 nsew signal bidirectional
rlabel metal4 s 21000 124946 25992 125200 6 vddio
port 44 nsew signal bidirectional
rlabel metal4 s 35113 124946 36043 125200 6 vddio
port 45 nsew signal bidirectional
rlabel metal5 s 35133 110200 36023 110454 6 vddio
port 46 nsew signal bidirectional
rlabel metal5 s 21003 110200 25993 110454 6 vddio
port 47 nsew signal bidirectional
rlabel metal5 s 35133 124946 36023 125200 6 vddio
port 48 nsew signal bidirectional
rlabel metal5 s 21003 124946 25993 125200 6 vddio
port 49 nsew signal bidirectional
rlabel metal3 s 36040 110299 40000 115079 6 vddio
port 50 nsew signal bidirectional
rlabel metal3 s 36040 120278 40000 125058 6 vddio
port 51 nsew signal bidirectional
rlabel metal4 s 93546 31963 93800 32653 6 vssa
port 53 nsew signal bidirectional
rlabel metal4 s 93546 28653 93800 28719 6 vssa
port 54 nsew signal bidirectional
rlabel metal4 s 93546 29435 93800 29671 6 vssa
port 55 nsew signal bidirectional
rlabel metal4 s 93546 30387 93800 30453 6 vssa
port 56 nsew signal bidirectional
rlabel metal4 s 78800 31963 79054 32653 6 vssa
port 57 nsew signal bidirectional
rlabel metal4 s 78800 30387 79054 30453 6 vssa
port 58 nsew signal bidirectional
rlabel metal4 s 78800 28653 79054 28719 6 vssa
port 59 nsew signal bidirectional
rlabel metal4 s 78800 29435 79054 29671 6 vssa
port 60 nsew signal bidirectional
rlabel metal5 s 93546 31983 93800 32631 6 vssa
port 61 nsew signal bidirectional
rlabel metal5 s 93546 28653 93800 30453 6 vssa
port 62 nsew signal bidirectional
rlabel metal5 s 78800 31983 79054 32631 6 vssa
port 63 nsew signal bidirectional
rlabel metal5 s 78800 28653 79054 30453 6 vssa
port 64 nsew signal bidirectional
rlabel metal3 s 78942 32648 83722 40000 6 vssa
port 65 nsew signal bidirectional
rlabel metal3 s 88921 33497 93701 39999 6 vssa
port 66 nsew signal bidirectional
rlabel metal4 s 255946 30753 256200 31683 6 vssd
port 68 nsew signal bidirectional
rlabel metal4 s 241200 30753 241454 31683 6 vssd
port 69 nsew signal bidirectional
rlabel metal5 s 255946 30773 256200 31663 6 vssd
port 70 nsew signal bidirectional
rlabel metal5 s 241200 30773 241454 31663 6 vssd
port 71 nsew signal bidirectional
rlabel metal3 s 251300 31680 256100 39600 6 vssd
port 72 nsew signal bidirectional
rlabel metal3 s 241260 31680 246048 39600 6 vssd
port 73 nsew signal bidirectional
rlabel metal4 s 333400 1002767 333654 1003697 6 vssio
port 75 nsew signal bidirectional
rlabel metal4 s 333400 1032757 333654 1037599 6 vssio
port 76 nsew signal bidirectional
rlabel metal4 s 348146 1032757 348400 1037599 6 vssio
port 77 nsew signal bidirectional
rlabel metal4 s 348146 1002767 348400 1003697 6 vssio
port 78 nsew signal bidirectional
rlabel metal5 s 333400 1002787 333654 1003677 6 vssio
port 79 nsew signal bidirectional
rlabel metal5 s 348146 1002787 348400 1003677 6 vssio
port 80 nsew signal bidirectional
rlabel metal3 s 343478 997600 348258 1002770 6 vssio
port 81 nsew signal bidirectional
rlabel metal3 s 333499 997600 338279 1002770 6 vssio
port 82 nsew signal bidirectional
rlabel metal4 s 348250 1032757 348400 1037599 6 vssio
port 83 nsew signal bidirectional
rlabel metal4 s 333526 1035920 333528 1035922 6 vssio
port 84 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 86 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 87 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 88 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 89 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 90 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 91 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 92 nsew signal input
rlabel metal2 s 675407 108931 675887 108987 6 mprj_io_enh[0]
port 93 nsew signal input
rlabel metal2 s 675407 109575 675887 109631 6 mprj_io_hldh_n[0]
port 94 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 95 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 96 nsew signal input
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 97 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 98 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 99 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 100 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 101 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 102 nsew signal tristate
rlabel metal2 s 675407 686611 675887 686667 6 mprj_analog_io[3]
port 103 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 104 nsew signal bidirectional
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 105 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 106 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 107 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 108 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 109 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 110 nsew signal input
rlabel metal2 s 675407 692131 675887 692187 6 mprj_io_enh[10]
port 111 nsew signal input
rlabel metal2 s 675407 692775 675887 692831 6 mprj_io_hldh_n[10]
port 112 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 113 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 114 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 115 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 116 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 117 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 118 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 119 nsew signal input
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 120 nsew signal tristate
rlabel metal2 s 675407 731611 675887 731667 6 mprj_analog_io[4]
port 121 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 122 nsew signal bidirectional
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 123 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 124 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 125 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 126 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 127 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 128 nsew signal input
rlabel metal2 s 675407 737131 675887 737187 6 mprj_io_enh[11]
port 129 nsew signal input
rlabel metal2 s 675407 737775 675887 737831 6 mprj_io_hldh_n[11]
port 130 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 131 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 132 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 133 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 134 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 135 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 136 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 137 nsew signal input
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 138 nsew signal tristate
rlabel metal2 s 675407 776611 675887 776667 6 mprj_analog_io[5]
port 139 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 140 nsew signal bidirectional
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 141 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 142 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 143 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 144 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 145 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 146 nsew signal input
rlabel metal2 s 675407 782131 675887 782187 6 mprj_io_enh[12]
port 147 nsew signal input
rlabel metal2 s 675407 782775 675887 782831 6 mprj_io_hldh_n[12]
port 148 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 149 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 150 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 151 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 152 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 153 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 154 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 155 nsew signal input
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 156 nsew signal tristate
rlabel metal2 s 675407 865811 675887 865867 6 mprj_analog_io[6]
port 157 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 158 nsew signal bidirectional
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 159 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 160 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 161 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 162 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 163 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 164 nsew signal input
rlabel metal2 s 675407 871331 675887 871387 6 mprj_io_enh[13]
port 165 nsew signal input
rlabel metal2 s 675407 871975 675887 872031 6 mprj_io_hldh_n[13]
port 166 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 167 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 168 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 169 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 170 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 171 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 172 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 173 nsew signal input
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 174 nsew signal tristate
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 176 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 194 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 212 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 230 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 247 nsew signal bidirectional
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 248 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 249 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 250 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 251 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 252 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 253 nsew signal input
rlabel metal2 s 675407 154131 675887 154187 6 mprj_io_enh[1]
port 254 nsew signal input
rlabel metal2 s 675407 154775 675887 154831 6 mprj_io_hldh_n[1]
port 255 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 256 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 257 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 258 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 259 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 260 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 261 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 262 nsew signal input
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 263 nsew signal tristate
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 264 nsew signal bidirectional
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 265 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 266 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 267 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 268 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 269 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 270 nsew signal input
rlabel metal2 s 675407 199131 675887 199187 6 mprj_io_enh[2]
port 271 nsew signal input
rlabel metal2 s 675407 199775 675887 199831 6 mprj_io_hldh_n[2]
port 272 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 273 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 274 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 275 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 276 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 277 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 278 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 279 nsew signal input
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 280 nsew signal tristate
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 281 nsew signal bidirectional
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 282 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 283 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 284 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 285 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 286 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 287 nsew signal input
rlabel metal2 s 675407 244331 675887 244387 6 mprj_io_enh[3]
port 288 nsew signal input
rlabel metal2 s 675407 244975 675887 245031 6 mprj_io_hldh_n[3]
port 289 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 290 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 291 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 292 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 293 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 294 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 295 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 296 nsew signal input
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 297 nsew signal tristate
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 298 nsew signal bidirectional
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 299 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 300 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 301 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 302 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 303 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 304 nsew signal input
rlabel metal2 s 675407 289331 675887 289387 6 mprj_io_enh[4]
port 305 nsew signal input
rlabel metal2 s 675407 289975 675887 290031 6 mprj_io_hldh_n[4]
port 306 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 307 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 308 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 309 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 310 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 311 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 312 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 313 nsew signal input
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 314 nsew signal tristate
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 315 nsew signal bidirectional
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 316 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 317 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 318 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 319 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 320 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 321 nsew signal input
rlabel metal2 s 675407 334331 675887 334387 6 mprj_io_enh[5]
port 322 nsew signal input
rlabel metal2 s 675407 334975 675887 335031 6 mprj_io_hldh_n[5]
port 323 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 324 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 325 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 326 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 327 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 328 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 329 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 330 nsew signal input
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 331 nsew signal tristate
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 332 nsew signal bidirectional
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 333 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 334 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 335 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 336 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 337 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 338 nsew signal input
rlabel metal2 s 675407 379531 675887 379587 6 mprj_io_enh[6]
port 339 nsew signal input
rlabel metal2 s 675407 380175 675887 380231 6 mprj_io_hldh_n[6]
port 340 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 341 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 342 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 343 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 344 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 345 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 346 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 347 nsew signal input
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 348 nsew signal tristate
rlabel metal2 s 675407 551211 675887 551267 6 mprj_analog_io[0]
port 349 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 350 nsew signal bidirectional
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 351 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 352 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 353 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 354 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 355 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 356 nsew signal input
rlabel metal2 s 675407 556731 675887 556787 6 mprj_io_enh[7]
port 357 nsew signal input
rlabel metal2 s 675407 557375 675887 557431 6 mprj_io_hldh_n[7]
port 358 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 359 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 360 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 361 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 362 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 363 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 364 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 365 nsew signal input
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 366 nsew signal tristate
rlabel metal2 s 675407 596411 675887 596467 6 mprj_analog_io[1]
port 367 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 368 nsew signal bidirectional
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 369 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 370 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 371 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 372 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 373 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 374 nsew signal input
rlabel metal2 s 675407 601931 675887 601987 6 mprj_io_enh[8]
port 375 nsew signal input
rlabel metal2 s 675407 602575 675887 602631 6 mprj_io_hldh_n[8]
port 376 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 377 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 378 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 379 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 380 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 381 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 382 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 383 nsew signal input
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 384 nsew signal tristate
rlabel metal2 s 675407 641411 675887 641467 6 mprj_analog_io[2]
port 385 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 386 nsew signal bidirectional
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 387 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 388 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 389 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 390 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 391 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 392 nsew signal input
rlabel metal2 s 675407 646931 675887 646987 6 mprj_io_enh[9]
port 393 nsew signal input
rlabel metal2 s 675407 647575 675887 647631 6 mprj_io_hldh_n[9]
port 394 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 395 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 396 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 397 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 398 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 399 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 400 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 401 nsew signal input
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 402 nsew signal tristate
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 404 nsew signal bidirectional
rlabel metal2 s 41713 667333 42193 667389 6 mprj_analog_io[21]
port 421 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 422 nsew signal bidirectional
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[28]
port 423 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[28]
port 424 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[28]
port 425 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[84]
port 426 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[85]
port 427 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[86]
port 428 nsew signal input
rlabel metal2 s 41713 661813 42193 661869 6 mprj_io_enh[28]
port 429 nsew signal input
rlabel metal2 s 41713 661169 42193 661225 6 mprj_io_hldh_n[28]
port 430 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[28]
port 431 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[28]
port 432 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[28]
port 433 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[28]
port 434 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[28]
port 435 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[28]
port 436 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[28]
port 437 nsew signal input
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[28]
port 438 nsew signal tristate
rlabel metal2 s 41713 624133 42193 624189 6 mprj_analog_io[22]
port 439 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 440 nsew signal bidirectional
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[29]
port 441 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[29]
port 442 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[29]
port 443 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[87]
port 444 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[88]
port 445 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[89]
port 446 nsew signal input
rlabel metal2 s 41713 618613 42193 618669 6 mprj_io_enh[29]
port 447 nsew signal input
rlabel metal2 s 41713 617969 42193 618025 6 mprj_io_hldh_n[29]
port 448 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[29]
port 449 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[29]
port 450 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[29]
port 451 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[29]
port 452 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[29]
port 453 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[29]
port 454 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[29]
port 455 nsew signal input
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[29]
port 456 nsew signal tristate
rlabel metal2 s 41713 580933 42193 580989 6 mprj_analog_io[23]
port 457 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 458 nsew signal bidirectional
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[30]
port 459 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[30]
port 460 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[30]
port 461 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[90]
port 462 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[91]
port 463 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[92]
port 464 nsew signal input
rlabel metal2 s 41713 575413 42193 575469 6 mprj_io_enh[30]
port 465 nsew signal input
rlabel metal2 s 41713 574769 42193 574825 6 mprj_io_hldh_n[30]
port 466 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[30]
port 467 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[30]
port 468 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[30]
port 469 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[30]
port 470 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[30]
port 471 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[30]
port 472 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[30]
port 473 nsew signal input
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[30]
port 474 nsew signal tristate
rlabel metal2 s 41713 537733 42193 537789 6 mprj_analog_io[24]
port 475 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 476 nsew signal bidirectional
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[31]
port 477 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[31]
port 478 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[31]
port 479 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[93]
port 480 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[94]
port 481 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[95]
port 482 nsew signal input
rlabel metal2 s 41713 532213 42193 532269 6 mprj_io_enh[31]
port 483 nsew signal input
rlabel metal2 s 41713 531569 42193 531625 6 mprj_io_hldh_n[31]
port 484 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[31]
port 485 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[31]
port 486 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[31]
port 487 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[31]
port 488 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[31]
port 489 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[31]
port 490 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[31]
port 491 nsew signal input
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[31]
port 492 nsew signal tristate
rlabel metal2 s 41713 410133 42193 410189 6 mprj_analog_io[25]
port 493 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 494 nsew signal bidirectional
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[32]
port 495 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[32]
port 496 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[32]
port 497 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[96]
port 498 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[97]
port 499 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[98]
port 500 nsew signal input
rlabel metal2 s 41713 404613 42193 404669 6 mprj_io_enh[32]
port 501 nsew signal input
rlabel metal2 s 41713 403969 42193 404025 6 mprj_io_hldh_n[32]
port 502 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[32]
port 503 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[32]
port 504 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[32]
port 505 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[32]
port 506 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[32]
port 507 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[32]
port 508 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[32]
port 509 nsew signal input
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[32]
port 510 nsew signal tristate
rlabel metal2 s 41713 366933 42193 366989 6 mprj_analog_io[26]
port 511 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 512 nsew signal bidirectional
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[33]
port 513 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[33]
port 514 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[33]
port 515 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[100]
port 516 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[101]
port 517 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[99]
port 518 nsew signal input
rlabel metal2 s 41713 361413 42193 361469 6 mprj_io_enh[33]
port 519 nsew signal input
rlabel metal2 s 41713 360769 42193 360825 6 mprj_io_hldh_n[33]
port 520 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[33]
port 521 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[33]
port 522 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[33]
port 523 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[33]
port 524 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[33]
port 525 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[33]
port 526 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[33]
port 527 nsew signal input
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[33]
port 528 nsew signal tristate
rlabel metal2 s 41713 323733 42193 323789 6 mprj_analog_io[27]
port 529 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 530 nsew signal bidirectional
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[34]
port 531 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[34]
port 532 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[34]
port 533 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[102]
port 534 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[103]
port 535 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[104]
port 536 nsew signal input
rlabel metal2 s 41713 318213 42193 318269 6 mprj_io_enh[34]
port 537 nsew signal input
rlabel metal2 s 41713 317569 42193 317625 6 mprj_io_hldh_n[34]
port 538 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[34]
port 539 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[34]
port 540 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[34]
port 541 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[34]
port 542 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[34]
port 543 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[34]
port 544 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[34]
port 545 nsew signal input
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[34]
port 546 nsew signal tristate
rlabel metal2 s 41713 280533 42193 280589 6 mprj_analog_io[28]
port 547 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 548 nsew signal bidirectional
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[35]
port 549 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[35]
port 550 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[35]
port 551 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[105]
port 552 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[106]
port 553 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[107]
port 554 nsew signal input
rlabel metal2 s 41713 275013 42193 275069 6 mprj_io_enh[35]
port 555 nsew signal input
rlabel metal2 s 41713 274369 42193 274425 6 mprj_io_hldh_n[35]
port 556 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[35]
port 557 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[35]
port 558 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[35]
port 559 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[35]
port 560 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[35]
port 561 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[35]
port 562 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[35]
port 563 nsew signal input
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[35]
port 564 nsew signal tristate
rlabel metal2 s 41713 237333 42193 237389 6 mprj_analog_io[29]
port 565 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 566 nsew signal bidirectional
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[36]
port 567 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[36]
port 568 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[36]
port 569 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[108]
port 570 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[109]
port 571 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[110]
port 572 nsew signal input
rlabel metal2 s 41713 231813 42193 231869 6 mprj_io_enh[36]
port 573 nsew signal input
rlabel metal2 s 41713 231169 42193 231225 6 mprj_io_hldh_n[36]
port 574 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[36]
port 575 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[36]
port 576 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[36]
port 577 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[36]
port 578 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[36]
port 579 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[36]
port 580 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[36]
port 581 nsew signal input
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[36]
port 582 nsew signal tristate
rlabel metal2 s 41713 194133 42193 194189 6 mprj_analog_io[30]
port 583 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 584 nsew signal bidirectional
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[37]
port 585 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[37]
port 586 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[37]
port 587 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[111]
port 588 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[112]
port 589 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[113]
port 590 nsew signal input
rlabel metal2 s 41713 188613 42193 188669 6 mprj_io_enh[37]
port 591 nsew signal input
rlabel metal2 s 41713 187969 42193 188025 6 mprj_io_hldh_n[37]
port 592 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[37]
port 593 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[37]
port 594 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[37]
port 595 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[37]
port 596 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[37]
port 597 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[37]
port 598 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[37]
port 599 nsew signal input
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[37]
port 600 nsew signal tristate
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 602 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 620 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 638 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 656 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 674 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 692 nsew signal bidirectional
rlabel metal2 s 41713 796933 42193 796989 6 mprj_analog_io[18]
port 709 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 710 nsew signal bidirectional
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[25]
port 711 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[25]
port 712 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[25]
port 713 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[75]
port 714 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[76]
port 715 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[77]
port 716 nsew signal input
rlabel metal2 s 41713 791413 42193 791469 6 mprj_io_enh[25]
port 717 nsew signal input
rlabel metal2 s 41713 790769 42193 790825 6 mprj_io_hldh_n[25]
port 718 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[25]
port 719 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[25]
port 720 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[25]
port 721 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[25]
port 722 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[25]
port 723 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[25]
port 724 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[25]
port 725 nsew signal input
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[25]
port 726 nsew signal tristate
rlabel metal2 s 41713 753733 42193 753789 6 mprj_analog_io[19]
port 727 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 728 nsew signal bidirectional
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[26]
port 729 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[26]
port 730 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[26]
port 731 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[78]
port 732 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[79]
port 733 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[80]
port 734 nsew signal input
rlabel metal2 s 41713 748213 42193 748269 6 mprj_io_enh[26]
port 735 nsew signal input
rlabel metal2 s 41713 747569 42193 747625 6 mprj_io_hldh_n[26]
port 736 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[26]
port 737 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[26]
port 738 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[26]
port 739 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[26]
port 740 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[26]
port 741 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[26]
port 742 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[26]
port 743 nsew signal input
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[26]
port 744 nsew signal tristate
rlabel metal2 s 41713 710533 42193 710589 6 mprj_analog_io[20]
port 745 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 746 nsew signal bidirectional
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[27]
port 747 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[27]
port 748 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[27]
port 749 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[81]
port 750 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[82]
port 751 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[83]
port 752 nsew signal input
rlabel metal2 s 41713 705013 42193 705069 6 mprj_io_enh[27]
port 753 nsew signal input
rlabel metal2 s 41713 704369 42193 704425 6 mprj_io_hldh_n[27]
port 754 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[27]
port 755 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[27]
port 756 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[27]
port 757 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[27]
port 758 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[27]
port 759 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[27]
port 760 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[27]
port 761 nsew signal input
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[27]
port 762 nsew signal tristate
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 763 nsew signal input
rlabel metal2 s 145091 39934 145143 40000 6 porb_h
port 764 nsew signal input
rlabel metal1 s 145091 39934 145143 40000 6 porb_h
port 765 nsew signal input
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 766 nsew signal input
rlabel metal3 s 141667 37971 141813 39199 6 resetb_core_h
port 767 nsew signal tristate
rlabel metal3 s 141667 38031 141813 39999 6 resetb_core_h
port 768 nsew signal tristate
rlabel metal3 s 141667 39934 141813 40000 6 resetb_core_h
port 769 nsew signal tristate
rlabel metal2 s 141667 39934 141813 40000 6 resetb_core_h
port 778 nsew signal tristate
rlabel metal4 s 679377 922346 680307 922600 6 vccd1
port 779 nsew signal bidirectional
rlabel metal4 s 679377 907600 680307 907854 6 vccd1
port 780 nsew signal bidirectional
rlabel metal5 s 679397 922346 680287 922600 6 vccd1
port 781 nsew signal bidirectional
rlabel metal5 s 679397 907600 680287 907854 6 vccd1
port 782 nsew signal bidirectional
rlabel metal3 s 678000 917700 679380 922500 6 vccd1
port 783 nsew signal bidirectional
rlabel metal3 s 678000 907660 679380 912448 6 vccd1
port 784 nsew signal bidirectional
rlabel metal4 s 680587 833207 681277 833399 6 vdda1
port 786 nsew signal bidirectional
rlabel metal4 s 680587 818400 681277 818592 6 vdda1
port 787 nsew signal bidirectional
rlabel metal5 s 680607 833207 681257 833399 6 vdda1
port 788 nsew signal bidirectional
rlabel metal5 s 680607 818400 681257 818592 6 vdda1
port 789 nsew signal bidirectional
rlabel metal3 s 677600 828521 680592 833301 6 vdda1
port 790 nsew signal bidirectional
rlabel metal3 s 677600 818542 680592 823322 6 vdda1
port 791 nsew signal bidirectional
rlabel metal4 s 575600 1004947 575854 1005637 6 vssa1
port 793 nsew signal bidirectional
rlabel metal4 s 575600 1008881 575854 1008947 6 vssa1
port 794 nsew signal bidirectional
rlabel metal4 s 575600 1007929 575854 1008165 6 vssa1
port 795 nsew signal bidirectional
rlabel metal4 s 575600 1007147 575854 1007213 6 vssa1
port 796 nsew signal bidirectional
rlabel metal4 s 590346 1004947 590600 1005637 6 vssa1
port 797 nsew signal bidirectional
rlabel metal4 s 590346 1007147 590600 1007213 6 vssa1
port 798 nsew signal bidirectional
rlabel metal4 s 590346 1008881 590600 1008947 6 vssa1
port 799 nsew signal bidirectional
rlabel metal4 s 590346 1007929 590600 1008165 6 vssa1
port 800 nsew signal bidirectional
rlabel metal5 s 575600 1004968 575854 1005616 6 vssa1
port 801 nsew signal bidirectional
rlabel metal5 s 575600 1007147 575854 1008947 6 vssa1
port 802 nsew signal bidirectional
rlabel metal5 s 590346 1004968 590600 1005616 6 vssa1
port 803 nsew signal bidirectional
rlabel metal5 s 590346 1007147 590600 1008947 6 vssa1
port 804 nsew signal bidirectional
rlabel metal3 s 585678 997600 590458 1004952 6 vssa1
port 805 nsew signal bidirectional
rlabel metal3 s 575699 997600 580479 1004102 6 vssa1
port 806 nsew signal bidirectional
rlabel metal4 s 685917 474546 686847 474800 6 vssd1
port 808 nsew signal bidirectional
rlabel metal4 s 685917 459800 686847 460054 6 vssd1
port 809 nsew signal bidirectional
rlabel metal5 s 685937 474546 686827 474800 6 vssd1
port 810 nsew signal bidirectional
rlabel metal5 s 685937 459800 686827 460054 6 vssd1
port 811 nsew signal bidirectional
rlabel metal3 s 678000 469900 685920 474700 6 vssd1
port 812 nsew signal bidirectional
rlabel metal3 s 678000 459860 685920 464648 6 vssd1
port 813 nsew signal bidirectional
rlabel metal4 s 37293 912000 38223 912254 6 vccd2
port 815 nsew signal bidirectional
rlabel metal4 s 37293 926746 38223 927000 6 vccd2
port 816 nsew signal bidirectional
rlabel metal5 s 37313 912000 38203 912254 6 vccd2
port 817 nsew signal bidirectional
rlabel metal5 s 37313 926746 38203 927000 6 vccd2
port 818 nsew signal bidirectional
rlabel metal3 s 38220 912100 39600 916900 6 vccd2
port 819 nsew signal bidirectional
rlabel metal3 s 38220 922151 39600 926939 6 vccd2
port 820 nsew signal bidirectional
rlabel metal4 s 36323 483000 37013 483192 6 vdda2
port 822 nsew signal bidirectional
rlabel metal4 s 36323 497807 37013 497999 6 vdda2
port 823 nsew signal bidirectional
rlabel metal5 s 36343 483000 36993 483192 6 vdda2
port 824 nsew signal bidirectional
rlabel metal5 s 36343 497807 36993 497999 6 vdda2
port 825 nsew signal bidirectional
rlabel metal3 s 37008 483099 40000 487879 6 vdda2
port 826 nsew signal bidirectional
rlabel metal3 s 37008 493078 40000 497858 6 vdda2
port 827 nsew signal bidirectional
rlabel metal4 s 31963 827600 32653 827854 6 vssa2
port 829 nsew signal bidirectional
rlabel metal4 s 28653 827600 28719 827854 6 vssa2
port 830 nsew signal bidirectional
rlabel metal4 s 29435 827600 29671 827854 6 vssa2
port 831 nsew signal bidirectional
rlabel metal4 s 30387 827600 30453 827854 6 vssa2
port 832 nsew signal bidirectional
rlabel metal4 s 31963 842346 32653 842600 6 vssa2
port 833 nsew signal bidirectional
rlabel metal4 s 30387 842346 30453 842600 6 vssa2
port 834 nsew signal bidirectional
rlabel metal4 s 28653 842346 28719 842600 6 vssa2
port 835 nsew signal bidirectional
rlabel metal4 s 29435 842346 29671 842600 6 vssa2
port 836 nsew signal bidirectional
rlabel metal5 s 31983 827600 32631 827854 6 vssa2
port 837 nsew signal bidirectional
rlabel metal5 s 28653 827600 30453 827854 6 vssa2
port 838 nsew signal bidirectional
rlabel metal5 s 31983 842346 32631 842600 6 vssa2
port 839 nsew signal bidirectional
rlabel metal5 s 28653 842346 30453 842600 6 vssa2
port 840 nsew signal bidirectional
rlabel metal3 s 32648 837678 40000 842458 6 vssa2
port 841 nsew signal bidirectional
rlabel metal3 s 33497 827699 39999 832479 6 vssa2
port 842 nsew signal bidirectional
rlabel metal4 s 30753 440800 31683 441054 6 vssd2
port 844 nsew signal bidirectional
rlabel metal4 s 30753 455546 31683 455800 6 vssd2
port 845 nsew signal bidirectional
rlabel metal5 s 30773 440800 31663 441054 6 vssd2
port 846 nsew signal bidirectional
rlabel metal5 s 30773 455546 31663 455800 6 vssd2
port 847 nsew signal bidirectional
rlabel metal3 s 31680 440900 39600 445700 6 vssd2
port 848 nsew signal bidirectional
rlabel metal3 s 31680 450951 39600 455739 6 vssd2
port 849 nsew signal bidirectional
rlabel metal3 579121 34830 583901 40000 1 vssio
port 75 n
rlabel metal3 569142 34830 573922 40000 1 vssio
port 75 n
rlabel metal5 80222 6811 92390 18976 1 vssa
port 53 n
rlabel metal5 243266 6167 254146 19620 1 vssd
port 68 n
rlabel metal5 570422 6811 582590 18976 1 vssio
port 75 n
rlabel metal5 624222 6811 636390 18976 1 vdda
port 35 n
rlabel metal5 697980 461866 711433 472746 1 vssd1
port 808 n
rlabel metal5 698624 819822 710789 831990 1 vdda1
port 786 n
rlabel metal5 697980 909666 711433 920546 1 vccd1
port 779 n
rlabel metal5 577010 1018624 589178 1030789 1 vssa1
port 793 n
rlabel metal5 334810 1018624 346978 1030789 1 vssio
port 75 n
rlabel metal5 6167 914054 19620 924934 1 vccd2
port 815 n
rlabel metal5 6811 829010 18976 841178 1 vssa2
port 829 n
rlabel metal5 6811 484410 18976 496578 1 vdda2
port 822 n
rlabel metal5 6167 442854 19620 453734 1 vssd2
port 844 n
rlabel metal5 6811 111610 18976 123778 1 vddio
port 42 n
rlabel metal5 6167 70054 19620 80934 1 vccd
port 28 n
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
