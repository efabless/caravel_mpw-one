magic
tech sky130A
magscale 1 2
timestamp 1605064459
<< viali >>
rect 1931 5496 1965 5530
rect 1547 5274 1581 5308
rect 1931 4682 1965 4716
rect 1547 4460 1581 4494
rect 1451 3868 1485 3902
<< metal1 >>
rect 556 5724 3148 5749
rect 556 5672 1298 5724
rect 1350 5672 1362 5724
rect 1414 5672 1426 5724
rect 1478 5672 1490 5724
rect 1542 5672 2162 5724
rect 2214 5672 2226 5724
rect 2278 5672 2290 5724
rect 2342 5672 2354 5724
rect 2406 5672 3148 5724
rect 556 5647 3148 5672
rect 764 5487 770 5539
rect 822 5527 828 5539
rect 1919 5530 1977 5536
rect 1919 5527 1931 5530
rect 822 5499 1931 5527
rect 822 5487 828 5499
rect 1919 5496 1931 5499
rect 1965 5496 1977 5530
rect 1919 5490 1977 5496
rect 1532 5305 1538 5317
rect 1493 5277 1538 5305
rect 1532 5265 1538 5277
rect 1590 5265 1596 5317
rect 556 4910 3148 4935
rect 556 4858 866 4910
rect 918 4858 930 4910
rect 982 4858 994 4910
rect 1046 4858 1058 4910
rect 1110 4858 1730 4910
rect 1782 4858 1794 4910
rect 1846 4858 1858 4910
rect 1910 4858 1922 4910
rect 1974 4858 2594 4910
rect 2646 4858 2658 4910
rect 2710 4858 2722 4910
rect 2774 4858 2786 4910
rect 2838 4858 3148 4910
rect 556 4833 3148 4858
rect 1532 4673 1538 4725
rect 1590 4713 1596 4725
rect 1919 4716 1977 4722
rect 1919 4713 1931 4716
rect 1590 4685 1931 4713
rect 1590 4673 1596 4685
rect 1919 4682 1931 4685
rect 1965 4682 1977 4716
rect 1919 4676 1977 4682
rect 1535 4494 1593 4500
rect 1535 4460 1547 4494
rect 1581 4491 1593 4494
rect 1628 4491 1634 4503
rect 1581 4463 1634 4491
rect 1581 4460 1593 4463
rect 1535 4454 1593 4460
rect 1628 4451 1634 4463
rect 1686 4451 1692 4503
rect 556 4096 3148 4121
rect 556 4044 1298 4096
rect 1350 4044 1362 4096
rect 1414 4044 1426 4096
rect 1478 4044 1490 4096
rect 1542 4044 2162 4096
rect 2214 4044 2226 4096
rect 2278 4044 2290 4096
rect 2342 4044 2354 4096
rect 2406 4044 3148 4096
rect 556 4019 3148 4044
rect 1439 3902 1497 3908
rect 1439 3868 1451 3902
rect 1485 3899 1497 3902
rect 1628 3899 1634 3911
rect 1485 3871 1634 3899
rect 1485 3868 1497 3871
rect 1439 3862 1497 3868
rect 1628 3859 1634 3871
rect 1686 3859 1692 3911
rect 556 3282 3148 3307
rect 556 3230 866 3282
rect 918 3230 930 3282
rect 982 3230 994 3282
rect 1046 3230 1058 3282
rect 1110 3230 1730 3282
rect 1782 3230 1794 3282
rect 1846 3230 1858 3282
rect 1910 3230 1922 3282
rect 1974 3230 2594 3282
rect 2646 3230 2658 3282
rect 2710 3230 2722 3282
rect 2774 3230 2786 3282
rect 2838 3230 3148 3282
rect 556 3205 3148 3230
<< via1 >>
rect 1298 5672 1350 5724
rect 1362 5672 1414 5724
rect 1426 5672 1478 5724
rect 1490 5672 1542 5724
rect 2162 5672 2214 5724
rect 2226 5672 2278 5724
rect 2290 5672 2342 5724
rect 2354 5672 2406 5724
rect 770 5487 822 5539
rect 1538 5308 1590 5317
rect 1538 5274 1547 5308
rect 1547 5274 1581 5308
rect 1581 5274 1590 5308
rect 1538 5265 1590 5274
rect 866 4858 918 4910
rect 930 4858 982 4910
rect 994 4858 1046 4910
rect 1058 4858 1110 4910
rect 1730 4858 1782 4910
rect 1794 4858 1846 4910
rect 1858 4858 1910 4910
rect 1922 4858 1974 4910
rect 2594 4858 2646 4910
rect 2658 4858 2710 4910
rect 2722 4858 2774 4910
rect 2786 4858 2838 4910
rect 1538 4673 1590 4725
rect 1634 4451 1686 4503
rect 1298 4044 1350 4096
rect 1362 4044 1414 4096
rect 1426 4044 1478 4096
rect 1490 4044 1542 4096
rect 2162 4044 2214 4096
rect 2226 4044 2278 4096
rect 2290 4044 2342 4096
rect 2354 4044 2406 4096
rect 1634 3859 1686 3911
rect 866 3230 918 3282
rect 930 3230 982 3282
rect 994 3230 1046 3282
rect 1058 3230 1110 3282
rect 1730 3230 1782 3282
rect 1794 3230 1846 3282
rect 1858 3230 1910 3282
rect 1922 3230 1974 3282
rect 2594 3230 2646 3282
rect 2658 3230 2710 3282
rect 2722 3230 2774 3282
rect 2786 3230 2838 3282
<< metal2 >>
rect 768 8364 824 9164
rect 782 5545 810 8364
rect 1272 5726 1568 5749
rect 1328 5724 1352 5726
rect 1408 5724 1432 5726
rect 1488 5724 1512 5726
rect 1350 5672 1352 5724
rect 1414 5672 1426 5724
rect 1488 5672 1490 5724
rect 1328 5670 1352 5672
rect 1408 5670 1432 5672
rect 1488 5670 1512 5672
rect 1272 5647 1568 5670
rect 2136 5726 2432 5749
rect 2192 5724 2216 5726
rect 2272 5724 2296 5726
rect 2352 5724 2376 5726
rect 2214 5672 2216 5724
rect 2278 5672 2290 5724
rect 2352 5672 2354 5724
rect 2192 5670 2216 5672
rect 2272 5670 2296 5672
rect 2352 5670 2376 5672
rect 2136 5647 2432 5670
rect 770 5539 822 5545
rect 770 5481 822 5487
rect 1538 5317 1590 5323
rect 1538 5259 1590 5265
rect 840 4912 1136 4935
rect 896 4910 920 4912
rect 976 4910 1000 4912
rect 1056 4910 1080 4912
rect 918 4858 920 4910
rect 982 4858 994 4910
rect 1056 4858 1058 4910
rect 896 4856 920 4858
rect 976 4856 1000 4858
rect 1056 4856 1080 4858
rect 840 4833 1136 4856
rect 1550 4731 1578 5259
rect 1704 4912 2000 4935
rect 1760 4910 1784 4912
rect 1840 4910 1864 4912
rect 1920 4910 1944 4912
rect 1782 4858 1784 4910
rect 1846 4858 1858 4910
rect 1920 4858 1922 4910
rect 1760 4856 1784 4858
rect 1840 4856 1864 4858
rect 1920 4856 1944 4858
rect 1704 4833 2000 4856
rect 2568 4912 2864 4935
rect 2624 4910 2648 4912
rect 2704 4910 2728 4912
rect 2784 4910 2808 4912
rect 2646 4858 2648 4910
rect 2710 4858 2722 4910
rect 2784 4858 2786 4910
rect 2624 4856 2648 4858
rect 2704 4856 2728 4858
rect 2784 4856 2808 4858
rect 2568 4833 2864 4856
rect 1538 4725 1590 4731
rect 1538 4667 1590 4673
rect 1634 4503 1686 4509
rect 1634 4445 1686 4451
rect 1272 4098 1568 4121
rect 1328 4096 1352 4098
rect 1408 4096 1432 4098
rect 1488 4096 1512 4098
rect 1350 4044 1352 4096
rect 1414 4044 1426 4096
rect 1488 4044 1490 4096
rect 1328 4042 1352 4044
rect 1408 4042 1432 4044
rect 1488 4042 1512 4044
rect 1272 4019 1568 4042
rect 1646 3917 1674 4445
rect 2136 4098 2432 4121
rect 2192 4096 2216 4098
rect 2272 4096 2296 4098
rect 2352 4096 2376 4098
rect 2214 4044 2216 4096
rect 2278 4044 2290 4096
rect 2352 4044 2354 4096
rect 2192 4042 2216 4044
rect 2272 4042 2296 4044
rect 2352 4042 2376 4044
rect 2136 4019 2432 4042
rect 1634 3911 1686 3917
rect 1634 3853 1686 3859
rect 840 3284 1136 3307
rect 896 3282 920 3284
rect 976 3282 1000 3284
rect 1056 3282 1080 3284
rect 918 3230 920 3282
rect 982 3230 994 3282
rect 1056 3230 1058 3282
rect 896 3228 920 3230
rect 976 3228 1000 3230
rect 1056 3228 1080 3230
rect 840 3205 1136 3228
rect 1704 3284 2000 3307
rect 1760 3282 1784 3284
rect 1840 3282 1864 3284
rect 1920 3282 1944 3284
rect 1782 3230 1784 3282
rect 1846 3230 1858 3282
rect 1920 3230 1922 3282
rect 1760 3228 1784 3230
rect 1840 3228 1864 3230
rect 1920 3228 1944 3230
rect 1704 3205 2000 3228
rect 2568 3284 2864 3307
rect 2624 3282 2648 3284
rect 2704 3282 2728 3284
rect 2784 3282 2808 3284
rect 2646 3230 2648 3282
rect 2710 3230 2722 3282
rect 2784 3230 2786 3282
rect 2624 3228 2648 3230
rect 2704 3228 2728 3230
rect 2784 3228 2808 3230
rect 2568 3205 2864 3228
rect 0 0 56 800
<< via2 >>
rect 1272 5724 1328 5726
rect 1352 5724 1408 5726
rect 1432 5724 1488 5726
rect 1512 5724 1568 5726
rect 1272 5672 1298 5724
rect 1298 5672 1328 5724
rect 1352 5672 1362 5724
rect 1362 5672 1408 5724
rect 1432 5672 1478 5724
rect 1478 5672 1488 5724
rect 1512 5672 1542 5724
rect 1542 5672 1568 5724
rect 1272 5670 1328 5672
rect 1352 5670 1408 5672
rect 1432 5670 1488 5672
rect 1512 5670 1568 5672
rect 2136 5724 2192 5726
rect 2216 5724 2272 5726
rect 2296 5724 2352 5726
rect 2376 5724 2432 5726
rect 2136 5672 2162 5724
rect 2162 5672 2192 5724
rect 2216 5672 2226 5724
rect 2226 5672 2272 5724
rect 2296 5672 2342 5724
rect 2342 5672 2352 5724
rect 2376 5672 2406 5724
rect 2406 5672 2432 5724
rect 2136 5670 2192 5672
rect 2216 5670 2272 5672
rect 2296 5670 2352 5672
rect 2376 5670 2432 5672
rect 840 4910 896 4912
rect 920 4910 976 4912
rect 1000 4910 1056 4912
rect 1080 4910 1136 4912
rect 840 4858 866 4910
rect 866 4858 896 4910
rect 920 4858 930 4910
rect 930 4858 976 4910
rect 1000 4858 1046 4910
rect 1046 4858 1056 4910
rect 1080 4858 1110 4910
rect 1110 4858 1136 4910
rect 840 4856 896 4858
rect 920 4856 976 4858
rect 1000 4856 1056 4858
rect 1080 4856 1136 4858
rect 1704 4910 1760 4912
rect 1784 4910 1840 4912
rect 1864 4910 1920 4912
rect 1944 4910 2000 4912
rect 1704 4858 1730 4910
rect 1730 4858 1760 4910
rect 1784 4858 1794 4910
rect 1794 4858 1840 4910
rect 1864 4858 1910 4910
rect 1910 4858 1920 4910
rect 1944 4858 1974 4910
rect 1974 4858 2000 4910
rect 1704 4856 1760 4858
rect 1784 4856 1840 4858
rect 1864 4856 1920 4858
rect 1944 4856 2000 4858
rect 2568 4910 2624 4912
rect 2648 4910 2704 4912
rect 2728 4910 2784 4912
rect 2808 4910 2864 4912
rect 2568 4858 2594 4910
rect 2594 4858 2624 4910
rect 2648 4858 2658 4910
rect 2658 4858 2704 4910
rect 2728 4858 2774 4910
rect 2774 4858 2784 4910
rect 2808 4858 2838 4910
rect 2838 4858 2864 4910
rect 2568 4856 2624 4858
rect 2648 4856 2704 4858
rect 2728 4856 2784 4858
rect 2808 4856 2864 4858
rect 1272 4096 1328 4098
rect 1352 4096 1408 4098
rect 1432 4096 1488 4098
rect 1512 4096 1568 4098
rect 1272 4044 1298 4096
rect 1298 4044 1328 4096
rect 1352 4044 1362 4096
rect 1362 4044 1408 4096
rect 1432 4044 1478 4096
rect 1478 4044 1488 4096
rect 1512 4044 1542 4096
rect 1542 4044 1568 4096
rect 1272 4042 1328 4044
rect 1352 4042 1408 4044
rect 1432 4042 1488 4044
rect 1512 4042 1568 4044
rect 2136 4096 2192 4098
rect 2216 4096 2272 4098
rect 2296 4096 2352 4098
rect 2376 4096 2432 4098
rect 2136 4044 2162 4096
rect 2162 4044 2192 4096
rect 2216 4044 2226 4096
rect 2226 4044 2272 4096
rect 2296 4044 2342 4096
rect 2342 4044 2352 4096
rect 2376 4044 2406 4096
rect 2406 4044 2432 4096
rect 2136 4042 2192 4044
rect 2216 4042 2272 4044
rect 2296 4042 2352 4044
rect 2376 4042 2432 4044
rect 840 3282 896 3284
rect 920 3282 976 3284
rect 1000 3282 1056 3284
rect 1080 3282 1136 3284
rect 840 3230 866 3282
rect 866 3230 896 3282
rect 920 3230 930 3282
rect 930 3230 976 3282
rect 1000 3230 1046 3282
rect 1046 3230 1056 3282
rect 1080 3230 1110 3282
rect 1110 3230 1136 3282
rect 840 3228 896 3230
rect 920 3228 976 3230
rect 1000 3228 1056 3230
rect 1080 3228 1136 3230
rect 1704 3282 1760 3284
rect 1784 3282 1840 3284
rect 1864 3282 1920 3284
rect 1944 3282 2000 3284
rect 1704 3230 1730 3282
rect 1730 3230 1760 3282
rect 1784 3230 1794 3282
rect 1794 3230 1840 3282
rect 1864 3230 1910 3282
rect 1910 3230 1920 3282
rect 1944 3230 1974 3282
rect 1974 3230 2000 3282
rect 1704 3228 1760 3230
rect 1784 3228 1840 3230
rect 1864 3228 1920 3230
rect 1944 3228 2000 3230
rect 2568 3282 2624 3284
rect 2648 3282 2704 3284
rect 2728 3282 2784 3284
rect 2808 3282 2864 3284
rect 2568 3230 2594 3282
rect 2594 3230 2624 3282
rect 2648 3230 2658 3282
rect 2658 3230 2704 3282
rect 2728 3230 2774 3282
rect 2774 3230 2784 3282
rect 2808 3230 2838 3282
rect 2838 3230 2864 3282
rect 2568 3228 2624 3230
rect 2648 3228 2704 3230
rect 2728 3228 2784 3230
rect 2808 3228 2864 3230
<< metal3 >>
rect 1260 5730 1580 5731
rect 1260 5666 1268 5730
rect 1332 5666 1348 5730
rect 1412 5666 1428 5730
rect 1492 5666 1508 5730
rect 1572 5666 1580 5730
rect 1260 5665 1580 5666
rect 2124 5730 2444 5731
rect 2124 5666 2132 5730
rect 2196 5666 2212 5730
rect 2276 5666 2292 5730
rect 2356 5666 2372 5730
rect 2436 5666 2444 5730
rect 2124 5665 2444 5666
rect 828 4916 1148 4917
rect 828 4852 836 4916
rect 900 4852 916 4916
rect 980 4852 996 4916
rect 1060 4852 1076 4916
rect 1140 4852 1148 4916
rect 828 4851 1148 4852
rect 1692 4916 2012 4917
rect 1692 4852 1700 4916
rect 1764 4852 1780 4916
rect 1844 4852 1860 4916
rect 1924 4852 1940 4916
rect 2004 4852 2012 4916
rect 1692 4851 2012 4852
rect 2556 4916 2876 4917
rect 2556 4852 2564 4916
rect 2628 4852 2644 4916
rect 2708 4852 2724 4916
rect 2788 4852 2804 4916
rect 2868 4852 2876 4916
rect 2556 4851 2876 4852
rect 1260 4102 1580 4103
rect 1260 4038 1268 4102
rect 1332 4038 1348 4102
rect 1412 4038 1428 4102
rect 1492 4038 1508 4102
rect 1572 4038 1580 4102
rect 1260 4037 1580 4038
rect 2124 4102 2444 4103
rect 2124 4038 2132 4102
rect 2196 4038 2212 4102
rect 2276 4038 2292 4102
rect 2356 4038 2372 4102
rect 2436 4038 2444 4102
rect 2124 4037 2444 4038
rect 3560 3862 4360 3982
rect 828 3288 1148 3289
rect 828 3224 836 3288
rect 900 3224 916 3288
rect 980 3224 996 3288
rect 1060 3224 1076 3288
rect 1140 3224 1148 3288
rect 828 3223 1148 3224
rect 1692 3288 2012 3289
rect 1692 3224 1700 3288
rect 1764 3224 1780 3288
rect 1844 3224 1860 3288
rect 1924 3224 1940 3288
rect 2004 3224 2012 3288
rect 1692 3223 2012 3224
rect 2556 3288 2876 3289
rect 2556 3224 2564 3288
rect 2628 3224 2644 3288
rect 2708 3224 2724 3288
rect 2788 3224 2804 3288
rect 2868 3224 2876 3288
rect 2556 3223 2876 3224
<< via3 >>
rect 1268 5726 1332 5730
rect 1268 5670 1272 5726
rect 1272 5670 1328 5726
rect 1328 5670 1332 5726
rect 1268 5666 1332 5670
rect 1348 5726 1412 5730
rect 1348 5670 1352 5726
rect 1352 5670 1408 5726
rect 1408 5670 1412 5726
rect 1348 5666 1412 5670
rect 1428 5726 1492 5730
rect 1428 5670 1432 5726
rect 1432 5670 1488 5726
rect 1488 5670 1492 5726
rect 1428 5666 1492 5670
rect 1508 5726 1572 5730
rect 1508 5670 1512 5726
rect 1512 5670 1568 5726
rect 1568 5670 1572 5726
rect 1508 5666 1572 5670
rect 2132 5726 2196 5730
rect 2132 5670 2136 5726
rect 2136 5670 2192 5726
rect 2192 5670 2196 5726
rect 2132 5666 2196 5670
rect 2212 5726 2276 5730
rect 2212 5670 2216 5726
rect 2216 5670 2272 5726
rect 2272 5670 2276 5726
rect 2212 5666 2276 5670
rect 2292 5726 2356 5730
rect 2292 5670 2296 5726
rect 2296 5670 2352 5726
rect 2352 5670 2356 5726
rect 2292 5666 2356 5670
rect 2372 5726 2436 5730
rect 2372 5670 2376 5726
rect 2376 5670 2432 5726
rect 2432 5670 2436 5726
rect 2372 5666 2436 5670
rect 836 4912 900 4916
rect 836 4856 840 4912
rect 840 4856 896 4912
rect 896 4856 900 4912
rect 836 4852 900 4856
rect 916 4912 980 4916
rect 916 4856 920 4912
rect 920 4856 976 4912
rect 976 4856 980 4912
rect 916 4852 980 4856
rect 996 4912 1060 4916
rect 996 4856 1000 4912
rect 1000 4856 1056 4912
rect 1056 4856 1060 4912
rect 996 4852 1060 4856
rect 1076 4912 1140 4916
rect 1076 4856 1080 4912
rect 1080 4856 1136 4912
rect 1136 4856 1140 4912
rect 1076 4852 1140 4856
rect 1700 4912 1764 4916
rect 1700 4856 1704 4912
rect 1704 4856 1760 4912
rect 1760 4856 1764 4912
rect 1700 4852 1764 4856
rect 1780 4912 1844 4916
rect 1780 4856 1784 4912
rect 1784 4856 1840 4912
rect 1840 4856 1844 4912
rect 1780 4852 1844 4856
rect 1860 4912 1924 4916
rect 1860 4856 1864 4912
rect 1864 4856 1920 4912
rect 1920 4856 1924 4912
rect 1860 4852 1924 4856
rect 1940 4912 2004 4916
rect 1940 4856 1944 4912
rect 1944 4856 2000 4912
rect 2000 4856 2004 4912
rect 1940 4852 2004 4856
rect 2564 4912 2628 4916
rect 2564 4856 2568 4912
rect 2568 4856 2624 4912
rect 2624 4856 2628 4912
rect 2564 4852 2628 4856
rect 2644 4912 2708 4916
rect 2644 4856 2648 4912
rect 2648 4856 2704 4912
rect 2704 4856 2708 4912
rect 2644 4852 2708 4856
rect 2724 4912 2788 4916
rect 2724 4856 2728 4912
rect 2728 4856 2784 4912
rect 2784 4856 2788 4912
rect 2724 4852 2788 4856
rect 2804 4912 2868 4916
rect 2804 4856 2808 4912
rect 2808 4856 2864 4912
rect 2864 4856 2868 4912
rect 2804 4852 2868 4856
rect 1268 4098 1332 4102
rect 1268 4042 1272 4098
rect 1272 4042 1328 4098
rect 1328 4042 1332 4098
rect 1268 4038 1332 4042
rect 1348 4098 1412 4102
rect 1348 4042 1352 4098
rect 1352 4042 1408 4098
rect 1408 4042 1412 4098
rect 1348 4038 1412 4042
rect 1428 4098 1492 4102
rect 1428 4042 1432 4098
rect 1432 4042 1488 4098
rect 1488 4042 1492 4098
rect 1428 4038 1492 4042
rect 1508 4098 1572 4102
rect 1508 4042 1512 4098
rect 1512 4042 1568 4098
rect 1568 4042 1572 4098
rect 1508 4038 1572 4042
rect 2132 4098 2196 4102
rect 2132 4042 2136 4098
rect 2136 4042 2192 4098
rect 2192 4042 2196 4098
rect 2132 4038 2196 4042
rect 2212 4098 2276 4102
rect 2212 4042 2216 4098
rect 2216 4042 2272 4098
rect 2272 4042 2276 4098
rect 2212 4038 2276 4042
rect 2292 4098 2356 4102
rect 2292 4042 2296 4098
rect 2296 4042 2352 4098
rect 2352 4042 2356 4098
rect 2292 4038 2356 4042
rect 2372 4098 2436 4102
rect 2372 4042 2376 4098
rect 2376 4042 2432 4098
rect 2432 4042 2436 4098
rect 2372 4038 2436 4042
rect 836 3284 900 3288
rect 836 3228 840 3284
rect 840 3228 896 3284
rect 896 3228 900 3284
rect 836 3224 900 3228
rect 916 3284 980 3288
rect 916 3228 920 3284
rect 920 3228 976 3284
rect 976 3228 980 3284
rect 916 3224 980 3228
rect 996 3284 1060 3288
rect 996 3228 1000 3284
rect 1000 3228 1056 3284
rect 1056 3228 1060 3284
rect 996 3224 1060 3228
rect 1076 3284 1140 3288
rect 1076 3228 1080 3284
rect 1080 3228 1136 3284
rect 1136 3228 1140 3284
rect 1076 3224 1140 3228
rect 1700 3284 1764 3288
rect 1700 3228 1704 3284
rect 1704 3228 1760 3284
rect 1760 3228 1764 3284
rect 1700 3224 1764 3228
rect 1780 3284 1844 3288
rect 1780 3228 1784 3284
rect 1784 3228 1840 3284
rect 1840 3228 1844 3284
rect 1780 3224 1844 3228
rect 1860 3284 1924 3288
rect 1860 3228 1864 3284
rect 1864 3228 1920 3284
rect 1920 3228 1924 3284
rect 1860 3224 1924 3228
rect 1940 3284 2004 3288
rect 1940 3228 1944 3284
rect 1944 3228 2000 3284
rect 2000 3228 2004 3284
rect 1940 3224 2004 3228
rect 2564 3284 2628 3288
rect 2564 3228 2568 3284
rect 2568 3228 2624 3284
rect 2624 3228 2628 3284
rect 2564 3224 2628 3228
rect 2644 3284 2708 3288
rect 2644 3228 2648 3284
rect 2648 3228 2704 3284
rect 2704 3228 2708 3284
rect 2644 3224 2708 3228
rect 2724 3284 2788 3288
rect 2724 3228 2728 3284
rect 2728 3228 2784 3284
rect 2784 3228 2788 3284
rect 2724 3224 2788 3228
rect 2804 3284 2868 3288
rect 2804 3228 2808 3284
rect 2808 3228 2864 3284
rect 2864 3228 2868 3284
rect 2804 3224 2868 3228
<< metal4 >>
rect 828 5358 1148 5749
rect 828 5122 870 5358
rect 1106 5122 1148 5358
rect 828 4916 1148 5122
rect 828 4852 836 4916
rect 900 4852 916 4916
rect 980 4852 996 4916
rect 1060 4852 1076 4916
rect 1140 4852 1148 4916
rect 828 4544 1148 4852
rect 828 4308 870 4544
rect 1106 4308 1148 4544
rect 828 3730 1148 4308
rect 828 3494 870 3730
rect 1106 3494 1148 3730
rect 828 3288 1148 3494
rect 828 3224 836 3288
rect 900 3224 916 3288
rect 980 3224 996 3288
rect 1060 3224 1076 3288
rect 1140 3224 1148 3288
rect 828 3205 1148 3224
rect 1260 5730 1580 5749
rect 1260 5666 1268 5730
rect 1332 5666 1348 5730
rect 1412 5666 1428 5730
rect 1492 5666 1508 5730
rect 1572 5666 1580 5730
rect 1260 4951 1580 5666
rect 1260 4715 1302 4951
rect 1538 4715 1580 4951
rect 1260 4137 1580 4715
rect 1260 4102 1302 4137
rect 1538 4102 1580 4137
rect 1260 4038 1268 4102
rect 1572 4038 1580 4102
rect 1260 3901 1302 4038
rect 1538 3901 1580 4038
rect 1260 3205 1580 3901
rect 1692 5358 2012 5749
rect 1692 5122 1734 5358
rect 1970 5122 2012 5358
rect 1692 4916 2012 5122
rect 1692 4852 1700 4916
rect 1764 4852 1780 4916
rect 1844 4852 1860 4916
rect 1924 4852 1940 4916
rect 2004 4852 2012 4916
rect 1692 4544 2012 4852
rect 1692 4308 1734 4544
rect 1970 4308 2012 4544
rect 1692 3730 2012 4308
rect 1692 3494 1734 3730
rect 1970 3494 2012 3730
rect 1692 3288 2012 3494
rect 1692 3224 1700 3288
rect 1764 3224 1780 3288
rect 1844 3224 1860 3288
rect 1924 3224 1940 3288
rect 2004 3224 2012 3288
rect 1692 3205 2012 3224
rect 2124 5730 2444 5749
rect 2124 5666 2132 5730
rect 2196 5666 2212 5730
rect 2276 5666 2292 5730
rect 2356 5666 2372 5730
rect 2436 5666 2444 5730
rect 2124 4951 2444 5666
rect 2124 4715 2166 4951
rect 2402 4715 2444 4951
rect 2124 4137 2444 4715
rect 2124 4102 2166 4137
rect 2402 4102 2444 4137
rect 2124 4038 2132 4102
rect 2436 4038 2444 4102
rect 2124 3901 2166 4038
rect 2402 3901 2444 4038
rect 2124 3205 2444 3901
rect 2556 5358 2876 5749
rect 2556 5122 2598 5358
rect 2834 5122 2876 5358
rect 2556 4916 2876 5122
rect 2556 4852 2564 4916
rect 2628 4852 2644 4916
rect 2708 4852 2724 4916
rect 2788 4852 2804 4916
rect 2868 4852 2876 4916
rect 2556 4544 2876 4852
rect 2556 4308 2598 4544
rect 2834 4308 2876 4544
rect 2556 3730 2876 4308
rect 2556 3494 2598 3730
rect 2834 3494 2876 3730
rect 2556 3288 2876 3494
rect 2556 3224 2564 3288
rect 2628 3224 2644 3288
rect 2708 3224 2724 3288
rect 2788 3224 2804 3288
rect 2868 3224 2876 3288
rect 2556 3205 2876 3224
<< via4 >>
rect 870 5122 1106 5358
rect 870 4308 1106 4544
rect 870 3494 1106 3730
rect 1302 4715 1538 4951
rect 1302 4102 1538 4137
rect 1302 4038 1332 4102
rect 1332 4038 1348 4102
rect 1348 4038 1412 4102
rect 1412 4038 1428 4102
rect 1428 4038 1492 4102
rect 1492 4038 1508 4102
rect 1508 4038 1538 4102
rect 1302 3901 1538 4038
rect 1734 5122 1970 5358
rect 1734 4308 1970 4544
rect 1734 3494 1970 3730
rect 2166 4715 2402 4951
rect 2166 4102 2402 4137
rect 2166 4038 2196 4102
rect 2196 4038 2212 4102
rect 2212 4038 2276 4102
rect 2276 4038 2292 4102
rect 2292 4038 2356 4102
rect 2356 4038 2372 4102
rect 2372 4038 2402 4102
rect 2166 3901 2402 4038
rect 2598 5122 2834 5358
rect 2598 4308 2834 4544
rect 2598 3494 2834 3730
<< metal5 >>
rect 556 5358 3148 5400
rect 556 5122 870 5358
rect 1106 5122 1734 5358
rect 1970 5122 2598 5358
rect 2834 5122 3148 5358
rect 556 5080 3148 5122
rect 556 4951 3148 4993
rect 556 4715 1302 4951
rect 1538 4715 2166 4951
rect 2402 4715 3148 4951
rect 556 4673 3148 4715
rect 556 4544 3148 4586
rect 556 4308 870 4544
rect 1106 4308 1734 4544
rect 1970 4308 2598 4544
rect 2834 4308 3148 4544
rect 556 4266 3148 4308
rect 556 4137 3148 4179
rect 556 3901 1302 4137
rect 1538 3901 2166 4137
rect 2402 3901 3148 4137
rect 556 3859 3148 3901
rect 556 3730 3148 3772
rect 556 3494 870 3730
rect 1106 3494 1734 3730
rect 1970 3494 2598 3730
rect 2834 3494 3148 3730
rect 556 3452 3148 3494
use sky130_fd_sc_hvl__conb_1  _1_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1604489734
transform 1 0 1228 0 -1 4070
box -66 -23 546 897
use sky130_fd_sc_hvl__schmittbuf_1  hystbuf1 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1604489734
transform 1 0 940 0 1 4070
box -66 -23 1122 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_0 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1604489734
transform 1 0 556 0 -1 4070
box -66 -23 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_0_4 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1604489734
transform 1 0 940 0 -1 4070
box -66 -23 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_0_6 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1604489734
transform 1 0 1132 0 -1 4070
box -66 -23 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_12 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1604489734
transform 1 0 1708 0 -1 4070
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_0
timestamp 1604489734
transform 1 0 556 0 1 4070
box -66 -23 450 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_20
timestamp 1604489734
transform 1 0 2476 0 -1 4070
box -66 -23 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_0_24
timestamp 1604489734
transform 1 0 2860 0 -1 4070
box -66 -23 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_15
timestamp 1604489734
transform 1 0 1996 0 1 4070
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_23
timestamp 1604489734
transform 1 0 2764 0 1 4070
box -66 -23 450 897
use sky130_fd_sc_hvl__fill_1  FILLER_0_26
timestamp 1604489734
transform 1 0 3052 0 -1 4070
box -66 -23 162 897
use sky130_fd_sc_hvl__schmittbuf_1  hystbuf2
timestamp 1604489734
transform 1 0 940 0 -1 5698
box -66 -23 1122 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_0
timestamp 1604489734
transform 1 0 556 0 -1 5698
box -66 -23 450 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_15
timestamp 1604489734
transform 1 0 1996 0 -1 5698
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_23
timestamp 1604489734
transform 1 0 2764 0 -1 5698
box -66 -23 450 897
<< labels >>
rlabel metal2 s 768 8364 824 9164 6 porb_h
port 0 nsew default tristate
rlabel metal2 s 0 0 56 800 6 vdd3v3
port 1 nsew default input
rlabel metal3 s 3560 3862 4360 3982 6 vss
port 2 nsew default input
rlabel metal5 s 556 3452 3148 3772 6 VPWR
port 3 nsew default input
rlabel metal5 s 556 3859 3148 4179 6 VGND
port 4 nsew default input
<< properties >>
string FIXED_BBOX 0 0 4360 9164
<< end >>
