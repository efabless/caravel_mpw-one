***  
* Most models come from here:

.lib ../../../sky130A-xyce/libs.tech/xyce/sky130.lib.spice tt

.include ./sky130_fd_io__condiode.spice
.include ./sky130_fd_pr__model__parasitic__diode_ps2nw.spice 
.include ./sky130_fd_pr__model__parasitic__diode_pw2dn.spice
.include ./sky130_fd_pr__model__parasitic__diode_ps2dn.spice


*.include ./sky130_fd_pr__model__parasitic__diode_ps2nw.model.spice 
*.include ./sky130_fd_pr__model__parasitic__diode_pw2dn.model.spice
*.include ./sky130_fd_pr__model__parasitic__diode_ps2dn.model.spice


***************************************

.include 	../NETLISTS/sky130_fd_io__top_xres4v2-extracted.spice

*** no space before the .include
*** removed subckts without any ports
*** converted calibre extracted netlist to spice with hs2ng
*** changed parasitic diodes to level=2.0
*** used sky130A-xyce PDK from MG

***************************************
Xsky130_fd_io__top_xres4v2 
+ VSS		; VSSD 
+ VDD3V3	; VDDIO 
+ VDD1V8	; VCCHIB 
+ VDD3V3	; VDDIO_Q 
+ ONE3V3	; ENABLE_H 
+ ONE3V3	; EN_VDDIO_SIG_H 
+ ZERO	 	; INP_SEL_H 
+ ONE1V8	; ENABLE_VDDIO 
+ PAD		; PAD 
+ ZERO		; PULLUP_H 
+ ONE3V3	; DISABLE_PULLUP_H
+ OPEN2		; PAD_A_ESD_H 
+ VSS		; VSSIO 
+ ONE3V3	; FILT_IN_H 
+ OPEN3		; TIE_LO_ESD 
+ ZERO		; XRES_H_N 
+ OPEN4		; TIE_HI_ESD 
+ OPEN5		; TIE_WEAK_HI_H 
+ VDD1V8	; VCCD 
+ VDD3V3	; VDDA
+ VDD3V3	; VSWITCH 
+ VSS		; VSSA 
+ OPEN6		; AMUXBUS_B 
+ OPEN7		; AMUXBUS_A 
+ VSS		; VSSIO_Q 
+ sky130_fd_io__top_xres4v2


vvss		VSS		0 		dc 	0
vvdd1v8		VDD1V8		0 		pwl	0 0 3u  1.8  1m 1.8
vvdd3v3		VDD3V3		0 		pwl	0 0 2u  3.3  1m 3.3

vzero		ZERO		0		dc	0
vone1v8		ONE1V8		0		pwl	0 0 5.5u 0 5.6u 1.8  1m 1.8
vone3v3		ONE3V3		0		pwl	0 0 5.5u 0 5.6u 3.3  1m 3.3

vout		OUT		0		pwl	0 0 8u 0  8.1u 1.8 11u 1.8 11.1u 0 15u 0
rload		PAD		0		1000K


.PRINT TRAN FORMAT=RAW v(pad) v(out) i(vvdd3v3) i(vvdd1v8) v(vdd3v3) v(vdd1v8) v(ONE1V8) v(ONE3V3) i(vone1v8) i(vone3v3) i(vout) i(rload)
.TRAN 10n 15u

.END
