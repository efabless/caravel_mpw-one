magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1260 -1260 1261 1261
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 8815304
string GDS_START 8809604
<< end >>
