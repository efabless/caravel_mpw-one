magic
tech sky130A
magscale 1 2
timestamp 1606520338
<< error_p >>
rect -2181 -1600 -2061 1600
rect -1941 -1600 -1821 1600
rect 1821 -1600 1941 1600
rect 2061 -1600 2181 1600
<< metal3 >>
rect -5943 1572 -2061 1600
rect -5943 -1572 -2145 1572
rect -2081 -1572 -2061 1572
rect -5943 -1600 -2061 -1572
rect -1941 1572 1941 1600
rect -1941 -1572 1857 1572
rect 1921 -1572 1941 1572
rect -1941 -1600 1941 -1572
rect 2061 1572 5943 1600
rect 2061 -1572 5859 1572
rect 5923 -1572 5943 1572
rect 2061 -1600 5943 -1572
<< via3 >>
rect -2145 -1572 -2081 1572
rect 1857 -1572 1921 1572
rect 5859 -1572 5923 1572
<< mimcap >>
rect -5843 1460 -2333 1500
rect -5843 -1460 -5803 1460
rect -2373 -1460 -2333 1460
rect -5843 -1500 -2333 -1460
rect -1841 1460 1669 1500
rect -1841 -1460 -1801 1460
rect 1629 -1460 1669 1460
rect -1841 -1500 1669 -1460
rect 2161 1460 5671 1500
rect 2161 -1460 2201 1460
rect 5631 -1460 5671 1460
rect 2161 -1500 5671 -1460
<< mimcapcontact >>
rect -5803 -1460 -2373 1460
rect -1801 -1460 1629 1460
rect 2201 -1460 5631 1460
<< metal4 >>
rect -2161 1572 -2065 1588
rect -5804 1460 -2372 1461
rect -5804 -1460 -5803 1460
rect -2373 -1460 -2372 1460
rect -5804 -1461 -2372 -1460
rect -2161 -1572 -2145 1572
rect -2081 -1572 -2065 1572
rect 1841 1572 1937 1588
rect -1802 1460 1630 1461
rect -1802 -1460 -1801 1460
rect 1629 -1460 1630 1460
rect -1802 -1461 1630 -1460
rect -2161 -1588 -2065 -1572
rect 1841 -1572 1857 1572
rect 1921 -1572 1937 1572
rect 5843 1572 5939 1588
rect 2200 1460 5632 1461
rect 2200 -1460 2201 1460
rect 5631 -1460 5632 1460
rect 2200 -1461 5632 -1460
rect 1841 -1588 1937 -1572
rect 5843 -1572 5859 1572
rect 5923 -1572 5939 1572
rect 5843 -1588 5939 -1572
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 2061 -1600 5771 1600
string parameters w 17.55 l 15.0 val 274.317 carea 1.00 cperi 0.17 nx 3 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 0
string library sky130
<< end >>
