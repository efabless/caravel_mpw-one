magic
tech sky130A
magscale 12 1
timestamp 1598774708
<< metal5 >>
rect 15 90 30 105
rect 0 75 45 90
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
