magic
tech sky130A
magscale 1 2
timestamp 1607547389
<< checkpaint >>
rect -1260 -1259 41262 5465
<< viali >>
rect 13471 2694 13505 2728
rect 14815 2694 14849 2728
rect 10495 1880 10529 1914
rect 36799 1880 36833 1914
rect 10975 1288 11009 1322
rect 37375 1066 37409 1100
<< metal1 >>
rect 960 4180 39936 4205
rect 960 4128 13947 4180
rect 13999 4128 26960 4180
rect 27012 4128 39936 4180
rect 960 4103 39936 4128
rect 960 3366 39936 3391
rect 960 3314 7440 3366
rect 7492 3314 20454 3366
rect 20506 3314 33467 3366
rect 33519 3314 39936 3366
rect 960 3289 39936 3314
rect 13456 2725 13462 2737
rect 13417 2697 13462 2725
rect 13456 2685 13462 2697
rect 13514 2685 13520 2737
rect 14512 2685 14518 2737
rect 14570 2725 14576 2737
rect 14803 2728 14861 2734
rect 14803 2725 14815 2728
rect 14570 2697 14815 2725
rect 14570 2685 14576 2697
rect 14803 2694 14815 2697
rect 14849 2694 14861 2728
rect 14803 2688 14861 2694
rect 960 2552 39936 2577
rect 960 2500 13947 2552
rect 13999 2500 26960 2552
rect 27012 2500 39936 2552
rect 960 2475 39936 2500
rect 14512 1985 14518 1997
rect 10498 1957 14518 1985
rect 10498 1920 10526 1957
rect 14512 1945 14518 1957
rect 14570 1945 14576 1997
rect 10483 1914 10541 1920
rect 10483 1880 10495 1914
rect 10529 1880 10541 1914
rect 10483 1874 10541 1880
rect 13456 1871 13462 1923
rect 13514 1911 13520 1923
rect 36787 1914 36845 1920
rect 36787 1911 36799 1914
rect 13514 1883 36799 1911
rect 13514 1871 13520 1883
rect 36787 1880 36799 1883
rect 36833 1880 36845 1914
rect 36787 1874 36845 1880
rect 960 1738 39936 1763
rect 960 1686 7440 1738
rect 7492 1686 20454 1738
rect 20506 1686 33467 1738
rect 33519 1686 39936 1738
rect 960 1661 39936 1686
rect 880 1279 886 1331
rect 938 1319 944 1331
rect 10963 1322 11021 1328
rect 10963 1319 10975 1322
rect 938 1291 10975 1319
rect 938 1279 944 1291
rect 10963 1288 10975 1291
rect 11009 1288 11021 1322
rect 10963 1282 11021 1288
rect 784 1057 790 1109
rect 842 1097 848 1109
rect 37363 1100 37421 1106
rect 37363 1097 37375 1100
rect 842 1069 37375 1097
rect 842 1057 848 1069
rect 37363 1066 37375 1069
rect 37409 1066 37421 1100
rect 37363 1060 37421 1066
rect 960 924 39936 949
rect 960 872 13947 924
rect 13999 872 26960 924
rect 27012 872 39936 924
rect 960 847 39936 872
rect 960 110 39936 135
rect 960 58 7440 110
rect 7492 58 20454 110
rect 20506 58 33467 110
rect 33519 58 39936 110
rect 960 33 39936 58
<< via1 >>
rect 13947 4128 13999 4180
rect 26960 4128 27012 4180
rect 7440 3314 7492 3366
rect 20454 3314 20506 3366
rect 33467 3314 33519 3366
rect 13462 2728 13514 2737
rect 13462 2694 13471 2728
rect 13471 2694 13505 2728
rect 13505 2694 13514 2728
rect 13462 2685 13514 2694
rect 14518 2685 14570 2737
rect 13947 2500 13999 2552
rect 26960 2500 27012 2552
rect 14518 1945 14570 1997
rect 13462 1871 13514 1923
rect 7440 1686 7492 1738
rect 20454 1686 20506 1738
rect 33467 1686 33519 1738
rect 886 1279 938 1331
rect 790 1057 842 1109
rect 13947 872 13999 924
rect 26960 872 27012 924
rect 7440 58 7492 110
rect 20454 58 20506 110
rect 33467 58 33519 110
<< metal2 >>
rect 788 3812 844 3821
rect 788 3747 844 3756
rect 802 1115 830 3747
rect 7436 3704 7497 4205
rect 13943 4180 14003 4205
rect 7436 3648 7438 3704
rect 7494 3648 7497 3704
rect 7436 3366 7497 3648
rect 7436 3314 7440 3366
rect 7492 3314 7497 3366
rect 7436 2247 7497 3314
rect 7436 2191 7438 2247
rect 7494 2191 7497 2247
rect 7436 1738 7497 2191
rect 7436 1686 7440 1738
rect 7492 1686 7497 1738
rect 886 1331 938 1337
rect 886 1273 938 1279
rect 790 1109 842 1115
rect 790 1051 842 1057
rect 788 852 844 861
rect 898 838 926 1273
rect 844 810 926 838
rect 788 787 844 796
rect 7436 789 7497 1686
rect 7436 733 7438 789
rect 7494 733 7497 789
rect 7436 110 7497 733
rect 7436 58 7440 110
rect 7492 58 7497 110
rect 7836 2698 7897 4154
rect 7836 2642 7838 2698
rect 7894 2642 7897 2698
rect 7836 1240 7897 2642
rect 7836 1184 7838 1240
rect 7894 1184 7897 1240
rect 7836 84 7897 1184
rect 8236 3098 8297 4154
rect 8236 3042 8238 3098
rect 8294 3042 8297 3098
rect 8236 1640 8297 3042
rect 13943 4128 13947 4180
rect 13999 4128 14003 4180
rect 13943 2975 14003 4128
rect 13943 2919 13945 2975
rect 14001 2919 14003 2975
rect 13462 2737 13514 2743
rect 13462 2679 13514 2685
rect 13474 1929 13502 2679
rect 13943 2552 14003 2919
rect 13943 2500 13947 2552
rect 13999 2500 14003 2552
rect 13462 1923 13514 1929
rect 13462 1865 13514 1871
rect 8236 1584 8238 1640
rect 8294 1584 8297 1640
rect 8236 84 8297 1584
rect 13943 1518 14003 2500
rect 13943 1462 13945 1518
rect 14001 1462 14003 1518
rect 13943 924 14003 1462
rect 13943 872 13947 924
rect 13999 872 14003 924
rect 7436 33 7497 58
rect 13943 33 14003 872
rect 14343 3426 14403 4154
rect 14343 3370 14345 3426
rect 14401 3370 14403 3426
rect 14343 1969 14403 3370
rect 14743 3826 14803 4154
rect 14743 3770 14745 3826
rect 14801 3770 14803 3826
rect 14518 2737 14570 2743
rect 14518 2679 14570 2685
rect 14530 2003 14558 2679
rect 14743 2369 14803 3770
rect 14743 2313 14745 2369
rect 14801 2313 14803 2369
rect 14343 1913 14345 1969
rect 14401 1913 14403 1969
rect 14518 1997 14570 2003
rect 14518 1939 14570 1945
rect 14343 84 14403 1913
rect 14743 84 14803 2313
rect 20450 3704 20510 4205
rect 26956 4180 27017 4205
rect 20450 3648 20452 3704
rect 20508 3648 20510 3704
rect 20450 3366 20510 3648
rect 20450 3314 20454 3366
rect 20506 3314 20510 3366
rect 20450 2247 20510 3314
rect 20450 2191 20452 2247
rect 20508 2191 20510 2247
rect 20450 1738 20510 2191
rect 20450 1686 20454 1738
rect 20506 1686 20510 1738
rect 20450 789 20510 1686
rect 20450 733 20452 789
rect 20508 733 20510 789
rect 20450 110 20510 733
rect 20450 58 20454 110
rect 20506 58 20510 110
rect 20850 2698 20910 4154
rect 20850 2642 20852 2698
rect 20908 2642 20910 2698
rect 20850 1240 20910 2642
rect 20850 1184 20852 1240
rect 20908 1184 20910 1240
rect 20850 84 20910 1184
rect 21250 3098 21310 4154
rect 21250 3042 21252 3098
rect 21308 3042 21310 3098
rect 21250 1640 21310 3042
rect 21250 1584 21252 1640
rect 21308 1584 21310 1640
rect 21250 84 21310 1584
rect 26956 4128 26960 4180
rect 27012 4128 27017 4180
rect 26956 2975 27017 4128
rect 26956 2919 26958 2975
rect 27014 2919 27017 2975
rect 26956 2552 27017 2919
rect 26956 2500 26960 2552
rect 27012 2500 27017 2552
rect 26956 1518 27017 2500
rect 26956 1462 26958 1518
rect 27014 1462 27017 1518
rect 26956 924 27017 1462
rect 26956 872 26960 924
rect 27012 872 27017 924
rect 20450 33 20510 58
rect 26956 33 27017 872
rect 27356 3426 27417 4154
rect 27356 3370 27358 3426
rect 27414 3370 27417 3426
rect 27356 1969 27417 3370
rect 27356 1913 27358 1969
rect 27414 1913 27417 1969
rect 27356 84 27417 1913
rect 27756 3826 27817 4154
rect 27756 3770 27758 3826
rect 27814 3770 27817 3826
rect 27756 2369 27817 3770
rect 27756 2313 27758 2369
rect 27814 2313 27817 2369
rect 27756 84 27817 2313
rect 33463 3704 33523 4205
rect 33463 3648 33465 3704
rect 33521 3648 33523 3704
rect 33463 3366 33523 3648
rect 33463 3314 33467 3366
rect 33519 3314 33523 3366
rect 33463 2247 33523 3314
rect 33463 2191 33465 2247
rect 33521 2191 33523 2247
rect 33463 1738 33523 2191
rect 33463 1686 33467 1738
rect 33519 1686 33523 1738
rect 33463 789 33523 1686
rect 33463 733 33465 789
rect 33521 733 33523 789
rect 33463 110 33523 733
rect 33463 58 33467 110
rect 33519 58 33523 110
rect 33863 2698 33923 4154
rect 33863 2642 33865 2698
rect 33921 2642 33923 2698
rect 33863 1240 33923 2642
rect 33863 1184 33865 1240
rect 33921 1184 33923 1240
rect 33863 84 33923 1184
rect 34263 3098 34323 4154
rect 34263 3042 34265 3098
rect 34321 3042 34323 3098
rect 34263 1640 34323 3042
rect 34263 1584 34265 1640
rect 34321 1584 34323 1640
rect 34263 84 34323 1584
rect 33463 33 33523 58
<< via2 >>
rect 788 3756 844 3812
rect 7438 3648 7494 3704
rect 7438 2191 7494 2247
rect 788 796 844 852
rect 7438 733 7494 789
rect 7838 2642 7894 2698
rect 7838 1184 7894 1240
rect 8238 3042 8294 3098
rect 13945 2919 14001 2975
rect 8238 1584 8294 1640
rect 13945 1462 14001 1518
rect 14345 3370 14401 3426
rect 14745 3770 14801 3826
rect 14745 2313 14801 2369
rect 14345 1913 14401 1969
rect 20452 3648 20508 3704
rect 20452 2191 20508 2247
rect 20452 733 20508 789
rect 20852 2642 20908 2698
rect 20852 1184 20908 1240
rect 21252 3042 21308 3098
rect 21252 1584 21308 1640
rect 26958 2919 27014 2975
rect 26958 1462 27014 1518
rect 27358 3370 27414 3426
rect 27358 1913 27414 1969
rect 27758 3770 27814 3826
rect 27758 2313 27814 2369
rect 33465 3648 33521 3704
rect 33465 2191 33521 2247
rect 33465 733 33521 789
rect 33865 2642 33921 2698
rect 33865 1184 33921 1240
rect 34265 3042 34321 3098
rect 34265 1584 34321 1640
<< metal3 >>
rect 0 3817 800 3844
rect 14740 3829 14806 3831
rect 27753 3829 27819 3831
rect 960 3826 39936 3829
rect 0 3812 849 3817
rect 0 3756 788 3812
rect 844 3756 849 3812
rect 960 3770 14745 3826
rect 14801 3770 27758 3826
rect 27814 3770 39936 3826
rect 960 3768 39936 3770
rect 14740 3765 14806 3768
rect 27753 3765 27819 3768
rect 0 3751 849 3756
rect 0 3724 800 3751
rect 7433 3706 7499 3709
rect 20447 3706 20513 3709
rect 33460 3706 33526 3709
rect 960 3704 39936 3706
rect 960 3648 7438 3704
rect 7494 3648 20452 3704
rect 20508 3648 33465 3704
rect 33521 3648 39936 3704
rect 960 3646 39936 3648
rect 7433 3643 7499 3646
rect 20447 3643 20513 3646
rect 33460 3643 33526 3646
rect 14340 3429 14406 3431
rect 27353 3429 27419 3431
rect 960 3426 39936 3429
rect 960 3370 14345 3426
rect 14401 3370 27358 3426
rect 27414 3370 39936 3426
rect 960 3368 39936 3370
rect 14340 3365 14406 3368
rect 27353 3365 27419 3368
rect 8233 3100 8299 3103
rect 21247 3100 21313 3103
rect 34260 3100 34326 3103
rect 960 3098 39936 3100
rect 960 3042 8238 3098
rect 8294 3042 21252 3098
rect 21308 3042 34265 3098
rect 34321 3042 39936 3098
rect 960 3040 39936 3042
rect 8233 3037 8299 3040
rect 21247 3037 21313 3040
rect 34260 3037 34326 3040
rect 13940 2978 14006 2980
rect 26953 2978 27019 2980
rect 960 2975 39936 2978
rect 960 2919 13945 2975
rect 14001 2919 26958 2975
rect 27014 2919 39936 2975
rect 960 2917 39936 2919
rect 13940 2914 14006 2917
rect 26953 2914 27019 2917
rect 7833 2700 7899 2703
rect 20847 2700 20913 2703
rect 33860 2700 33926 2703
rect 960 2698 39936 2700
rect 960 2642 7838 2698
rect 7894 2642 20852 2698
rect 20908 2642 33865 2698
rect 33921 2642 39936 2698
rect 960 2640 39936 2642
rect 7833 2637 7899 2640
rect 20847 2637 20913 2640
rect 33860 2637 33926 2640
rect 14740 2371 14806 2374
rect 27753 2371 27819 2374
rect 960 2369 39936 2371
rect 960 2313 14745 2369
rect 14801 2313 27758 2369
rect 27814 2313 39936 2369
rect 960 2311 39936 2313
rect 14740 2308 14806 2311
rect 27753 2308 27819 2311
rect 7433 2249 7499 2252
rect 20447 2249 20513 2252
rect 33460 2249 33526 2252
rect 960 2247 39936 2249
rect 960 2191 7438 2247
rect 7494 2191 20452 2247
rect 20508 2191 33465 2247
rect 33521 2191 39936 2247
rect 960 2189 39936 2191
rect 7433 2186 7499 2189
rect 20447 2186 20513 2189
rect 33460 2186 33526 2189
rect 14340 1971 14406 1974
rect 27353 1971 27419 1974
rect 960 1969 39936 1971
rect 960 1913 14345 1969
rect 14401 1913 27358 1969
rect 27414 1913 39936 1969
rect 960 1911 39936 1913
rect 14340 1908 14406 1911
rect 27353 1908 27419 1911
rect 8233 1643 8299 1645
rect 21247 1643 21313 1645
rect 34260 1643 34326 1645
rect 960 1640 39936 1643
rect 960 1584 8238 1640
rect 8294 1584 21252 1640
rect 21308 1584 34265 1640
rect 34321 1584 39936 1640
rect 960 1582 39936 1584
rect 8233 1579 8299 1582
rect 21247 1579 21313 1582
rect 34260 1579 34326 1582
rect 13940 1520 14006 1523
rect 26953 1520 27019 1523
rect 960 1518 39936 1520
rect 960 1462 13945 1518
rect 14001 1462 26958 1518
rect 27014 1462 39936 1518
rect 960 1460 39936 1462
rect 13940 1457 14006 1460
rect 26953 1457 27019 1460
rect 7833 1243 7899 1245
rect 20847 1243 20913 1245
rect 33860 1243 33926 1245
rect 960 1240 39936 1243
rect 960 1184 7838 1240
rect 7894 1184 20852 1240
rect 20908 1184 33865 1240
rect 33921 1184 39936 1240
rect 960 1182 39936 1184
rect 7833 1179 7899 1182
rect 20847 1179 20913 1182
rect 33860 1179 33926 1182
rect 0 857 800 884
rect 0 852 849 857
rect 0 796 788 852
rect 844 796 849 852
rect 0 791 849 796
rect 7433 792 7499 794
rect 20447 792 20513 794
rect 33460 792 33526 794
rect 0 764 800 791
rect 960 789 39936 792
rect 960 733 7438 789
rect 7494 733 20452 789
rect 20508 733 33465 789
rect 33521 733 39936 789
rect 960 731 39936 733
rect 7433 728 7499 731
rect 20447 728 20513 731
rect 33460 728 33526 731
use sky130_fd_sc_hvl__decap_8  FILLER_3_388
timestamp 1607547389
transform 1 0 38208 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_396
timestamp 1607547389
transform 1 0 38976 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_2  FILLER_3_404
timestamp 1607547389
transform 1 0 39744 0 1 2526
box -66 -23 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_392
timestamp 1607547389
transform 1 0 38592 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_4_400
timestamp 1607547389
transform 1 0 39360 0 -1 4154
box -66 -23 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_4_404
timestamp 1607547389
transform 1 0 39744 0 -1 4154
box -66 -23 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_372
timestamp 1607547389
transform 1 0 36672 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_380
timestamp 1607547389
transform 1 0 37440 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_368
timestamp 1607547389
transform 1 0 36288 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_376
timestamp 1607547389
transform 1 0 37056 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_384
timestamp 1607547389
transform 1 0 37824 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_356
timestamp 1607547389
transform 1 0 35136 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_364
timestamp 1607547389
transform 1 0 35904 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_352
timestamp 1607547389
transform 1 0 34752 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_360
timestamp 1607547389
transform 1 0 35520 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_332
timestamp 1607547389
transform 1 0 32832 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_340
timestamp 1607547389
transform 1 0 33600 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_348
timestamp 1607547389
transform 1 0 34368 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_336
timestamp 1607547389
transform 1 0 33216 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_344
timestamp 1607547389
transform 1 0 33984 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_316
timestamp 1607547389
transform 1 0 31296 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_324
timestamp 1607547389
transform 1 0 32064 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_320
timestamp 1607547389
transform 1 0 31680 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_328
timestamp 1607547389
transform 1 0 32448 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_300
timestamp 1607547389
transform 1 0 29760 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_308
timestamp 1607547389
transform 1 0 30528 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_296
timestamp 1607547389
transform 1 0 29376 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_304
timestamp 1607547389
transform 1 0 30144 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_312
timestamp 1607547389
transform 1 0 30912 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_276
timestamp 1607547389
transform 1 0 27456 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_284
timestamp 1607547389
transform 1 0 28224 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_292
timestamp 1607547389
transform 1 0 28992 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_280
timestamp 1607547389
transform 1 0 27840 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_288
timestamp 1607547389
transform 1 0 28608 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_260
timestamp 1607547389
transform 1 0 25920 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_268
timestamp 1607547389
transform 1 0 26688 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_264
timestamp 1607547389
transform 1 0 26304 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_272
timestamp 1607547389
transform 1 0 27072 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_244
timestamp 1607547389
transform 1 0 24384 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_252
timestamp 1607547389
transform 1 0 25152 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_240
timestamp 1607547389
transform 1 0 24000 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_248
timestamp 1607547389
transform 1 0 24768 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_256
timestamp 1607547389
transform 1 0 25536 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_228
timestamp 1607547389
transform 1 0 22848 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_236
timestamp 1607547389
transform 1 0 23616 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_224
timestamp 1607547389
transform 1 0 22464 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_232
timestamp 1607547389
transform 1 0 23232 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_204
timestamp 1607547389
transform 1 0 20544 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_212
timestamp 1607547389
transform 1 0 21312 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_220
timestamp 1607547389
transform 1 0 22080 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_208
timestamp 1607547389
transform 1 0 20928 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_216
timestamp 1607547389
transform 1 0 21696 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_188
timestamp 1607547389
transform 1 0 19008 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_196
timestamp 1607547389
transform 1 0 19776 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_184
timestamp 1607547389
transform 1 0 18624 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_192
timestamp 1607547389
transform 1 0 19392 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_200
timestamp 1607547389
transform 1 0 20160 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_172
timestamp 1607547389
transform 1 0 17472 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_180
timestamp 1607547389
transform 1 0 18240 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_168
timestamp 1607547389
transform 1 0 17088 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_176
timestamp 1607547389
transform 1 0 17856 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_148
timestamp 1607547389
transform 1 0 15168 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_156
timestamp 1607547389
transform 1 0 15936 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_164
timestamp 1607547389
transform 1 0 16704 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_152
timestamp 1607547389
transform 1 0 15552 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_160
timestamp 1607547389
transform 1 0 16320 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__conb_1  mprj2_logic_high_hvl
timestamp 1607547389
transform 1 0 14688 0 1 2526
box -66 -23 546 897
use sky130_fd_sc_hvl__conb_1  mprj_logic_high_hvl
timestamp 1607547389
transform 1 0 13344 0 1 2526
box -66 -23 546 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_134
timestamp 1607547389
transform 1 0 13824 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_1  FILLER_3_142
timestamp 1607547389
transform 1 0 14592 0 1 2526
box -66 -23 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_136
timestamp 1607547389
transform 1 0 14016 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_144
timestamp 1607547389
transform 1 0 14784 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_112
timestamp 1607547389
transform 1 0 11712 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_120
timestamp 1607547389
transform 1 0 12480 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_1  FILLER_3_128
timestamp 1607547389
transform 1 0 13248 0 1 2526
box -66 -23 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_112
timestamp 1607547389
transform 1 0 11712 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_120
timestamp 1607547389
transform 1 0 12480 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_128
timestamp 1607547389
transform 1 0 13248 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_96
timestamp 1607547389
transform 1 0 10176 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_104
timestamp 1607547389
transform 1 0 10944 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_96
timestamp 1607547389
transform 1 0 10176 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_104
timestamp 1607547389
transform 1 0 10944 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_80
timestamp 1607547389
transform 1 0 8640 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_88
timestamp 1607547389
transform 1 0 9408 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_80
timestamp 1607547389
transform 1 0 8640 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_88
timestamp 1607547389
transform 1 0 9408 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_56
timestamp 1607547389
transform 1 0 6336 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_64
timestamp 1607547389
transform 1 0 7104 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_72
timestamp 1607547389
transform 1 0 7872 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_56
timestamp 1607547389
transform 1 0 6336 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_64
timestamp 1607547389
transform 1 0 7104 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_72
timestamp 1607547389
transform 1 0 7872 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_40
timestamp 1607547389
transform 1 0 4800 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_48
timestamp 1607547389
transform 1 0 5568 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_40
timestamp 1607547389
transform 1 0 4800 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_48
timestamp 1607547389
transform 1 0 5568 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_24
timestamp 1607547389
transform 1 0 3264 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_32
timestamp 1607547389
transform 1 0 4032 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_24
timestamp 1607547389
transform 1 0 3264 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_32
timestamp 1607547389
transform 1 0 4032 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_0
timestamp 1607547389
transform 1 0 960 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_8
timestamp 1607547389
transform 1 0 1728 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_16
timestamp 1607547389
transform 1 0 2496 0 1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_0
timestamp 1607547389
transform 1 0 960 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_8
timestamp 1607547389
transform 1 0 1728 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_16
timestamp 1607547389
transform 1 0 2496 0 -1 4154
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_405
timestamp 1607547389
transform 1 0 39840 0 1 898
box -66 -23 162 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_405
timestamp 1607547389
transform 1 0 39840 0 -1 2526
box -66 -23 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_392
timestamp 1607547389
transform 1 0 38592 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_400
timestamp 1607547389
transform 1 0 39360 0 -1 898
box -66 -23 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_0_404
timestamp 1607547389
transform 1 0 39744 0 -1 898
box -66 -23 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_389
timestamp 1607547389
transform 1 0 38304 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_397
timestamp 1607547389
transform 1 0 39072 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_389
timestamp 1607547389
transform 1 0 38304 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_397
timestamp 1607547389
transform 1 0 39072 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  mprj_logic_high_lv
timestamp 1607547389
transform 1 0 36672 0 1 898
box -66 -23 1698 1651
use sky130_fd_sc_hvl__decap_8  FILLER_0_368
timestamp 1607547389
transform 1 0 36288 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_376
timestamp 1607547389
transform 1 0 37056 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_384
timestamp 1607547389
transform 1 0 37824 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_2  FILLER_1_370
timestamp 1607547389
transform 1 0 36480 0 1 898
box -66 -23 258 897
use sky130_fd_sc_hvl__fill_2  FILLER_2_370
timestamp 1607547389
transform 1 0 36480 0 -1 2526
box -66 -23 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_352
timestamp 1607547389
transform 1 0 34752 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_360
timestamp 1607547389
transform 1 0 35520 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_354
timestamp 1607547389
transform 1 0 34944 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_362
timestamp 1607547389
transform 1 0 35712 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_354
timestamp 1607547389
transform 1 0 34944 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_362
timestamp 1607547389
transform 1 0 35712 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_336
timestamp 1607547389
transform 1 0 33216 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_344
timestamp 1607547389
transform 1 0 33984 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_338
timestamp 1607547389
transform 1 0 33408 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_346
timestamp 1607547389
transform 1 0 34176 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_338
timestamp 1607547389
transform 1 0 33408 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_346
timestamp 1607547389
transform 1 0 34176 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_320
timestamp 1607547389
transform 1 0 31680 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_328
timestamp 1607547389
transform 1 0 32448 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_314
timestamp 1607547389
transform 1 0 31104 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_322
timestamp 1607547389
transform 1 0 31872 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_330
timestamp 1607547389
transform 1 0 32640 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_314
timestamp 1607547389
transform 1 0 31104 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_322
timestamp 1607547389
transform 1 0 31872 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_330
timestamp 1607547389
transform 1 0 32640 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_296
timestamp 1607547389
transform 1 0 29376 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_304
timestamp 1607547389
transform 1 0 30144 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_312
timestamp 1607547389
transform 1 0 30912 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_298
timestamp 1607547389
transform 1 0 29568 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_306
timestamp 1607547389
transform 1 0 30336 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_298
timestamp 1607547389
transform 1 0 29568 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_306
timestamp 1607547389
transform 1 0 30336 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_280
timestamp 1607547389
transform 1 0 27840 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_288
timestamp 1607547389
transform 1 0 28608 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_282
timestamp 1607547389
transform 1 0 28032 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_290
timestamp 1607547389
transform 1 0 28800 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_282
timestamp 1607547389
transform 1 0 28032 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_290
timestamp 1607547389
transform 1 0 28800 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_264
timestamp 1607547389
transform 1 0 26304 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_272
timestamp 1607547389
transform 1 0 27072 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_258
timestamp 1607547389
transform 1 0 25728 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_266
timestamp 1607547389
transform 1 0 26496 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_274
timestamp 1607547389
transform 1 0 27264 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_258
timestamp 1607547389
transform 1 0 25728 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_266
timestamp 1607547389
transform 1 0 26496 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_274
timestamp 1607547389
transform 1 0 27264 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_240
timestamp 1607547389
transform 1 0 24000 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_248
timestamp 1607547389
transform 1 0 24768 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_256
timestamp 1607547389
transform 1 0 25536 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_242
timestamp 1607547389
transform 1 0 24192 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_250
timestamp 1607547389
transform 1 0 24960 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_242
timestamp 1607547389
transform 1 0 24192 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_250
timestamp 1607547389
transform 1 0 24960 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_224
timestamp 1607547389
transform 1 0 22464 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_232
timestamp 1607547389
transform 1 0 23232 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_226
timestamp 1607547389
transform 1 0 22656 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_234
timestamp 1607547389
transform 1 0 23424 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_226
timestamp 1607547389
transform 1 0 22656 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_234
timestamp 1607547389
transform 1 0 23424 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_208
timestamp 1607547389
transform 1 0 20928 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_216
timestamp 1607547389
transform 1 0 21696 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_210
timestamp 1607547389
transform 1 0 21120 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_218
timestamp 1607547389
transform 1 0 21888 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_210
timestamp 1607547389
transform 1 0 21120 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_218
timestamp 1607547389
transform 1 0 21888 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_184
timestamp 1607547389
transform 1 0 18624 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_192
timestamp 1607547389
transform 1 0 19392 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_200
timestamp 1607547389
transform 1 0 20160 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_186
timestamp 1607547389
transform 1 0 18816 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_194
timestamp 1607547389
transform 1 0 19584 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_202
timestamp 1607547389
transform 1 0 20352 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_186
timestamp 1607547389
transform 1 0 18816 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_194
timestamp 1607547389
transform 1 0 19584 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_202
timestamp 1607547389
transform 1 0 20352 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_168
timestamp 1607547389
transform 1 0 17088 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_176
timestamp 1607547389
transform 1 0 17856 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_170
timestamp 1607547389
transform 1 0 17280 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_178
timestamp 1607547389
transform 1 0 18048 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_170
timestamp 1607547389
transform 1 0 17280 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_178
timestamp 1607547389
transform 1 0 18048 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_152
timestamp 1607547389
transform 1 0 15552 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_160
timestamp 1607547389
transform 1 0 16320 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_154
timestamp 1607547389
transform 1 0 15744 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_162
timestamp 1607547389
transform 1 0 16512 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_154
timestamp 1607547389
transform 1 0 15744 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_162
timestamp 1607547389
transform 1 0 16512 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_136
timestamp 1607547389
transform 1 0 14016 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_144
timestamp 1607547389
transform 1 0 14784 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_130
timestamp 1607547389
transform 1 0 13440 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_138
timestamp 1607547389
transform 1 0 14208 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_146
timestamp 1607547389
transform 1 0 14976 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_130
timestamp 1607547389
transform 1 0 13440 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_138
timestamp 1607547389
transform 1 0 14208 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_146
timestamp 1607547389
transform 1 0 14976 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_112
timestamp 1607547389
transform 1 0 11712 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_120
timestamp 1607547389
transform 1 0 12480 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_128
timestamp 1607547389
transform 1 0 13248 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_114
timestamp 1607547389
transform 1 0 11904 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_122
timestamp 1607547389
transform 1 0 12672 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_114
timestamp 1607547389
transform 1 0 11904 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_122
timestamp 1607547389
transform 1 0 12672 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  mprj2_logic_high_lv
timestamp 1607547389
transform 1 0 10272 0 1 898
box -66 -23 1698 1651
use sky130_fd_sc_hvl__decap_8  FILLER_0_96
timestamp 1607547389
transform 1 0 10176 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_104
timestamp 1607547389
transform 1 0 10944 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_96
timestamp 1607547389
transform 1 0 10176 0 1 898
box -66 -23 162 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_96
timestamp 1607547389
transform 1 0 10176 0 -1 2526
box -66 -23 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_80
timestamp 1607547389
transform 1 0 8640 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_88
timestamp 1607547389
transform 1 0 9408 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_80
timestamp 1607547389
transform 1 0 8640 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_88
timestamp 1607547389
transform 1 0 9408 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_80
timestamp 1607547389
transform 1 0 8640 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_88
timestamp 1607547389
transform 1 0 9408 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_56
timestamp 1607547389
transform 1 0 6336 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_64
timestamp 1607547389
transform 1 0 7104 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_72
timestamp 1607547389
transform 1 0 7872 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_56
timestamp 1607547389
transform 1 0 6336 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_64
timestamp 1607547389
transform 1 0 7104 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_72
timestamp 1607547389
transform 1 0 7872 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_56
timestamp 1607547389
transform 1 0 6336 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_64
timestamp 1607547389
transform 1 0 7104 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_72
timestamp 1607547389
transform 1 0 7872 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_40
timestamp 1607547389
transform 1 0 4800 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_48
timestamp 1607547389
transform 1 0 5568 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_40
timestamp 1607547389
transform 1 0 4800 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_48
timestamp 1607547389
transform 1 0 5568 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_40
timestamp 1607547389
transform 1 0 4800 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_48
timestamp 1607547389
transform 1 0 5568 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_24
timestamp 1607547389
transform 1 0 3264 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_32
timestamp 1607547389
transform 1 0 4032 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_24
timestamp 1607547389
transform 1 0 3264 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_32
timestamp 1607547389
transform 1 0 4032 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_24
timestamp 1607547389
transform 1 0 3264 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_32
timestamp 1607547389
transform 1 0 4032 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_0
timestamp 1607547389
transform 1 0 960 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_8
timestamp 1607547389
transform 1 0 1728 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_16
timestamp 1607547389
transform 1 0 2496 0 -1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_0
timestamp 1607547389
transform 1 0 960 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_8
timestamp 1607547389
transform 1 0 1728 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_16
timestamp 1607547389
transform 1 0 2496 0 1 898
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_0
timestamp 1607547389
transform 1 0 960 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_8
timestamp 1607547389
transform 1 0 1728 0 -1 2526
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_16
timestamp 1607547389
transform 1 0 2496 0 -1 2526
box -66 -23 834 897
<< labels >>
rlabel metal3 s 0 764 800 884 4 mprj2_vdd_logic1
port 1 nsew
rlabel metal3 s 0 3724 800 3844 4 mprj_vdd_logic1
port 2 nsew
rlabel metal2 s 33463 33 33523 4205 4 vccd
port 3 nsew
rlabel metal2 s 20450 33 20510 4205 4 vccd
port 3 nsew
rlabel metal2 s 7437 33 7497 4205 4 vccd
port 3 nsew
rlabel metal3 s 960 3646 39936 3706 4 vccd
port 3 nsew
rlabel metal3 s 960 2189 39936 2249 4 vccd
port 3 nsew
rlabel metal3 s 960 732 39936 792 4 vccd
port 3 nsew
rlabel metal2 s 26957 33 27017 4205 4 vssd
port 4 nsew
rlabel metal2 s 13943 33 14003 4205 4 vssd
port 4 nsew
rlabel metal3 s 960 2918 39936 2978 4 vssd
port 4 nsew
rlabel metal3 s 960 1460 39936 1520 4 vssd
port 4 nsew
rlabel metal2 s 33863 84 33923 4154 4 vdda1
port 5 nsew
rlabel metal2 s 20850 84 20910 4154 4 vdda1
port 5 nsew
rlabel metal2 s 7837 84 7897 4154 4 vdda1
port 5 nsew
rlabel metal3 s 960 2640 39936 2700 4 vdda1
port 5 nsew
rlabel metal3 s 960 1183 39936 1243 4 vdda1
port 5 nsew
rlabel metal2 s 27357 84 27417 4154 4 vssa1
port 6 nsew
rlabel metal2 s 14343 84 14403 4154 4 vssa1
port 6 nsew
rlabel metal3 s 960 3369 39936 3429 4 vssa1
port 6 nsew
rlabel metal3 s 960 1911 39936 1971 4 vssa1
port 6 nsew
rlabel metal2 s 34263 84 34323 4154 4 vdda2
port 7 nsew
rlabel metal2 s 21250 84 21310 4154 4 vdda2
port 7 nsew
rlabel metal2 s 8237 84 8297 4154 4 vdda2
port 7 nsew
rlabel metal3 s 960 3040 39936 3100 4 vdda2
port 7 nsew
rlabel metal3 s 960 1583 39936 1643 4 vdda2
port 7 nsew
rlabel metal2 s 27757 84 27817 4154 4 vssa2
port 8 nsew
rlabel metal2 s 14743 84 14803 4154 4 vssa2
port 8 nsew
rlabel metal3 s 960 3769 39936 3829 4 vssa2
port 8 nsew
rlabel metal3 s 960 2311 39936 2371 4 vssa2
port 8 nsew
<< properties >>
string FIXED_BBOX 0 1 40002 4205
<< end >>
