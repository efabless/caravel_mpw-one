magic
tech sky130A
magscale 12 1
timestamp 1598768719
<< metal5 >>
rect 0 100 35 105
rect 0 95 40 100
rect 0 85 45 95
rect 0 70 15 85
rect 30 70 45 85
rect 0 60 45 70
rect 0 55 40 60
rect 0 50 35 55
rect 0 35 30 50
rect 0 30 35 35
rect 0 25 40 30
rect 0 15 45 25
rect 0 0 15 15
rect 30 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
