magic
tech sky130A
magscale 1 2
timestamp 1602626460
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_61 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602619247
transform 0 -1 39547 -1 0 78134
box -143 -543 16134 39593
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602619247
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_0
timestamp 1602619247
transform -1 0 73400 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_1
timestamp 1602619247
transform -1 0 124200 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_2
timestamp 1602619247
transform -1 0 175000 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_4
timestamp 1602619247
transform -1 0 276600 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_3
timestamp 1602619247
transform -1 0 225800 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_5
timestamp 1602619247
transform -1 0 327400 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_6
timestamp 1602619247
transform -1 0 378200 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_7
timestamp 1602619247
transform -1 0 429000 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_8
timestamp 1602619247
transform -1 0 479800 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_21
timestamp 1602619247
transform 0 1 600058 1 0 54143
box -143 -543 16134 39593
use sky130_fd_io__corner_bus_overlay  sky130_fd_io__corner_bus_overlay_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602619247
transform 0 1 599792 -1 0 40000
box 0 0 40000 40733
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_9
timestamp 1602619247
transform -1 0 530600 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_10
timestamp 1602619247
transform -1 0 581400 0 -1 39593
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_60
timestamp 1602619247
transform 0 -1 39547 -1 0 175734
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_59
timestamp 1602619247
transform 0 -1 39547 -1 0 126934
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_19
timestamp 1602619247
transform 0 1 600058 1 0 102943
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_18
timestamp 1602619247
transform 0 1 600058 1 0 200543
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_20
timestamp 1602619247
transform 0 1 600058 1 0 151743
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_53
timestamp 1602619247
transform 0 -1 39547 -1 0 273334
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_54
timestamp 1602619247
transform 0 -1 39547 -1 0 224534
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_17
timestamp 1602619247
transform 0 1 600058 1 0 298143
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_16
timestamp 1602619247
transform 0 1 600058 1 0 249343
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_55
timestamp 1602619247
transform 0 -1 39547 -1 0 322134
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_56
timestamp 1602619247
transform 0 -1 39547 -1 0 419734
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_57
timestamp 1602619247
transform 0 -1 39547 -1 0 370934
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_14
timestamp 1602619247
transform 0 1 600058 1 0 395743
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_15
timestamp 1602619247
transform 0 1 600058 1 0 346943
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_48
timestamp 1602619247
transform 0 -1 39547 -1 0 523534
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_58
timestamp 1602619247
transform 0 -1 39547 -1 0 468534
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_13
timestamp 1602619247
transform 0 1 600058 1 0 493343
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_12
timestamp 1602619247
transform 0 1 600058 1 0 444543
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_49
timestamp 1602619247
transform 0 -1 39547 -1 0 572334
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_50
timestamp 1602619247
transform 0 -1 39547 -1 0 619134
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_11
timestamp 1602619247
transform 0 1 600058 1 0 542143
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_22
timestamp 1602619247
transform 0 1 600058 1 0 595143
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_51
timestamp 1602619247
transform 0 -1 39547 -1 0 716734
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_52
timestamp 1602619247
transform 0 -1 39547 -1 0 667934
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_24
timestamp 1602619247
transform 0 1 600058 1 0 692743
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_23
timestamp 1602619247
transform 0 1 600058 1 0 643943
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_43
timestamp 1602619247
transform 0 -1 39547 -1 0 765534
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_42
timestamp 1602619247
transform 0 -1 39547 -1 0 814334
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_25
timestamp 1602619247
transform 0 1 600058 1 0 741543
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_31
timestamp 1602619247
transform 0 1 600058 1 0 790343
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_46
timestamp 1602619247
transform 0 -1 39547 -1 0 911934
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_44
timestamp 1602619247
transform 0 -1 39547 -1 0 863134
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_29
timestamp 1602619247
transform 0 1 600058 1 0 887943
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_32
timestamp 1602619247
transform 0 1 600058 1 0 839143
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_47
timestamp 1602619247
transform 0 -1 39547 -1 0 1006534
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_45
timestamp 1602619247
transform 0 -1 39547 -1 0 960734
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_27
timestamp 1602619247
transform 0 1 600058 1 0 985543
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_30
timestamp 1602619247
transform 0 1 600058 1 0 936743
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_41
timestamp 1602619247
transform 1 0 58205 0 1 1023084
box -143 -543 16134 39593
use sky130_fd_io__corner_bus_overlay  sky130_fd_io__corner_bus_overlay_1
timestamp 1602619247
transform 0 -1 39813 1 0 1022677
box 0 0 40000 40733
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_39
timestamp 1602619247
transform 1 0 159805 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_40
timestamp 1602619247
transform 1 0 109005 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_38
timestamp 1602619247
transform 1 0 210605 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_37
timestamp 1602619247
transform 1 0 261405 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_35
timestamp 1602619247
transform 1 0 363005 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_36
timestamp 1602619247
transform 1 0 312205 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_34
timestamp 1602619247
transform 1 0 413805 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_33
timestamp 1602619247
transform 1 0 464605 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_28
timestamp 1602619247
transform 1 0 515405 0 1 1023084
box -143 -543 16134 39593
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_1
timestamp 1602619247
transform 1 0 599605 0 1 1021877
box 0 0 40000 40800
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_26
timestamp 1602619247
transform 1 0 566205 0 1 1023084
box -143 -543 16134 39593
use bump_pad  bump_pad_3
array 0 1 100000 0 1 100000
timestamp 1602626256
transform 1 0 468644 0 1 471210
box -24800 -24800 25000 24800
use bump_pad  bump_pad_2
array 0 1 100000 0 1 100000
timestamp 1602626256
transform 1 0 68644 0 1 471210
box -24800 -24800 25000 24800
use bump_pad  bump_pad_1
array 0 5 100000 0 3 100000
timestamp 1602626256
transform 1 0 68644 0 1 671210
box -24800 -24800 25000 24800
use bump_pad  bump_pad_0
array 0 5 100000 0 3 100000
timestamp 1602626256
transform 1 0 68644 0 1 71210
box -24800 -24800 25000 24800
<< end >>
