magic
tech sky130A
magscale 1 2
timestamp 1621450687
<< viali >>
rect 1133 425 1167 459
<< metal1 >>
rect 0 1114 1564 1136
rect 0 1062 174 1114
rect 226 1062 574 1114
rect 626 1062 974 1114
rect 1026 1062 1374 1114
rect 1426 1062 1564 1114
rect 0 1040 1564 1062
rect 0 570 1564 592
rect 0 518 374 570
rect 426 518 774 570
rect 826 518 1174 570
rect 1226 518 1564 570
rect 0 496 1564 518
rect 14 416 20 468
rect 72 456 78 468
rect 1121 459 1179 465
rect 1121 456 1133 459
rect 72 428 1133 456
rect 72 416 78 428
rect 1121 425 1133 428
rect 1167 425 1179 459
rect 1121 419 1179 425
rect 0 26 1564 48
rect 0 -26 174 26
rect 226 -26 574 26
rect 626 -26 974 26
rect 1026 -26 1374 26
rect 1426 -26 1564 26
rect 0 -48 1564 -26
<< via1 >>
rect 174 1062 226 1114
rect 574 1062 626 1114
rect 974 1062 1026 1114
rect 1374 1062 1426 1114
rect 374 518 426 570
rect 774 518 826 570
rect 1174 518 1226 570
rect 20 416 72 468
rect 174 -26 226 26
rect 574 -26 626 26
rect 974 -26 1026 26
rect 1374 -26 1426 26
<< metal2 >>
rect 160 1114 240 1136
rect 160 1080 174 1114
rect 226 1080 240 1114
rect 160 1024 172 1080
rect 228 1024 240 1080
rect 18 912 74 921
rect 18 847 74 856
rect 32 474 60 847
rect 20 468 72 474
rect 20 410 72 416
rect 160 180 240 1024
rect 160 124 172 180
rect 228 124 240 180
rect 160 26 240 124
rect 160 -26 174 26
rect 226 -26 240 26
rect 160 -48 240 -26
rect 360 630 440 1136
rect 360 574 372 630
rect 428 574 440 630
rect 360 570 440 574
rect 360 518 374 570
rect 426 518 440 570
rect 360 -48 440 518
rect 560 1114 640 1136
rect 560 1080 574 1114
rect 626 1080 640 1114
rect 560 1024 572 1080
rect 628 1024 640 1080
rect 560 180 640 1024
rect 560 124 572 180
rect 628 124 640 180
rect 560 26 640 124
rect 560 -26 574 26
rect 626 -26 640 26
rect 560 -48 640 -26
rect 760 630 840 1136
rect 760 574 772 630
rect 828 574 840 630
rect 760 570 840 574
rect 760 518 774 570
rect 826 518 840 570
rect 760 -48 840 518
rect 960 1114 1040 1136
rect 960 1080 974 1114
rect 1026 1080 1040 1114
rect 960 1024 972 1080
rect 1028 1024 1040 1080
rect 960 180 1040 1024
rect 960 124 972 180
rect 1028 124 1040 180
rect 960 26 1040 124
rect 960 -26 974 26
rect 1026 -26 1040 26
rect 960 -48 1040 -26
rect 1160 630 1240 1136
rect 1160 574 1172 630
rect 1228 574 1240 630
rect 1160 570 1240 574
rect 1160 518 1174 570
rect 1226 518 1240 570
rect 1160 -48 1240 518
rect 1360 1114 1440 1136
rect 1360 1080 1374 1114
rect 1426 1080 1440 1114
rect 1360 1024 1372 1080
rect 1428 1024 1440 1080
rect 1360 180 1440 1024
rect 1360 124 1372 180
rect 1428 124 1440 180
rect 1360 26 1440 124
rect 1360 -26 1374 26
rect 1426 -26 1440 26
rect 1360 -48 1440 -26
<< via2 >>
rect 172 1062 174 1080
rect 174 1062 226 1080
rect 226 1062 228 1080
rect 172 1024 228 1062
rect 18 856 74 912
rect 172 124 228 180
rect 372 574 428 630
rect 572 1062 574 1080
rect 574 1062 626 1080
rect 626 1062 628 1080
rect 572 1024 628 1062
rect 572 124 628 180
rect 772 574 828 630
rect 972 1062 974 1080
rect 974 1062 1026 1080
rect 1026 1062 1028 1080
rect 972 1024 1028 1062
rect 972 124 1028 180
rect 1172 574 1228 630
rect 1372 1062 1374 1080
rect 1374 1062 1426 1080
rect 1426 1062 1428 1080
rect 1372 1024 1428 1062
rect 1372 124 1428 180
<< metal3 >>
rect 0 1080 1564 1092
rect 0 1024 172 1080
rect 228 1024 572 1080
rect 628 1024 972 1080
rect 1028 1024 1372 1080
rect 1428 1024 1564 1080
rect 0 1012 1564 1024
rect 13 914 79 917
rect 800 914 1600 944
rect 13 912 1600 914
rect 13 856 18 912
rect 74 856 1600 912
rect 13 854 1600 856
rect 13 851 79 854
rect 800 824 1600 854
rect 0 630 1564 642
rect 0 574 372 630
rect 428 574 772 630
rect 828 574 1172 630
rect 1228 574 1564 630
rect 0 562 1564 574
rect 0 180 1564 192
rect 0 124 172 180
rect 228 124 572 180
rect 628 124 972 180
rect 1028 124 1372 180
rect 1428 124 1564 180
rect 0 112 1564 124
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 0 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1618914159
transform 1 0 0 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 276 0 -1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1618914159
transform 1 0 276 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  gpio_logic_high $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform -1 0 1196 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 828 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_5
timestamp 1618914159
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 1196 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 920 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618914159
transform -1 0 1564 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618914159
transform -1 0 1564 0 1 544
box -38 -48 314 592
<< labels >>
rlabel metal3 s 800 824 1600 944 6 gpio_logic1
port 0 nsew signal tristate
rlabel metal2 s 1360 -48 1440 1136 6 vccd1
port 1 nsew power bidirectional
rlabel metal2 s 960 -48 1040 1136 6 vccd1
port 2 nsew power bidirectional
rlabel metal2 s 560 -48 640 1136 6 vccd1
port 3 nsew power bidirectional
rlabel metal2 s 160 -48 240 1136 6 vccd1
port 4 nsew power bidirectional
rlabel metal3 s 0 1012 1564 1092 6 vccd1
port 5 nsew power bidirectional
rlabel metal3 s 0 112 1564 192 6 vccd1
port 6 nsew power bidirectional
rlabel metal2 s 1160 -48 1240 1136 6 vssd1
port 7 nsew ground bidirectional
rlabel metal2 s 760 -48 840 1136 6 vssd1
port 8 nsew ground bidirectional
rlabel metal2 s 360 -48 440 1136 6 vssd1
port 9 nsew ground bidirectional
rlabel metal3 s 0 562 1564 642 6 vssd1
port 10 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1600 1600
<< end >>
