magic
tech sky130A
magscale 12 1
timestamp 1598768325
<< metal5 >>
rect 10 100 35 105
rect 5 95 40 100
rect 0 85 45 95
rect 0 35 15 85
rect 30 35 45 85
rect 0 10 45 35
rect 5 5 45 10
rect 10 0 45 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
