magic
tech sky130A
magscale 12 1
timestamp 1598766505
<< metal5 >>
rect 0 90 15 105
rect 60 90 75 105
rect 0 75 30 90
rect 45 75 75 90
rect 0 60 75 75
rect 0 0 15 60
rect 30 45 45 60
rect 60 0 75 60
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
