magic
tech sky130A
magscale 12 1
timestamp 1598765560
<< metal5 >>
rect 0 60 15 105
rect 30 60 45 105
rect 0 45 45 60
rect 0 0 15 45
rect 30 0 45 45
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
