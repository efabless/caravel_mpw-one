magic
tech sky130A
timestamp 1584566829
use seal_ring_corner_abstract seal_ring_corner_abstract_0
timestamp 1584566221
transform 1 0 0 0 1 0
box 0 0 160716 265712
use seal_ring_corner_abstract seal_ring_corner_abstract_3
timestamp 1584566221
transform -1 0 321432 0 1 0
box 0 0 160716 265712
use seal_ring_corner_abstract seal_ring_corner_abstract_1
timestamp 1584566221
transform 1 0 0 0 -1 531424
box 0 0 160716 265712
use seal_ring_corner_abstract seal_ring_corner_abstract_2
timestamp 1584566221
transform -1 0 321432 0 -1 531424
box 0 0 160716 265712
<< properties >>
string LEFview no_prefix
string GDS_FILE advSeal_6um_gen.gds
string GDS_START 0
string FIXED_BBOX 0 0 321432 531424
<< end >>
