magic
tech sky130A
magscale 1 2
timestamp 1622497372
<< viali >>
rect 16773 221 16807 255
<< metal1 >>
rect 0 1114 19964 1136
rect 0 1062 174 1114
rect 226 1062 8174 1114
rect 8226 1062 16174 1114
rect 16226 1062 19964 1114
rect 0 1040 19964 1062
rect 0 570 19964 592
rect 0 518 4174 570
rect 4226 518 12174 570
rect 12226 518 19964 570
rect 0 496 19964 518
rect 16758 252 16764 264
rect 16719 224 16764 252
rect 16758 212 16764 224
rect 16816 212 16822 264
rect 0 26 19964 48
rect 0 -26 174 26
rect 226 -26 8174 26
rect 8226 -26 16174 26
rect 16226 -26 19964 26
rect 0 -48 19964 -26
<< via1 >>
rect 174 1062 226 1114
rect 8174 1062 8226 1114
rect 16174 1062 16226 1114
rect 4174 518 4226 570
rect 12174 518 12226 570
rect 16764 255 16816 264
rect 16764 221 16773 255
rect 16773 221 16807 255
rect 16807 221 16816 255
rect 16764 212 16816 221
rect 174 -26 226 26
rect 8174 -26 8226 26
rect 16174 -26 16226 26
<< metal2 >>
rect 170 1114 230 1136
rect 170 1062 174 1114
rect 226 1062 230 1114
rect 170 380 230 1062
rect 4170 940 4230 1136
rect 4170 884 4172 940
rect 4228 884 4230 940
rect 3146 776 3202 785
rect 3146 711 3202 720
rect 170 324 172 380
rect 228 324 230 380
rect 170 26 230 324
rect 3160 241 3188 711
rect 4170 570 4230 884
rect 4170 518 4174 570
rect 4226 518 4230 570
rect 3146 232 3202 241
rect 3146 167 3202 176
rect 170 -26 174 26
rect 226 -26 230 26
rect 170 -48 230 -26
rect 4170 -48 4230 518
rect 8170 1114 8230 1136
rect 8170 1062 8174 1114
rect 8226 1062 8230 1114
rect 8170 380 8230 1062
rect 8170 324 8172 380
rect 8228 324 8230 380
rect 8170 26 8230 324
rect 8170 -26 8174 26
rect 8226 -26 8230 26
rect 8170 -48 8230 -26
rect 12170 940 12230 1136
rect 12170 884 12172 940
rect 12228 884 12230 940
rect 12170 570 12230 884
rect 12170 518 12174 570
rect 12226 518 12230 570
rect 12170 -48 12230 518
rect 16170 1114 16230 1136
rect 16170 1062 16174 1114
rect 16226 1062 16230 1114
rect 16170 380 16230 1062
rect 16170 324 16172 380
rect 16228 324 16230 380
rect 16170 26 16230 324
rect 16764 264 16816 270
rect 16762 232 16764 241
rect 16816 232 16818 241
rect 16762 167 16818 176
rect 16170 -26 16174 26
rect 16226 -26 16230 26
rect 16170 -48 16230 -26
<< via2 >>
rect 4172 884 4228 940
rect 3146 720 3202 776
rect 172 324 228 380
rect 3146 176 3202 232
rect 8172 324 8228 380
rect 12172 884 12228 940
rect 16172 324 16228 380
rect 16762 212 16764 232
rect 16764 212 16816 232
rect 16816 212 16818 232
rect 16762 176 16818 212
<< metal3 >>
rect 4167 942 4233 945
rect 12167 942 12233 945
rect 0 940 19964 942
rect 0 884 4172 940
rect 4228 884 12172 940
rect 12228 884 19964 940
rect 0 882 19964 884
rect 4167 879 4233 882
rect 12167 879 12233 882
rect 0 778 800 808
rect 3141 778 3207 781
rect 0 776 3207 778
rect 0 720 3146 776
rect 3202 720 3207 776
rect 0 718 3207 720
rect 0 688 800 718
rect 3141 715 3207 718
rect 167 382 233 385
rect 8167 382 8233 385
rect 16167 382 16233 385
rect 0 380 19964 382
rect 0 324 172 380
rect 228 324 8172 380
rect 8228 324 16172 380
rect 16228 324 19964 380
rect 0 322 19964 324
rect 167 319 233 322
rect 8167 319 8233 322
rect 16167 319 16233 322
rect 3141 234 3207 237
rect 16757 234 16823 237
rect 3141 232 16823 234
rect 3141 176 3146 232
rect 3202 176 16762 232
rect 16818 176 16823 232
rect 3141 174 16823 176
rect 3141 171 3207 174
rect 16757 171 16823 174
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 0 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1618914159
transform 1 0 0 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 276 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1618914159
transform 1 0 276 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1618914159
transform 1 0 1380 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1618914159
transform 1 0 1380 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 2668 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_11
timestamp 1618914159
transform 1 0 2668 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 2484 0 -1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1618914159
transform 1 0 2760 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1618914159
transform 1 0 2484 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 1618914159
transform 1 0 2760 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1618914159
transform 1 0 3864 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 1618914159
transform 1 0 3864 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_5
timestamp 1618914159
transform 1 0 5336 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_12
timestamp 1618914159
transform 1 0 5336 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 4968 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1618914159
transform 1 0 5428 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_54
timestamp 1618914159
transform 1 0 4968 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_59
timestamp 1618914159
transform 1 0 5428 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1618914159
transform 1 0 6532 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_71
timestamp 1618914159
transform 1 0 6532 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_6
timestamp 1618914159
transform 1 0 8004 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_13
timestamp 1618914159
transform 1 0 8004 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1618914159
transform 1 0 7636 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1618914159
transform 1 0 8096 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1618914159
transform 1 0 7636 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_88
timestamp 1618914159
transform 1 0 8096 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1618914159
transform 1 0 9200 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_100
timestamp 1618914159
transform 1 0 9200 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1618914159
transform 1 0 10304 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_112
timestamp 1618914159
transform 1 0 10304 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_7
timestamp 1618914159
transform 1 0 10672 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_14
timestamp 1618914159
transform 1 0 10672 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1618914159
transform 1 0 10764 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1618914159
transform 1 0 10764 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_129
timestamp 1618914159
transform 1 0 11868 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1618914159
transform 1 0 12972 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1618914159
transform 1 0 11868 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1618914159
transform 1 0 12972 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_8
timestamp 1618914159
transform 1 0 13340 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_15
timestamp 1618914159
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1618914159
transform 1 0 13432 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_146
timestamp 1618914159
transform 1 0 13432 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_158
timestamp 1618914159
transform 1 0 14536 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_158
timestamp 1618914159
transform 1 0 14536 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_9
timestamp 1618914159
transform 1 0 16008 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16
timestamp 1618914159
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1618914159
transform 1 0 15640 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_175 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 16100 0 -1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_170
timestamp 1618914159
transform 1 0 15640 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_175
timestamp 1618914159
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  inst $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 16744 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_181 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 16652 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_185
timestamp 1618914159
transform 1 0 17020 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_187
timestamp 1618914159
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_10
timestamp 1618914159
transform 1 0 18676 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1618914159
transform 1 0 18676 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1618914159
transform 1 0 18124 0 -1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 18768 0 -1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1618914159
transform 1 0 18308 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_204
timestamp 1618914159
transform 1 0 18768 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618914159
transform -1 0 19964 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618914159
transform -1 0 19964 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_212
timestamp 1618914159
transform 1 0 19504 0 -1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_212
timestamp 1618914159
transform 1 0 19504 0 1 544
box -38 -48 222 592
<< labels >>
rlabel metal3 s 0 688 800 808 6 HI
port 0 nsew signal tristate
rlabel metal2 s 16170 -48 16230 1136 6 vccd2
port 1 nsew power bidirectional
rlabel metal2 s 8170 -48 8230 1136 6 vccd2
port 2 nsew power bidirectional
rlabel metal2 s 170 -48 230 1136 6 vccd2
port 3 nsew power bidirectional
rlabel metal3 s 0 322 19964 382 6 vccd2
port 4 nsew power bidirectional
rlabel metal2 s 12170 -48 12230 1136 6 vssd2
port 5 nsew ground bidirectional
rlabel metal2 s 4170 -48 4230 1136 6 vssd2
port 6 nsew ground bidirectional
rlabel metal3 s 0 882 19964 942 6 vssd2
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 1400
<< end >>
