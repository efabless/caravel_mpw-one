* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 VPWR VGND
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[1] la_data_in_mprj[20]
+ la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23] la_data_in_mprj[24]
+ la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27] la_data_in_mprj[28]
+ la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31] la_data_in_mprj[32]
+ la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35] la_data_in_mprj[36]
+ la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39] la_data_in_mprj[3] la_data_in_mprj[40]
+ la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43] la_data_in_mprj[44]
+ la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47] la_data_in_mprj[48]
+ la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51] la_data_in_mprj[52]
+ la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55] la_data_in_mprj[56]
+ la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59] la_data_in_mprj[5] la_data_in_mprj[60]
+ la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63] la_data_in_mprj[64]
+ la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67] la_data_in_mprj[68]
+ la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71] la_data_in_mprj[72]
+ la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75] la_data_in_mprj[76]
+ la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79] la_data_in_mprj[7] la_data_in_mprj[80]
+ la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83] la_data_in_mprj[84]
+ la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87] la_data_in_mprj[88]
+ la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91] la_data_in_mprj[92]
+ la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95] la_data_in_mprj[96]
+ la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99] la_data_in_mprj[9] la_data_out_core[0]
+ la_data_out_core[100] la_data_out_core[101] la_data_out_core[102] la_data_out_core[103]
+ la_data_out_core[104] la_data_out_core[105] la_data_out_core[106] la_data_out_core[107]
+ la_data_out_core[108] la_data_out_core[109] la_data_out_core[10] la_data_out_core[110]
+ la_data_out_core[111] la_data_out_core[112] la_data_out_core[113] la_data_out_core[114]
+ la_data_out_core[115] la_data_out_core[116] la_data_out_core[117] la_data_out_core[118]
+ la_data_out_core[119] la_data_out_core[11] la_data_out_core[120] la_data_out_core[121]
+ la_data_out_core[122] la_data_out_core[123] la_data_out_core[124] la_data_out_core[125]
+ la_data_out_core[126] la_data_out_core[127] la_data_out_core[12] la_data_out_core[13]
+ la_data_out_core[14] la_data_out_core[15] la_data_out_core[16] la_data_out_core[17]
+ la_data_out_core[18] la_data_out_core[19] la_data_out_core[1] la_data_out_core[20]
+ la_data_out_core[21] la_data_out_core[22] la_data_out_core[23] la_data_out_core[24]
+ la_data_out_core[25] la_data_out_core[26] la_data_out_core[27] la_data_out_core[28]
+ la_data_out_core[29] la_data_out_core[2] la_data_out_core[30] la_data_out_core[31]
+ la_data_out_core[32] la_data_out_core[33] la_data_out_core[34] la_data_out_core[35]
+ la_data_out_core[36] la_data_out_core[37] la_data_out_core[38] la_data_out_core[39]
+ la_data_out_core[3] la_data_out_core[40] la_data_out_core[41] la_data_out_core[42]
+ la_data_out_core[43] la_data_out_core[44] la_data_out_core[45] la_data_out_core[46]
+ la_data_out_core[47] la_data_out_core[48] la_data_out_core[49] la_data_out_core[4]
+ la_data_out_core[50] la_data_out_core[51] la_data_out_core[52] la_data_out_core[53]
+ la_data_out_core[54] la_data_out_core[55] la_data_out_core[56] la_data_out_core[57]
+ la_data_out_core[58] la_data_out_core[59] la_data_out_core[5] la_data_out_core[60]
+ la_data_out_core[61] la_data_out_core[62] la_data_out_core[63] la_data_out_core[64]
+ la_data_out_core[65] la_data_out_core[66] la_data_out_core[67] la_data_out_core[68]
+ la_data_out_core[69] la_data_out_core[6] la_data_out_core[70] la_data_out_core[71]
+ la_data_out_core[72] la_data_out_core[73] la_data_out_core[74] la_data_out_core[75]
+ la_data_out_core[76] la_data_out_core[77] la_data_out_core[78] la_data_out_core[79]
+ la_data_out_core[7] la_data_out_core[80] la_data_out_core[81] la_data_out_core[82]
+ la_data_out_core[83] la_data_out_core[84] la_data_out_core[85] la_data_out_core[86]
+ la_data_out_core[87] la_data_out_core[88] la_data_out_core[89] la_data_out_core[8]
+ la_data_out_core[90] la_data_out_core[91] la_data_out_core[92] la_data_out_core[93]
+ la_data_out_core[94] la_data_out_core[95] la_data_out_core[96] la_data_out_core[97]
+ la_data_out_core[98] la_data_out_core[99] la_data_out_core[9] la_data_out_mprj[0]
+ la_data_out_mprj[100] la_data_out_mprj[101] la_data_out_mprj[102] la_data_out_mprj[103]
+ la_data_out_mprj[104] la_data_out_mprj[105] la_data_out_mprj[106] la_data_out_mprj[107]
+ la_data_out_mprj[108] la_data_out_mprj[109] la_data_out_mprj[10] la_data_out_mprj[110]
+ la_data_out_mprj[111] la_data_out_mprj[112] la_data_out_mprj[113] la_data_out_mprj[114]
+ la_data_out_mprj[115] la_data_out_mprj[116] la_data_out_mprj[117] la_data_out_mprj[118]
+ la_data_out_mprj[119] la_data_out_mprj[11] la_data_out_mprj[120] la_data_out_mprj[121]
+ la_data_out_mprj[122] la_data_out_mprj[123] la_data_out_mprj[124] la_data_out_mprj[125]
+ la_data_out_mprj[126] la_data_out_mprj[127] la_data_out_mprj[12] la_data_out_mprj[13]
+ la_data_out_mprj[14] la_data_out_mprj[15] la_data_out_mprj[16] la_data_out_mprj[17]
+ la_data_out_mprj[18] la_data_out_mprj[19] la_data_out_mprj[1] la_data_out_mprj[20]
+ la_data_out_mprj[21] la_data_out_mprj[22] la_data_out_mprj[23] la_data_out_mprj[24]
+ la_data_out_mprj[25] la_data_out_mprj[26] la_data_out_mprj[27] la_data_out_mprj[28]
+ la_data_out_mprj[29] la_data_out_mprj[2] la_data_out_mprj[30] la_data_out_mprj[31]
+ la_data_out_mprj[32] la_data_out_mprj[33] la_data_out_mprj[34] la_data_out_mprj[35]
+ la_data_out_mprj[36] la_data_out_mprj[37] la_data_out_mprj[38] la_data_out_mprj[39]
+ la_data_out_mprj[3] la_data_out_mprj[40] la_data_out_mprj[42] la_data_out_mprj[43]
+ la_data_out_mprj[44] la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47]
+ la_data_out_mprj[48] la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50]
+ la_data_out_mprj[51] la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54]
+ la_data_out_mprj[55] la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58]
+ la_data_out_mprj[59] la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61]
+ la_data_out_mprj[62] la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65]
+ la_data_out_mprj[66] la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69]
+ la_data_out_mprj[6] la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72]
+ la_data_out_mprj[73] la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76]
+ la_data_out_mprj[77] la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7]
+ la_data_out_mprj[80] la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83]
+ la_data_out_mprj[84] la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87]
+ la_data_out_mprj[88] la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90]
+ la_data_out_mprj[91] la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94]
+ la_data_out_mprj[95] la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98]
+ la_data_out_mprj[99] la_data_out_mprj[9] la_oen_core[0] la_oen_core[100] la_oen_core[101]
+ la_oen_core[102] la_oen_core[103] la_oen_core[104] la_oen_core[105] la_oen_core[106]
+ la_oen_core[107] la_oen_core[108] la_oen_core[109] la_oen_core[10] la_oen_core[110]
+ la_oen_core[111] la_oen_core[112] la_oen_core[113] la_oen_core[114] la_oen_core[115]
+ la_oen_core[116] la_oen_core[117] la_oen_core[118] la_oen_core[119] la_oen_core[11]
+ la_oen_core[120] la_oen_core[121] la_oen_core[122] la_oen_core[123] la_oen_core[124]
+ la_oen_core[125] la_oen_core[126] la_oen_core[127] la_oen_core[12] la_oen_core[13]
+ la_oen_core[14] la_oen_core[15] la_oen_core[16] la_oen_core[17] la_oen_core[18]
+ la_oen_core[19] la_oen_core[1] la_oen_core[20] la_oen_core[21] la_oen_core[22] la_oen_core[23]
+ la_oen_core[24] la_oen_core[25] la_oen_core[26] la_oen_core[27] la_oen_core[28]
+ la_oen_core[29] la_oen_core[2] la_oen_core[30] la_oen_core[31] la_oen_core[32] la_oen_core[33]
+ la_oen_core[34] la_oen_core[35] la_oen_core[36] la_oen_core[37] la_oen_core[38]
+ la_oen_core[39] la_oen_core[3] la_oen_core[40] la_oen_core[41] la_oen_core[42] la_oen_core[43]
+ la_oen_core[44] la_oen_core[45] la_oen_core[46] la_oen_core[47] la_oen_core[48]
+ la_oen_core[49] la_oen_core[4] la_oen_core[50] la_oen_core[51] la_oen_core[52] la_oen_core[53]
+ la_oen_core[54] la_oen_core[55] la_oen_core[56] la_oen_core[57] la_oen_core[58]
+ la_oen_core[59] la_oen_core[5] la_oen_core[60] la_oen_core[61] la_oen_core[62] la_oen_core[63]
+ la_oen_core[64] la_oen_core[65] la_oen_core[66] la_oen_core[67] la_oen_core[68]
+ la_oen_core[69] la_oen_core[6] la_oen_core[70] la_oen_core[71] la_oen_core[72] la_oen_core[73]
+ la_oen_core[74] la_oen_core[75] la_oen_core[76] la_oen_core[77] la_oen_core[78]
+ la_oen_core[79] la_oen_core[7] la_oen_core[80] la_oen_core[81] la_oen_core[82] la_oen_core[83]
+ la_oen_core[84] la_oen_core[85] la_oen_core[86] la_oen_core[87] la_oen_core[88]
+ la_oen_core[89] la_oen_core[8] la_oen_core[90] la_oen_core[91] la_oen_core[92] la_oen_core[93]
+ la_oen_core[94] la_oen_core[95] la_oen_core[96] la_oen_core[97] la_oen_core[98]
+ la_oen_core[99] la_oen_core[9] la_oen_mprj[0] la_oen_mprj[100] la_oen_mprj[101]
+ la_oen_mprj[102] la_oen_mprj[103] la_oen_mprj[104] la_oen_mprj[105] la_oen_mprj[106]
+ la_oen_mprj[107] la_oen_mprj[108] la_oen_mprj[109] la_oen_mprj[10] la_oen_mprj[110]
+ la_oen_mprj[111] la_oen_mprj[112] la_oen_mprj[113] la_oen_mprj[114] la_oen_mprj[115]
+ la_oen_mprj[116] la_oen_mprj[117] la_oen_mprj[118] la_oen_mprj[119] la_oen_mprj[11]
+ la_oen_mprj[120] la_oen_mprj[121] la_oen_mprj[122] la_oen_mprj[123] la_oen_mprj[124]
+ la_oen_mprj[125] la_oen_mprj[126] la_oen_mprj[127] la_oen_mprj[12] la_oen_mprj[13]
+ la_oen_mprj[14] la_oen_mprj[15] la_oen_mprj[16] la_oen_mprj[17] la_oen_mprj[18]
+ la_oen_mprj[19] la_oen_mprj[1] la_oen_mprj[20] la_oen_mprj[21] la_oen_mprj[22] la_oen_mprj[23]
+ la_oen_mprj[24] la_oen_mprj[25] la_oen_mprj[26] la_oen_mprj[27] la_oen_mprj[28]
+ la_oen_mprj[29] la_oen_mprj[2] la_oen_mprj[30] la_oen_mprj[31] la_oen_mprj[32] la_oen_mprj[33]
+ la_oen_mprj[34] la_oen_mprj[35] la_oen_mprj[36] la_oen_mprj[37] la_oen_mprj[38]
+ la_oen_mprj[39] la_oen_mprj[3] la_oen_mprj[40] la_oen_mprj[41] la_oen_mprj[42] la_oen_mprj[43]
+ la_oen_mprj[44] la_oen_mprj[45] la_oen_mprj[46] la_oen_mprj[47] la_oen_mprj[48]
+ la_oen_mprj[49] la_oen_mprj[4] la_oen_mprj[50] la_oen_mprj[51] la_oen_mprj[52] la_oen_mprj[53]
+ la_oen_mprj[54] la_oen_mprj[55] la_oen_mprj[56] la_oen_mprj[57] la_oen_mprj[58]
+ la_oen_mprj[59] la_oen_mprj[5] la_oen_mprj[60] la_oen_mprj[61] la_oen_mprj[62] la_oen_mprj[63]
+ la_oen_mprj[64] la_oen_mprj[65] la_oen_mprj[66] la_oen_mprj[67] la_oen_mprj[68]
+ la_oen_mprj[69] la_oen_mprj[6] la_oen_mprj[70] la_oen_mprj[71] la_oen_mprj[72] la_oen_mprj[73]
+ la_oen_mprj[74] la_oen_mprj[75] la_oen_mprj[76] la_oen_mprj[77] la_oen_mprj[78]
+ la_oen_mprj[79] la_oen_mprj[7] la_oen_mprj[80] la_oen_mprj[81] la_oen_mprj[82] la_oen_mprj[84]
+ la_oen_mprj[85] la_oen_mprj[86] la_oen_mprj[87] la_oen_mprj[88] la_oen_mprj[89]
+ la_oen_mprj[8] la_oen_mprj[90] la_oen_mprj[91] la_oen_mprj[92] la_oen_mprj[93] la_oen_mprj[94]
+ la_oen_mprj[95] la_oen_mprj[96] la_oen_mprj[97] la_oen_mprj[98] la_oen_mprj[99]
+ la_oen_mprj[9] mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12]
+ mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16]
+ mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20]
+ mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24]
+ mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28]
+ mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3]
+ mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8]
+ mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12]
+ mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16]
+ mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20]
+ mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24]
+ mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28]
+ mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3]
+ mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8]
+ mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_o_core[0] mprj_dat_o_core[10]
+ mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14]
+ mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18]
+ mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22]
+ mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26]
+ mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30]
+ mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6]
+ mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10]
+ mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14]
+ mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18]
+ mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22]
+ mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26]
+ mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30]
+ mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6]
+ mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_sel_o_core[0] mprj_sel_o_core[1]
+ mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2]
+ mprj_sel_o_user[3] mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user
+ user1_vcc_powergood user1_vdd_powergood user2_vcc_powergood user2_vdd_powergood
+ user_clock user_clock2 user_reset user_resetn VPWR VGND
XFILLER_3_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[299\] VGND VGND VPWR VPWR mprj_logic_high\[299\]/HI mprj_logic_high\[299\]/LO
+ sky130_fd_sc_hd__conb_1
X_501_ la_data_out_mprj[30] VGND VGND VPWR VPWR _501_/Y sky130_fd_sc_hd__inv_2
X_432_ mprj_adr_o_core[25] VGND VGND VPWR VPWR _432_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_363_ la_oen_mprj[95] VGND VGND VPWR VPWR _363_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[36\] _507_/Y la_buf\[36\]/TE VGND VGND VPWR VPWR la_data_in_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_6_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] mprj_logic_high\[355\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[25\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[76\] _344_/Y mprj_logic_high\[278\]/HI VGND VGND VPWR VPWR
+ la_oen_core[76] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[214\] VGND VGND VPWR VPWR mprj_logic_high\[214\]/HI mprj_logic_high\[214\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[24\] _463_/Y mprj_dat_buf\[24\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_20_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high\[306\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_415_ mprj_adr_o_core[8] VGND VGND VPWR VPWR _415_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_346_ la_oen_mprj[78] VGND VGND VPWR VPWR _346_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high\[329\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[75\] VGND VGND VPWR VPWR la_buf\[1\]/TE mprj_logic_high\[75\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[164\] VGND VGND VPWR VPWR la_buf\[90\]/TE mprj_logic_high\[164\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[331\] VGND VGND VPWR VPWR mprj_logic_high\[331\]/HI mprj_logic_high\[331\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[429\] VGND VGND VPWR VPWR mprj_logic_high\[429\]/HI mprj_logic_high\[429\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[41\]_TE la_buf\[41\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[26\]_TE mprj_logic_high\[228\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] mprj_logic_high\[422\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[92\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[64\]_TE la_buf\[64\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high\[251\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[109\] _377_/Y mprj_logic_high\[311\]/HI VGND VGND VPWR
+ VPWR la_oen_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_18_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[39\] _638_/Y mprj_logic_high\[241\]/HI VGND VGND VPWR VPWR
+ la_oen_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_16_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[281\] VGND VGND VPWR VPWR mprj_logic_high\[281\]/HI mprj_logic_high\[281\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[379\] VGND VGND VPWR VPWR mprj_logic_high\[379\]/HI mprj_logic_high\[379\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[13\]_TE mprj_dat_buf\[13\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__402__A mprj_we_o_core VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y VGND VGND VPWR VPWR la_data_in_mprj[62]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[87\]_TE la_buf\[87\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[38\] VGND VGND VPWR VPWR mprj_adr_buf\[28\]/TE mprj_logic_high\[38\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[127\] VGND VGND VPWR VPWR la_buf\[53\]/TE mprj_logic_high\[127\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_594_ la_data_out_mprj[123] VGND VGND VPWR VPWR _594_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xla_buf\[66\] _537_/Y la_buf\[66\]/TE VGND VGND VPWR VPWR la_data_in_core[66] sky130_fd_sc_hd__einvp_8
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[122\] _593_/Y la_buf\[122\]/TE VGND VGND VPWR VPWR la_data_in_core[122] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[70\]_B mprj_logic_high\[400\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] mprj_logic_high\[385\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[55\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[61\]_B mprj_logic_high\[391\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[244\] VGND VGND VPWR VPWR mprj_logic_high\[244\]/HI mprj_logic_high\[244\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[52\]_B mprj_logic_high\[382\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[411\] VGND VGND VPWR VPWR mprj_logic_high\[411\]/HI mprj_logic_high\[411\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_646_ la_oen_mprj[47] VGND VGND VPWR VPWR _646_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_577_ la_data_out_mprj[106] VGND VGND VPWR VPWR _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[6\]_A _445_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y VGND VGND VPWR VPWR la_data_in_mprj[25]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[43\]_B mprj_logic_high\[373\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[112\]_TE la_buf\[112\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[27\]_TE mprj_adr_buf\[27\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[95\]_A user_to_mprj_in_gates\[95\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[34\]_B mprj_logic_high\[364\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__500__A la_data_out_mprj[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_500_ la_data_out_mprj[29] VGND VGND VPWR VPWR _500_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_431_ mprj_adr_o_core[24] VGND VGND VPWR VPWR _431_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[194\] VGND VGND VPWR VPWR la_buf\[120\]/TE mprj_logic_high\[194\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[3\] _602_/Y mprj_logic_high\[205\]/HI VGND VGND VPWR VPWR
+ la_oen_core[3] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[21\] _620_/Y mprj_logic_high\[223\]/HI VGND VGND VPWR VPWR
+ la_oen_core[21] sky130_fd_sc_hd__einvp_8
X_362_ la_oen_mprj[94] VGND VGND VPWR VPWR _362_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[361\] VGND VGND VPWR VPWR mprj_logic_high\[361\]/HI mprj_logic_high\[361\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[122\]_A _593_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[29\] _500_/Y la_buf\[29\]/TE VGND VGND VPWR VPWR la_data_in_core[29] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[86\]_A user_to_mprj_in_gates\[86\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_B mprj_logic_high\[355\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__410__A mprj_adr_o_core[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[10\]_A user_to_mprj_in_gates\[10\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_629_ la_oen_mprj[30] VGND VGND VPWR VPWR _629_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[124\]_A user_to_mprj_in_gates\[124\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] mprj_logic_high\[348\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[18\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[113\]_A _584_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[77\]_A user_to_mprj_in_gates\[77\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[16\]_B mprj_logic_high\[346\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[50\]_A _521_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_B mprj_logic_high\[430\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high\[284\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[115\]_A user_to_mprj_in_gates\[115\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[104\]_A _575_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[68\]_A user_to_mprj_in_gates\[68\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[41\]_A _512_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[20\] VGND VGND VPWR VPWR mprj_adr_buf\[10\]/TE mprj_logic_high\[20\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[69\] _337_/Y mprj_logic_high\[271\]/HI VGND VGND VPWR VPWR
+ la_oen_core[69] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[17\] _456_/Y mprj_dat_buf\[17\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[17]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[207\] VGND VGND VPWR VPWR mprj_logic_high\[207\]/HI mprj_logic_high\[207\]/LO
+ sky130_fd_sc_hd__conb_1
X_414_ mprj_adr_o_core[7] VGND VGND VPWR VPWR _414_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[106\]_A user_to_mprj_in_gates\[106\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_345_ la_oen_mprj[77] VGND VGND VPWR VPWR _345_/Y sky130_fd_sc_hd__inv_2
XANTENNA__405__A mprj_sel_o_core[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[59\]_A user_to_mprj_in_gates\[59\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[32\]_A _503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[12\] _419_/Y mprj_adr_buf\[12\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[12]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[126] sky130_fd_sc_hd__inv_8
XFILLER_2_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y VGND VGND VPWR VPWR la_data_in_mprj[92]
+ sky130_fd_sc_hd__inv_8
XFILLER_2_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[99\]_A _570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[23\]_A _494_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[68\] VGND VGND VPWR VPWR mprj_dat_buf\[26\]/TE mprj_logic_high\[68\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[157\] VGND VGND VPWR VPWR la_buf\[83\]/TE mprj_logic_high\[157\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[14\]_A _485_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[324\] VGND VGND VPWR VPWR mprj_logic_high\[324\]/HI mprj_logic_high\[324\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[96\] _567_/Y la_buf\[96\]/TE VGND VGND VPWR VPWR la_data_in_core[96] sky130_fd_sc_hd__einvp_8
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] mprj_logic_high\[415\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[85\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[92\]_A _360_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[274\] VGND VGND VPWR VPWR mprj_logic_high\[274\]/HI mprj_logic_high\[274\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[83\]_A _351_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[441\] VGND VGND VPWR VPWR mprj_logic_high\[441\]/HI mprj_logic_high\[441\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[7\] _478_/Y la_buf\[7\]/TE VGND VGND VPWR VPWR la_data_in_core[7] sky130_fd_sc_hd__einvp_8
Xla_buf\[11\] _482_/Y la_buf\[11\]/TE VGND VGND VPWR VPWR la_data_in_core[11] sky130_fd_sc_hd__einvp_8
XFILLER_3_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[4\] _411_/Y mprj_adr_buf\[4\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y VGND VGND VPWR VPWR la_data_in_mprj[55]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high\[319\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[74\]_A _342_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] mprj_logic_high\[441\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[111\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[31\]_TE la_buf\[31\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[65\]_A _333_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high\[218\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__503__A la_data_out_mprj[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[121\] _389_/Y mprj_logic_high\[323\]/HI VGND VGND VPWR
+ VPWR la_oen_core[121] sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[2\] _405_/Y mprj_sel_buf\[2\]/TE VGND VGND VPWR VPWR mprj_sel_o_user[2]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[51\] _650_/Y mprj_logic_high\[253\]/HI VGND VGND VPWR VPWR
+ la_oen_core[51] sky130_fd_sc_hd__einvp_8
XFILLER_5_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[391\] VGND VGND VPWR VPWR mprj_logic_high\[391\]/HI mprj_logic_high\[391\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_593_ la_data_out_mprj[122] VGND VGND VPWR VPWR _593_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[59\] _530_/Y la_buf\[59\]/TE VGND VGND VPWR VPWR la_data_in_core[59] sky130_fd_sc_hd__einvp_8
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[56\]_A _655_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__413__A mprj_adr_o_core[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[115\] _586_/Y la_buf\[115\]/TE VGND VGND VPWR VPWR la_data_in_core[115] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[54\]_TE la_buf\[54\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] mprj_logic_high\[378\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[48\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[39\]_TE mprj_logic_high\[241\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[47\]_A _646_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[38\]_A _637_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[50\] VGND VGND VPWR VPWR mprj_dat_buf\[8\]/TE mprj_logic_high\[50\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[99\] _367_/Y mprj_logic_high\[301\]/HI VGND VGND VPWR VPWR
+ la_oen_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_5_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[237\] VGND VGND VPWR VPWR mprj_logic_high\[237\]/HI mprj_logic_high\[237\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[404\] VGND VGND VPWR VPWR mprj_logic_high\[404\]/HI mprj_logic_high\[404\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj2_vdd_pwrgood mprj2_pwrgood/A VGND VGND VPWR VPWR user2_vdd_powergood sky130_fd_sc_hd__buf_8
XANTENNA_la_buf\[77\]_TE la_buf\[77\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_645_ la_oen_mprj[46] VGND VGND VPWR VPWR _645_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_576_ la_data_out_mprj[105] VGND VGND VPWR VPWR _576_/Y sky130_fd_sc_hd__inv_2
XANTENNA__408__A mprj_adr_o_core[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[29\]_A _628_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y VGND VGND VPWR VPWR la_data_in_mprj[18]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[25\]_A _432_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[26\]_TE mprj_dat_buf\[26\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[5\]_TE mprj_logic_high\[207\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[2\]_A _601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_A _423_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[98\] VGND VGND VPWR VPWR la_buf\[24\]/TE mprj_logic_high\[98\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_430_ mprj_adr_o_core[23] VGND VGND VPWR VPWR _430_/Y sky130_fd_sc_hd__inv_2
X_361_ la_oen_mprj[93] VGND VGND VPWR VPWR _361_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[187\] VGND VGND VPWR VPWR la_buf\[113\]/TE mprj_logic_high\[187\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[14\] _613_/Y mprj_logic_high\[216\]/HI VGND VGND VPWR VPWR
+ la_oen_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_14_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[354\] VGND VGND VPWR VPWR mprj_logic_high\[354\]/HI mprj_logic_high\[354\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_628_ la_oen_mprj[29] VGND VGND VPWR VPWR _628_/Y sky130_fd_sc_hd__inv_2
X_559_ la_data_out_mprj[88] VGND VGND VPWR VPWR _559_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__601__A la_oen_mprj[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[13\] VGND VGND VPWR VPWR mprj_adr_buf\[3\]/TE mprj_logic_high\[13\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__511__A la_data_out_mprj[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[102\] VGND VGND VPWR VPWR la_buf\[28\]/TE mprj_logic_high\[102\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_413_ mprj_adr_o_core[6] VGND VGND VPWR VPWR _413_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[41\] _512_/Y la_buf\[41\]/TE VGND VGND VPWR VPWR la_data_in_core[41] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[102\]_TE la_buf\[102\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_344_ la_oen_mprj[76] VGND VGND VPWR VPWR _344_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[17\]_TE mprj_adr_buf\[17\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__421__A mprj_adr_o_core[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[119] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[29\]_A _468_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y VGND VGND VPWR VPWR la_data_in_mprj[85]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] mprj_logic_high\[360\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[30\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[1\]_A _408_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__331__A la_oen_mprj[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[5\]_TE mprj_dat_buf\[5\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_TE la_buf\[125\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__506__A la_data_out_mprj[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[81\] _349_/Y mprj_logic_high\[283\]/HI VGND VGND VPWR VPWR
+ la_oen_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_3_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[317\] VGND VGND VPWR VPWR mprj_logic_high\[317\]/HI mprj_logic_high\[317\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xla_buf\[89\] _560_/Y la_buf\[89\]/TE VGND VGND VPWR VPWR la_data_in_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[72\]_TE mprj_logic_high\[274\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__416__A mprj_adr_o_core[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] mprj_logic_high\[408\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[78\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj2_pwrgood_A mprj2_pwrgood/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high\[297\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[80\] VGND VGND VPWR VPWR la_buf\[6\]/TE mprj_logic_high\[80\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[267\] VGND VGND VPWR VPWR mprj_logic_high\[267\]/HI mprj_logic_high\[267\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[434\] VGND VGND VPWR VPWR mprj_logic_high\[434\]/HI mprj_logic_high\[434\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[7\]_A _478_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y VGND VGND VPWR VPWR la_data_in_mprj[48]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] mprj_logic_high\[434\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[104\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[1\]_B mprj_logic_high\[331\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[114\] _382_/Y mprj_logic_high\[316\]/HI VGND VGND VPWR
+ VPWR la_oen_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_0_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[44\] _643_/Y mprj_logic_high\[246\]/HI VGND VGND VPWR VPWR
+ la_oen_core[44] sky130_fd_sc_hd__einvp_8
X_592_ la_data_out_mprj[121] VGND VGND VPWR VPWR _592_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[384\] VGND VGND VPWR VPWR mprj_logic_high\[384\]/HI mprj_logic_high\[384\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[108\] _579_/Y la_buf\[108\]/TE VGND VGND VPWR VPWR la_data_in_core[108] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[101] sky130_fd_sc_hd__inv_8
XFILLER_0_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[5\]_A user_to_mprj_in_gates\[5\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__604__A la_oen_mprj[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[0\] _439_/Y mprj_dat_buf\[0\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__514__A la_data_out_mprj[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[43\] VGND VGND VPWR VPWR mprj_dat_buf\[1\]/TE mprj_logic_high\[43\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[132\] VGND VGND VPWR VPWR la_buf\[58\]/TE mprj_logic_high\[132\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[107\]_TE mprj_logic_high\[309\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_644_ la_oen_mprj[45] VGND VGND VPWR VPWR _644_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[71\] _542_/Y la_buf\[71\]/TE VGND VGND VPWR VPWR la_data_in_core[71] sky130_fd_sc_hd__einvp_8
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_575_ la_data_out_mprj[104] VGND VGND VPWR VPWR _575_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__424__A mprj_adr_o_core[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[21\]_TE la_buf\[21\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] mprj_logic_high\[390\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[60\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__334__A la_oen_mprj[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__509__A la_data_out_mprj[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_360_ la_oen_mprj[92] VGND VGND VPWR VPWR _360_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[347\] VGND VGND VPWR VPWR mprj_logic_high\[347\]/HI mprj_logic_high\[347\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[44\]_TE la_buf\[44\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high\[231\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_627_ la_oen_mprj[28] VGND VGND VPWR VPWR _627_/Y sky130_fd_sc_hd__inv_2
XANTENNA__419__A mprj_adr_o_core[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_558_ la_data_out_mprj[87] VGND VGND VPWR VPWR _558_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y VGND VGND VPWR VPWR la_data_in_mprj[30]
+ sky130_fd_sc_hd__inv_8
X_489_ la_data_out_mprj[18] VGND VGND VPWR VPWR _489_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[8\] VGND VGND VPWR VPWR mprj_sel_buf\[2\]/TE mprj_logic_high\[8\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[67\]_TE la_buf\[67\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[297\] VGND VGND VPWR VPWR mprj_logic_high\[297\]/HI mprj_logic_high\[297\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_412_ mprj_adr_o_core[5] VGND VGND VPWR VPWR _412_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ la_oen_mprj[75] VGND VGND VPWR VPWR _343_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[34\] _505_/Y la_buf\[34\]/TE VGND VGND VPWR VPWR la_data_in_core[34] sky130_fd_sc_hd__einvp_8
XFILLER_6_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y VGND VGND VPWR VPWR la_data_in_mprj[78]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] mprj_logic_high\[353\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[23\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__612__A la_oen_mprj[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__522__A la_data_out_mprj[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[74\] _342_/Y mprj_logic_high\[276\]/HI VGND VGND VPWR VPWR
+ la_oen_core[74] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[212\] VGND VGND VPWR VPWR mprj_logic_high\[212\]/HI mprj_logic_high\[212\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[22\] _461_/Y mprj_dat_buf\[22\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__432__A mprj_adr_o_core[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__607__A la_oen_mprj[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[91\]_B mprj_logic_high\[421\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__342__A la_oen_mprj[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__517__A la_data_out_mprj[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[73\] VGND VGND VPWR VPWR mprj_dat_buf\[31\]/TE mprj_logic_high\[73\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[162\] VGND VGND VPWR VPWR la_buf\[88\]/TE mprj_logic_high\[162\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[82\]_B mprj_logic_high\[412\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[427\] VGND VGND VPWR VPWR mprj_logic_high\[427\]/HI mprj_logic_high\[427\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__427__A mprj_adr_o_core[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[73\]_B mprj_logic_high\[403\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] mprj_logic_high\[420\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[90\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[115\]_TE la_buf\[115\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__337__A la_oen_mprj[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[64\]_B mprj_logic_high\[394\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[62\]_TE mprj_logic_high\[264\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[107\] _375_/Y mprj_logic_high\[309\]/HI VGND VGND VPWR
+ VPWR la_oen_core[107] sky130_fd_sc_hd__einvp_8
X_660_ la_oen_mprj[61] VGND VGND VPWR VPWR _660_/Y sky130_fd_sc_hd__inv_2
X_591_ la_data_out_mprj[120] VGND VGND VPWR VPWR _591_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[37\] _636_/Y mprj_logic_high\[239\]/HI VGND VGND VPWR VPWR
+ la_oen_core[37] sky130_fd_sc_hd__einvp_8
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[377\] VGND VGND VPWR VPWR mprj_logic_high\[377\]/HI mprj_logic_high\[377\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[55\]_B mprj_logic_high\[385\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_1728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[40\]_A user_to_mprj_in_gates\[40\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y VGND VGND VPWR VPWR la_data_in_mprj[60]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[9\]_A _448_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[46\]_B mprj_logic_high\[376\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[80\]_A _551_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high\[287\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__620__A la_oen_mprj[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[31\]_A user_to_mprj_in_gates\[31\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[98\]_A user_to_mprj_in_gates\[98\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_B mprj_logic_high\[367\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_A _542_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[121\]_B mprj_logic_high\[451\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[36\] VGND VGND VPWR VPWR mprj_adr_buf\[26\]/TE mprj_logic_high\[36\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[125\] VGND VGND VPWR VPWR la_buf\[51\]/TE mprj_logic_high\[125\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__530__A la_data_out_mprj[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[22\]_A user_to_mprj_in_gates\[22\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_643_ la_oen_mprj[44] VGND VGND VPWR VPWR _643_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[64\] _535_/Y la_buf\[64\]/TE VGND VGND VPWR VPWR la_data_in_core[64] sky130_fd_sc_hd__einvp_8
X_574_ la_data_out_mprj[103] VGND VGND VPWR VPWR _574_/Y sky130_fd_sc_hd__inv_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[125\]_A _596_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[89\]_A user_to_mprj_in_gates\[89\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[28\]_B mprj_logic_high\[358\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[62\]_A _533_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B mprj_logic_high\[442\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[28\] _435_/Y mprj_adr_buf\[28\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[28]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[120\] _591_/Y la_buf\[120\]/TE VGND VGND VPWR VPWR la_data_in_core[120] sky130_fd_sc_hd__einvp_8
XFILLER_4_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__440__A mprj_dat_o_core[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[13\]_A user_to_mprj_in_gates\[13\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] mprj_logic_high\[383\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[53\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[127\]_A user_to_mprj_in_gates\[127\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__615__A la_oen_mprj[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[116\]_A _587_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[19\]_B mprj_logic_high\[349\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[53\]_A _524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B mprj_logic_high\[433\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__350__A la_oen_mprj[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[118\]_A user_to_mprj_in_gates\[118\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__525__A la_data_out_mprj[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[107\]_A _578_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[44\]_A _515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[242\] VGND VGND VPWR VPWR mprj_logic_high\[242\]/HI mprj_logic_high\[242\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_626_ la_oen_mprj[27] VGND VGND VPWR VPWR _626_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_557_ la_data_out_mprj[86] VGND VGND VPWR VPWR _557_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[109\]_A user_to_mprj_in_gates\[109\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__435__A mprj_adr_o_core[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_488_ la_data_out_mprj[17] VGND VGND VPWR VPWR _488_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y VGND VGND VPWR VPWR la_data_in_mprj[23]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[35\]_A _506_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[120\]_A _388_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__345__A la_oen_mprj[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_A _497_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[111\]_A _379_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_411_ mprj_adr_o_core[4] VGND VGND VPWR VPWR _411_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[192\] VGND VGND VPWR VPWR la_buf\[118\]/TE mprj_logic_high\[192\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[1\] _600_/Y mprj_logic_high\[203\]/HI VGND VGND VPWR VPWR
+ la_oen_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_15_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_342_ la_oen_mprj[74] VGND VGND VPWR VPWR _342_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[11\]_TE la_buf\[11\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[457\] VGND VGND VPWR VPWR mprj_logic_high\[457\]/HI mprj_logic_high\[457\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[17\]_A _488_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[27\] _498_/Y la_buf\[27\]/TE VGND VGND VPWR VPWR la_data_in_core[27] sky130_fd_sc_hd__einvp_8
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[102\]_A _370_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_609_ la_oen_mprj[10] VGND VGND VPWR VPWR _609_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] mprj_logic_high\[346\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[16\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] mprj_logic_high\[457\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[127\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[34\]_TE la_buf\[34\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high\[221\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[95\]_A _363_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[67\] _335_/Y mprj_logic_high\[269\]/HI VGND VGND VPWR VPWR
+ la_oen_core[67] sky130_fd_sc_hd__einvp_8
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[15\] _454_/Y mprj_dat_buf\[15\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[205\] VGND VGND VPWR VPWR mprj_logic_high\[205\]/HI mprj_logic_high\[205\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[86\]_A _354_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[2\]_TE la_buf\[2\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[10\] _417_/Y mprj_adr_buf\[10\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[124] sky130_fd_sc_hd__inv_8
XFILLER_2_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[10\]_A _609_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y VGND VGND VPWR VPWR la_data_in_mprj[90]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[57\]_TE la_buf\[57\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[77\]_A _345_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__623__A la_oen_mprj[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[68\]_A _336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[66\] VGND VGND VPWR VPWR mprj_dat_buf\[24\]/TE mprj_logic_high\[66\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[155\] VGND VGND VPWR VPWR la_buf\[81\]/TE mprj_logic_high\[155\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__533__A la_data_out_mprj[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[322\] VGND VGND VPWR VPWR mprj_logic_high\[322\]/HI mprj_logic_high\[322\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[94\] _565_/Y la_buf\[94\]/TE VGND VGND VPWR VPWR la_data_in_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_19_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[59\]_A _658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__443__A mprj_dat_o_core[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] mprj_logic_high\[413\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[83\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__618__A la_oen_mprj[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high\[210\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__353__A la_oen_mprj[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_590_ la_data_out_mprj[119] VGND VGND VPWR VPWR _590_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__528__A la_data_out_mprj[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[272\] VGND VGND VPWR VPWR mprj_logic_high\[272\]/HI mprj_logic_high\[272\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xla_buf\[5\] _476_/Y la_buf\[5\]/TE VGND VGND VPWR VPWR la_data_in_core[5] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[2\] _409_/Y mprj_adr_buf\[2\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__438__A mprj_adr_o_core[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y VGND VGND VPWR VPWR la_data_in_mprj[53]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[10\]_A _449_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[28\]_A _435_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__348__A la_oen_mprj[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[5\]_A _604_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[19\]_A _426_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[29\] VGND VGND VPWR VPWR mprj_adr_buf\[19\]/TE mprj_logic_high\[29\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_sel_buf\[0\] _403_/Y mprj_sel_buf\[0\]/TE VGND VGND VPWR VPWR mprj_sel_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[118\] VGND VGND VPWR VPWR la_buf\[44\]/TE mprj_logic_high\[118\]/LO
+ sky130_fd_sc_hd__conb_1
X_642_ la_oen_mprj[43] VGND VGND VPWR VPWR _642_/Y sky130_fd_sc_hd__inv_2
X_573_ la_data_out_mprj[102] VGND VGND VPWR VPWR _573_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[105\]_TE la_buf\[105\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[57\] _528_/Y la_buf\[57\]/TE VGND VGND VPWR VPWR la_data_in_core[57] sky130_fd_sc_hd__einvp_8
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[113\] _584_/Y la_buf\[113\]/TE VGND VGND VPWR VPWR la_data_in_core[113] sky130_fd_sc_hd__einvp_8
XFILLER_4_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] mprj_logic_high\[376\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[46\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high\[254\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__631__A la_oen_mprj[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[8\]_TE mprj_dat_buf\[8\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] mprj_logic_high\[338\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[8\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[97\] _365_/Y mprj_logic_high\[299\]/HI VGND VGND VPWR VPWR
+ la_oen_core[97] sky130_fd_sc_hd__einvp_8
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__541__A la_data_out_mprj[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[235\] VGND VGND VPWR VPWR mprj_logic_high\[235\]/HI mprj_logic_high\[235\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[402\] VGND VGND VPWR VPWR mprj_logic_high\[402\]/HI mprj_logic_high\[402\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[90\]_TE la_buf\[90\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_625_ la_oen_mprj[26] VGND VGND VPWR VPWR _625_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high\[277\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_556_ la_data_out_mprj[85] VGND VGND VPWR VPWR _556_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_487_ la_data_out_mprj[16] VGND VGND VPWR VPWR _487_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y VGND VGND VPWR VPWR la_data_in_mprj[16]
+ sky130_fd_sc_hd__inv_8
XANTENNA__451__A mprj_dat_o_core[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__626__A la_oen_mprj[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[4\]_A _411_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__361__A la_oen_mprj[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high\[300\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[96\] VGND VGND VPWR VPWR la_buf\[22\]/TE mprj_logic_high\[96\]/LO
+ sky130_fd_sc_hd__conb_1
X_410_ mprj_adr_o_core[3] VGND VGND VPWR VPWR _410_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__536__A la_data_out_mprj[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[12\] _611_/Y mprj_logic_high\[214\]/HI VGND VGND VPWR VPWR
+ la_oen_core[12] sky130_fd_sc_hd__einvp_8
X_341_ la_oen_mprj[73] VGND VGND VPWR VPWR _341_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[185\] VGND VGND VPWR VPWR la_buf\[111\]/TE mprj_logic_high\[185\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y VGND VGND VPWR VPWR la_data_in_mprj[8]
+ sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[352\] VGND VGND VPWR VPWR mprj_logic_high\[352\]/HI mprj_logic_high\[352\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_stb_buf _401_/Y mprj_stb_buf/TE VGND VGND VPWR VPWR mprj_stb_o_user sky130_fd_sc_hd__einvp_8
XFILLER_20_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_608_ la_oen_mprj[9] VGND VGND VPWR VPWR _608_/Y sky130_fd_sc_hd__inv_2
XANTENNA__446__A mprj_dat_o_core[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_539_ la_data_out_mprj[68] VGND VGND VPWR VPWR _539_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__356__A la_oen_mprj[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[11\] VGND VGND VPWR VPWR mprj_adr_buf\[1\]/TE mprj_logic_high\[11\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[100\] VGND VGND VPWR VPWR la_buf\[26\]/TE mprj_logic_high\[100\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk_buf_A _398_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[30\]_TE mprj_adr_buf\[30\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[117] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y VGND VGND VPWR VPWR la_data_in_mprj[83]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[4\]_B mprj_logic_high\[334\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[59\] VGND VGND VPWR VPWR mprj_dat_buf\[17\]/TE mprj_logic_high\[59\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[148\] VGND VGND VPWR VPWR la_buf\[74\]/TE mprj_logic_high\[148\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[315\] VGND VGND VPWR VPWR mprj_logic_high\[315\]/HI mprj_logic_high\[315\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[87\] _558_/Y la_buf\[87\]/TE VGND VGND VPWR VPWR la_data_in_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_1_1803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[24\]_TE la_buf\[24\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] mprj_logic_high\[406\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[76\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[8\]_A user_to_mprj_in_gates\[8\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__634__A la_oen_mprj[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[265\] VGND VGND VPWR VPWR mprj_logic_high\[265\]/HI mprj_logic_high\[265\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__544__A la_data_out_mprj[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[47\]_TE la_buf\[47\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[432\] VGND VGND VPWR VPWR mprj_logic_high\[432\]/HI mprj_logic_high\[432\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y VGND VGND VPWR VPWR la_data_in_mprj[46]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__454__A mprj_dat_o_core[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__629__A la_oen_mprj[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] mprj_logic_high\[432\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[102\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__364__A la_oen_mprj[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[112\] _380_/Y mprj_logic_high\[314\]/HI VGND VGND VPWR
+ VPWR la_oen_core[112] sky130_fd_sc_hd__einvp_8
X_641_ la_oen_mprj[42] VGND VGND VPWR VPWR _641_/Y sky130_fd_sc_hd__inv_2
XANTENNA__539__A la_data_out_mprj[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[42\] _641_/Y mprj_logic_high\[244\]/HI VGND VGND VPWR VPWR
+ la_oen_core[42] sky130_fd_sc_hd__einvp_8
X_572_ la_data_out_mprj[101] VGND VGND VPWR VPWR _572_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[382\] VGND VGND VPWR VPWR mprj_logic_high\[382\]/HI mprj_logic_high\[382\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xla_buf\[106\] _577_/Y la_buf\[106\]/TE VGND VGND VPWR VPWR la_data_in_core[106] sky130_fd_sc_hd__einvp_8
XFILLER_7_1820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__449__A mprj_dat_o_core[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] mprj_logic_high\[369\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[39\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__359__A la_oen_mprj[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[41\] VGND VGND VPWR VPWR mprj_adr_buf\[31\]/TE mprj_logic_high\[41\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[130\] VGND VGND VPWR VPWR la_buf\[56\]/TE mprj_logic_high\[130\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[228\] VGND VGND VPWR VPWR mprj_logic_high\[228\]/HI mprj_logic_high\[228\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high\[322\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_624_ la_oen_mprj[25] VGND VGND VPWR VPWR _624_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_555_ la_data_out_mprj[84] VGND VGND VPWR VPWR _555_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_486_ la_data_out_mprj[15] VGND VGND VPWR VPWR _486_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_we_buf _402_/Y mprj_we_buf/TE VGND VGND VPWR VPWR mprj_we_o_user sky130_fd_sc_hd__einvp_8
XFILLER_13_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_pwrgood mprj_pwrgood/A VGND VGND VPWR VPWR user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_7_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__642__A la_oen_mprj[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[89\] VGND VGND VPWR VPWR la_buf\[15\]/TE mprj_logic_high\[89\]/LO
+ sky130_fd_sc_hd__conb_1
X_340_ la_oen_mprj[72] VGND VGND VPWR VPWR _340_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[178\] VGND VGND VPWR VPWR la_buf\[104\]/TE mprj_logic_high\[178\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__552__A la_data_out_mprj[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[345\] VGND VGND VPWR VPWR mprj_logic_high\[345\]/HI mprj_logic_high\[345\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[42\]_TE mprj_logic_high\[244\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_607_ la_oen_mprj[8] VGND VGND VPWR VPWR _607_/Y sky130_fd_sc_hd__inv_2
X_538_ la_data_out_mprj[67] VGND VGND VPWR VPWR _538_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_469_ mprj_dat_o_core[30] VGND VGND VPWR VPWR _469_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__462__A mprj_dat_o_core[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[118\]_TE la_buf\[118\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[6\] VGND VGND VPWR VPWR mprj_sel_buf\[0\]/TE mprj_logic_high\[6\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__637__A la_oen_mprj[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[94\]_B mprj_logic_high\[424\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__372__A la_oen_mprj[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_TE la_buf\[80\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[65\]_TE mprj_logic_high\[267\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__547__A la_data_out_mprj[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[295\] VGND VGND VPWR VPWR mprj_logic_high\[295\]/HI mprj_logic_high\[295\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_we_buf_A _402_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[85\]_B mprj_logic_high\[415\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[32\] _503_/Y la_buf\[32\]/TE VGND VGND VPWR VPWR la_data_in_core[32] sky130_fd_sc_hd__einvp_8
XFILLER_11_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[70\]_A user_to_mprj_in_gates\[70\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y VGND VGND VPWR VPWR la_data_in_mprj[76]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__457__A mprj_dat_o_core[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] mprj_logic_high\[351\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[21\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[76\]_B mprj_logic_high\[406\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high\[290\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[9\] _448_/Y mprj_dat_buf\[9\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[61\]_A user_to_mprj_in_gates\[61\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__367__A la_oen_mprj[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[67\]_B mprj_logic_high\[397\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[72\] _340_/Y mprj_logic_high\[274\]/HI VGND VGND VPWR VPWR
+ la_oen_core[72] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[210\] VGND VGND VPWR VPWR mprj_logic_high\[210\]/HI mprj_logic_high\[210\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[20\] _459_/Y mprj_dat_buf\[20\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[20]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[308\] VGND VGND VPWR VPWR mprj_logic_high\[308\]/HI mprj_logic_high\[308\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[52\]_A user_to_mprj_in_gates\[52\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[58\]_B mprj_logic_high\[388\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[92\]_A _563_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[43\]_A user_to_mprj_in_gates\[43\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] mprj_logic_high\[399\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[69\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[49\]_B mprj_logic_high\[379\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[83\]_A _554_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__650__A la_oen_mprj[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[34\]_A user_to_mprj_in_gates\[34\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[20\]_TE mprj_adr_buf\[20\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[71\] VGND VGND VPWR VPWR mprj_dat_buf\[29\]/TE mprj_logic_high\[71\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[74\]_A _545_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_B mprj_logic_high\[454\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[258\] VGND VGND VPWR VPWR mprj_logic_high\[258\]/HI mprj_logic_high\[258\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[160\] VGND VGND VPWR VPWR la_buf\[86\]/TE mprj_logic_high\[160\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__560__A la_data_out_mprj[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[425\] VGND VGND VPWR VPWR mprj_logic_high\[425\]/HI mprj_logic_high\[425\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[25\]_A user_to_mprj_in_gates\[25\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y VGND VGND VPWR VPWR la_data_in_mprj[39]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[65\]_A _536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_B mprj_logic_high\[445\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__470__A mprj_dat_o_core[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[16\]_A user_to_mprj_in_gates\[16\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__645__A la_oen_mprj[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[119\]_A _590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[56\]_A _527_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_B mprj_logic_high\[436\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__380__A la_oen_mprj[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[105\] _373_/Y mprj_logic_high\[307\]/HI VGND VGND VPWR
+ VPWR la_oen_core[105] sky130_fd_sc_hd__einvp_8
X_640_ la_oen_mprj[41] VGND VGND VPWR VPWR _640_/Y sky130_fd_sc_hd__inv_2
X_571_ la_data_out_mprj[100] VGND VGND VPWR VPWR _571_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[35\] _634_/Y mprj_logic_high\[237\]/HI VGND VGND VPWR VPWR
+ la_oen_core[35] sky130_fd_sc_hd__einvp_8
XANTENNA__555__A la_data_out_mprj[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[14\]_TE la_buf\[14\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[375\] VGND VGND VPWR VPWR mprj_logic_high\[375\]/HI mprj_logic_high\[375\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[47\]_A _518_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__465__A mprj_dat_o_core[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[38\]_A _509_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[123\]_A _391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[37\]_TE la_buf\[37\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__375__A la_oen_mprj[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[29\]_A _500_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[34\] VGND VGND VPWR VPWR mprj_adr_buf\[24\]/TE mprj_logic_high\[34\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[114\]_A _382_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[123\] VGND VGND VPWR VPWR la_buf\[49\]/TE mprj_logic_high\[123\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_623_ la_oen_mprj[24] VGND VGND VPWR VPWR _623_/Y sky130_fd_sc_hd__inv_2
X_554_ la_data_out_mprj[83] VGND VGND VPWR VPWR _554_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[62\] _533_/Y la_buf\[62\]/TE VGND VGND VPWR VPWR la_data_in_core[62] sky130_fd_sc_hd__einvp_8
XFILLER_18_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_485_ la_data_out_mprj[14] VGND VGND VPWR VPWR _485_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[5\]_TE la_buf\[5\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[26\] _433_/Y mprj_adr_buf\[26\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[105\]_A _373_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[40\]_A _639_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] mprj_logic_high\[381\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[51\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[31\]_A _630_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_A _366_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[240\] VGND VGND VPWR VPWR mprj_logic_high\[240\]/HI mprj_logic_high\[240\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[338\] VGND VGND VPWR VPWR mprj_logic_high\[338\]/HI mprj_logic_high\[338\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[22\]_A _621_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_606_ la_oen_mprj[7] VGND VGND VPWR VPWR _606_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[89\]_A _357_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_537_ la_data_out_mprj[66] VGND VGND VPWR VPWR _537_/Y sky130_fd_sc_hd__inv_2
X_468_ mprj_dat_o_core[29] VGND VGND VPWR VPWR _468_/Y sky130_fd_sc_hd__inv_2
X_399_ caravel_clk2 VGND VGND VPWR VPWR _399_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y VGND VGND VPWR VPWR la_data_in_mprj[21]
+ sky130_fd_sc_hd__inv_8
XFILLER_16_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] mprj_logic_high\[429\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[99\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[13\]_A _612_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__653__A la_oen_mprj[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[110\]_TE mprj_logic_high\[312\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[190\] VGND VGND VPWR VPWR la_buf\[116\]/TE mprj_logic_high\[190\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[288\] VGND VGND VPWR VPWR mprj_logic_high\[288\]/HI mprj_logic_high\[288\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__563__A la_data_out_mprj[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[455\] VGND VGND VPWR VPWR mprj_logic_high\[455\]/HI mprj_logic_high\[455\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[25\] _496_/Y la_buf\[25\]/TE VGND VGND VPWR VPWR la_data_in_core[25] sky130_fd_sc_hd__einvp_8
XFILLER_13_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y VGND VGND VPWR VPWR la_data_in_mprj[69]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__473__A la_data_out_mprj[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] mprj_logic_high\[344\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[14\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] mprj_logic_high\[455\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[125\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__648__A la_oen_mprj[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[31\]_A _470_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__383__A la_oen_mprj[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[32\]_TE mprj_logic_high\[234\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[65\] _333_/Y mprj_logic_high\[267\]/HI VGND VGND VPWR VPWR
+ la_oen_core[65] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[13\] _452_/Y mprj_dat_buf\[13\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[13]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[203\] VGND VGND VPWR VPWR mprj_logic_high\[203\]/HI mprj_logic_high\[203\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__558__A la_data_out_mprj[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[108\]_TE la_buf\[108\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[22\]_A _461_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[7\]_TE mprj_adr_buf\[7\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[122] sky130_fd_sc_hd__inv_8
XFILLER_2_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__468__A mprj_dat_o_core[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[70\]_TE la_buf\[70\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[13\]_A _452_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[55\]_TE mprj_logic_high\[257\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__378__A la_oen_mprj[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[8\]_A _607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[64\] VGND VGND VPWR VPWR mprj_dat_buf\[22\]/TE mprj_logic_high\[64\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[153\] VGND VGND VPWR VPWR la_buf\[79\]/TE mprj_logic_high\[153\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[320\] VGND VGND VPWR VPWR mprj_logic_high\[320\]/HI mprj_logic_high\[320\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[418\] VGND VGND VPWR VPWR mprj_logic_high\[418\]/HI mprj_logic_high\[418\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[92\] _563_/Y la_buf\[92\]/TE VGND VGND VPWR VPWR la_data_in_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_0_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[93\]_TE la_buf\[93\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high\[280\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A VGND VGND VPWR VPWR user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_1_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] mprj_logic_high\[411\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[81\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_570_ la_data_out_mprj[99] VGND VGND VPWR VPWR _570_/Y sky130_fd_sc_hd__inv_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[28\] _627_/Y mprj_logic_high\[230\]/HI VGND VGND VPWR VPWR
+ la_oen_core[28] sky130_fd_sc_hd__einvp_8
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[0\]_A _471_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[368\] VGND VGND VPWR VPWR mprj_logic_high\[368\]/HI mprj_logic_high\[368\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[270\] VGND VGND VPWR VPWR mprj_logic_high\[270\]/HI mprj_logic_high\[270\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__571__A la_data_out_mprj[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[3\] _474_/Y la_buf\[3\]/TE VGND VGND VPWR VPWR la_data_in_core[3] sky130_fd_sc_hd__einvp_8
XFILLER_10_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[0\] _407_/Y mprj_adr_buf\[0\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y VGND VGND VPWR VPWR la_data_in_mprj[51]
+ sky130_fd_sc_hd__inv_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__481__A la_data_out_mprj[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__656__A la_oen_mprj[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[7\]_A _414_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__391__A la_oen_mprj[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[27\] VGND VGND VPWR VPWR mprj_adr_buf\[17\]/TE mprj_logic_high\[27\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[116\] VGND VGND VPWR VPWR la_buf\[42\]/TE mprj_logic_high\[116\]/LO
+ sky130_fd_sc_hd__conb_1
X_622_ la_oen_mprj[23] VGND VGND VPWR VPWR _622_/Y sky130_fd_sc_hd__inv_2
XANTENNA__566__A la_data_out_mprj[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_553_ la_data_out_mprj[82] VGND VGND VPWR VPWR _553_/Y sky130_fd_sc_hd__inv_2
X_484_ la_data_out_mprj[13] VGND VGND VPWR VPWR _484_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[55\] _526_/Y la_buf\[55\]/TE VGND VGND VPWR VPWR la_data_in_core[55] sky130_fd_sc_hd__einvp_8
XFILLER_9_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[19\] _426_/Y mprj_adr_buf\[19\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[19]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[111\] _582_/Y la_buf\[111\]/TE VGND VGND VPWR VPWR la_data_in_core[111] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y VGND VGND VPWR VPWR la_data_in_mprj[99]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__476__A la_data_out_mprj[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] mprj_logic_high\[374\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[44\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] mprj_logic_high\[336\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[6\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__386__A la_oen_mprj[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[95\] _363_/Y mprj_logic_high\[297\]/HI VGND VGND VPWR VPWR
+ la_oen_core[95] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[233\] VGND VGND VPWR VPWR mprj_logic_high\[233\]/HI mprj_logic_high\[233\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[400\] VGND VGND VPWR VPWR mprj_logic_high\[400\]/HI mprj_logic_high\[400\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_605_ la_oen_mprj[6] VGND VGND VPWR VPWR _605_/Y sky130_fd_sc_hd__inv_2
X_536_ la_data_out_mprj[65] VGND VGND VPWR VPWR _536_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_467_ mprj_dat_o_core[28] VGND VGND VPWR VPWR _467_/Y sky130_fd_sc_hd__inv_2
X_398_ caravel_clk VGND VGND VPWR VPWR _398_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y VGND VGND VPWR VPWR la_data_in_mprj[14]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[27\]_TE la_buf\[27\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[7\]_B mprj_logic_high\[337\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[94\] VGND VGND VPWR VPWR la_buf\[20\]/TE mprj_logic_high\[94\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[10\] _609_/Y mprj_logic_high\[212\]/HI VGND VGND VPWR VPWR
+ la_oen_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[183\] VGND VGND VPWR VPWR la_buf\[109\]/TE mprj_logic_high\[183\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y VGND VGND VPWR VPWR la_data_in_mprj[6]
+ sky130_fd_sc_hd__inv_8
XFILLER_11_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[448\] VGND VGND VPWR VPWR mprj_logic_high\[448\]/HI mprj_logic_high\[448\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[350\] VGND VGND VPWR VPWR mprj_logic_high\[350\]/HI mprj_logic_high\[350\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[18\] _489_/Y la_buf\[18\]/TE VGND VGND VPWR VPWR la_data_in_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_2_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_519_ la_data_out_mprj[48] VGND VGND VPWR VPWR _519_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] mprj_logic_high\[448\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[118\]/Y sky130_fd_sc_hd__nand2_4
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[58\] _657_/Y mprj_logic_high\[260\]/HI VGND VGND VPWR VPWR
+ la_oen_core[58] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[398\] VGND VGND VPWR VPWR mprj_logic_high\[398\]/HI mprj_logic_high\[398\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__574__A la_data_out_mprj[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[115] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y VGND VGND VPWR VPWR la_data_in_mprj[81]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high\[302\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__484__A la_data_out_mprj[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__659__A la_oen_mprj[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__394__A la_oen_mprj[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[57\] VGND VGND VPWR VPWR mprj_dat_buf\[15\]/TE mprj_logic_high\[57\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[146\] VGND VGND VPWR VPWR la_buf\[72\]/TE mprj_logic_high\[146\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[313\] VGND VGND VPWR VPWR mprj_logic_high\[313\]/HI mprj_logic_high\[313\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__569__A la_data_out_mprj[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[85\] _556_/Y la_buf\[85\]/TE VGND VGND VPWR VPWR la_data_in_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_5_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high\[325\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__479__A la_data_out_mprj[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] mprj_logic_high\[404\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[74\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[22\]_TE mprj_logic_high\[224\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__389__A la_oen_mprj[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[263\] VGND VGND VPWR VPWR mprj_logic_high\[263\]/HI mprj_logic_high\[263\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[430\] VGND VGND VPWR VPWR mprj_logic_high\[430\]/HI mprj_logic_high\[430\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[60\]_TE la_buf\[60\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[45\]_TE mprj_logic_high\[247\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y VGND VGND VPWR VPWR la_data_in_mprj[44]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_sel_buf\[1\]_A _404_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] mprj_logic_high\[430\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[100\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[83\]_TE la_buf\[83\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[68\]_TE mprj_logic_high\[270\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[110\] _378_/Y mprj_logic_high\[312\]/HI VGND VGND VPWR
+ VPWR la_oen_core[110] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[109\] VGND VGND VPWR VPWR la_buf\[35\]/TE mprj_logic_high\[109\]/LO
+ sky130_fd_sc_hd__conb_1
X_621_ la_oen_mprj[22] VGND VGND VPWR VPWR _621_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[40\] _639_/Y mprj_logic_high\[242\]/HI VGND VGND VPWR VPWR
+ la_oen_core[40] sky130_fd_sc_hd__einvp_8
XFILLER_18_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_552_ la_data_out_mprj[81] VGND VGND VPWR VPWR _552_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_483_ la_data_out_mprj[12] VGND VGND VPWR VPWR _483_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[380\] VGND VGND VPWR VPWR mprj_logic_high\[380\]/HI mprj_logic_high\[380\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__582__A la_data_out_mprj[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[48\] _519_/Y la_buf\[48\]/TE VGND VGND VPWR VPWR la_data_in_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[2\]_A _441_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[104\] _575_/Y la_buf\[104\]/TE VGND VGND VPWR VPWR la_data_in_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] mprj_logic_high\[367\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[37\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__492__A la_data_out_mprj[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[91\]_A user_to_mprj_in_gates\[91\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[30\]_B mprj_logic_high\[360\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[97\]_B mprj_logic_high\[427\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[88\] _356_/Y mprj_logic_high\[290\]/HI VGND VGND VPWR VPWR
+ la_oen_core[88] sky130_fd_sc_hd__einvp_8
XFILLER_2_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[21\]_B mprj_logic_high\[351\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[226\] VGND VGND VPWR VPWR mprj_logic_high\[226\]/HI mprj_logic_high\[226\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[82\]_A user_to_mprj_in_gates\[82\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__577__A la_data_out_mprj[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_604_ la_oen_mprj[5] VGND VGND VPWR VPWR _604_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_535_ la_data_out_mprj[64] VGND VGND VPWR VPWR _535_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[88\]_B mprj_logic_high\[418\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_466_ mprj_dat_o_core[27] VGND VGND VPWR VPWR _466_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_397_ user_resetn VGND VGND VPWR VPWR user_reset sky130_fd_sc_hd__inv_2
XFILLER_13_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[31\] _438_/Y mprj_adr_buf\[31\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_16_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[120\]_A user_to_mprj_in_gates\[120\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[73\]_A user_to_mprj_in_gates\[73\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[12\]_B mprj_logic_high\[342\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_1759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__487__A la_data_out_mprj[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[79\]_B mprj_logic_high\[409\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[111\]_A user_to_mprj_in_gates\[111\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[100\]_A _571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[64\]_A user_to_mprj_in_gates\[64\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__397__A user_resetn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[23\]_TE mprj_adr_buf\[23\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[87\] VGND VGND VPWR VPWR la_buf\[13\]/TE mprj_logic_high\[87\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[176\] VGND VGND VPWR VPWR la_buf\[102\]/TE mprj_logic_high\[176\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[343\] VGND VGND VPWR VPWR mprj_logic_high\[343\]/HI mprj_logic_high\[343\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[102\]_A user_to_mprj_in_gates\[102\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[55\]_A user_to_mprj_in_gates\[55\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_A _566_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_518_ la_data_out_mprj[47] VGND VGND VPWR VPWR _518_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_449_ mprj_dat_o_core[10] VGND VGND VPWR VPWR _449_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[46\]_A user_to_mprj_in_gates\[46\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[4\] VGND VGND VPWR VPWR mprj_stb_buf/TE mprj_logic_high\[4\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[86\]_A _557_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[37\]_A user_to_mprj_in_gates\[37\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[10\]_A _481_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[17\]_TE la_buf\[17\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[293\] VGND VGND VPWR VPWR mprj_logic_high\[293\]/HI mprj_logic_high\[293\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[77\]_A _548_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_B mprj_logic_high\[457\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__590__A la_data_out_mprj[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[30\] _501_/Y la_buf\[30\]/TE VGND VGND VPWR VPWR la_data_in_core[30] sky130_fd_sc_hd__einvp_8
XFILLER_6_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[28\]_A user_to_mprj_in_gates\[28\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[108] sky130_fd_sc_hd__inv_8
XFILLER_6_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y VGND VGND VPWR VPWR la_data_in_mprj[74]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[118\]_B mprj_logic_high\[448\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[68\]_A _539_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[19\]_A user_to_mprj_in_gates\[19\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[7\] _446_/Y mprj_dat_buf\[7\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[109\]_B mprj_logic_high\[439\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[59\]_A _530_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[139\] VGND VGND VPWR VPWR la_buf\[65\]/TE mprj_logic_high\[139\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[70\] _338_/Y mprj_logic_high\[272\]/HI VGND VGND VPWR VPWR
+ la_oen_core[70] sky130_fd_sc_hd__einvp_8
XFILLER_0_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[306\] VGND VGND VPWR VPWR mprj_logic_high\[306\]/HI mprj_logic_high\[306\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[78\] _549_/Y la_buf\[78\]/TE VGND VGND VPWR VPWR la_data_in_core[78] sky130_fd_sc_hd__einvp_8
XFILLER_5_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__585__A la_data_out_mprj[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[8\]_TE la_buf\[8\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[70\]_A _338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] mprj_logic_high\[397\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[67\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__495__A la_data_out_mprj[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[61\]_A _660_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[126\]_A _394_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[256\] VGND VGND VPWR VPWR mprj_logic_high\[256\]/HI mprj_logic_high\[256\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[52\]_A _651_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_A _385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[423\] VGND VGND VPWR VPWR mprj_logic_high\[423\]/HI mprj_logic_high\[423\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y VGND VGND VPWR VPWR la_data_in_mprj[37]
+ sky130_fd_sc_hd__inv_8
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[43\]_A _642_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[108\]_A _376_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high\[315\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[34\]_A _633_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[103\] _371_/Y mprj_logic_high\[305\]/HI VGND VGND VPWR
+ VPWR la_oen_core[103] sky130_fd_sc_hd__einvp_8
X_620_ la_oen_mprj[21] VGND VGND VPWR VPWR _620_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_adr_buf\[30\]_A _437_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_551_ la_data_out_mprj[80] VGND VGND VPWR VPWR _551_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[33\] _632_/Y mprj_logic_high\[235\]/HI VGND VGND VPWR VPWR
+ la_oen_core[33] sky130_fd_sc_hd__einvp_8
X_482_ la_data_out_mprj[11] VGND VGND VPWR VPWR _482_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[373\] VGND VGND VPWR VPWR mprj_logic_high\[373\]/HI mprj_logic_high\[373\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high\[214\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[25\]_A _624_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[21\]_A _428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj2_vdd_pwrgood_A mprj2_pwrgood/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_A _615_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[12\]_A _419_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[50\]_TE la_buf\[50\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high\[237\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[32\] VGND VGND VPWR VPWR mprj_adr_buf\[22\]/TE mprj_logic_high\[32\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[29\] _468_/Y mprj_dat_buf\[29\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[29]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[121\] VGND VGND VPWR VPWR la_buf\[47\]/TE mprj_logic_high\[121\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[219\] VGND VGND VPWR VPWR mprj_logic_high\[219\]/HI mprj_logic_high\[219\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_603_ la_oen_mprj[4] VGND VGND VPWR VPWR _603_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[60\] _531_/Y la_buf\[60\]/TE VGND VGND VPWR VPWR la_data_in_core[60] sky130_fd_sc_hd__einvp_8
X_534_ la_data_out_mprj[63] VGND VGND VPWR VPWR _534_/Y sky130_fd_sc_hd__inv_2
XANTENNA__593__A la_data_out_mprj[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_465_ mprj_dat_o_core[26] VGND VGND VPWR VPWR _465_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_396_ caravel_rstn VGND VGND VPWR VPWR _396_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[24\] _431_/Y mprj_adr_buf\[24\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[73\]_TE la_buf\[73\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[58\]_TE mprj_logic_high\[260\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[169\] VGND VGND VPWR VPWR la_buf\[95\]/TE mprj_logic_high\[169\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[1\]_TE mprj_logic_high\[203\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[336\] VGND VGND VPWR VPWR mprj_logic_high\[336\]/HI mprj_logic_high\[336\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__588__A la_data_out_mprj[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[96\]_TE la_buf\[96\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[25\]_A _464_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_517_ la_data_out_mprj[46] VGND VGND VPWR VPWR _517_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_448_ mprj_dat_o_core[9] VGND VGND VPWR VPWR _448_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_379_ la_oen_mprj[111] VGND VGND VPWR VPWR _379_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] mprj_logic_high\[427\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[97\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__498__A la_data_out_mprj[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[16\]_A _455_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[286\] VGND VGND VPWR VPWR mprj_logic_high\[286\]/HI mprj_logic_high\[286\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[453\] VGND VGND VPWR VPWR mprj_logic_high\[453\]/HI mprj_logic_high\[453\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[23\] _494_/Y la_buf\[23\]/TE VGND VGND VPWR VPWR la_data_in_core[23] sky130_fd_sc_hd__einvp_8
XFILLER_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y VGND VGND VPWR VPWR la_data_in_mprj[67]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] mprj_logic_high\[342\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[12\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[13\]_TE mprj_adr_buf\[13\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] mprj_logic_high\[453\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[123\]/Y sky130_fd_sc_hd__nand2_4
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[63\] _331_/Y mprj_logic_high\[265\]/HI VGND VGND VPWR VPWR
+ la_oen_core[63] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[11\] _450_/Y mprj_dat_buf\[11\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[11]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[201\] VGND VGND VPWR VPWR la_buf\[127\]/TE mprj_logic_high\[201\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_mprj_dat_buf\[1\]_TE mprj_dat_buf\[1\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[3\]_A _474_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[121\]_TE la_buf\[121\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[127\] _598_/Y la_buf\[127\]/TE VGND VGND VPWR VPWR la_data_in_core[127] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[120] sky130_fd_sc_hd__inv_8
XFILLER_3_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[62\] VGND VGND VPWR VPWR mprj_dat_buf\[20\]/TE mprj_logic_high\[62\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[151\] VGND VGND VPWR VPWR la_buf\[77\]/TE mprj_logic_high\[151\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[249\] VGND VGND VPWR VPWR mprj_logic_high\[249\]/HI mprj_logic_high\[249\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[416\] VGND VGND VPWR VPWR mprj_logic_high\[416\]/HI mprj_logic_high\[416\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__596__A la_data_out_mprj[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[90\] _561_/Y la_buf\[90\]/TE VGND VGND VPWR VPWR la_data_in_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_1_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high\[293\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[1\]_A user_to_mprj_in_gates\[1\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_550_ la_data_out_mprj[79] VGND VGND VPWR VPWR _550_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[8\] _607_/Y mprj_logic_high\[210\]/HI VGND VGND VPWR VPWR
+ la_oen_core[8] sky130_fd_sc_hd__einvp_8
X_481_ la_data_out_mprj[10] VGND VGND VPWR VPWR _481_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[199\] VGND VGND VPWR VPWR la_buf\[125\]/TE mprj_logic_high\[199\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[26\] _625_/Y mprj_logic_high\[228\]/HI VGND VGND VPWR VPWR
+ la_oen_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_12_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[366\] VGND VGND VPWR VPWR mprj_logic_high\[366\]/HI mprj_logic_high\[366\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[1\] _472_/Y la_buf\[1\]/TE VGND VGND VPWR VPWR la_data_in_core[1] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[25\] VGND VGND VPWR VPWR mprj_adr_buf\[15\]/TE mprj_logic_high\[25\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[114\] VGND VGND VPWR VPWR la_buf\[40\]/TE mprj_logic_high\[114\]/LO
+ sky130_fd_sc_hd__conb_1
X_602_ la_oen_mprj[3] VGND VGND VPWR VPWR _602_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_533_ la_data_out_mprj[62] VGND VGND VPWR VPWR _533_/Y sky130_fd_sc_hd__inv_2
X_464_ mprj_dat_o_core[25] VGND VGND VPWR VPWR _464_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[53\] _524_/Y la_buf\[53\]/TE VGND VGND VPWR VPWR la_data_in_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_395_ la_oen_mprj[127] VGND VGND VPWR VPWR _395_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[17\] _424_/Y mprj_adr_buf\[17\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y VGND VGND VPWR VPWR la_data_in_mprj[97]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high\[305\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] mprj_logic_high\[372\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[42\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] mprj_logic_high\[334\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[4\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[93\] _361_/Y mprj_logic_high\[295\]/HI VGND VGND VPWR VPWR
+ la_oen_core[93] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[231\] VGND VGND VPWR VPWR mprj_logic_high\[231\]/HI mprj_logic_high\[231\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[329\] VGND VGND VPWR VPWR mprj_logic_high\[329\]/HI mprj_logic_high\[329\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high\[328\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_516_ la_data_out_mprj[45] VGND VGND VPWR VPWR _516_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_447_ mprj_dat_o_core[8] VGND VGND VPWR VPWR _447_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_378_ la_oen_mprj[110] VGND VGND VPWR VPWR _378_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y VGND VGND VPWR VPWR la_data_in_mprj[12]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[40\]_TE la_buf\[40\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[25\]_TE mprj_logic_high\[227\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[92\] VGND VGND VPWR VPWR la_buf\[18\]/TE mprj_logic_high\[92\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y VGND VGND VPWR VPWR la_data_in_mprj[4]
+ sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[181\] VGND VGND VPWR VPWR la_buf\[107\]/TE mprj_logic_high\[181\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[279\] VGND VGND VPWR VPWR mprj_logic_high\[279\]/HI mprj_logic_high\[279\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[446\] VGND VGND VPWR VPWR mprj_logic_high\[446\]/HI mprj_logic_high\[446\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[63\]_TE la_buf\[63\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[16\] _487_/Y la_buf\[16\]/TE VGND VGND VPWR VPWR la_data_in_core[16] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[48\]_TE mprj_logic_high\[250\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__599__A la_oen_mprj[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[9\] _416_/Y mprj_adr_buf\[9\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] mprj_logic_high\[446\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[116\]/Y sky130_fd_sc_hd__nand2_4
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[86\]_TE la_buf\[86\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[126\] _394_/Y mprj_logic_high\[328\]/HI VGND VGND VPWR
+ VPWR la_oen_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_0_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[56\] _655_/Y mprj_logic_high\[258\]/HI VGND VGND VPWR VPWR
+ la_oen_core[56] sky130_fd_sc_hd__einvp_8
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[396\] VGND VGND VPWR VPWR mprj_logic_high\[396\]/HI mprj_logic_high\[396\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[113] sky130_fd_sc_hd__inv_8
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[60\]_B mprj_logic_high\[390\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[55\] VGND VGND VPWR VPWR mprj_dat_buf\[13\]/TE mprj_logic_high\[55\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[144\] VGND VGND VPWR VPWR la_buf\[70\]/TE mprj_logic_high\[144\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[51\]_B mprj_logic_high\[381\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[409\] VGND VGND VPWR VPWR mprj_logic_high\[409\]/HI mprj_logic_high\[409\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[311\] VGND VGND VPWR VPWR mprj_logic_high\[311\]/HI mprj_logic_high\[311\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[83\] _554_/Y la_buf\[83\]/TE VGND VGND VPWR VPWR la_data_in_core[83] sky130_fd_sc_hd__einvp_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[5\]_A _444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[42\]_B mprj_logic_high\[372\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] mprj_logic_high\[402\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[72\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[94\]_A user_to_mprj_in_gates\[94\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[33\]_B mprj_logic_high\[363\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[111\]_TE la_buf\[111\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[26\]_TE mprj_adr_buf\[26\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_480_ la_data_out_mprj[9] VGND VGND VPWR VPWR _480_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[19\] _618_/Y mprj_logic_high\[221\]/HI VGND VGND VPWR VPWR
+ la_oen_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[261\] VGND VGND VPWR VPWR mprj_logic_high\[261\]/HI mprj_logic_high\[261\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[359\] VGND VGND VPWR VPWR mprj_logic_high\[359\]/HI mprj_logic_high\[359\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[121\]_A _592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[85\]_A user_to_mprj_in_gates\[85\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[24\]_B mprj_logic_high\[354\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__400__A mprj_cyc_o_core VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y VGND VGND VPWR VPWR la_data_in_mprj[42]
+ sky130_fd_sc_hd__inv_8
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[123\]_A user_to_mprj_in_gates\[123\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[112\]_A _583_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[76\]_A user_to_mprj_in_gates\[76\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[15\]_B mprj_logic_high\[345\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[114\]_A user_to_mprj_in_gates\[114\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[103\]_A _574_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[67\]_A user_to_mprj_in_gates\[67\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[40\]_A _511_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[18\] VGND VGND VPWR VPWR mprj_adr_buf\[8\]/TE mprj_logic_high\[18\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high\[283\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[107\] VGND VGND VPWR VPWR la_buf\[33\]/TE mprj_logic_high\[107\]/LO
+ sky130_fd_sc_hd__conb_1
X_601_ la_oen_mprj[2] VGND VGND VPWR VPWR _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_532_ la_data_out_mprj[61] VGND VGND VPWR VPWR _532_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_463_ mprj_dat_o_core[24] VGND VGND VPWR VPWR _463_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_394_ la_oen_mprj[126] VGND VGND VPWR VPWR _394_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[46\] _517_/Y la_buf\[46\]/TE VGND VGND VPWR VPWR la_data_in_core[46] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[105\]_A user_to_mprj_in_gates\[105\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[58\]_A user_to_mprj_in_gates\[58\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[31\]_A _502_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[102\] _573_/Y la_buf\[102\]/TE VGND VGND VPWR VPWR la_data_in_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_1_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[98\]_A _569_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] mprj_logic_high\[365\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[35\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[49\]_A user_to_mprj_in_gates\[49\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[22\]_A _493_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[89\]_A _560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[86\] _354_/Y mprj_logic_high\[288\]/HI VGND VGND VPWR VPWR
+ la_oen_core[86] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[13\]_A _484_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[224\] VGND VGND VPWR VPWR mprj_logic_high\[224\]/HI mprj_logic_high\[224\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_18_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_515_ la_data_out_mprj[44] VGND VGND VPWR VPWR _515_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_446_ mprj_dat_o_core[7] VGND VGND VPWR VPWR _446_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_377_ la_oen_mprj[109] VGND VGND VPWR VPWR _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[91\]_A _359_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[85\] VGND VGND VPWR VPWR la_buf\[11\]/TE mprj_logic_high\[85\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[174\] VGND VGND VPWR VPWR la_buf\[100\]/TE mprj_logic_high\[174\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[341\] VGND VGND VPWR VPWR mprj_logic_high\[341\]/HI mprj_logic_high\[341\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_A _350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[439\] VGND VGND VPWR VPWR mprj_logic_high\[439\]/HI mprj_logic_high\[439\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_429_ mprj_adr_o_core[22] VGND VGND VPWR VPWR _429_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[73\]_A _341_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[2\] VGND VGND VPWR VPWR mprj_clk2_buf/TE mprj_logic_high\[2\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] mprj_logic_high\[439\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[109\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high\[318\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[64\]_A _332_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[119\] _387_/Y mprj_logic_high\[321\]/HI VGND VGND VPWR
+ VPWR la_oen_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[49\] _648_/Y mprj_logic_high\[251\]/HI VGND VGND VPWR VPWR
+ la_oen_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_5_1787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[291\] VGND VGND VPWR VPWR mprj_logic_high\[291\]/HI mprj_logic_high\[291\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[389\] VGND VGND VPWR VPWR mprj_logic_high\[389\]/HI mprj_logic_high\[389\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[30\]_TE la_buf\[30\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high\[217\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[55\]_A _654_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__403__A mprj_sel_o_core[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[106] sky130_fd_sc_hd__inv_8
XFILLER_19_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y VGND VGND VPWR VPWR la_data_in_mprj[72]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_A _645_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[5\] _444_/Y mprj_dat_buf\[5\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[53\]_TE la_buf\[53\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[38\]_TE mprj_logic_high\[240\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[37\]_A _636_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[48\] VGND VGND VPWR VPWR mprj_dat_buf\[6\]/TE mprj_logic_high\[48\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[137\] VGND VGND VPWR VPWR la_buf\[63\]/TE mprj_logic_high\[137\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[304\] VGND VGND VPWR VPWR mprj_logic_high\[304\]/HI mprj_logic_high\[304\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[76\] _547_/Y la_buf\[76\]/TE VGND VGND VPWR VPWR la_data_in_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_1_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[28\]_A _627_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[24\]_A _431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[76\]_TE la_buf\[76\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] mprj_logic_high\[395\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[65\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[19\]_A _618_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[1\]_A _600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[15\]_A _422_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high\[206\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[254\] VGND VGND VPWR VPWR mprj_logic_high\[254\]/HI mprj_logic_high\[254\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[421\] VGND VGND VPWR VPWR mprj_logic_high\[421\]/HI mprj_logic_high\[421\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[99\]_TE la_buf\[99\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y VGND VGND VPWR VPWR la_data_in_mprj[35]
+ sky130_fd_sc_hd__inv_8
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__501__A la_data_out_mprj[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _369_/Y mprj_logic_high\[303\]/HI VGND VGND VPWR
+ VPWR la_oen_core[101] sky130_fd_sc_hd__einvp_8
X_600_ la_oen_mprj[1] VGND VGND VPWR VPWR _600_/Y sky130_fd_sc_hd__inv_2
X_531_ la_data_out_mprj[60] VGND VGND VPWR VPWR _531_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[31\] _630_/Y mprj_logic_high\[233\]/HI VGND VGND VPWR VPWR
+ la_oen_core[31] sky130_fd_sc_hd__einvp_8
X_462_ mprj_dat_o_core[23] VGND VGND VPWR VPWR _462_/Y sky130_fd_sc_hd__inv_2
X_393_ la_oen_mprj[125] VGND VGND VPWR VPWR _393_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[371\] VGND VGND VPWR VPWR mprj_logic_high\[371\]/HI mprj_logic_high\[371\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[39\] _510_/Y la_buf\[39\]/TE VGND VGND VPWR VPWR la_data_in_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_16_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__411__A mprj_adr_o_core[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[28\]_A _467_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] mprj_logic_high\[358\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[28\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[101\]_TE la_buf\[101\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[0\]_A _407_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[19\]_A _458_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[30\] VGND VGND VPWR VPWR mprj_adr_buf\[20\]/TE mprj_logic_high\[30\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[79\] _347_/Y mprj_logic_high\[281\]/HI VGND VGND VPWR VPWR
+ la_oen_core[79] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[27\] _466_/Y mprj_dat_buf\[27\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[27]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[217\] VGND VGND VPWR VPWR mprj_logic_high\[217\]/HI mprj_logic_high\[217\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_mprj_dat_buf\[4\]_TE mprj_dat_buf\[4\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_514_ la_data_out_mprj[43] VGND VGND VPWR VPWR _514_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[124\]_TE la_buf\[124\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_445_ mprj_dat_o_core[6] VGND VGND VPWR VPWR _445_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_376_ la_oen_mprj[108] VGND VGND VPWR VPWR _376_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__406__A mprj_sel_o_core[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[22\] _429_/Y mprj_adr_buf\[22\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high\[273\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[78\] VGND VGND VPWR VPWR la_buf\[4\]/TE mprj_logic_high\[78\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[167\] VGND VGND VPWR VPWR la_buf\[93\]/TE mprj_logic_high\[167\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[334\] VGND VGND VPWR VPWR mprj_logic_high\[334\]/HI mprj_logic_high\[334\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[6\]_A _477_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high\[296\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_428_ mprj_adr_o_core[21] VGND VGND VPWR VPWR _428_/Y sky130_fd_sc_hd__inv_2
X_359_ la_oen_mprj[91] VGND VGND VPWR VPWR _359_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] mprj_logic_high\[425\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[95\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[0\]_B mprj_logic_high\[330\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[284\] VGND VGND VPWR VPWR mprj_logic_high\[284\]/HI mprj_logic_high\[284\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[451\] VGND VGND VPWR VPWR mprj_logic_high\[451\]/HI mprj_logic_high\[451\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[21\] _492_/Y la_buf\[21\]/TE VGND VGND VPWR VPWR la_data_in_core[21] sky130_fd_sc_hd__einvp_8
XFILLER_20_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[4\]_A user_to_mprj_in_gates\[4\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y VGND VGND VPWR VPWR la_data_in_mprj[65]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] mprj_logic_high\[340\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[10\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] mprj_logic_high\[451\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[121\]/Y sky130_fd_sc_hd__nand2_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__504__A la_data_out_mprj[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[61\] _660_/Y mprj_logic_high\[263\]/HI VGND VGND VPWR VPWR
+ la_oen_core[61] sky130_fd_sc_hd__einvp_8
XFILLER_5_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xla_buf\[69\] _540_/Y la_buf\[69\]/TE VGND VGND VPWR VPWR la_data_in_core[69] sky130_fd_sc_hd__einvp_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__414__A mprj_adr_o_core[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[125\] _596_/Y la_buf\[125\]/TE VGND VGND VPWR VPWR la_data_in_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_6_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high\[308\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] mprj_logic_high\[388\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[58\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[20\]_TE la_buf\[20\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[60\] VGND VGND VPWR VPWR mprj_dat_buf\[18\]/TE mprj_logic_high\[60\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[247\] VGND VGND VPWR VPWR mprj_logic_high\[247\]/HI mprj_logic_high\[247\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[414\] VGND VGND VPWR VPWR mprj_logic_high\[414\]/HI mprj_logic_high\[414\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__409__A mprj_adr_o_core[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y VGND VGND VPWR VPWR la_data_in_mprj[28]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_TE la_buf\[43\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[28\]_TE mprj_logic_high\[230\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_530_ la_data_out_mprj[59] VGND VGND VPWR VPWR _530_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[6\] _605_/Y mprj_logic_high\[208\]/HI VGND VGND VPWR VPWR
+ la_oen_core[6] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[197\] VGND VGND VPWR VPWR la_buf\[123\]/TE mprj_logic_high\[197\]/LO
+ sky130_fd_sc_hd__conb_1
X_461_ mprj_dat_o_core[22] VGND VGND VPWR VPWR _461_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[24\] _623_/Y mprj_logic_high\[226\]/HI VGND VGND VPWR VPWR
+ la_oen_core[24] sky130_fd_sc_hd__einvp_8
X_392_ la_oen_mprj[124] VGND VGND VPWR VPWR _392_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[364\] VGND VGND VPWR VPWR mprj_logic_high\[364\]/HI mprj_logic_high\[364\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[66\]_TE la_buf\[66\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_659_ la_oen_mprj[60] VGND VGND VPWR VPWR _659_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[15\]_TE mprj_dat_buf\[15\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__602__A la_oen_mprj[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[89\]_TE la_buf\[89\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__512__A VPWR VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[23\] VGND VGND VPWR VPWR mprj_adr_buf\[13\]/TE mprj_logic_high\[23\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[112\] VGND VGND VPWR VPWR la_buf\[38\]/TE mprj_logic_high\[112\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_513_ la_data_out_mprj[42] VGND VGND VPWR VPWR _513_/Y sky130_fd_sc_hd__inv_2
X_444_ mprj_dat_o_core[5] VGND VGND VPWR VPWR _444_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[51\] _522_/Y la_buf\[51\]/TE VGND VGND VPWR VPWR la_data_in_core[51] sky130_fd_sc_hd__einvp_8
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_375_ la_oen_mprj[107] VGND VGND VPWR VPWR _375_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__422__A mprj_adr_o_core[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[15\] _422_/Y mprj_adr_buf\[15\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y VGND VGND VPWR VPWR la_data_in_mprj[95]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] mprj_logic_high\[370\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[40\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[90\]_B mprj_logic_high\[420\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__332__A la_oen_mprj[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] mprj_logic_high\[332\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[2\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__507__A la_data_out_mprj[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[81\]_B mprj_logic_high\[411\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[91\] _359_/Y mprj_logic_high\[293\]/HI VGND VGND VPWR VPWR
+ la_oen_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_3_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[327\] VGND VGND VPWR VPWR mprj_logic_high\[327\]/HI mprj_logic_high\[327\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[99\] _570_/Y la_buf\[99\]/TE VGND VGND VPWR VPWR la_data_in_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_19_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_427_ mprj_adr_o_core[20] VGND VGND VPWR VPWR _427_/Y sky130_fd_sc_hd__inv_2
XANTENNA__417__A mprj_adr_o_core[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_358_ la_oen_mprj[90] VGND VGND VPWR VPWR _358_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[72\]_B mprj_logic_high\[402\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y VGND VGND VPWR VPWR la_data_in_mprj[10]
+ sky130_fd_sc_hd__inv_8
XFILLER_13_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] mprj_logic_high\[418\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[88\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[63\]_B mprj_logic_high\[393\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[114\]_TE la_buf\[114\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[29\]_TE mprj_adr_buf\[29\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[90\] VGND VGND VPWR VPWR la_buf\[16\]/TE mprj_logic_high\[90\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y VGND VGND VPWR VPWR la_data_in_mprj[2]
+ sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[277\] VGND VGND VPWR VPWR mprj_logic_high\[277\]/HI mprj_logic_high\[277\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[444\] VGND VGND VPWR VPWR mprj_logic_high\[444\]/HI mprj_logic_high\[444\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[54\]_B mprj_logic_high\[384\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xla_buf\[14\] _485_/Y la_buf\[14\]/TE VGND VGND VPWR VPWR la_data_in_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_3_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[61\]_TE mprj_logic_high\[263\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[7\] _414_/Y mprj_adr_buf\[7\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_20_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y VGND VGND VPWR VPWR la_data_in_mprj[58]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[8\]_A _447_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[45\]_B mprj_logic_high\[375\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__610__A la_oen_mprj[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] mprj_logic_high\[444\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[114\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[30\]_A user_to_mprj_in_gates\[30\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[36\]_B mprj_logic_high\[366\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[97\]_A user_to_mprj_in_gates\[97\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_B mprj_logic_high\[450\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[70\]_A _541_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high\[286\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[124\] _392_/Y mprj_logic_high\[326\]/HI VGND VGND VPWR
+ VPWR la_oen_core[124] sky130_fd_sc_hd__einvp_8
XANTENNA__520__A la_data_out_mprj[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[54\] _653_/Y mprj_logic_high\[256\]/HI VGND VGND VPWR VPWR
+ la_oen_core[54] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[21\]_A user_to_mprj_in_gates\[21\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[394\] VGND VGND VPWR VPWR mprj_logic_high\[394\]/HI mprj_logic_high\[394\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[124\]_A _595_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[88\]_A user_to_mprj_in_gates\[88\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[111\]_B mprj_logic_high\[441\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_B mprj_logic_high\[357\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[61\]_A _532_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[118\] _589_/Y la_buf\[118\]/TE VGND VGND VPWR VPWR la_data_in_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[111] sky130_fd_sc_hd__inv_8
XANTENNA__430__A mprj_adr_o_core[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[12\]_A user_to_mprj_in_gates\[12\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[126\]_A user_to_mprj_in_gates\[126\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[115\]_A _586_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__605__A la_oen_mprj[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[79\]_A user_to_mprj_in_gates\[79\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[102\]_B mprj_logic_high\[432\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_B mprj_logic_high\[348\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[52\]_A _523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__340__A la_oen_mprj[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[117\]_A user_to_mprj_in_gates\[117\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[53\] VGND VGND VPWR VPWR mprj_dat_buf\[11\]/TE mprj_logic_high\[53\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__515__A la_data_out_mprj[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[106\]_A _577_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[43\]_A _514_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[142\] VGND VGND VPWR VPWR la_buf\[68\]/TE mprj_logic_high\[142\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[407\] VGND VGND VPWR VPWR mprj_logic_high\[407\]/HI mprj_logic_high\[407\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[81\] _552_/Y la_buf\[81\]/TE VGND VGND VPWR VPWR la_data_in_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_5_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[108\]_A user_to_mprj_in_gates\[108\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__425__A mprj_adr_o_core[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[34\]_A _505_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] mprj_logic_high\[400\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[70\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_clk_buf _398_/Y mprj_clk_buf/TE VGND VGND VPWR VPWR user_clock sky130_fd_sc_hd__einvp_8
XFILLER_17_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__335__A la_oen_mprj[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[25\]_A _496_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[110\]_A _378_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_460_ mprj_dat_o_core[21] VGND VGND VPWR VPWR _460_/Y sky130_fd_sc_hd__inv_2
X_391_ la_oen_mprj[123] VGND VGND VPWR VPWR _391_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[17\] _616_/Y mprj_logic_high\[219\]/HI VGND VGND VPWR VPWR
+ la_oen_core[17] sky130_fd_sc_hd__einvp_8
XFILLER_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[357\] VGND VGND VPWR VPWR mprj_logic_high\[357\]/HI mprj_logic_high\[357\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[16\]_A _487_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[101\]_A _369_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_658_ la_oen_mprj[59] VGND VGND VPWR VPWR _658_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_589_ la_data_out_mprj[118] VGND VGND VPWR VPWR _589_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y VGND VGND VPWR VPWR la_data_in_mprj[40]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[10\]_TE la_buf\[10\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high\[321\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_A _362_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[16\] VGND VGND VPWR VPWR mprj_adr_buf\[6\]/TE mprj_logic_high\[16\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[105\] VGND VGND VPWR VPWR la_buf\[31\]/TE mprj_logic_high\[105\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_512_ VPWR VGND VGND VPWR VPWR _512_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[33\]_TE la_buf\[33\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_443_ mprj_dat_o_core[4] VGND VGND VPWR VPWR _443_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high\[220\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_374_ la_oen_mprj[106] VGND VGND VPWR VPWR _374_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_A _353_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xla_buf\[44\] _515_/Y la_buf\[44\]/TE VGND VGND VPWR VPWR la_data_in_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[100\] _571_/Y la_buf\[100\]/TE VGND VGND VPWR VPWR la_data_in_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_1_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y VGND VGND VPWR VPWR la_data_in_mprj[88]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] mprj_logic_high\[363\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[33\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[76\]_A _344_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[1\]_TE la_buf\[1\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__613__A la_oen_mprj[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[56\]_TE la_buf\[56\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[67\]_A _335_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__523__A la_data_out_mprj[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[84\] _352_/Y mprj_logic_high\[286\]/HI VGND VGND VPWR VPWR
+ la_oen_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_2_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[222\] VGND VGND VPWR VPWR mprj_logic_high\[222\]/HI mprj_logic_high\[222\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_426_ mprj_adr_o_core[19] VGND VGND VPWR VPWR _426_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[58\]_A _657_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_357_ la_oen_mprj[89] VGND VGND VPWR VPWR _357_/Y sky130_fd_sc_hd__inv_2
XANTENNA__433__A mprj_adr_o_core[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[79\]_TE la_buf\[79\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__608__A la_oen_mprj[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[49\]_A _648_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__343__A la_oen_mprj[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[83\] VGND VGND VPWR VPWR la_buf\[9\]/TE mprj_logic_high\[83\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__518__A la_data_out_mprj[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[7\]_TE mprj_logic_high\[209\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[172\] VGND VGND VPWR VPWR la_buf\[98\]/TE mprj_logic_high\[172\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[437\] VGND VGND VPWR VPWR mprj_logic_high\[437\]/HI mprj_logic_high\[437\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__428__A mprj_adr_o_core[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_409_ mprj_adr_o_core[2] VGND VGND VPWR VPWR _409_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[27\]_A _434_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[0\] VGND VGND VPWR VPWR mprj_rstn_buf/TE mprj_logic_high\[0\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_mprj_sel_buf\[2\]_TE mprj_sel_buf\[2\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] mprj_logic_high\[437\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[107\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__338__A la_oen_mprj[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[4\]_A _603_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[18\]_A _425_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[117\] _385_/Y mprj_logic_high\[319\]/HI VGND VGND VPWR
+ VPWR la_oen_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_5_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[47\] _646_/Y mprj_logic_high\[249\]/HI VGND VGND VPWR VPWR
+ la_oen_core[47] sky130_fd_sc_hd__einvp_8
XFILLER_5_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[387\] VGND VGND VPWR VPWR mprj_logic_high\[387\]/HI mprj_logic_high\[387\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[104] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y VGND VGND VPWR VPWR la_data_in_mprj[70]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[104\]_TE la_buf\[104\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[19\]_TE mprj_adr_buf\[19\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__621__A la_oen_mprj[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[3\] _442_/Y mprj_dat_buf\[3\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[51\]_TE mprj_logic_high\[253\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[46\] VGND VGND VPWR VPWR mprj_dat_buf\[4\]/TE mprj_logic_high\[46\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[135\] VGND VGND VPWR VPWR la_buf\[61\]/TE mprj_logic_high\[135\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__531__A la_data_out_mprj[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[7\]_TE mprj_dat_buf\[7\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[302\] VGND VGND VPWR VPWR mprj_logic_high\[302\]/HI mprj_logic_high\[302\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[74\] _545_/Y la_buf\[74\]/TE VGND VGND VPWR VPWR la_data_in_core[74] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[127\]_TE la_buf\[127\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__441__A mprj_dat_o_core[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] mprj_logic_high\[393\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[63\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high\[276\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__616__A la_oen_mprj[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[3\]_A _410_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__351__A VPWR VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_390_ la_oen_mprj[122] VGND VGND VPWR VPWR _390_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__526__A la_data_out_mprj[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[252\] VGND VGND VPWR VPWR mprj_logic_high\[252\]/HI mprj_logic_high\[252\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high\[299\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_657_ la_oen_mprj[58] VGND VGND VPWR VPWR _657_/Y sky130_fd_sc_hd__inv_2
X_588_ la_data_out_mprj[117] VGND VGND VPWR VPWR _588_/Y sky130_fd_sc_hd__inv_2
XANTENNA__436__A mprj_adr_o_core[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y VGND VGND VPWR VPWR la_data_in_mprj[33]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__346__A la_oen_mprj[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_511_ la_data_out_mprj[40] VGND VGND VPWR VPWR _511_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_442_ mprj_dat_o_core[3] VGND VGND VPWR VPWR _442_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_373_ la_oen_mprj[105] VGND VGND VPWR VPWR _373_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[37\] _508_/Y la_buf\[37\]/TE VGND VGND VPWR VPWR la_data_in_core[37] sky130_fd_sc_hd__einvp_8
XFILLER_10_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_A _480_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] mprj_logic_high\[356\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[26\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[3\]_B mprj_logic_high\[333\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[77\] _345_/Y mprj_logic_high\[279\]/HI VGND VGND VPWR VPWR
+ la_oen_core[77] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[25\] _464_/Y mprj_dat_buf\[25\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[25]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[215\] VGND VGND VPWR VPWR mprj_logic_high\[215\]/HI mprj_logic_high\[215\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_425_ mprj_adr_o_core[18] VGND VGND VPWR VPWR _425_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_356_ la_oen_mprj[88] VGND VGND VPWR VPWR _356_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[20\] _427_/Y mprj_adr_buf\[20\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XFILLER_10_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high\[311\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[7\]_A user_to_mprj_in_gates\[7\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__624__A la_oen_mprj[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_TE la_buf\[23\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[76\] VGND VGND VPWR VPWR la_buf\[2\]/TE mprj_logic_high\[76\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__534__A la_data_out_mprj[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[165\] VGND VGND VPWR VPWR la_buf\[91\]/TE mprj_logic_high\[165\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[332\] VGND VGND VPWR VPWR mprj_logic_high\[332\]/HI mprj_logic_high\[332\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_408_ mprj_adr_o_core[1] VGND VGND VPWR VPWR _408_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__444__A mprj_dat_o_core[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_339_ la_oen_mprj[71] VGND VGND VPWR VPWR _339_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[46\]_TE la_buf\[46\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] mprj_logic_high\[423\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[93\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__619__A la_oen_mprj[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__354__A la_oen_mprj[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__529__A la_data_out_mprj[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[282\] VGND VGND VPWR VPWR mprj_logic_high\[282\]/HI mprj_logic_high\[282\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[69\]_TE la_buf\[69\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__439__A mprj_dat_o_core[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y VGND VGND VPWR VPWR la_data_in_mprj[63]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[18\]_TE mprj_dat_buf\[18\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__349__A la_oen_mprj[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[39\] VGND VGND VPWR VPWR mprj_adr_buf\[29\]/TE mprj_logic_high\[39\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[128\] VGND VGND VPWR VPWR la_buf\[54\]/TE mprj_logic_high\[128\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[67\] _538_/Y la_buf\[67\]/TE VGND VGND VPWR VPWR la_data_in_core[67] sky130_fd_sc_hd__einvp_8
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[123\] _594_/Y la_buf\[123\]/TE VGND VGND VPWR VPWR la_data_in_core[123] sky130_fd_sc_hd__einvp_8
XFILLER_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] mprj_logic_high\[386\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[56\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__632__A la_oen_mprj[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__542__A la_data_out_mprj[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[245\] VGND VGND VPWR VPWR mprj_logic_high\[245\]/HI mprj_logic_high\[245\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[412\] VGND VGND VPWR VPWR mprj_logic_high\[412\]/HI mprj_logic_high\[412\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_656_ la_oen_mprj[57] VGND VGND VPWR VPWR _656_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_587_ la_data_out_mprj[116] VGND VGND VPWR VPWR _587_/Y sky130_fd_sc_hd__inv_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y VGND VGND VPWR VPWR la_data_in_mprj[26]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__452__A mprj_dat_o_core[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[41\]_TE mprj_logic_high\[243\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__627__A la_oen_mprj[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_B mprj_logic_high\[423\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__362__A la_oen_mprj[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[117\]_TE la_buf\[117\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_510_ la_data_out_mprj[39] VGND VGND VPWR VPWR _510_/Y sky130_fd_sc_hd__inv_2
X_441_ mprj_dat_o_core[2] VGND VGND VPWR VPWR _441_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[195\] VGND VGND VPWR VPWR la_buf\[121\]/TE mprj_logic_high\[195\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__537__A la_data_out_mprj[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[4\] _603_/Y mprj_logic_high\[206\]/HI VGND VGND VPWR VPWR
+ la_oen_core[4] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[22\] _621_/Y mprj_logic_high\[224\]/HI VGND VGND VPWR VPWR
+ la_oen_core[22] sky130_fd_sc_hd__einvp_8
X_372_ la_oen_mprj[104] VGND VGND VPWR VPWR _372_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[362\] VGND VGND VPWR VPWR mprj_logic_high\[362\]/HI mprj_logic_high\[362\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B mprj_logic_high\[414\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[64\]_TE mprj_logic_high\[266\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_639_ la_oen_mprj[40] VGND VGND VPWR VPWR _639_/Y sky130_fd_sc_hd__inv_2
XANTENNA__447__A mprj_dat_o_core[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] mprj_logic_high\[349\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[19\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[75\]_B mprj_logic_high\[405\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[60\]_A user_to_mprj_in_gates\[60\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__357__A la_oen_mprj[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[66\]_B mprj_logic_high\[396\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high\[289\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[21\] VGND VGND VPWR VPWR mprj_adr_buf\[11\]/TE mprj_logic_high\[21\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[110\] VGND VGND VPWR VPWR la_buf\[36\]/TE mprj_logic_high\[110\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[51\]_A user_to_mprj_in_gates\[51\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[18\] _457_/Y mprj_dat_buf\[18\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[18]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[208\] VGND VGND VPWR VPWR mprj_logic_high\[208\]/HI mprj_logic_high\[208\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_424_ mprj_adr_o_core[17] VGND VGND VPWR VPWR _424_/Y sky130_fd_sc_hd__inv_2
X_355_ la_oen_mprj[87] VGND VGND VPWR VPWR _355_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_B mprj_logic_high\[387\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[91\]_A _562_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[13\] _420_/Y mprj_adr_buf\[13\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[13]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[127] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y VGND VGND VPWR VPWR la_data_in_mprj[93]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_buffers\[42\]_A user_to_mprj_in_gates\[42\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[48\]_B mprj_logic_high\[378\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[82\]_A _553_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__640__A la_oen_mprj[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] mprj_logic_high\[330\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[0\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[33\]_A user_to_mprj_in_gates\[33\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[69\] VGND VGND VPWR VPWR mprj_dat_buf\[27\]/TE mprj_logic_high\[69\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[123\]_B mprj_logic_high\[453\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[39\]_B mprj_logic_high\[369\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[73\]_A _544_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[158\] VGND VGND VPWR VPWR la_buf\[84\]/TE mprj_logic_high\[158\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__550__A la_data_out_mprj[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[325\] VGND VGND VPWR VPWR mprj_logic_high\[325\]/HI mprj_logic_high\[325\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[24\]_A user_to_mprj_in_gates\[24\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[97\] _568_/Y la_buf\[97\]/TE VGND VGND VPWR VPWR la_data_in_core[97] sky130_fd_sc_hd__einvp_8
XFILLER_4_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[127\]_A _598_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_407_ mprj_adr_o_core[0] VGND VGND VPWR VPWR _407_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_338_ la_oen_mprj[70] VGND VGND VPWR VPWR _338_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[114\]_B mprj_logic_high\[444\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[64\]_A _535_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__460__A mprj_dat_o_core[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] mprj_logic_high\[416\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[86\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[15\]_A user_to_mprj_in_gates\[15\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__635__A la_oen_mprj[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[118\]_A _589_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[105\]_B mprj_logic_high\[435\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[55\]_A _526_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__370__A la_oen_mprj[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y VGND VGND VPWR VPWR la_data_in_mprj[0]
+ sky130_fd_sc_hd__inv_8
XANTENNA__545__A la_data_out_mprj[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[109\]_A _580_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[275\] VGND VGND VPWR VPWR mprj_logic_high\[275\]/HI mprj_logic_high\[275\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[46\]_A _517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[442\] VGND VGND VPWR VPWR mprj_logic_high\[442\]/HI mprj_logic_high\[442\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[12\] _483_/Y la_buf\[12\]/TE VGND VGND VPWR VPWR la_data_in_core[12] sky130_fd_sc_hd__einvp_8
Xla_buf\[8\] _479_/Y la_buf\[8\]/TE VGND VGND VPWR VPWR la_data_in_core[8] sky130_fd_sc_hd__einvp_8
XFILLER_10_1731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[5\] _412_/Y mprj_adr_buf\[5\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y VGND VGND VPWR VPWR la_data_in_mprj[56]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[13\]_TE la_buf\[13\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__455__A mprj_dat_o_core[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[37\]_A _508_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[122\]_A _390_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] mprj_logic_high\[442\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[112\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__365__A la_oen_mprj[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[28\]_A _499_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[113\]_A _381_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[122\] _390_/Y mprj_logic_high\[324\]/HI VGND VGND VPWR
+ VPWR la_oen_core[122] sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[3\] _406_/Y mprj_sel_buf\[3\]/TE VGND VGND VPWR VPWR mprj_sel_o_user[3]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[52\] _651_/Y mprj_logic_high\[254\]/HI VGND VGND VPWR VPWR
+ la_oen_core[52] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[36\]_TE la_buf\[36\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[392\] VGND VGND VPWR VPWR mprj_logic_high\[392\]/HI mprj_logic_high\[392\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[19\]_A _490_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[116\] _587_/Y la_buf\[116\]/TE VGND VGND VPWR VPWR la_data_in_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_10_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[104\]_A _372_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk2_buf_A _399_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] mprj_logic_high\[379\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[49\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[4\]_TE la_buf\[4\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[30\]_A _629_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[59\]_TE la_buf\[59\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_A _365_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[51\] VGND VGND VPWR VPWR mprj_dat_buf\[9\]/TE mprj_logic_high\[51\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[238\] VGND VGND VPWR VPWR mprj_logic_high\[238\]/HI mprj_logic_high\[238\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[140\] VGND VGND VPWR VPWR la_buf\[66\]/TE mprj_logic_high\[140\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[21\]_A _620_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[405\] VGND VGND VPWR VPWR mprj_logic_high\[405\]/HI mprj_logic_high\[405\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_655_ la_oen_mprj[56] VGND VGND VPWR VPWR _655_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[88\]_A _356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_586_ la_data_out_mprj[115] VGND VGND VPWR VPWR _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y VGND VGND VPWR VPWR VPWR
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_oen_buffers\[12\]_A _611_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[79\]_A _347_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__643__A la_oen_mprj[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[99\] VGND VGND VPWR VPWR la_buf\[25\]/TE mprj_logic_high\[99\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_440_ mprj_dat_o_core[1] VGND VGND VPWR VPWR _440_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[188\] VGND VGND VPWR VPWR la_buf\[114\]/TE mprj_logic_high\[188\]/LO
+ sky130_fd_sc_hd__conb_1
X_371_ la_oen_mprj[103] VGND VGND VPWR VPWR _371_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[15\] _614_/Y mprj_logic_high\[217\]/HI VGND VGND VPWR VPWR
+ la_oen_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_9_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__553__A la_data_out_mprj[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[355\] VGND VGND VPWR VPWR mprj_logic_high\[355\]/HI mprj_logic_high\[355\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_638_ la_oen_mprj[39] VGND VGND VPWR VPWR _638_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_569_ la_data_out_mprj[98] VGND VGND VPWR VPWR _569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__463__A mprj_dat_o_core[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__638__A la_oen_mprj[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[30\]_A _469_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__373__A la_oen_mprj[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[14\] VGND VGND VPWR VPWR mprj_adr_buf\[4\]/TE mprj_logic_high\[14\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[103\] VGND VGND VPWR VPWR la_buf\[29\]/TE mprj_logic_high\[103\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__548__A la_data_out_mprj[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_423_ mprj_adr_o_core[16] VGND VGND VPWR VPWR _423_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_A _460_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[42\] _513_/Y la_buf\[42\]/TE VGND VGND VPWR VPWR la_data_in_core[42] sky130_fd_sc_hd__einvp_8
X_354_ la_oen_mprj[86] VGND VGND VPWR VPWR _354_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[31\]_TE mprj_logic_high\[233\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y VGND VGND VPWR VPWR la_data_in_mprj[86]
+ sky130_fd_sc_hd__inv_8
XANTENNA__458__A mprj_dat_o_core[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[107\]_TE la_buf\[107\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] mprj_logic_high\[361\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[31\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[12\]_A _451_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[6\]_TE mprj_adr_buf\[6\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__368__A la_oen_mprj[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[7\]_A _606_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_TE mprj_logic_high\[256\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[82\] _350_/Y mprj_logic_high\[284\]/HI VGND VGND VPWR VPWR
+ la_oen_core[82] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[318\] VGND VGND VPWR VPWR mprj_logic_high\[318\]/HI mprj_logic_high\[318\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[30\] _469_/Y mprj_dat_buf\[30\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[220\] VGND VGND VPWR VPWR mprj_logic_high\[220\]/HI mprj_logic_high\[220\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_406_ mprj_sel_o_core[3] VGND VGND VPWR VPWR _406_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_337_ la_oen_mprj[69] VGND VGND VPWR VPWR _337_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] mprj_logic_high\[409\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[79\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[92\]_TE la_buf\[92\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high\[279\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__651__A la_oen_mprj[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_cyc_buf_TE mprj_cyc_buf/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[81\] VGND VGND VPWR VPWR la_buf\[7\]/TE mprj_logic_high\[81\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[170\] VGND VGND VPWR VPWR la_buf\[96\]/TE mprj_logic_high\[170\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[268\] VGND VGND VPWR VPWR mprj_logic_high\[268\]/HI mprj_logic_high\[268\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__561__A la_data_out_mprj[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[435\] VGND VGND VPWR VPWR mprj_logic_high\[435\]/HI mprj_logic_high\[435\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y VGND VGND VPWR VPWR la_data_in_mprj[49]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__471__A la_data_out_mprj[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] mprj_logic_high\[435\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[105\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__646__A la_oen_mprj[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[6\]_A _413_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__381__A la_oen_mprj[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[115\] _383_/Y mprj_logic_high\[317\]/HI VGND VGND VPWR
+ VPWR la_oen_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_0_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[45\] _644_/Y mprj_logic_high\[247\]/HI VGND VGND VPWR VPWR
+ la_oen_core[45] sky130_fd_sc_hd__einvp_8
XFILLER_17_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[385\] VGND VGND VPWR VPWR mprj_logic_high\[385\]/HI mprj_logic_high\[385\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__556__A la_data_out_mprj[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[109\] _580_/Y la_buf\[109\]/TE VGND VGND VPWR VPWR la_data_in_core[109] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[102] sky130_fd_sc_hd__inv_8
XFILLER_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__466__A mprj_dat_o_core[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[1\] _440_/Y mprj_dat_buf\[1\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__376__A la_oen_mprj[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[44\] VGND VGND VPWR VPWR mprj_dat_buf\[2\]/TE mprj_logic_high\[44\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[133\] VGND VGND VPWR VPWR la_buf\[59\]/TE mprj_logic_high\[133\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[300\] VGND VGND VPWR VPWR mprj_logic_high\[300\]/HI mprj_logic_high\[300\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_654_ la_oen_mprj[55] VGND VGND VPWR VPWR _654_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[72\] _543_/Y la_buf\[72\]/TE VGND VGND VPWR VPWR la_data_in_core[72] sky130_fd_sc_hd__einvp_8
X_585_ la_data_out_mprj[114] VGND VGND VPWR VPWR _585_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] mprj_logic_high\[391\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[61\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[26\]_TE la_buf\[26\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[6\]_B mprj_logic_high\[336\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_370_ la_oen_mprj[102] VGND VGND VPWR VPWR _370_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[348\] VGND VGND VPWR VPWR mprj_logic_high\[348\]/HI mprj_logic_high\[348\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[250\] VGND VGND VPWR VPWR mprj_logic_high\[250\]/HI mprj_logic_high\[250\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_637_ la_oen_mprj[38] VGND VGND VPWR VPWR _637_/Y sky130_fd_sc_hd__inv_2
X_568_ la_data_out_mprj[97] VGND VGND VPWR VPWR _568_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y VGND VGND VPWR VPWR la_data_in_mprj[31]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[49\]_TE la_buf\[49\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_499_ la_data_out_mprj[28] VGND VGND VPWR VPWR _499_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[9\] VGND VGND VPWR VPWR mprj_sel_buf\[3\]/TE mprj_logic_high\[9\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__654__A la_oen_mprj[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[298\] VGND VGND VPWR VPWR mprj_logic_high\[298\]/HI mprj_logic_high\[298\]/LO
+ sky130_fd_sc_hd__conb_1
X_422_ mprj_adr_o_core[15] VGND VGND VPWR VPWR _422_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__564__A la_data_out_mprj[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_353_ la_oen_mprj[85] VGND VGND VPWR VPWR _353_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xla_buf\[35\] _506_/Y la_buf\[35\]/TE VGND VGND VPWR VPWR la_data_in_core[35] sky130_fd_sc_hd__einvp_8
XFILLER_6_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y VGND VGND VPWR VPWR la_data_in_mprj[79]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__474__A la_data_out_mprj[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] mprj_logic_high\[354\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[24\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__649__A la_oen_mprj[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__384__A la_oen_mprj[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[75\] _343_/Y mprj_logic_high\[277\]/HI VGND VGND VPWR VPWR
+ la_oen_core[75] sky130_fd_sc_hd__einvp_8
XFILLER_2_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[213\] VGND VGND VPWR VPWR mprj_logic_high\[213\]/HI mprj_logic_high\[213\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[23\] _462_/Y mprj_dat_buf\[23\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__559__A la_data_out_mprj[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ mprj_sel_o_core[2] VGND VGND VPWR VPWR _405_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_336_ la_oen_mprj[68] VGND VGND VPWR VPWR _336_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__469__A mprj_dat_o_core[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high\[324\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__379__A la_oen_mprj[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[21\]_TE mprj_logic_high\[223\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[74\] VGND VGND VPWR VPWR la_buf\[0\]/TE mprj_logic_high\[74\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[163\] VGND VGND VPWR VPWR la_buf\[89\]/TE mprj_logic_high\[163\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[428\] VGND VGND VPWR VPWR mprj_logic_high\[428\]/HI mprj_logic_high\[428\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[330\] VGND VGND VPWR VPWR mprj_logic_high\[330\]/HI mprj_logic_high\[330\]/LO
+ sky130_fd_sc_hd__conb_1
Xpowergood_check mprj2_pwrgood/A mprj_vdd_pwrgood/A powergood_check/VPWR powergood_check/VGND
+ mgmt_protect_hv
XFILLER_15_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] mprj_logic_high\[421\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[91\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[44\]_TE mprj_logic_high\[246\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[0\]_A _403_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[108\] _376_/Y mprj_logic_high\[310\]/HI VGND VGND VPWR
+ VPWR la_oen_core[108] sky130_fd_sc_hd__einvp_8
XFILLER_5_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[38\] _637_/Y mprj_logic_high\[240\]/HI VGND VGND VPWR VPWR
+ la_oen_core[38] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[280\] VGND VGND VPWR VPWR mprj_logic_high\[280\]/HI mprj_logic_high\[280\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[378\] VGND VGND VPWR VPWR mprj_logic_high\[378\]/HI mprj_logic_high\[378\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__572__A la_data_out_mprj[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[82\]_TE la_buf\[82\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[1\]_A _440_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[67\]_TE mprj_logic_high\[269\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y VGND VGND VPWR VPWR la_data_in_mprj[61]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__482__A la_data_out_mprj[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[90\]_A user_to_mprj_in_gates\[90\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__657__A la_oen_mprj[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[96\]_B mprj_logic_high\[426\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__392__A la_oen_mprj[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[37\] VGND VGND VPWR VPWR mprj_adr_buf\[27\]/TE mprj_logic_high\[37\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[126\] VGND VGND VPWR VPWR la_buf\[52\]/TE mprj_logic_high\[126\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[81\]_A user_to_mprj_in_gates\[81\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[20\]_B mprj_logic_high\[350\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__567__A la_data_out_mprj[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_653_ la_oen_mprj[54] VGND VGND VPWR VPWR _653_/Y sky130_fd_sc_hd__inv_2
X_584_ la_data_out_mprj[113] VGND VGND VPWR VPWR _584_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[65\] _536_/Y la_buf\[65\]/TE VGND VGND VPWR VPWR la_data_in_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[87\]_B mprj_logic_high\[417\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[29\] _436_/Y mprj_adr_buf\[29\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[29]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[121\] _592_/Y la_buf\[121\]/TE VGND VGND VPWR VPWR la_data_in_core[121] sky130_fd_sc_hd__einvp_8
XFILLER_4_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[72\]_A user_to_mprj_in_gates\[72\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_B mprj_logic_high\[341\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__477__A la_data_out_mprj[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] mprj_logic_high\[384\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[54\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[78\]_B mprj_logic_high\[408\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[110\]_A user_to_mprj_in_gates\[110\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[63\]_A user_to_mprj_in_gates\[63\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__387__A la_oen_mprj[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[69\]_B mprj_logic_high\[399\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[243\] VGND VGND VPWR VPWR mprj_logic_high\[243\]/HI mprj_logic_high\[243\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[101\]_A user_to_mprj_in_gates\[101\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[410\] VGND VGND VPWR VPWR mprj_logic_high\[410\]/HI mprj_logic_high\[410\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[54\]_A user_to_mprj_in_gates\[54\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_636_ la_oen_mprj[37] VGND VGND VPWR VPWR _636_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_567_ la_data_out_mprj[96] VGND VGND VPWR VPWR _567_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_498_ la_data_out_mprj[27] VGND VGND VPWR VPWR _498_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[94\]_A _565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y VGND VGND VPWR VPWR la_data_in_mprj[24]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[45\]_A user_to_mprj_in_gates\[45\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[85\]_A _556_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[36\]_A user_to_mprj_in_gates\[36\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[193\] VGND VGND VPWR VPWR la_buf\[119\]/TE mprj_logic_high\[193\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[2\] _601_/Y mprj_logic_high\[204\]/HI VGND VGND VPWR VPWR
+ la_oen_core[2] sky130_fd_sc_hd__einvp_8
X_421_ mprj_adr_o_core[14] VGND VGND VPWR VPWR _421_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[20\] _619_/Y mprj_logic_high\[222\]/HI VGND VGND VPWR VPWR
+ la_oen_core[20] sky130_fd_sc_hd__einvp_8
X_352_ la_oen_mprj[84] VGND VGND VPWR VPWR _352_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[126\]_B mprj_logic_high\[456\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[76\]_A _547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[458\] VGND VGND VPWR VPWR mprj_pwrgood/A mprj_logic_high\[458\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[360\] VGND VGND VPWR VPWR mprj_logic_high\[360\]/HI mprj_logic_high\[360\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__580__A la_data_out_mprj[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[28\] _499_/Y la_buf\[28\]/TE VGND VGND VPWR VPWR la_data_in_core[28] sky130_fd_sc_hd__einvp_8
XFILLER_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[27\]_A user_to_mprj_in_gates\[27\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[16\]_TE la_buf\[16\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_619_ la_oen_mprj[20] VGND VGND VPWR VPWR _619_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[67\]_A _538_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_B mprj_logic_high\[447\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] mprj_logic_high\[347\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[17\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__490__A la_data_out_mprj[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[18\]_A user_to_mprj_in_gates\[18\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[58\]_A _529_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_B mprj_logic_high\[438\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[68\] _336_/Y mprj_logic_high\[270\]/HI VGND VGND VPWR VPWR
+ la_oen_core[68] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[16\] _455_/Y mprj_dat_buf\[16\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[39\]_TE la_buf\[39\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[206\] VGND VGND VPWR VPWR mprj_logic_high\[206\]/HI mprj_logic_high\[206\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__575__A la_data_out_mprj[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[49\]_A _520_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_404_ mprj_sel_o_core[1] VGND VGND VPWR VPWR _404_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ la_oen_mprj[67] VGND VGND VPWR VPWR _335_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[11\] _418_/Y mprj_adr_buf\[11\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[11]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[125] sky130_fd_sc_hd__inv_8
XFILLER_2_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y VGND VGND VPWR VPWR la_data_in_mprj[91]
+ sky130_fd_sc_hd__inv_8
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__485__A la_data_out_mprj[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[7\]_TE la_buf\[7\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_A _659_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[125\]_A _393_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__395__A la_oen_mprj[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[67\] VGND VGND VPWR VPWR mprj_dat_buf\[25\]/TE mprj_logic_high\[67\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[156\] VGND VGND VPWR VPWR la_buf\[82\]/TE mprj_logic_high\[156\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[51\]_A _650_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[116\]_A _384_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[323\] VGND VGND VPWR VPWR mprj_logic_high\[323\]/HI mprj_logic_high\[323\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[95\] _566_/Y la_buf\[95\]/TE VGND VGND VPWR VPWR la_data_in_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_8_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[107\]_A _375_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[42\]_A _641_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] mprj_logic_high\[414\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[84\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[33\]_A _632_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[273\] VGND VGND VPWR VPWR mprj_logic_high\[273\]/HI mprj_logic_high\[273\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[440\] VGND VGND VPWR VPWR mprj_logic_high\[440\]/HI mprj_logic_high\[440\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[112\]_TE mprj_logic_high\[314\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[6\] _477_/Y la_buf\[6\]/TE VGND VGND VPWR VPWR la_data_in_core[6] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[24\]_A _623_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[10\] _481_/Y la_buf\[10\]/TE VGND VGND VPWR VPWR la_data_in_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_4_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[3\] _410_/Y mprj_adr_buf\[3\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_we_buf_TE mprj_we_buf/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[20\]_A _427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y VGND VGND VPWR VPWR la_data_in_mprj[54]
+ sky130_fd_sc_hd__inv_8
XFILLER_16_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high\[213\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[15\]_A _614_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] mprj_logic_high\[440\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[110\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[11\]_A _418_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[120\] _388_/Y mprj_logic_high\[322\]/HI VGND VGND VPWR
+ VPWR la_oen_core[120] sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[1\] _404_/Y mprj_sel_buf\[1\]/TE VGND VGND VPWR VPWR mprj_sel_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[119\] VGND VGND VPWR VPWR la_buf\[45\]/TE mprj_logic_high\[119\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[50\] _649_/Y mprj_logic_high\[252\]/HI VGND VGND VPWR VPWR
+ la_oen_core[50] sky130_fd_sc_hd__einvp_8
X_652_ la_oen_mprj[53] VGND VGND VPWR VPWR _652_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[390\] VGND VGND VPWR VPWR mprj_logic_high\[390\]/HI mprj_logic_high\[390\]/LO
+ sky130_fd_sc_hd__conb_1
X_583_ la_data_out_mprj[112] VGND VGND VPWR VPWR _583_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__583__A la_data_out_mprj[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[58\] _529_/Y la_buf\[58\]/TE VGND VGND VPWR VPWR la_data_in_core[58] sky130_fd_sc_hd__einvp_8
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[34\]_TE mprj_logic_high\[236\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xla_buf\[114\] _585_/Y la_buf\[114\]/TE VGND VGND VPWR VPWR la_data_in_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_10_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] mprj_logic_high\[377\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[47\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__493__A la_data_out_mprj[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[9\]_TE mprj_adr_buf\[9\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] mprj_logic_high\[339\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[9\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[72\]_TE la_buf\[72\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[57\]_TE mprj_logic_high\[259\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[98\] _366_/Y mprj_logic_high\[300\]/HI VGND VGND VPWR VPWR
+ la_oen_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_5_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[236\] VGND VGND VPWR VPWR mprj_logic_high\[236\]/HI mprj_logic_high\[236\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[403\] VGND VGND VPWR VPWR mprj_logic_high\[403\]/HI mprj_logic_high\[403\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__578__A la_data_out_mprj[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[24\]_A _463_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_635_ la_oen_mprj[36] VGND VGND VPWR VPWR _635_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_566_ la_data_out_mprj[95] VGND VGND VPWR VPWR _566_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_497_ la_data_out_mprj[26] VGND VGND VPWR VPWR _497_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[0\]_TE mprj_logic_high\[202\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y VGND VGND VPWR VPWR la_data_in_mprj[17]
+ sky130_fd_sc_hd__inv_8
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_TE la_buf\[95\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__488__A la_data_out_mprj[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[15\]_A _454_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__398__A caravel_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[97\] VGND VGND VPWR VPWR la_buf\[23\]/TE mprj_logic_high\[97\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_420_ mprj_adr_o_core[13] VGND VGND VPWR VPWR _420_/Y sky130_fd_sc_hd__inv_2
X_351_ VPWR VGND VGND VPWR VPWR _351_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[13\] _612_/Y mprj_logic_high\[215\]/HI VGND VGND VPWR VPWR
+ la_oen_core[13] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y VGND VGND VPWR VPWR la_data_in_mprj[9]
+ sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[186\] VGND VGND VPWR VPWR la_buf\[112\]/TE mprj_logic_high\[186\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[353\] VGND VGND VPWR VPWR mprj_logic_high\[353\]/HI mprj_logic_high\[353\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_618_ la_oen_mprj[19] VGND VGND VPWR VPWR _618_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_549_ la_data_out_mprj[78] VGND VGND VPWR VPWR _549_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[12\] VGND VGND VPWR VPWR mprj_adr_buf\[2\]/TE mprj_logic_high\[12\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[101\] VGND VGND VPWR VPWR la_buf\[27\]/TE mprj_logic_high\[101\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_403_ mprj_sel_o_core[0] VGND VGND VPWR VPWR _403_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[2\]_A _473_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_334_ la_oen_mprj[66] VGND VGND VPWR VPWR _334_/Y sky130_fd_sc_hd__inv_2
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[40\] _511_/Y la_buf\[40\]/TE VGND VGND VPWR VPWR la_data_in_core[40] sky130_fd_sc_hd__einvp_8
XANTENNA__591__A la_data_out_mprj[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[118] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y VGND VGND VPWR VPWR la_data_in_mprj[84]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[0\]_TE mprj_dat_buf\[0\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[120\]_TE la_buf\[120\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[9\]_A _416_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[149\] VGND VGND VPWR VPWR la_buf\[75\]/TE mprj_logic_high\[149\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[80\] _348_/Y mprj_logic_high\[282\]/HI VGND VGND VPWR VPWR
+ la_oen_core[80] sky130_fd_sc_hd__einvp_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[316\] VGND VGND VPWR VPWR mprj_logic_high\[316\]/HI mprj_logic_high\[316\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__586__A la_data_out_mprj[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[88\] _559_/Y la_buf\[88\]/TE VGND VGND VPWR VPWR la_data_in_core[88] sky130_fd_sc_hd__einvp_8
XFILLER_15_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[0\]_A user_to_mprj_in_gates\[0\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] mprj_logic_high\[407\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[77\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__496__A la_data_out_mprj[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high\[292\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[29\]_TE la_buf\[29\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[266\] VGND VGND VPWR VPWR mprj_logic_high\[266\]/HI mprj_logic_high\[266\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[433\] VGND VGND VPWR VPWR mprj_logic_high\[433\]/HI mprj_logic_high\[433\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y VGND VGND VPWR VPWR la_data_in_mprj[47]
+ sky130_fd_sc_hd__inv_8
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] mprj_logic_high\[433\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[103\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_clk2_buf _399_/Y mprj_clk2_buf/TE VGND VGND VPWR VPWR user_clock2 sky130_fd_sc_hd__einvp_8
XFILLER_1_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[113\] _381_/Y mprj_logic_high\[315\]/HI VGND VGND VPWR
+ VPWR la_oen_core[113] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[9\]_B mprj_logic_high\[339\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[43\] _642_/Y mprj_logic_high\[245\]/HI VGND VGND VPWR VPWR
+ la_oen_core[43] sky130_fd_sc_hd__einvp_8
X_651_ la_oen_mprj[52] VGND VGND VPWR VPWR _651_/Y sky130_fd_sc_hd__inv_2
X_582_ la_data_out_mprj[111] VGND VGND VPWR VPWR _582_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[383\] VGND VGND VPWR VPWR mprj_logic_high\[383\]/HI mprj_logic_high\[383\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[107\] _578_/Y la_buf\[107\]/TE VGND VGND VPWR VPWR la_data_in_core[107] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[100] sky130_fd_sc_hd__inv_8
XFILLER_0_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high\[304\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[42\] VGND VGND VPWR VPWR mprj_dat_buf\[0\]/TE mprj_logic_high\[42\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[131\] VGND VGND VPWR VPWR la_buf\[57\]/TE mprj_logic_high\[131\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[229\] VGND VGND VPWR VPWR mprj_logic_high\[229\]/HI mprj_logic_high\[229\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_634_ la_oen_mprj[35] VGND VGND VPWR VPWR _634_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[70\] _541_/Y la_buf\[70\]/TE VGND VGND VPWR VPWR la_data_in_core[70] sky130_fd_sc_hd__einvp_8
XANTENNA__594__A la_data_out_mprj[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_565_ la_data_out_mprj[94] VGND VGND VPWR VPWR _565_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_496_ la_data_out_mprj[25] VGND VGND VPWR VPWR _496_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high\[327\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[24\]_TE mprj_logic_high\[226\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_350_ la_oen_mprj[82] VGND VGND VPWR VPWR _350_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[179\] VGND VGND VPWR VPWR la_buf\[105\]/TE mprj_logic_high\[179\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[346\] VGND VGND VPWR VPWR mprj_logic_high\[346\]/HI mprj_logic_high\[346\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__589__A la_data_out_mprj[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_617_ la_oen_mprj[18] VGND VGND VPWR VPWR _617_/Y sky130_fd_sc_hd__inv_2
X_548_ la_data_out_mprj[77] VGND VGND VPWR VPWR _548_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_479_ la_data_out_mprj[8] VGND VGND VPWR VPWR _479_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[62\]_TE la_buf\[62\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high\[249\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[7\] VGND VGND VPWR VPWR mprj_sel_buf\[1\]/TE mprj_logic_high\[7\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__499__A la_data_out_mprj[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[296\] VGND VGND VPWR VPWR mprj_logic_high\[296\]/HI mprj_logic_high\[296\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_402_ mprj_we_o_core VGND VGND VPWR VPWR _402_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_333_ la_oen_mprj[65] VGND VGND VPWR VPWR _333_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[85\]_TE la_buf\[85\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[33\] _504_/Y la_buf\[33\]/TE VGND VGND VPWR VPWR la_data_in_core[33] sky130_fd_sc_hd__einvp_8
XFILLER_6_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y VGND VGND VPWR VPWR la_data_in_mprj[77]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] mprj_logic_high\[352\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[22\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[3\]_A _406_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[50\]_B mprj_logic_high\[380\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[211\] VGND VGND VPWR VPWR mprj_logic_high\[211\]/HI mprj_logic_high\[211\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[73\] _341_/Y mprj_logic_high\[275\]/HI VGND VGND VPWR VPWR
+ la_oen_core[73] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[21\] _460_/Y mprj_dat_buf\[21\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[21]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[309\] VGND VGND VPWR VPWR mprj_logic_high\[309\]/HI mprj_logic_high\[309\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[4\]_A _443_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[41\]_B mprj_logic_high\[371\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[93\]_A user_to_mprj_in_gates\[93\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[32\]_B mprj_logic_high\[362\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[99\]_B mprj_logic_high\[429\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[72\] VGND VGND VPWR VPWR mprj_dat_buf\[30\]/TE mprj_logic_high\[72\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[161\] VGND VGND VPWR VPWR la_buf\[87\]/TE mprj_logic_high\[161\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[259\] VGND VGND VPWR VPWR mprj_logic_high\[259\]/HI mprj_logic_high\[259\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[120\]_A _591_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[426\] VGND VGND VPWR VPWR mprj_logic_high\[426\]/HI mprj_logic_high\[426\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[84\]_A user_to_mprj_in_gates\[84\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[23\]_B mprj_logic_high\[353\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__597__A la_data_out_mprj[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[110\]_TE la_buf\[110\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[122\]_A user_to_mprj_in_gates\[122\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[111\]_A _582_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[75\]_A user_to_mprj_in_gates\[75\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B mprj_logic_high\[344\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[113\]_A user_to_mprj_in_gates\[113\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[102\]_A _573_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[66\]_A user_to_mprj_in_gates\[66\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _374_/Y mprj_logic_high\[308\]/HI VGND VGND VPWR
+ VPWR la_oen_core[106] sky130_fd_sc_hd__einvp_8
X_650_ la_oen_mprj[51] VGND VGND VPWR VPWR _650_/Y sky130_fd_sc_hd__inv_2
X_581_ la_data_out_mprj[110] VGND VGND VPWR VPWR _581_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[36\] _635_/Y mprj_logic_high\[238\]/HI VGND VGND VPWR VPWR
+ la_oen_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[376\] VGND VGND VPWR VPWR mprj_logic_high\[376\]/HI mprj_logic_high\[376\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[104\]_A user_to_mprj_in_gates\[104\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[57\]_A user_to_mprj_in_gates\[57\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[30\]_A _501_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high\[282\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[19\]_TE la_buf\[19\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[97\]_A _568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[48\]_A user_to_mprj_in_gates\[48\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[21\]_A _492_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_A _559_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[35\] VGND VGND VPWR VPWR mprj_adr_buf\[25\]/TE mprj_logic_high\[35\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[39\]_A user_to_mprj_in_gates\[39\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[124\] VGND VGND VPWR VPWR la_buf\[50\]/TE mprj_logic_high\[124\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[12\]_A _483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_633_ la_oen_mprj[34] VGND VGND VPWR VPWR _633_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[63\] _534_/Y la_buf\[63\]/TE VGND VGND VPWR VPWR la_data_in_core[63] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[79\]_A _550_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_564_ la_data_out_mprj[93] VGND VGND VPWR VPWR _564_/Y sky130_fd_sc_hd__inv_2
X_495_ la_data_out_mprj[24] VGND VGND VPWR VPWR _495_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[27\] _434_/Y mprj_adr_buf\[27\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] mprj_logic_high\[382\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[52\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[90\]_A _358_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[81\]_A _349_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[339\] VGND VGND VPWR VPWR mprj_logic_high\[339\]/HI mprj_logic_high\[339\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[241\] VGND VGND VPWR VPWR mprj_logic_high\[241\]/HI mprj_logic_high\[241\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_616_ la_oen_mprj[17] VGND VGND VPWR VPWR _616_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_547_ la_data_out_mprj[76] VGND VGND VPWR VPWR _547_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_478_ la_data_out_mprj[7] VGND VGND VPWR VPWR _478_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y VGND VGND VPWR VPWR la_data_in_mprj[22]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_oen_buffers\[72\]_A _340_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[63\]_A _331_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_401_ mprj_stb_o_core VGND VGND VPWR VPWR _401_/Y sky130_fd_sc_hd__inv_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[191\] VGND VGND VPWR VPWR la_buf\[117\]/TE mprj_logic_high\[191\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[0\] _599_/Y mprj_logic_high\[202\]/HI VGND VGND VPWR VPWR
+ la_oen_core[0] sky130_fd_sc_hd__einvp_8
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[289\] VGND VGND VPWR VPWR mprj_logic_high\[289\]/HI mprj_logic_high\[289\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_332_ la_oen_mprj[64] VGND VGND VPWR VPWR _332_/Y sky130_fd_sc_hd__inv_2
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[456\] VGND VGND VPWR VPWR mprj_logic_high\[456\]/HI mprj_logic_high\[456\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high\[317\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_A _653_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[119\]_A _387_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[26\] _497_/Y la_buf\[26\]/TE VGND VGND VPWR VPWR la_data_in_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] mprj_logic_high\[345\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[15\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[45\]_A _644_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high\[216\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] mprj_logic_high\[456\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[126\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_A _635_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[66\] _334_/Y mprj_logic_high\[268\]/HI VGND VGND VPWR VPWR
+ la_oen_core[66] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[14\] _453_/Y mprj_dat_buf\[14\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[14]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[204\] VGND VGND VPWR VPWR mprj_logic_high\[204\]/HI mprj_logic_high\[204\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[52\]_TE la_buf\[52\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[37\]_TE mprj_logic_high\[239\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[27\]_A _626_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[123] sky130_fd_sc_hd__inv_8
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[23\]_A _430_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[0\]_A _599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[18\]_A _617_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[14\]_A _421_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[75\]_TE la_buf\[75\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[65\] VGND VGND VPWR VPWR mprj_dat_buf\[23\]/TE mprj_logic_high\[65\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[154\] VGND VGND VPWR VPWR la_buf\[80\]/TE mprj_logic_high\[154\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[321\] VGND VGND VPWR VPWR mprj_logic_high\[321\]/HI mprj_logic_high\[321\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[419\] VGND VGND VPWR VPWR mprj_logic_high\[419\]/HI mprj_logic_high\[419\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[93\] _564_/Y la_buf\[93\]/TE VGND VGND VPWR VPWR la_data_in_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high\[205\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[98\]_TE la_buf\[98\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] mprj_logic_high\[412\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[82\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_580_ la_data_out_mprj[109] VGND VGND VPWR VPWR _580_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[29\] _628_/Y mprj_logic_high\[231\]/HI VGND VGND VPWR VPWR
+ la_oen_core[29] sky130_fd_sc_hd__einvp_8
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[271\] VGND VGND VPWR VPWR mprj_logic_high\[271\]/HI mprj_logic_high\[271\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[369\] VGND VGND VPWR VPWR mprj_logic_high\[369\]/HI mprj_logic_high\[369\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[4\] _475_/Y la_buf\[4\]/TE VGND VGND VPWR VPWR la_data_in_core[4] sky130_fd_sc_hd__einvp_8
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__401__A mprj_stb_o_core VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[1\] _408_/Y mprj_adr_buf\[1\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[27\]_A _466_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y VGND VGND VPWR VPWR la_data_in_mprj[52]
+ sky130_fd_sc_hd__inv_8
XFILLER_16_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[18\]_A _457_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[100\]_TE la_buf\[100\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[28\] VGND VGND VPWR VPWR mprj_adr_buf\[18\]/TE mprj_logic_high\[28\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[117\] VGND VGND VPWR VPWR la_buf\[43\]/TE mprj_logic_high\[117\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_632_ la_oen_mprj[33] VGND VGND VPWR VPWR _632_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_563_ la_data_out_mprj[92] VGND VGND VPWR VPWR _563_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[56\] _527_/Y la_buf\[56\]/TE VGND VGND VPWR VPWR la_data_in_core[56] sky130_fd_sc_hd__einvp_8
X_494_ la_data_out_mprj[23] VGND VGND VPWR VPWR _494_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xla_buf\[112\] _583_/Y la_buf\[112\]/TE VGND VGND VPWR VPWR la_data_in_core[112] sky130_fd_sc_hd__einvp_8
XFILLER_5_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[3\]_TE mprj_dat_buf\[3\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] mprj_logic_high\[375\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[45\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[123\]_TE la_buf\[123\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] mprj_logic_high\[337\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[7\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[70\]_TE mprj_logic_high\[272\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[96\] _364_/Y mprj_logic_high\[298\]/HI VGND VGND VPWR VPWR
+ la_oen_core[96] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[234\] VGND VGND VPWR VPWR mprj_logic_high\[234\]/HI mprj_logic_high\[234\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[401\] VGND VGND VPWR VPWR mprj_logic_high\[401\]/HI mprj_logic_high\[401\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[5\]_A _476_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_615_ la_oen_mprj[16] VGND VGND VPWR VPWR _615_/Y sky130_fd_sc_hd__inv_2
X_546_ la_data_out_mprj[75] VGND VGND VPWR VPWR _546_/Y sky130_fd_sc_hd__inv_2
X_477_ la_data_out_mprj[6] VGND VGND VPWR VPWR _477_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y VGND VGND VPWR VPWR la_data_in_mprj[15]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high\[295\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj2_pwrgood mprj2_pwrgood/A VGND VGND VPWR VPWR user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_8_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[95\] VGND VGND VPWR VPWR la_buf\[21\]/TE mprj_logic_high\[95\]/LO
+ sky130_fd_sc_hd__conb_1
X_400_ mprj_cyc_o_core VGND VGND VPWR VPWR _400_/Y sky130_fd_sc_hd__inv_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[11\] _610_/Y mprj_logic_high\[213\]/HI VGND VGND VPWR VPWR
+ la_oen_core[11] sky130_fd_sc_hd__einvp_8
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ la_oen_mprj[63] VGND VGND VPWR VPWR _331_/Y sky130_fd_sc_hd__inv_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y VGND VGND VPWR VPWR la_data_in_mprj[7]
+ sky130_fd_sc_hd__inv_8
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[184\] VGND VGND VPWR VPWR la_buf\[110\]/TE mprj_logic_high\[184\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[449\] VGND VGND VPWR VPWR mprj_logic_high\[449\]/HI mprj_logic_high\[449\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[351\] VGND VGND VPWR VPWR mprj_logic_high\[351\]/HI mprj_logic_high\[351\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[19\] _490_/Y la_buf\[19\]/TE VGND VGND VPWR VPWR la_data_in_core[19] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[3\]_A user_to_mprj_in_gates\[3\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_529_ la_data_out_mprj[58] VGND VGND VPWR VPWR _529_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_vdd_pwrgood_A mprj_vdd_pwrgood/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] mprj_logic_high\[449\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[119\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[10\] VGND VGND VPWR VPWR mprj_adr_buf\[0\]/TE mprj_logic_high\[10\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[59\] _658_/Y mprj_logic_high\[261\]/HI VGND VGND VPWR VPWR
+ la_oen_core[59] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[399\] VGND VGND VPWR VPWR mprj_logic_high\[399\]/HI mprj_logic_high\[399\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__404__A mprj_sel_o_core[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[116] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y VGND VGND VPWR VPWR la_data_in_mprj[82]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_rstn_buf_A _396_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[105\]_TE mprj_logic_high\[307\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[58\] VGND VGND VPWR VPWR mprj_dat_buf\[16\]/TE mprj_logic_high\[58\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[147\] VGND VGND VPWR VPWR la_buf\[73\]/TE mprj_logic_high\[147\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[314\] VGND VGND VPWR VPWR mprj_logic_high\[314\]/HI mprj_logic_high\[314\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[86\] _557_/Y la_buf\[86\]/TE VGND VGND VPWR VPWR la_data_in_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_1_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] mprj_logic_high\[405\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[75\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[42\]_TE la_buf\[42\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high\[229\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[264\] VGND VGND VPWR VPWR mprj_logic_high\[264\]/HI mprj_logic_high\[264\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[431\] VGND VGND VPWR VPWR mprj_logic_high\[431\]/HI mprj_logic_high\[431\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y VGND VGND VPWR VPWR la_data_in_mprj[45]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[65\]_TE la_buf\[65\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] mprj_logic_high\[431\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[101\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[14\]_TE mprj_dat_buf\[14\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__502__A la_data_out_mprj[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[111\] _379_/Y mprj_logic_high\[313\]/HI VGND VGND VPWR
+ VPWR la_oen_core[111] sky130_fd_sc_hd__einvp_8
X_631_ la_oen_mprj[32] VGND VGND VPWR VPWR _631_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[41\] _640_/Y mprj_logic_high\[243\]/HI VGND VGND VPWR VPWR
+ la_oen_core[41] sky130_fd_sc_hd__einvp_8
XFILLER_2_1820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_562_ la_data_out_mprj[91] VGND VGND VPWR VPWR _562_/Y sky130_fd_sc_hd__inv_2
X_493_ la_data_out_mprj[22] VGND VGND VPWR VPWR _493_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[381\] VGND VGND VPWR VPWR mprj_logic_high\[381\]/HI mprj_logic_high\[381\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[88\]_TE la_buf\[88\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[49\] _520_/Y la_buf\[49\]/TE VGND VGND VPWR VPWR la_data_in_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__412__A mprj_adr_o_core[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[105\] _576_/Y la_buf\[105\]/TE VGND VGND VPWR VPWR la_data_in_core[105] sky130_fd_sc_hd__einvp_8
XFILLER_0_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] mprj_logic_high\[368\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[38\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[40\] VGND VGND VPWR VPWR mprj_adr_buf\[30\]/TE mprj_logic_high\[40\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[80\]_B mprj_logic_high\[410\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[89\] _357_/Y mprj_logic_high\[291\]/HI VGND VGND VPWR VPWR
+ la_oen_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[227\] VGND VGND VPWR VPWR mprj_logic_high\[227\]/HI mprj_logic_high\[227\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_614_ la_oen_mprj[15] VGND VGND VPWR VPWR _614_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_545_ la_data_out_mprj[74] VGND VGND VPWR VPWR _545_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__407__A mprj_adr_o_core[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_476_ la_data_out_mprj[5] VGND VGND VPWR VPWR _476_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[71\]_B mprj_logic_high\[401\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[62\]_B mprj_logic_high\[392\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ la_oen_mprj[62] VGND VGND VPWR VPWR _330_/Y sky130_fd_sc_hd__inv_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[88\] VGND VGND VPWR VPWR la_buf\[14\]/TE mprj_logic_high\[88\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[177\] VGND VGND VPWR VPWR la_buf\[103\]/TE mprj_logic_high\[177\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[344\] VGND VGND VPWR VPWR mprj_logic_high\[344\]/HI mprj_logic_high\[344\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[53\]_B mprj_logic_high\[383\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[113\]_TE la_buf\[113\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[28\]_TE mprj_adr_buf\[28\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_528_ la_data_out_mprj[57] VGND VGND VPWR VPWR _528_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[7\]_A _446_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_459_ mprj_dat_o_core[20] VGND VGND VPWR VPWR _459_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[44\]_B mprj_logic_high\[374\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[5\] VGND VGND VPWR VPWR mprj_we_buf/TE mprj_logic_high\[5\]/LO sky130_fd_sc_hd__conb_1
XANTENNA__600__A la_oen_mprj[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_TE mprj_logic_high\[262\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[96\]_A user_to_mprj_in_gates\[96\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[35\]_B mprj_logic_high\[365\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__510__A la_data_out_mprj[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[20\]_A user_to_mprj_in_gates\[20\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[294\] VGND VGND VPWR VPWR mprj_logic_high\[294\]/HI mprj_logic_high\[294\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[123\]_A _594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[31\] _502_/Y la_buf\[31\]/TE VGND VGND VPWR VPWR la_data_in_core[31] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[87\]_A user_to_mprj_in_gates\[87\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[26\]_B mprj_logic_high\[356\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_B mprj_logic_high\[440\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[60\]_A _531_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high\[285\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__420__A mprj_adr_o_core[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[109] sky130_fd_sc_hd__inv_8
XFILLER_19_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y VGND VGND VPWR VPWR la_data_in_mprj[75]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[11\]_A user_to_mprj_in_gates\[11\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] mprj_logic_high\[350\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[20\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[125\]_A user_to_mprj_in_gates\[125\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[114\]_A _585_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[17\]_B mprj_logic_high\[347\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[78\]_A user_to_mprj_in_gates\[78\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_B mprj_logic_high\[431\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[51\]_A _522_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__330__A la_oen_mprj[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[8\] _447_/Y mprj_dat_buf\[8\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[116\]_A user_to_mprj_in_gates\[116\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[105\]_A _576_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__505__A la_data_out_mprj[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[69\]_A user_to_mprj_in_gates\[69\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[42\]_A _513_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[71\] _339_/Y mprj_logic_high\[273\]/HI VGND VGND VPWR VPWR
+ la_oen_core[71] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[307\] VGND VGND VPWR VPWR mprj_logic_high\[307\]/HI mprj_logic_high\[307\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[79\] _550_/Y la_buf\[79\]/TE VGND VGND VPWR VPWR la_data_in_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_16_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[107\]_A user_to_mprj_in_gates\[107\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__415__A mprj_adr_o_core[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[33\]_A _504_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] mprj_logic_high\[398\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[68\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_A _495_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[70\] VGND VGND VPWR VPWR mprj_dat_buf\[28\]/TE mprj_logic_high\[70\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[257\] VGND VGND VPWR VPWR mprj_logic_high\[257\]/HI mprj_logic_high\[257\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[15\]_A _486_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[424\] VGND VGND VPWR VPWR mprj_logic_high\[424\]/HI mprj_logic_high\[424\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[100\]_A _368_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y VGND VGND VPWR VPWR la_data_in_mprj[38]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[93\]_A _361_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[104\] _372_/Y mprj_logic_high\[306\]/HI VGND VGND VPWR
+ VPWR la_oen_core[104] sky130_fd_sc_hd__einvp_8
X_630_ la_oen_mprj[31] VGND VGND VPWR VPWR _630_/Y sky130_fd_sc_hd__inv_2
X_561_ la_data_out_mprj[90] VGND VGND VPWR VPWR _561_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[34\] _633_/Y mprj_logic_high\[236\]/HI VGND VGND VPWR VPWR
+ la_oen_core[34] sky130_fd_sc_hd__einvp_8
X_492_ la_data_out_mprj[21] VGND VGND VPWR VPWR _492_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[374\] VGND VGND VPWR VPWR mprj_logic_high\[374\]/HI mprj_logic_high\[374\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high\[320\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[84\]_A _352_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[32\]_TE la_buf\[32\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[75\]_A _343_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[17\]_TE mprj_logic_high\[219\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__603__A la_oen_mprj[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[66\]_A _334_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[0\]_TE la_buf\[0\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[33\] VGND VGND VPWR VPWR mprj_adr_buf\[23\]/TE mprj_logic_high\[33\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__513__A la_data_out_mprj[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[122\] VGND VGND VPWR VPWR la_buf\[48\]/TE mprj_logic_high\[122\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_613_ la_oen_mprj[14] VGND VGND VPWR VPWR _613_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[55\]_TE la_buf\[55\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[61\] _532_/Y la_buf\[61\]/TE VGND VGND VPWR VPWR la_data_in_core[61] sky130_fd_sc_hd__einvp_8
X_544_ la_data_out_mprj[73] VGND VGND VPWR VPWR _544_/Y sky130_fd_sc_hd__inv_2
X_475_ la_data_out_mprj[4] VGND VGND VPWR VPWR _475_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[57\]_A _656_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[25\] _432_/Y mprj_adr_buf\[25\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__423__A mprj_adr_o_core[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] mprj_logic_high\[380\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[50\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[48\]_A _647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__333__A la_oen_mprj[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[78\]_TE la_buf\[78\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__508__A la_data_out_mprj[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[39\]_A _638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[337\] VGND VGND VPWR VPWR mprj_logic_high\[337\]/HI mprj_logic_high\[337\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[27\]_TE mprj_dat_buf\[27\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__418__A mprj_adr_o_core[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_527_ la_data_out_mprj[56] VGND VGND VPWR VPWR _527_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[6\]_TE mprj_logic_high\[208\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_458_ mprj_dat_o_core[19] VGND VGND VPWR VPWR _458_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_389_ la_oen_mprj[121] VGND VGND VPWR VPWR _389_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y VGND VGND VPWR VPWR la_data_in_mprj[20]
+ sky130_fd_sc_hd__inv_8
XFILLER_5_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] mprj_logic_high\[428\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[98\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[26\]_A _433_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[3\]_A _602_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[17\]_A _424_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[287\] VGND VGND VPWR VPWR mprj_logic_high\[287\]/HI mprj_logic_high\[287\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[454\] VGND VGND VPWR VPWR mprj_logic_high\[454\]/HI mprj_logic_high\[454\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[24\] _495_/Y la_buf\[24\]/TE VGND VGND VPWR VPWR la_data_in_core[24] sky130_fd_sc_hd__einvp_8
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y VGND VGND VPWR VPWR la_data_in_mprj[68]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] mprj_logic_high\[343\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[13\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__611__A la_oen_mprj[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] mprj_logic_high\[454\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[124\]/Y sky130_fd_sc_hd__nand2_4
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[103\]_TE la_buf\[103\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__521__A la_data_out_mprj[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[64\] _332_/Y mprj_logic_high\[266\]/HI VGND VGND VPWR VPWR
+ la_oen_core[64] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[202\] VGND VGND VPWR VPWR mprj_logic_high\[202\]/HI mprj_logic_high\[202\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[12\] _451_/Y mprj_dat_buf\[12\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_cyc_buf_A _400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[50\]_TE mprj_logic_high\[252\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__431__A mprj_adr_o_core[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[121] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[6\]_TE mprj_dat_buf\[6\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[126\]_TE la_buf\[126\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__606__A la_oen_mprj[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[2\]_A _409_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__341__A la_oen_mprj[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[73\]_TE mprj_logic_high\[275\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__516__A la_data_out_mprj[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[63\] VGND VGND VPWR VPWR mprj_dat_buf\[21\]/TE mprj_logic_high\[63\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[152\] VGND VGND VPWR VPWR la_buf\[78\]/TE mprj_logic_high\[152\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[417\] VGND VGND VPWR VPWR mprj_logic_high\[417\]/HI mprj_logic_high\[417\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[91\] _562_/Y la_buf\[91\]/TE VGND VGND VPWR VPWR la_data_in_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_1_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__426__A mprj_adr_o_core[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] mprj_logic_high\[410\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[80\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high\[298\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__336__A la_oen_mprj[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_560_ la_data_out_mprj[89] VGND VGND VPWR VPWR _560_/Y sky130_fd_sc_hd__inv_2
X_491_ la_data_out_mprj[20] VGND VGND VPWR VPWR _491_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[9\] _608_/Y mprj_logic_high\[211\]/HI VGND VGND VPWR VPWR
+ la_oen_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_13_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[27\] _626_/Y mprj_logic_high\[229\]/HI VGND VGND VPWR VPWR
+ la_oen_core[27] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[367\] VGND VGND VPWR VPWR mprj_logic_high\[367\]/HI mprj_logic_high\[367\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[2\] _473_/Y la_buf\[2\]/TE VGND VGND VPWR VPWR la_data_in_core[2] sky130_fd_sc_hd__einvp_8
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[8\]_A _479_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y VGND VGND VPWR VPWR la_data_in_mprj[50]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[2\]_B mprj_logic_high\[332\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[26\] VGND VGND VPWR VPWR mprj_adr_buf\[16\]/TE mprj_logic_high\[26\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[115\] VGND VGND VPWR VPWR la_buf\[41\]/TE mprj_logic_high\[115\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_612_ la_oen_mprj[13] VGND VGND VPWR VPWR _612_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_543_ la_data_out_mprj[72] VGND VGND VPWR VPWR _543_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_474_ la_data_out_mprj[3] VGND VGND VPWR VPWR _474_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[54\] _525_/Y la_buf\[54\]/TE VGND VGND VPWR VPWR la_data_in_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_13_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[18\] _425_/Y mprj_adr_buf\[18\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[110\] _581_/Y la_buf\[110\]/TE VGND VGND VPWR VPWR la_data_in_core[110] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y VGND VGND VPWR VPWR la_data_in_mprj[98]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[6\]_A user_to_mprj_in_gates\[6\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] mprj_logic_high\[373\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[43\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__614__A la_oen_mprj[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] mprj_logic_high\[335\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[5\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[108\]_TE mprj_logic_high\[310\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__524__A la_data_out_mprj[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[94\] _362_/Y mprj_logic_high\[296\]/HI VGND VGND VPWR VPWR
+ la_oen_core[94] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[232\] VGND VGND VPWR VPWR mprj_logic_high\[232\]/HI mprj_logic_high\[232\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[22\]_TE la_buf\[22\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_526_ la_data_out_mprj[55] VGND VGND VPWR VPWR _526_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_457_ mprj_dat_o_core[18] VGND VGND VPWR VPWR _457_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_388_ la_oen_mprj[120] VGND VGND VPWR VPWR _388_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__434__A mprj_adr_o_core[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y VGND VGND VPWR VPWR la_data_in_mprj[13]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__609__A la_oen_mprj[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__344__A la_oen_mprj[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[45\]_TE la_buf\[45\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__519__A la_data_out_mprj[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[93\] VGND VGND VPWR VPWR la_buf\[19\]/TE mprj_logic_high\[93\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_1780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y VGND VGND VPWR VPWR la_data_in_mprj[5]
+ sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[182\] VGND VGND VPWR VPWR la_buf\[108\]/TE mprj_logic_high\[182\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[447\] VGND VGND VPWR VPWR mprj_logic_high\[447\]/HI mprj_logic_high\[447\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[17\] _488_/Y la_buf\[17\]/TE VGND VGND VPWR VPWR la_data_in_core[17] sky130_fd_sc_hd__einvp_8
XFILLER_6_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__429__A mprj_adr_o_core[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_509_ la_data_out_mprj[38] VGND VGND VPWR VPWR _509_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[68\]_TE la_buf\[68\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] mprj_logic_high\[447\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[117\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__339__A la_oen_mprj[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[127\] _395_/Y mprj_logic_high\[329\]/HI VGND VGND VPWR
+ VPWR la_oen_core[127] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[57\] _656_/Y mprj_logic_high\[259\]/HI VGND VGND VPWR VPWR
+ la_oen_core[57] sky130_fd_sc_hd__einvp_8
XFILLER_5_1820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[397\] VGND VGND VPWR VPWR mprj_logic_high\[397\]/HI mprj_logic_high\[397\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[114] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y VGND VGND VPWR VPWR la_data_in_mprj[80]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__622__A la_oen_mprj[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[56\] VGND VGND VPWR VPWR mprj_dat_buf\[14\]/TE mprj_logic_high\[56\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__532__A la_data_out_mprj[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[145\] VGND VGND VPWR VPWR la_buf\[71\]/TE mprj_logic_high\[145\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[312\] VGND VGND VPWR VPWR mprj_logic_high\[312\]/HI mprj_logic_high\[312\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xla_buf\[84\] _555_/Y la_buf\[84\]/TE VGND VGND VPWR VPWR la_data_in_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_5_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__442__A mprj_dat_o_core[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] mprj_logic_high\[403\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[73\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__617__A la_oen_mprj[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[92\]_B mprj_logic_high\[422\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__352__A la_oen_mprj[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high\[242\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_490_ la_data_out_mprj[19] VGND VGND VPWR VPWR _490_/Y sky130_fd_sc_hd__inv_2
XANTENNA__527__A la_data_out_mprj[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[262\] VGND VGND VPWR VPWR mprj_logic_high\[262\]/HI mprj_logic_high\[262\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_gates\[83\]_B mprj_logic_high\[413\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[116\]_TE la_buf\[116\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__437__A mprj_adr_o_core[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y VGND VGND VPWR VPWR la_data_in_mprj[43]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[74\]_B mprj_logic_high\[404\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[63\]_TE mprj_logic_high\[265\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__347__A la_oen_mprj[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[65\]_B mprj_logic_high\[395\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_1739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[19\] VGND VGND VPWR VPWR mprj_adr_buf\[9\]/TE mprj_logic_high\[19\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[108\] VGND VGND VPWR VPWR la_buf\[34\]/TE mprj_logic_high\[108\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[50\]_A user_to_mprj_in_gates\[50\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_611_ la_oen_mprj[12] VGND VGND VPWR VPWR _611_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_542_ la_data_out_mprj[71] VGND VGND VPWR VPWR _542_/Y sky130_fd_sc_hd__inv_2
X_473_ la_data_out_mprj[2] VGND VGND VPWR VPWR _473_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[47\] _518_/Y la_buf\[47\]/TE VGND VGND VPWR VPWR la_data_in_core[47] sky130_fd_sc_hd__einvp_8
XFILLER_9_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[56\]_B mprj_logic_high\[386\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[90\]_A _561_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high\[288\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[103\] _574_/Y la_buf\[103\]/TE VGND VGND VPWR VPWR la_data_in_core[103] sky130_fd_sc_hd__einvp_8
XFILLER_7_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[41\]_A user_to_mprj_in_gates\[41\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] mprj_logic_high\[366\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[36\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[47\]_B mprj_logic_high\[377\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[81\]_A _552_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__630__A la_oen_mprj[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[32\]_A user_to_mprj_in_gates\[32\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[99\]_A user_to_mprj_in_gates\[99\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[38\]_B mprj_logic_high\[368\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[122\]_B mprj_logic_high\[452\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[72\]_A _543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__540__A la_data_out_mprj[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[87\] _355_/Y mprj_logic_high\[289\]/HI VGND VGND VPWR VPWR
+ la_oen_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_11_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[225\] VGND VGND VPWR VPWR mprj_logic_high\[225\]/HI mprj_logic_high\[225\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[23\]_A user_to_mprj_in_gates\[23\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_525_ la_data_out_mprj[54] VGND VGND VPWR VPWR _525_/Y sky130_fd_sc_hd__inv_2
X_456_ mprj_dat_o_core[17] VGND VGND VPWR VPWR _456_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[126\]_A _597_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_387_ la_oen_mprj[119] VGND VGND VPWR VPWR _387_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[113\]_B mprj_logic_high\[443\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_B mprj_logic_high\[359\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[30\] _437_/Y mprj_adr_buf\[30\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[63\]_A _534_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__450__A mprj_dat_o_core[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[14\]_A user_to_mprj_in_gates\[14\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[117\]_A _588_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__625__A la_oen_mprj[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_B mprj_logic_high\[434\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[54\]_A _525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__360__A la_oen_mprj[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_stb_buf_A _401_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[119\]_A user_to_mprj_in_gates\[119\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[86\] VGND VGND VPWR VPWR la_buf\[12\]/TE mprj_logic_high\[86\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[108\]_A _579_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[175\] VGND VGND VPWR VPWR la_buf\[101\]/TE mprj_logic_high\[175\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__535__A la_data_out_mprj[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[45\]_A _516_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[342\] VGND VGND VPWR VPWR mprj_logic_high\[342\]/HI mprj_logic_high\[342\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_508_ la_data_out_mprj[37] VGND VGND VPWR VPWR _508_/Y sky130_fd_sc_hd__inv_2
X_439_ mprj_dat_o_core[0] VGND VGND VPWR VPWR _439_/Y sky130_fd_sc_hd__inv_2
XANTENNA__445__A mprj_dat_o_core[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[36\]_A _507_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[3\] VGND VGND VPWR VPWR mprj_cyc_buf/TE mprj_logic_high\[3\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[121\]_A _389_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[12\]_TE la_buf\[12\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__355__A la_oen_mprj[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[27\]_A _498_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[112\]_A _380_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[292\] VGND VGND VPWR VPWR mprj_logic_high\[292\]/HI mprj_logic_high\[292\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[18\]_A _489_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[103\]_A _371_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[107] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y VGND VGND VPWR VPWR la_data_in_mprj[73]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[35\]_TE la_buf\[35\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _445_/Y mprj_dat_buf\[6\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[96\]_A _364_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[3\]_TE la_buf\[3\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[49\] VGND VGND VPWR VPWR mprj_dat_buf\[7\]/TE mprj_logic_high\[49\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[138\] VGND VGND VPWR VPWR la_buf\[64\]/TE mprj_logic_high\[138\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[20\]_A _619_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[305\] VGND VGND VPWR VPWR mprj_logic_high\[305\]/HI mprj_logic_high\[305\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[58\]_TE la_buf\[58\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[77\] _548_/Y la_buf\[77\]/TE VGND VGND VPWR VPWR la_data_in_core[77] sky130_fd_sc_hd__einvp_8
XFILLER_5_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_A _355_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[11\]_A _610_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] mprj_logic_high\[396\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[66\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[78\]_A _346_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__633__A la_oen_mprj[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[69\]_A _337_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__543__A la_data_out_mprj[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[255\] VGND VGND VPWR VPWR mprj_logic_high\[255\]/HI mprj_logic_high\[255\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[422\] VGND VGND VPWR VPWR mprj_logic_high\[422\]/HI mprj_logic_high\[422\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high\[211\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y VGND VGND VPWR VPWR la_data_in_mprj[36]
+ sky130_fd_sc_hd__inv_8
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__453__A mprj_dat_o_core[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__628__A la_oen_mprj[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__363__A la_oen_mprj[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[102\] _370_/Y mprj_logic_high\[304\]/HI VGND VGND VPWR
+ VPWR la_oen_core[102] sky130_fd_sc_hd__einvp_8
X_610_ la_oen_mprj[11] VGND VGND VPWR VPWR _610_/Y sky130_fd_sc_hd__inv_2
XANTENNA__538__A la_data_out_mprj[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_541_ la_data_out_mprj[70] VGND VGND VPWR VPWR _541_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[32\] _631_/Y mprj_logic_high\[234\]/HI VGND VGND VPWR VPWR
+ la_oen_core[32] sky130_fd_sc_hd__einvp_8
X_472_ la_data_out_mprj[1] VGND VGND VPWR VPWR _472_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[20\]_A _459_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[372\] VGND VGND VPWR VPWR mprj_logic_high\[372\]/HI mprj_logic_high\[372\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__448__A mprj_dat_o_core[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[11\]_A _450_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] mprj_logic_high\[359\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[29\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high\[232\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[29\]_A _436_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__358__A la_oen_mprj[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[6\]_A _605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[106\]_TE la_buf\[106\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[31\] VGND VGND VPWR VPWR mprj_adr_buf\[21\]/TE mprj_logic_high\[31\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[28\] _467_/Y mprj_dat_buf\[28\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[28]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[120\] VGND VGND VPWR VPWR la_buf\[46\]/TE mprj_logic_high\[120\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[218\] VGND VGND VPWR VPWR mprj_logic_high\[218\]/HI mprj_logic_high\[218\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_524_ la_data_out_mprj[53] VGND VGND VPWR VPWR _524_/Y sky130_fd_sc_hd__inv_2
X_455_ mprj_dat_o_core[16] VGND VGND VPWR VPWR _455_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[53\]_TE mprj_logic_high\[255\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_386_ la_oen_mprj[118] VGND VGND VPWR VPWR _386_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[23\] _430_/Y mprj_adr_buf\[23\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[9\]_TE mprj_dat_buf\[9\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__641__A la_oen_mprj[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[91\]_TE la_buf\[91\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[76\]_TE mprj_logic_high\[278\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[79\] VGND VGND VPWR VPWR la_buf\[5\]/TE mprj_logic_high\[79\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[168\] VGND VGND VPWR VPWR la_buf\[94\]/TE mprj_logic_high\[168\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__551__A la_data_out_mprj[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[335\] VGND VGND VPWR VPWR mprj_logic_high\[335\]/HI mprj_logic_high\[335\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_507_ la_data_out_mprj[36] VGND VGND VPWR VPWR _507_/Y sky130_fd_sc_hd__inv_2
X_438_ mprj_adr_o_core[31] VGND VGND VPWR VPWR _438_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_369_ la_oen_mprj[101] VGND VGND VPWR VPWR _369_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__461__A mprj_dat_o_core[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] mprj_logic_high\[426\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[96\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high\[301\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__636__A la_oen_mprj[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[5\]_A _412_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__371__A la_oen_mprj[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__546__A la_data_out_mprj[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[285\] VGND VGND VPWR VPWR mprj_logic_high\[285\]/HI mprj_logic_high\[285\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[452\] VGND VGND VPWR VPWR mprj_logic_high\[452\]/HI mprj_logic_high\[452\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[22\] _493_/Y la_buf\[22\]/TE VGND VGND VPWR VPWR la_data_in_core[22] sky130_fd_sc_hd__einvp_8
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y VGND VGND VPWR VPWR la_data_in_mprj[66]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_stb_buf_TE mprj_stb_buf/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__456__A mprj_dat_o_core[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] mprj_logic_high\[341\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[11\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] mprj_logic_high\[452\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[122\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__366__A la_oen_mprj[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[31\]_TE mprj_adr_buf\[31\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[62\] _330_/Y mprj_logic_high\[264\]/HI VGND VGND VPWR VPWR
+ la_oen_core[62] sky130_fd_sc_hd__einvp_8
XFILLER_0_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[10\] _449_/Y mprj_dat_buf\[10\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[10]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[200\] VGND VGND VPWR VPWR la_buf\[126\]/TE mprj_logic_high\[200\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[126\] _597_/Y la_buf\[126\]/TE VGND VGND VPWR VPWR la_data_in_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_6_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] mprj_logic_high\[389\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[59\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[5\]_B mprj_logic_high\[335\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[61\] VGND VGND VPWR VPWR mprj_dat_buf\[19\]/TE mprj_logic_high\[61\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[150\] VGND VGND VPWR VPWR la_buf\[76\]/TE mprj_logic_high\[150\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[25\]_TE la_buf\[25\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[248\] VGND VGND VPWR VPWR mprj_logic_high\[248\]/HI mprj_logic_high\[248\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[415\] VGND VGND VPWR VPWR mprj_logic_high\[415\]/HI mprj_logic_high\[415\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y VGND VGND VPWR VPWR la_data_in_mprj[29]
+ sky130_fd_sc_hd__inv_8
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__644__A la_oen_mprj[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[48\]_TE la_buf\[48\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_540_ la_data_out_mprj[69] VGND VGND VPWR VPWR _540_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_471_ la_data_out_mprj[0] VGND VGND VPWR VPWR _471_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[7\] _606_/Y mprj_logic_high\[209\]/HI VGND VGND VPWR VPWR
+ la_oen_core[7] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[198\] VGND VGND VPWR VPWR la_buf\[124\]/TE mprj_logic_high\[198\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[25\] _624_/Y mprj_logic_high\[227\]/HI VGND VGND VPWR VPWR
+ la_oen_core[25] sky130_fd_sc_hd__einvp_8
XFILLER_9_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__554__A la_data_out_mprj[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[365\] VGND VGND VPWR VPWR mprj_logic_high\[365\]/HI mprj_logic_high\[365\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[0\] _471_/Y la_buf\[0\]/TE VGND VGND VPWR VPWR la_data_in_core[0] sky130_fd_sc_hd__einvp_8
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__464__A mprj_dat_o_core[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__639__A la_oen_mprj[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__374__A la_oen_mprj[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[24\] VGND VGND VPWR VPWR mprj_adr_buf\[14\]/TE mprj_logic_high\[24\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[113\] VGND VGND VPWR VPWR la_buf\[39\]/TE mprj_logic_high\[113\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__549__A la_data_out_mprj[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_523_ la_data_out_mprj[52] VGND VGND VPWR VPWR _523_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_454_ mprj_dat_o_core[15] VGND VGND VPWR VPWR _454_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[52\] _523_/Y la_buf\[52\]/TE VGND VGND VPWR VPWR la_data_in_core[52] sky130_fd_sc_hd__einvp_8
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_385_ la_oen_mprj[117] VGND VGND VPWR VPWR _385_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[16\] _423_/Y mprj_adr_buf\[16\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y VGND VGND VPWR VPWR la_data_in_mprj[96]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__459__A mprj_dat_o_core[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_rstn_buf _396_/Y mprj_rstn_buf/TE VGND VGND VPWR VPWR user_resetn sky130_fd_sc_hd__einvp_8
XFILLER_3_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] mprj_logic_high\[371\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[41\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] mprj_logic_high\[333\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[3\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__369__A la_oen_mprj[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[121\]_TE mprj_logic_high\[323\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[92\] _360_/Y mprj_logic_high\[294\]/HI VGND VGND VPWR VPWR
+ la_oen_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_2_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[328\] VGND VGND VPWR VPWR mprj_logic_high\[328\]/HI mprj_logic_high\[328\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[230\] VGND VGND VPWR VPWR mprj_logic_high\[230\]/HI mprj_logic_high\[230\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[20\]_TE mprj_logic_high\[222\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_506_ la_data_out_mprj[35] VGND VGND VPWR VPWR _506_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_437_ mprj_adr_o_core[30] VGND VGND VPWR VPWR _437_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_368_ la_oen_mprj[100] VGND VGND VPWR VPWR _368_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y VGND VGND VPWR VPWR la_data_in_mprj[11]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] mprj_logic_high\[419\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[89\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__652__A la_oen_mprj[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[43\]_TE mprj_logic_high\[245\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_cyc_buf _400_/Y mprj_cyc_buf/TE VGND VGND VPWR VPWR mprj_cyc_o_user sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[91\] VGND VGND VPWR VPWR la_buf\[17\]/TE mprj_logic_high\[91\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y VGND VGND VPWR VPWR la_data_in_mprj[3]
+ sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[278\] VGND VGND VPWR VPWR mprj_logic_high\[278\]/HI mprj_logic_high\[278\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[180\] VGND VGND VPWR VPWR la_buf\[106\]/TE mprj_logic_high\[180\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__562__A la_data_out_mprj[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[445\] VGND VGND VPWR VPWR mprj_logic_high\[445\]/HI mprj_logic_high\[445\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[119\]_TE la_buf\[119\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[15\] _486_/Y la_buf\[15\]/TE VGND VGND VPWR VPWR la_data_in_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_13_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_A _439_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[8\] _415_/Y mprj_adr_buf\[8\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y VGND VGND VPWR VPWR la_data_in_mprj[59]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__472__A la_data_out_mprj[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[81\]_TE la_buf\[81\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[66\]_TE mprj_logic_high\[268\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] mprj_logic_high\[445\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[115\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__647__A la_oen_mprj[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[95\]_B mprj_logic_high\[425\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__382__A la_oen_mprj[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_clk2_buf_TE mprj_clk2_buf/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[30\]_TE mprj_dat_buf\[30\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[125\] _393_/Y mprj_logic_high\[327\]/HI VGND VGND VPWR
+ VPWR la_oen_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_0_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[55\] _654_/Y mprj_logic_high\[257\]/HI VGND VGND VPWR VPWR
+ la_oen_core[55] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[80\]_A user_to_mprj_in_gates\[80\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__557__A la_data_out_mprj[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[395\] VGND VGND VPWR VPWR mprj_logic_high\[395\]/HI mprj_logic_high\[395\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[86\]_B mprj_logic_high\[416\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high\[291\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xla_buf\[119\] _590_/Y la_buf\[119\]/TE VGND VGND VPWR VPWR la_data_in_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_3_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[112] sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_buffers\[71\]_A user_to_mprj_in_gates\[71\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[10\]_B mprj_logic_high\[340\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__467__A mprj_dat_o_core[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[77\]_B mprj_logic_high\[407\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[62\]_A user_to_mprj_in_gates\[62\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__377__A la_oen_mprj[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[68\]_B mprj_logic_high\[398\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[54\] VGND VGND VPWR VPWR mprj_dat_buf\[12\]/TE mprj_logic_high\[54\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[143\] VGND VGND VPWR VPWR la_buf\[69\]/TE mprj_logic_high\[143\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[100\]_A user_to_mprj_in_gates\[100\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[408\] VGND VGND VPWR VPWR mprj_logic_high\[408\]/HI mprj_logic_high\[408\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[310\] VGND VGND VPWR VPWR mprj_logic_high\[310\]/HI mprj_logic_high\[310\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[53\]_A user_to_mprj_in_gates\[53\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[82\] _553_/Y la_buf\[82\]/TE VGND VGND VPWR VPWR la_data_in_core[82] sky130_fd_sc_hd__einvp_8
XFILLER_16_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[59\]_B mprj_logic_high\[389\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[93\]_A _564_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[44\]_A user_to_mprj_in_gates\[44\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] mprj_logic_high\[401\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[71\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[84\]_A _555_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__660__A la_oen_mprj[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[35\]_A user_to_mprj_in_gates\[35\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_470_ mprj_dat_o_core[31] VGND VGND VPWR VPWR _470_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[18\] _617_/Y mprj_logic_high\[220\]/HI VGND VGND VPWR VPWR
+ la_oen_core[18] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[125\]_B mprj_logic_high\[455\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[260\] VGND VGND VPWR VPWR mprj_logic_high\[260\]/HI mprj_logic_high\[260\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[75\]_A _546_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[358\] VGND VGND VPWR VPWR mprj_logic_high\[358\]/HI mprj_logic_high\[358\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__570__A la_data_out_mprj[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[26\]_A user_to_mprj_in_gates\[26\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_599_ la_oen_mprj[0] VGND VGND VPWR VPWR _599_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y VGND VGND VPWR VPWR la_data_in_mprj[41]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[116\]_B mprj_logic_high\[446\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[66\]_A _537_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__480__A la_data_out_mprj[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[17\]_A user_to_mprj_in_gates\[17\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[15\]_TE la_buf\[15\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__655__A la_oen_mprj[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[107\]_B mprj_logic_high\[437\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[57\]_A _528_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__390__A la_oen_mprj[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[17\] VGND VGND VPWR VPWR mprj_adr_buf\[7\]/TE mprj_logic_high\[17\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[106\] VGND VGND VPWR VPWR la_buf\[32\]/TE mprj_logic_high\[106\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_522_ la_data_out_mprj[51] VGND VGND VPWR VPWR _522_/Y sky130_fd_sc_hd__inv_2
XANTENNA__565__A la_data_out_mprj[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_453_ mprj_dat_o_core[14] VGND VGND VPWR VPWR _453_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[45\] _516_/Y la_buf\[45\]/TE VGND VGND VPWR VPWR la_data_in_core[45] sky130_fd_sc_hd__einvp_8
X_384_ la_oen_mprj[116] VGND VGND VPWR VPWR _384_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[48\]_A _519_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[101\] _572_/Y la_buf\[101\]/TE VGND VGND VPWR VPWR la_data_in_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y VGND VGND VPWR VPWR la_data_in_mprj[89]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[38\]_TE la_buf\[38\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__475__A la_data_out_mprj[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] mprj_logic_high\[364\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[34\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[39\]_A _510_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[124\]_A _392_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__385__A la_oen_mprj[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[6\]_TE la_buf\[6\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[115\]_A _383_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[50\]_A _649_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[85\] _353_/Y mprj_logic_high\[287\]/HI VGND VGND VPWR VPWR
+ la_oen_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_2_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[223\] VGND VGND VPWR VPWR mprj_logic_high\[223\]/HI mprj_logic_high\[223\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_505_ la_data_out_mprj[34] VGND VGND VPWR VPWR _505_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_436_ mprj_adr_o_core[29] VGND VGND VPWR VPWR _436_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_367_ la_oen_mprj[99] VGND VGND VPWR VPWR _367_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[106\]_A _374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[41\]_A _640_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[32\]_A _631_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[99\]_A _367_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[84\] VGND VGND VPWR VPWR la_buf\[10\]/TE mprj_logic_high\[84\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[173\] VGND VGND VPWR VPWR la_buf\[99\]/TE mprj_logic_high\[173\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[340\] VGND VGND VPWR VPWR mprj_logic_high\[340\]/HI mprj_logic_high\[340\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[438\] VGND VGND VPWR VPWR mprj_logic_high\[438\]/HI mprj_logic_high\[438\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[23\]_A _622_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_419_ mprj_adr_o_core[12] VGND VGND VPWR VPWR _419_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high\[313\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_A _613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[1\] VGND VGND VPWR VPWR mprj_clk_buf/TE mprj_logic_high\[1\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] mprj_logic_high\[438\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[108\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[10\]_A _417_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high\[212\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[118\] _386_/Y mprj_logic_high\[320\]/HI VGND VGND VPWR
+ VPWR la_oen_core[118] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[48\] _647_/Y mprj_logic_high\[250\]/HI VGND VGND VPWR VPWR
+ la_oen_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_1_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[388\] VGND VGND VPWR VPWR mprj_logic_high\[388\]/HI mprj_logic_high\[388\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[290\] VGND VGND VPWR VPWR mprj_logic_high\[290\]/HI mprj_logic_high\[290\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__573__A la_data_out_mprj[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[105] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y VGND VGND VPWR VPWR la_data_in_mprj[71]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__483__A la_data_out_mprj[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[33\]_TE mprj_logic_high\[235\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[4\] _443_/Y mprj_dat_buf\[4\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__658__A la_oen_mprj[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[109\]_TE la_buf\[109\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__393__A la_oen_mprj[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[47\] VGND VGND VPWR VPWR mprj_dat_buf\[5\]/TE mprj_logic_high\[47\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[136\] VGND VGND VPWR VPWR la_buf\[62\]/TE mprj_logic_high\[136\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[303\] VGND VGND VPWR VPWR mprj_logic_high\[303\]/HI mprj_logic_high\[303\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__568__A la_data_out_mprj[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[71\]_TE la_buf\[71\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[23\]_A _462_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[75\] _546_/Y la_buf\[75\]/TE VGND VGND VPWR VPWR la_data_in_core[75] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[56\]_TE mprj_logic_high\[258\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__478__A la_data_out_mprj[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] mprj_logic_high\[394\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[64\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[14\]_A _453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[94\]_TE la_buf\[94\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__388__A la_oen_mprj[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[79\]_TE mprj_logic_high\[281\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[9\]_A _608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[253\] VGND VGND VPWR VPWR mprj_logic_high\[253\]/HI mprj_logic_high\[253\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[420\] VGND VGND VPWR VPWR mprj_logic_high\[420\]/HI mprj_logic_high\[420\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_598_ la_data_out_mprj[127] VGND VGND VPWR VPWR _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y VGND VGND VPWR VPWR la_data_in_mprj[34]
+ sky130_fd_sc_hd__inv_8
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[100\] _368_/Y mprj_logic_high\[302\]/HI VGND VGND VPWR
+ VPWR la_oen_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_18_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[30\] _629_/Y mprj_logic_high\[232\]/HI VGND VGND VPWR VPWR
+ la_oen_core[30] sky130_fd_sc_hd__einvp_8
X_521_ la_data_out_mprj[50] VGND VGND VPWR VPWR _521_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_452_ mprj_dat_o_core[13] VGND VGND VPWR VPWR _452_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[1\]_A _472_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_383_ la_oen_mprj[115] VGND VGND VPWR VPWR _383_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[370\] VGND VGND VPWR VPWR mprj_logic_high\[370\]/HI mprj_logic_high\[370\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__581__A la_data_out_mprj[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[38\] _509_/Y la_buf\[38\]/TE VGND VGND VPWR VPWR la_data_in_core[38] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] mprj_logic_high\[357\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[27\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__491__A la_data_out_mprj[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[8\]_A _415_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[78\] _346_/Y mprj_logic_high\[280\]/HI VGND VGND VPWR VPWR
+ la_oen_core[78] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[26\] _465_/Y mprj_dat_buf\[26\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[26]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[216\] VGND VGND VPWR VPWR mprj_logic_high\[216\]/HI mprj_logic_high\[216\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__576__A la_data_out_mprj[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_504_ la_data_out_mprj[33] VGND VGND VPWR VPWR _504_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_435_ mprj_adr_o_core[28] VGND VGND VPWR VPWR _435_/Y sky130_fd_sc_hd__inv_2
X_366_ la_oen_mprj[98] VGND VGND VPWR VPWR _366_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[21\] _428_/Y mprj_adr_buf\[21\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__486__A la_data_out_mprj[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__396__A caravel_rstn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[77\] VGND VGND VPWR VPWR la_buf\[3\]/TE mprj_logic_high\[77\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[166\] VGND VGND VPWR VPWR la_buf\[92\]/TE mprj_logic_high\[166\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[28\]_TE la_buf\[28\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[333\] VGND VGND VPWR VPWR mprj_logic_high\[333\]/HI mprj_logic_high\[333\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_418_ mprj_adr_o_core[11] VGND VGND VPWR VPWR _418_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_349_ la_oen_mprj[81] VGND VGND VPWR VPWR _349_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_1808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] mprj_logic_high\[424\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[94\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[8\]_B mprj_logic_high\[338\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[283\] VGND VGND VPWR VPWR mprj_logic_high\[283\]/HI mprj_logic_high\[283\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[450\] VGND VGND VPWR VPWR mprj_logic_high\[450\]/HI mprj_logic_high\[450\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xla_buf\[20\] _491_/Y la_buf\[20\]/TE VGND VGND VPWR VPWR la_data_in_core[20] sky130_fd_sc_hd__einvp_8
XFILLER_10_1830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y VGND VGND VPWR VPWR la_data_in_mprj[64]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] mprj_logic_high\[450\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[120\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[129\] VGND VGND VPWR VPWR la_buf\[55\]/TE mprj_logic_high\[129\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[60\] _659_/Y mprj_logic_high\[262\]/HI VGND VGND VPWR VPWR
+ la_oen_core[60] sky130_fd_sc_hd__einvp_8
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high\[303\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[68\] _539_/Y la_buf\[68\]/TE VGND VGND VPWR VPWR la_data_in_core[68] sky130_fd_sc_hd__einvp_8
XANTENNA__584__A la_data_out_mprj[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xla_buf\[124\] _595_/Y la_buf\[124\]/TE VGND VGND VPWR VPWR la_data_in_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] mprj_logic_high\[387\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[57\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__494__A la_data_out_mprj[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high\[326\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[246\] VGND VGND VPWR VPWR mprj_logic_high\[246\]/HI mprj_logic_high\[246\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[413\] VGND VGND VPWR VPWR mprj_logic_high\[413\]/HI mprj_logic_high\[413\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__579__A la_data_out_mprj[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[23\]_TE mprj_logic_high\[225\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_597_ la_data_out_mprj[126] VGND VGND VPWR VPWR _597_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y VGND VGND VPWR VPWR la_data_in_mprj[27]
+ sky130_fd_sc_hd__inv_8
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__489__A la_data_out_mprj[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[61\]_TE la_buf\[61\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__399__A caravel_clk2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high\[248\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_520_ la_data_out_mprj[49] VGND VGND VPWR VPWR _520_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[5\] _604_/Y mprj_logic_high\[207\]/HI VGND VGND VPWR VPWR
+ la_oen_core[5] sky130_fd_sc_hd__einvp_8
X_451_ mprj_dat_o_core[12] VGND VGND VPWR VPWR _451_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[196\] VGND VGND VPWR VPWR la_buf\[122\]/TE mprj_logic_high\[196\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[23\] _622_/Y mprj_logic_high\[225\]/HI VGND VGND VPWR VPWR
+ la_oen_core[23] sky130_fd_sc_hd__einvp_8
XFILLER_0_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_382_ la_oen_mprj[114] VGND VGND VPWR VPWR _382_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[363\] VGND VGND VPWR VPWR mprj_logic_high\[363\]/HI mprj_logic_high\[363\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[10\]_TE mprj_dat_buf\[10\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_649_ la_oen_mprj[50] VGND VGND VPWR VPWR _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[84\]_TE la_buf\[84\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[69\]_TE mprj_logic_high\[271\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[2\]_A _405_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[22\] VGND VGND VPWR VPWR mprj_adr_buf\[12\]/TE mprj_logic_high\[22\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[209\] VGND VGND VPWR VPWR mprj_logic_high\[209\]/HI mprj_logic_high\[209\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[111\] VGND VGND VPWR VPWR la_buf\[37\]/TE mprj_logic_high\[111\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[19\] _458_/Y mprj_dat_buf\[19\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[19]
+ sky130_fd_sc_hd__einvp_8
X_503_ la_data_out_mprj[32] VGND VGND VPWR VPWR _503_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_434_ mprj_adr_o_core[27] VGND VGND VPWR VPWR _434_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[50\] _521_/Y la_buf\[50\]/TE VGND VGND VPWR VPWR la_data_in_core[50] sky130_fd_sc_hd__einvp_8
XANTENNA__592__A la_data_out_mprj[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_365_ la_oen_mprj[97] VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[3\]_A _442_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[14\] _421_/Y mprj_adr_buf\[14\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[40\]_B mprj_logic_high\[370\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y VGND VGND VPWR VPWR la_data_in_mprj[94]
+ sky130_fd_sc_hd__inv_8
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[92\]_A user_to_mprj_in_gates\[92\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] mprj_logic_high\[331\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[1\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[31\]_B mprj_logic_high\[361\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[98\]_B mprj_logic_high\[428\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[159\] VGND VGND VPWR VPWR la_buf\[85\]/TE mprj_logic_high\[159\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[90\] _358_/Y mprj_logic_high\[292\]/HI VGND VGND VPWR VPWR
+ la_oen_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[326\] VGND VGND VPWR VPWR mprj_logic_high\[326\]/HI mprj_logic_high\[326\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[83\]_A user_to_mprj_in_gates\[83\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[22\]_B mprj_logic_high\[352\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xla_buf\[98\] _569_/Y la_buf\[98\]/TE VGND VGND VPWR VPWR la_data_in_core[98] sky130_fd_sc_hd__einvp_8
XANTENNA__587__A la_data_out_mprj[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[89\]_B mprj_logic_high\[419\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_417_ mprj_adr_o_core[10] VGND VGND VPWR VPWR _417_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_348_ la_oen_mprj[80] VGND VGND VPWR VPWR _348_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[121\]_A user_to_mprj_in_gates\[121\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[110\]_A _581_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[74\]_A user_to_mprj_in_gates\[74\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[13\]_B mprj_logic_high\[343\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] mprj_logic_high\[417\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[87\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__497__A la_data_out_mprj[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[112\]_A user_to_mprj_in_gates\[112\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[101\]_A _572_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[65\]_A user_to_mprj_in_gates\[65\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y VGND VGND VPWR VPWR la_data_in_mprj[1]
+ sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[276\] VGND VGND VPWR VPWR mprj_logic_high\[276\]/HI mprj_logic_high\[276\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[443\] VGND VGND VPWR VPWR mprj_logic_high\[443\]/HI mprj_logic_high\[443\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_in_buffers\[103\]_A user_to_mprj_in_gates\[103\]/Y VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[9\] _480_/Y la_buf\[9\]/TE VGND VGND VPWR VPWR la_data_in_core[9] sky130_fd_sc_hd__einvp_8
Xla_buf\[13\] _484_/Y la_buf\[13\]/TE VGND VGND VPWR VPWR la_data_in_core[13] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[56\]_A user_to_mprj_in_gates\[56\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[6\] _413_/Y mprj_adr_buf\[6\]/TE VGND VGND VPWR VPWR mprj_adr_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y VGND VGND VPWR VPWR la_data_in_mprj[57]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[96\]_A _567_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[47\]_A user_to_mprj_in_gates\[47\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[20\]_A _491_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] mprj_logic_high\[443\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[113\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[18\]_TE la_buf\[18\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[87\]_A _558_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[38\]_A user_to_mprj_in_gates\[38\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[11\]_A _482_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[123\] _391_/Y mprj_logic_high\[325\]/HI VGND VGND VPWR
+ VPWR la_oen_core[123] sky130_fd_sc_hd__einvp_8
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[53\] _652_/Y mprj_logic_high\[255\]/HI VGND VGND VPWR VPWR
+ la_oen_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_5_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[393\] VGND VGND VPWR VPWR mprj_logic_high\[393\]/HI mprj_logic_high\[393\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_la_buf\[78\]_A _549_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[29\]_A user_to_mprj_in_gates\[29\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xla_buf\[117\] _588_/Y la_buf\[117\]/TE VGND VGND VPWR VPWR la_data_in_core[117] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[110] sky130_fd_sc_hd__inv_8
XFILLER_6_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[119\]_B mprj_logic_high\[449\]/HI VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[69\]_A _540_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_TE la_buf\[9\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[52\] VGND VGND VPWR VPWR mprj_dat_buf\[10\]/TE mprj_logic_high\[52\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[80\]_A _348_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[141\] VGND VGND VPWR VPWR la_buf\[67\]/TE mprj_logic_high\[141\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[239\] VGND VGND VPWR VPWR mprj_logic_high\[239\]/HI mprj_logic_high\[239\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[406\] VGND VGND VPWR VPWR mprj_logic_high\[406\]/HI mprj_logic_high\[406\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[80\] _551_/Y la_buf\[80\]/TE VGND VGND VPWR VPWR la_data_in_core[80] sky130_fd_sc_hd__einvp_8
XANTENNA__595__A la_data_out_mprj[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_596_ la_data_out_mprj[125] VGND VGND VPWR VPWR _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[71\]_A _339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[62\]_A _330_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[127\]_A _395_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_450_ mprj_dat_o_core[11] VGND VGND VPWR VPWR _450_/Y sky130_fd_sc_hd__inv_2
X_381_ la_oen_mprj[113] VGND VGND VPWR VPWR _381_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[189\] VGND VGND VPWR VPWR la_buf\[115\]/TE mprj_logic_high\[189\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[16\] _615_/Y mprj_logic_high\[218\]/HI VGND VGND VPWR VPWR
+ la_oen_core[16] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[356\] VGND VGND VPWR VPWR mprj_logic_high\[356\]/HI mprj_logic_high\[356\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_user_to_mprj_oen_buffers\[118\]_A _386_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[53\]_A _652_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_648_ la_oen_mprj[49] VGND VGND VPWR VPWR _648_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_579_ la_data_out_mprj[108] VGND VGND VPWR VPWR _579_/Y sky130_fd_sc_hd__inv_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[114\]_TE mprj_logic_high\[316\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[109\]_A _377_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[44\]_A _643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high\[215\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[35\]_A _634_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[15\] VGND VGND VPWR VPWR mprj_adr_buf\[5\]/TE mprj_logic_high\[15\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[104\] VGND VGND VPWR VPWR la_buf\[30\]/TE mprj_logic_high\[104\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_mprj_adr_buf\[31\]_A _438_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_502_ la_data_out_mprj[31] VGND VGND VPWR VPWR _502_/Y sky130_fd_sc_hd__inv_2
X_433_ mprj_adr_o_core[26] VGND VGND VPWR VPWR _433_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xla_buf\[43\] _514_/Y la_buf\[43\]/TE VGND VGND VPWR VPWR la_data_in_core[43] sky130_fd_sc_hd__einvp_8
X_364_ la_oen_mprj[96] VGND VGND VPWR VPWR _364_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[26\]_A _625_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[22\]_A _429_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y VGND VGND VPWR VPWR la_data_in_mprj[87]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[51\]_TE la_buf\[51\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] mprj_logic_high\[362\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[32\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high\[238\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[17\]_A _616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[13\]_A _420_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[83\] _351_/Y mprj_logic_high\[285\]/HI VGND VGND VPWR VPWR
+ la_oen_core[83] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[31\] _470_/Y mprj_dat_buf\[31\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[319\] VGND VGND VPWR VPWR mprj_logic_high\[319\]/HI mprj_logic_high\[319\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[221\] VGND VGND VPWR VPWR mprj_logic_high\[221\]/HI mprj_logic_high\[221\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[74\]_TE la_buf\[74\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[59\]_TE mprj_logic_high\[261\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_416_ mprj_adr_o_core[9] VGND VGND VPWR VPWR _416_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_347_ la_oen_mprj[79] VGND VGND VPWR VPWR _347_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high\[204\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[97\]_TE la_buf\[97\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[82\] VGND VGND VPWR VPWR la_buf\[8\]/TE mprj_logic_high\[82\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[171\] VGND VGND VPWR VPWR la_buf\[97\]/TE mprj_logic_high\[171\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[269\] VGND VGND VPWR VPWR mprj_logic_high\[269\]/HI mprj_logic_high\[269\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[436\] VGND VGND VPWR VPWR mprj_logic_high\[436\]/HI mprj_logic_high\[436\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__598__A la_data_out_mprj[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[26\]_A _465_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[17\]_A _456_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] mprj_logic_high\[436\]/HI VGND
+ VGND VPWR VPWR user_to_mprj_in_gates\[106\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[116\] _384_/Y mprj_logic_high\[318\]/HI VGND VGND VPWR
+ VPWR la_oen_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_5_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[46\] _645_/Y mprj_logic_high\[248\]/HI VGND VGND VPWR VPWR
+ la_oen_core[46] sky130_fd_sc_hd__einvp_8
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[386\] VGND VGND VPWR VPWR mprj_logic_high\[386\]/HI mprj_logic_high\[386\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_TE mprj_adr_buf\[14\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y VGND VGND VPWR VPWR
+ la_data_in_mprj[103] sky130_fd_sc_hd__inv_8
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[2\] _441_/Y mprj_dat_buf\[2\]/TE VGND VGND VPWR VPWR mprj_dat_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[2\]_TE mprj_dat_buf\[2\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[122\]_TE la_buf\[122\]/TE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmprj_logic_high\[45\] VGND VGND VPWR VPWR mprj_dat_buf\[3\]/TE mprj_logic_high\[45\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[134\] VGND VGND VPWR VPWR la_buf\[60\]/TE mprj_logic_high\[134\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[301\] VGND VGND VPWR VPWR mprj_logic_high\[301\]/HI mprj_logic_high\[301\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[4\]_A _475_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xla_buf\[73\] _544_/Y la_buf\[73\]/TE VGND VGND VPWR VPWR la_data_in_core[73] sky130_fd_sc_hd__einvp_8
X_595_ la_data_out_mprj[124] VGND VGND VPWR VPWR _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] mprj_logic_high\[392\]/HI VGND VGND
+ VPWR VPWR user_to_mprj_in_gates\[62\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_380_ la_oen_mprj[112] VGND VGND VPWR VPWR _380_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high\[294\]/HI VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[251\] VGND VGND VPWR VPWR mprj_logic_high\[251\]/HI mprj_logic_high\[251\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[349\] VGND VGND VPWR VPWR mprj_logic_high\[349\]/HI mprj_logic_high\[349\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_647_ la_oen_mprj[48] VGND VGND VPWR VPWR _647_/Y sky130_fd_sc_hd__inv_2
X_578_ la_data_out_mprj[107] VGND VGND VPWR VPWR _578_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[2\]_A user_to_mprj_in_gates\[2\]/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y VGND VGND VPWR VPWR la_data_in_mprj[32]
+ sky130_fd_sc_hd__inv_8
XFILLER_13_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

