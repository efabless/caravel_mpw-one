* NGSPICE file created from caravel.ext - technology: sky130A

* Black-box entry subcircuit for gpio_control_block abstract view
.subckt gpio_control_block mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en
+ pad_gpio_ana_pol pad_gpio_ana_sel pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover
+ pad_gpio_ib_mode_sel pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel
+ pad_gpio_vtrip_sel resetn serial_clock serial_data_in serial_data_out user_gpio_in
+ user_gpio_oeb user_gpio_out zero vccd vssd vccd1 vssd1
.ends

* Black-box entry subcircuit for chip_io abstract view
.subckt chip_io clock clock_core por flash_clk flash_clk_core flash_clk_ieb_core flash_clk_oeb_core
+ flash_csb flash_csb_core flash_csb_ieb_core flash_csb_oeb_core flash_io0 flash_io0_di_core
+ flash_io0_do_core flash_io0_ieb_core flash_io0_oeb_core flash_io1 flash_io1_di_core
+ flash_io1_do_core flash_io1_ieb_core flash_io1_oeb_core gpio gpio_in_core gpio_inenb_core
+ gpio_mode0_core gpio_mode1_core gpio_out_core gpio_outenb_core mprj_io[0] mprj_io_analog_en[0]
+ mprj_io_analog_pol[0] mprj_io_analog_sel[0] mprj_io_dm[0] mprj_io_dm[1] mprj_io_dm[2]
+ mprj_io_enh[0] mprj_io_hldh_n[0] mprj_io_holdover[0] mprj_io_ib_mode_sel[0] mprj_io_inp_dis[0]
+ mprj_io_oeb[0] mprj_io_out[0] mprj_io_slow_sel[0] mprj_io_vtrip_sel[0] mprj_io_in[0]
+ mprj_analog_io[3] mprj_io[10] mprj_io_analog_en[10] mprj_io_analog_pol[10] mprj_io_analog_sel[10]
+ mprj_io_dm[30] mprj_io_dm[31] mprj_io_dm[32] mprj_io_enh[10] mprj_io_hldh_n[10]
+ mprj_io_holdover[10] mprj_io_ib_mode_sel[10] mprj_io_inp_dis[10] mprj_io_oeb[10]
+ mprj_io_out[10] mprj_io_slow_sel[10] mprj_io_vtrip_sel[10] mprj_io_in[10] mprj_analog_io[4]
+ mprj_io[11] mprj_io_analog_en[11] mprj_io_analog_pol[11] mprj_io_analog_sel[11]
+ mprj_io_dm[33] mprj_io_dm[34] mprj_io_dm[35] mprj_io_enh[11] mprj_io_hldh_n[11]
+ mprj_io_holdover[11] mprj_io_ib_mode_sel[11] mprj_io_inp_dis[11] mprj_io_oeb[11]
+ mprj_io_out[11] mprj_io_slow_sel[11] mprj_io_vtrip_sel[11] mprj_io_in[11] mprj_analog_io[5]
+ mprj_io[12] mprj_io_analog_en[12] mprj_io_analog_pol[12] mprj_io_analog_sel[12]
+ mprj_io_dm[36] mprj_io_dm[37] mprj_io_dm[38] mprj_io_enh[12] mprj_io_hldh_n[12]
+ mprj_io_holdover[12] mprj_io_ib_mode_sel[12] mprj_io_inp_dis[12] mprj_io_oeb[12]
+ mprj_io_out[12] mprj_io_slow_sel[12] mprj_io_vtrip_sel[12] mprj_io_in[12] mprj_analog_io[6]
+ mprj_io[13] mprj_io_analog_en[13] mprj_io_analog_pol[13] mprj_io_analog_sel[13]
+ mprj_io_dm[39] mprj_io_dm[40] mprj_io_dm[41] mprj_io_enh[13] mprj_io_hldh_n[13]
+ mprj_io_holdover[13] mprj_io_ib_mode_sel[13] mprj_io_inp_dis[13] mprj_io_oeb[13]
+ mprj_io_out[13] mprj_io_slow_sel[13] mprj_io_vtrip_sel[13] mprj_io_in[13] mprj_analog_io[7]
+ mprj_io[14] mprj_io_analog_en[14] mprj_io_analog_pol[14] mprj_io_analog_sel[14]
+ mprj_io_dm[42] mprj_io_dm[43] mprj_io_dm[44] mprj_io_enh[14] mprj_io_hldh_n[14]
+ mprj_io_holdover[14] mprj_io_ib_mode_sel[14] mprj_io_inp_dis[14] mprj_io_oeb[14]
+ mprj_io_out[14] mprj_io_slow_sel[14] mprj_io_vtrip_sel[14] mprj_io_in[14] mprj_analog_io[8]
+ mprj_io[15] mprj_io_analog_en[15] mprj_io_analog_pol[15] mprj_io_analog_sel[15]
+ mprj_io_dm[45] mprj_io_dm[46] mprj_io_dm[47] mprj_io_enh[15] mprj_io_hldh_n[15]
+ mprj_io_holdover[15] mprj_io_ib_mode_sel[15] mprj_io_inp_dis[15] mprj_io_oeb[15]
+ mprj_io_out[15] mprj_io_slow_sel[15] mprj_io_vtrip_sel[15] mprj_io_in[15] mprj_analog_io[9]
+ mprj_io[16] mprj_io_analog_en[16] mprj_io_analog_pol[16] mprj_io_analog_sel[16]
+ mprj_io_dm[48] mprj_io_dm[49] mprj_io_dm[50] mprj_io_enh[16] mprj_io_hldh_n[16]
+ mprj_io_holdover[16] mprj_io_ib_mode_sel[16] mprj_io_inp_dis[16] mprj_io_oeb[16]
+ mprj_io_out[16] mprj_io_slow_sel[16] mprj_io_vtrip_sel[16] mprj_io_in[16] mprj_analog_io[10]
+ mprj_io[17] mprj_io_analog_en[17] mprj_io_analog_pol[17] mprj_io_analog_sel[17]
+ mprj_io_dm[51] mprj_io_dm[52] mprj_io_dm[53] mprj_io_enh[17] mprj_io_hldh_n[17]
+ mprj_io_holdover[17] mprj_io_ib_mode_sel[17] mprj_io_inp_dis[17] mprj_io_oeb[17]
+ mprj_io_out[17] mprj_io_slow_sel[17] mprj_io_vtrip_sel[17] mprj_io_in[17] mprj_io[1]
+ mprj_io_analog_en[1] mprj_io_analog_pol[1] mprj_io_analog_sel[1] mprj_io_dm[3] mprj_io_dm[4]
+ mprj_io_dm[5] mprj_io_enh[1] mprj_io_hldh_n[1] mprj_io_holdover[1] mprj_io_ib_mode_sel[1]
+ mprj_io_inp_dis[1] mprj_io_oeb[1] mprj_io_out[1] mprj_io_slow_sel[1] mprj_io_vtrip_sel[1]
+ mprj_io_in[1] mprj_io[2] mprj_io_analog_en[2] mprj_io_analog_pol[2] mprj_io_analog_sel[2]
+ mprj_io_dm[6] mprj_io_dm[7] mprj_io_dm[8] mprj_io_enh[2] mprj_io_hldh_n[2] mprj_io_holdover[2]
+ mprj_io_ib_mode_sel[2] mprj_io_inp_dis[2] mprj_io_oeb[2] mprj_io_out[2] mprj_io_slow_sel[2]
+ mprj_io_vtrip_sel[2] mprj_io_in[2] mprj_io[3] mprj_io_analog_en[3] mprj_io_analog_pol[3]
+ mprj_io_analog_sel[3] mprj_io_dm[10] mprj_io_dm[11] mprj_io_dm[9] mprj_io_enh[3]
+ mprj_io_hldh_n[3] mprj_io_holdover[3] mprj_io_ib_mode_sel[3] mprj_io_inp_dis[3]
+ mprj_io_oeb[3] mprj_io_out[3] mprj_io_slow_sel[3] mprj_io_vtrip_sel[3] mprj_io_in[3]
+ mprj_io[4] mprj_io_analog_en[4] mprj_io_analog_pol[4] mprj_io_analog_sel[4] mprj_io_dm[12]
+ mprj_io_dm[13] mprj_io_dm[14] mprj_io_enh[4] mprj_io_hldh_n[4] mprj_io_holdover[4]
+ mprj_io_ib_mode_sel[4] mprj_io_inp_dis[4] mprj_io_oeb[4] mprj_io_out[4] mprj_io_slow_sel[4]
+ mprj_io_vtrip_sel[4] mprj_io_in[4] mprj_io[5] mprj_io_analog_en[5] mprj_io_analog_pol[5]
+ mprj_io_analog_sel[5] mprj_io_dm[15] mprj_io_dm[16] mprj_io_dm[17] mprj_io_enh[5]
+ mprj_io_hldh_n[5] mprj_io_holdover[5] mprj_io_ib_mode_sel[5] mprj_io_inp_dis[5]
+ mprj_io_oeb[5] mprj_io_out[5] mprj_io_slow_sel[5] mprj_io_vtrip_sel[5] mprj_io_in[5]
+ mprj_io[6] mprj_io_analog_en[6] mprj_io_analog_pol[6] mprj_io_analog_sel[6] mprj_io_dm[18]
+ mprj_io_dm[19] mprj_io_dm[20] mprj_io_enh[6] mprj_io_hldh_n[6] mprj_io_holdover[6]
+ mprj_io_ib_mode_sel[6] mprj_io_inp_dis[6] mprj_io_oeb[6] mprj_io_out[6] mprj_io_slow_sel[6]
+ mprj_io_vtrip_sel[6] mprj_io_in[6] mprj_analog_io[0] mprj_io[7] mprj_io_analog_en[7]
+ mprj_io_analog_pol[7] mprj_io_analog_sel[7] mprj_io_dm[21] mprj_io_dm[22] mprj_io_dm[23]
+ mprj_io_enh[7] mprj_io_hldh_n[7] mprj_io_holdover[7] mprj_io_ib_mode_sel[7] mprj_io_inp_dis[7]
+ mprj_io_oeb[7] mprj_io_out[7] mprj_io_slow_sel[7] mprj_io_vtrip_sel[7] mprj_io_in[7]
+ mprj_analog_io[1] mprj_io[8] mprj_io_analog_en[8] mprj_io_analog_pol[8] mprj_io_analog_sel[8]
+ mprj_io_dm[24] mprj_io_dm[25] mprj_io_dm[26] mprj_io_enh[8] mprj_io_hldh_n[8] mprj_io_holdover[8]
+ mprj_io_ib_mode_sel[8] mprj_io_inp_dis[8] mprj_io_oeb[8] mprj_io_out[8] mprj_io_slow_sel[8]
+ mprj_io_vtrip_sel[8] mprj_io_in[8] mprj_analog_io[2] mprj_io[9] mprj_io_analog_en[9]
+ mprj_io_analog_pol[9] mprj_io_analog_sel[9] mprj_io_dm[27] mprj_io_dm[28] mprj_io_dm[29]
+ mprj_io_enh[9] mprj_io_hldh_n[9] mprj_io_holdover[9] mprj_io_ib_mode_sel[9] mprj_io_inp_dis[9]
+ mprj_io_oeb[9] mprj_io_out[9] mprj_io_slow_sel[9] mprj_io_vtrip_sel[9] mprj_io_in[9]
+ mprj_analog_io[11] mprj_io[18] mprj_io_analog_en[18] mprj_io_analog_pol[18] mprj_io_analog_sel[18]
+ mprj_io_dm[54] mprj_io_dm[55] mprj_io_dm[56] mprj_io_enh[18] mprj_io_hldh_n[18]
+ mprj_io_holdover[18] mprj_io_ib_mode_sel[18] mprj_io_inp_dis[18] mprj_io_oeb[18]
+ mprj_io_out[18] mprj_io_slow_sel[18] mprj_io_vtrip_sel[18] mprj_io_in[18] mprj_analog_io[21]
+ mprj_io[28] mprj_io_analog_en[28] mprj_io_analog_pol[28] mprj_io_analog_sel[28]
+ mprj_io_dm[84] mprj_io_dm[85] mprj_io_dm[86] mprj_io_enh[28] mprj_io_hldh_n[28]
+ mprj_io_holdover[28] mprj_io_ib_mode_sel[28] mprj_io_inp_dis[28] mprj_io_oeb[28]
+ mprj_io_out[28] mprj_io_slow_sel[28] mprj_io_vtrip_sel[28] mprj_io_in[28] mprj_analog_io[22]
+ mprj_io[29] mprj_io_analog_en[29] mprj_io_analog_pol[29] mprj_io_analog_sel[29]
+ mprj_io_dm[87] mprj_io_dm[88] mprj_io_dm[89] mprj_io_enh[29] mprj_io_hldh_n[29]
+ mprj_io_holdover[29] mprj_io_ib_mode_sel[29] mprj_io_inp_dis[29] mprj_io_oeb[29]
+ mprj_io_out[29] mprj_io_slow_sel[29] mprj_io_vtrip_sel[29] mprj_io_in[29] mprj_analog_io[23]
+ mprj_io[30] mprj_io_analog_en[30] mprj_io_analog_pol[30] mprj_io_analog_sel[30]
+ mprj_io_dm[90] mprj_io_dm[91] mprj_io_dm[92] mprj_io_enh[30] mprj_io_hldh_n[30]
+ mprj_io_holdover[30] mprj_io_ib_mode_sel[30] mprj_io_inp_dis[30] mprj_io_oeb[30]
+ mprj_io_out[30] mprj_io_slow_sel[30] mprj_io_vtrip_sel[30] mprj_io_in[30] mprj_analog_io[24]
+ mprj_io[31] mprj_io_analog_en[31] mprj_io_analog_pol[31] mprj_io_analog_sel[31]
+ mprj_io_dm[93] mprj_io_dm[94] mprj_io_dm[95] mprj_io_enh[31] mprj_io_hldh_n[31]
+ mprj_io_holdover[31] mprj_io_ib_mode_sel[31] mprj_io_inp_dis[31] mprj_io_oeb[31]
+ mprj_io_out[31] mprj_io_slow_sel[31] mprj_io_vtrip_sel[31] mprj_io_in[31] mprj_analog_io[25]
+ mprj_io[32] mprj_io_analog_en[32] mprj_io_analog_pol[32] mprj_io_analog_sel[32]
+ mprj_io_dm[96] mprj_io_dm[97] mprj_io_dm[98] mprj_io_enh[32] mprj_io_hldh_n[32]
+ mprj_io_holdover[32] mprj_io_ib_mode_sel[32] mprj_io_inp_dis[32] mprj_io_oeb[32]
+ mprj_io_out[32] mprj_io_slow_sel[32] mprj_io_vtrip_sel[32] mprj_io_in[32] mprj_analog_io[26]
+ mprj_io[33] mprj_io_analog_en[33] mprj_io_analog_pol[33] mprj_io_analog_sel[33]
+ mprj_io_dm[100] mprj_io_dm[101] mprj_io_dm[99] mprj_io_enh[33] mprj_io_hldh_n[33]
+ mprj_io_holdover[33] mprj_io_ib_mode_sel[33] mprj_io_inp_dis[33] mprj_io_oeb[33]
+ mprj_io_out[33] mprj_io_slow_sel[33] mprj_io_vtrip_sel[33] mprj_io_in[33] mprj_analog_io[27]
+ mprj_io[34] mprj_io_analog_en[34] mprj_io_analog_pol[34] mprj_io_analog_sel[34]
+ mprj_io_dm[102] mprj_io_dm[103] mprj_io_dm[104] mprj_io_enh[34] mprj_io_hldh_n[34]
+ mprj_io_holdover[34] mprj_io_ib_mode_sel[34] mprj_io_inp_dis[34] mprj_io_oeb[34]
+ mprj_io_out[34] mprj_io_slow_sel[34] mprj_io_vtrip_sel[34] mprj_io_in[34] mprj_analog_io[28]
+ mprj_io[35] mprj_io_analog_en[35] mprj_io_analog_pol[35] mprj_io_analog_sel[35]
+ mprj_io_dm[105] mprj_io_dm[106] mprj_io_dm[107] mprj_io_enh[35] mprj_io_hldh_n[35]
+ mprj_io_holdover[35] mprj_io_ib_mode_sel[35] mprj_io_inp_dis[35] mprj_io_oeb[35]
+ mprj_io_out[35] mprj_io_slow_sel[35] mprj_io_vtrip_sel[35] mprj_io_in[35] mprj_analog_io[29]
+ mprj_io[36] mprj_io_analog_en[36] mprj_io_analog_pol[36] mprj_io_analog_sel[36]
+ mprj_io_dm[108] mprj_io_dm[109] mprj_io_dm[110] mprj_io_enh[36] mprj_io_hldh_n[36]
+ mprj_io_holdover[36] mprj_io_ib_mode_sel[36] mprj_io_inp_dis[36] mprj_io_oeb[36]
+ mprj_io_out[36] mprj_io_slow_sel[36] mprj_io_vtrip_sel[36] mprj_io_in[36] mprj_analog_io[30]
+ mprj_io[37] mprj_io_analog_en[37] mprj_io_analog_pol[37] mprj_io_analog_sel[37]
+ mprj_io_dm[111] mprj_io_dm[112] mprj_io_dm[113] mprj_io_enh[37] mprj_io_hldh_n[37]
+ mprj_io_holdover[37] mprj_io_ib_mode_sel[37] mprj_io_inp_dis[37] mprj_io_oeb[37]
+ mprj_io_out[37] mprj_io_slow_sel[37] mprj_io_vtrip_sel[37] mprj_io_in[37] mprj_analog_io[12]
+ mprj_io[19] mprj_io_analog_en[19] mprj_io_analog_pol[19] mprj_io_analog_sel[19]
+ mprj_io_dm[57] mprj_io_dm[58] mprj_io_dm[59] mprj_io_enh[19] mprj_io_hldh_n[19]
+ mprj_io_holdover[19] mprj_io_ib_mode_sel[19] mprj_io_inp_dis[19] mprj_io_oeb[19]
+ mprj_io_out[19] mprj_io_slow_sel[19] mprj_io_vtrip_sel[19] mprj_io_in[19] mprj_analog_io[13]
+ mprj_io[20] mprj_io_analog_en[20] mprj_io_analog_pol[20] mprj_io_analog_sel[20]
+ mprj_io_dm[60] mprj_io_dm[61] mprj_io_dm[62] mprj_io_enh[20] mprj_io_hldh_n[20]
+ mprj_io_holdover[20] mprj_io_ib_mode_sel[20] mprj_io_inp_dis[20] mprj_io_oeb[20]
+ mprj_io_out[20] mprj_io_slow_sel[20] mprj_io_vtrip_sel[20] mprj_io_in[20] mprj_analog_io[14]
+ mprj_io[21] mprj_io_analog_en[21] mprj_io_analog_pol[21] mprj_io_analog_sel[21]
+ mprj_io_dm[63] mprj_io_dm[64] mprj_io_dm[65] mprj_io_enh[21] mprj_io_hldh_n[21]
+ mprj_io_holdover[21] mprj_io_ib_mode_sel[21] mprj_io_inp_dis[21] mprj_io_oeb[21]
+ mprj_io_out[21] mprj_io_slow_sel[21] mprj_io_vtrip_sel[21] mprj_io_in[21] mprj_analog_io[15]
+ mprj_io[22] mprj_io_analog_en[22] mprj_io_analog_pol[22] mprj_io_analog_sel[22]
+ mprj_io_dm[66] mprj_io_dm[67] mprj_io_dm[68] mprj_io_enh[22] mprj_io_hldh_n[22]
+ mprj_io_holdover[22] mprj_io_ib_mode_sel[22] mprj_io_inp_dis[22] mprj_io_oeb[22]
+ mprj_io_out[22] mprj_io_slow_sel[22] mprj_io_vtrip_sel[22] mprj_io_in[22] mprj_analog_io[16]
+ mprj_io[23] mprj_io_analog_en[23] mprj_io_analog_pol[23] mprj_io_analog_sel[23]
+ mprj_io_dm[69] mprj_io_dm[70] mprj_io_dm[71] mprj_io_enh[23] mprj_io_hldh_n[23]
+ mprj_io_holdover[23] mprj_io_ib_mode_sel[23] mprj_io_inp_dis[23] mprj_io_oeb[23]
+ mprj_io_out[23] mprj_io_slow_sel[23] mprj_io_vtrip_sel[23] mprj_io_in[23] mprj_analog_io[17]
+ mprj_io[24] mprj_io_analog_en[24] mprj_io_analog_pol[24] mprj_io_analog_sel[24]
+ mprj_io_dm[72] mprj_io_dm[73] mprj_io_dm[74] mprj_io_enh[24] mprj_io_hldh_n[24]
+ mprj_io_holdover[24] mprj_io_ib_mode_sel[24] mprj_io_inp_dis[24] mprj_io_oeb[24]
+ mprj_io_out[24] mprj_io_slow_sel[24] mprj_io_vtrip_sel[24] mprj_io_in[24] mprj_analog_io[18]
+ mprj_io[25] mprj_io_analog_en[25] mprj_io_analog_pol[25] mprj_io_analog_sel[25]
+ mprj_io_dm[75] mprj_io_dm[76] mprj_io_dm[77] mprj_io_enh[25] mprj_io_hldh_n[25]
+ mprj_io_holdover[25] mprj_io_ib_mode_sel[25] mprj_io_inp_dis[25] mprj_io_oeb[25]
+ mprj_io_out[25] mprj_io_slow_sel[25] mprj_io_vtrip_sel[25] mprj_io_in[25] mprj_analog_io[19]
+ mprj_io[26] mprj_io_analog_en[26] mprj_io_analog_pol[26] mprj_io_analog_sel[26]
+ mprj_io_dm[78] mprj_io_dm[79] mprj_io_dm[80] mprj_io_enh[26] mprj_io_hldh_n[26]
+ mprj_io_holdover[26] mprj_io_ib_mode_sel[26] mprj_io_inp_dis[26] mprj_io_oeb[26]
+ mprj_io_out[26] mprj_io_slow_sel[26] mprj_io_vtrip_sel[26] mprj_io_in[26] mprj_analog_io[20]
+ mprj_io[27] mprj_io_analog_en[27] mprj_io_analog_pol[27] mprj_io_analog_sel[27]
+ mprj_io_dm[81] mprj_io_dm[82] mprj_io_dm[83] mprj_io_enh[27] mprj_io_hldh_n[27]
+ mprj_io_holdover[27] mprj_io_ib_mode_sel[27] mprj_io_inp_dis[27] mprj_io_oeb[27]
+ mprj_io_out[27] mprj_io_slow_sel[27] mprj_io_vtrip_sel[27] mprj_io_in[27] resetb
+ porb_h resetb_core_h vccd vccd1 vccd1_pad vccd2 vccd2_pad vccd_pad vdda vdda1 vdda1_pad
+ vdda2 vdda2_pad vdda_pad vddio vddio_pad vssa vssa1 vssa1_pad vssa2 vssa2_pad vssa_pad
+ vssd vssd1 vssd1_pad vssd2 vssd2_pad vssd_pad vssio vssio_pad vssio_pad2 vddio_pad2
+ vssa1_pad2 vdda1_pad2
.ends

* Black-box entry subcircuit for mgmt_core abstract view
.subckt mgmt_core clock core_clk core_rstn flash_clk flash_clk_ieb flash_clk_oeb flash_csb
+ flash_csb_ieb flash_csb_oeb flash_io0_di flash_io0_do flash_io0_ieb flash_io0_oeb
+ flash_io1_di flash_io1_do flash_io1_ieb flash_io1_oeb gpio_in_pad gpio_inenb_pad
+ gpio_mode0_pad gpio_mode1_pad gpio_out_pad gpio_outenb_pad jtag_out jtag_outenb
+ la_input[0] la_input[100] la_input[101] la_input[102] la_input[103] la_input[104]
+ la_input[105] la_input[106] la_input[107] la_input[108] la_input[109] la_input[10]
+ la_input[110] la_input[111] la_input[112] la_input[113] la_input[114] la_input[115]
+ la_input[116] la_input[117] la_input[118] la_input[119] la_input[11] la_input[120]
+ la_input[121] la_input[122] la_input[123] la_input[124] la_input[125] la_input[126]
+ la_input[127] la_input[12] la_input[13] la_input[14] la_input[15] la_input[16] la_input[17]
+ la_input[18] la_input[19] la_input[1] la_input[20] la_input[21] la_input[22] la_input[23]
+ la_input[24] la_input[25] la_input[26] la_input[27] la_input[28] la_input[29] la_input[2]
+ la_input[30] la_input[31] la_input[32] la_input[33] la_input[34] la_input[35] la_input[36]
+ la_input[37] la_input[38] la_input[39] la_input[3] la_input[40] la_input[41] la_input[42]
+ la_input[43] la_input[44] la_input[45] la_input[46] la_input[47] la_input[48] la_input[49]
+ la_input[4] la_input[50] la_input[51] la_input[52] la_input[53] la_input[54] la_input[55]
+ la_input[56] la_input[57] la_input[58] la_input[59] la_input[5] la_input[60] la_input[61]
+ la_input[62] la_input[63] la_input[64] la_input[65] la_input[66] la_input[67] la_input[68]
+ la_input[69] la_input[6] la_input[70] la_input[71] la_input[72] la_input[73] la_input[74]
+ la_input[75] la_input[76] la_input[77] la_input[78] la_input[79] la_input[7] la_input[80]
+ la_input[81] la_input[82] la_input[83] la_input[84] la_input[85] la_input[86] la_input[87]
+ la_input[88] la_input[89] la_input[8] la_input[90] la_input[91] la_input[92] la_input[93]
+ la_input[94] la_input[95] la_input[96] la_input[97] la_input[98] la_input[99] la_input[9]
+ la_oen[0] la_oen[100] la_oen[101] la_oen[102] la_oen[103] la_oen[104] la_oen[105]
+ la_oen[106] la_oen[107] la_oen[108] la_oen[109] la_oen[10] la_oen[110] la_oen[111]
+ la_oen[112] la_oen[113] la_oen[114] la_oen[115] la_oen[116] la_oen[117] la_oen[118]
+ la_oen[119] la_oen[11] la_oen[120] la_oen[121] la_oen[122] la_oen[123] la_oen[124]
+ la_oen[125] la_oen[126] la_oen[127] la_oen[12] la_oen[13] la_oen[14] la_oen[15]
+ la_oen[16] la_oen[17] la_oen[18] la_oen[19] la_oen[1] la_oen[20] la_oen[21] la_oen[22]
+ la_oen[23] la_oen[24] la_oen[25] la_oen[26] la_oen[27] la_oen[28] la_oen[29] la_oen[2]
+ la_oen[30] la_oen[31] la_oen[32] la_oen[33] la_oen[34] la_oen[35] la_oen[36] la_oen[37]
+ la_oen[38] la_oen[39] la_oen[3] la_oen[40] la_oen[41] la_oen[42] la_oen[43] la_oen[44]
+ la_oen[45] la_oen[46] la_oen[47] la_oen[48] la_oen[49] la_oen[4] la_oen[50] la_oen[51]
+ la_oen[52] la_oen[53] la_oen[54] la_oen[55] la_oen[56] la_oen[57] la_oen[58] la_oen[59]
+ la_oen[5] la_oen[60] la_oen[61] la_oen[62] la_oen[63] la_oen[64] la_oen[65] la_oen[66]
+ la_oen[67] la_oen[68] la_oen[69] la_oen[6] la_oen[70] la_oen[71] la_oen[72] la_oen[73]
+ la_oen[74] la_oen[75] la_oen[76] la_oen[77] la_oen[78] la_oen[79] la_oen[7] la_oen[80]
+ la_oen[81] la_oen[82] la_oen[83] la_oen[84] la_oen[85] la_oen[86] la_oen[87] la_oen[88]
+ la_oen[89] la_oen[8] la_oen[90] la_oen[91] la_oen[92] la_oen[93] la_oen[94] la_oen[95]
+ la_oen[96] la_oen[97] la_oen[98] la_oen[99] la_oen[9] la_output[0] la_output[100]
+ la_output[101] la_output[102] la_output[103] la_output[104] la_output[105] la_output[106]
+ la_output[107] la_output[108] la_output[109] la_output[10] la_output[110] la_output[111]
+ la_output[112] la_output[113] la_output[114] la_output[115] la_output[116] la_output[117]
+ la_output[118] la_output[119] la_output[11] la_output[120] la_output[121] la_output[122]
+ la_output[123] la_output[124] la_output[125] la_output[126] la_output[127] la_output[12]
+ la_output[13] la_output[14] la_output[15] la_output[16] la_output[17] la_output[18]
+ la_output[19] la_output[1] la_output[20] la_output[21] la_output[22] la_output[23]
+ la_output[24] la_output[25] la_output[26] la_output[27] la_output[28] la_output[29]
+ la_output[2] la_output[30] la_output[31] la_output[32] la_output[33] la_output[34]
+ la_output[35] la_output[36] la_output[37] la_output[38] la_output[39] la_output[3]
+ la_output[40] la_output[41] la_output[42] la_output[43] la_output[44] la_output[45]
+ la_output[46] la_output[47] la_output[48] la_output[49] la_output[4] la_output[50]
+ la_output[51] la_output[52] la_output[53] la_output[54] la_output[55] la_output[56]
+ la_output[57] la_output[58] la_output[59] la_output[5] la_output[60] la_output[61]
+ la_output[62] la_output[63] la_output[64] la_output[65] la_output[66] la_output[67]
+ la_output[68] la_output[69] la_output[6] la_output[70] la_output[71] la_output[72]
+ la_output[73] la_output[74] la_output[75] la_output[76] la_output[77] la_output[78]
+ la_output[79] la_output[7] la_output[80] la_output[81] la_output[82] la_output[83]
+ la_output[84] la_output[85] la_output[86] la_output[87] la_output[88] la_output[89]
+ la_output[8] la_output[90] la_output[91] la_output[92] la_output[93] la_output[94]
+ la_output[95] la_output[96] la_output[97] la_output[98] la_output[99] la_output[9]
+ mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13] mask_rev[14] mask_rev[15]
+ mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1] mask_rev[20] mask_rev[21]
+ mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27] mask_rev[28]
+ mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3] mask_rev[4] mask_rev[5]
+ mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] mgmt_addr[0] mgmt_addr[1] mgmt_addr[2]
+ mgmt_addr[3] mgmt_addr[4] mgmt_addr[5] mgmt_addr[6] mgmt_addr[7] mgmt_addr_ro[0]
+ mgmt_addr_ro[1] mgmt_addr_ro[2] mgmt_addr_ro[3] mgmt_addr_ro[4] mgmt_addr_ro[5]
+ mgmt_addr_ro[6] mgmt_addr_ro[7] mgmt_ena[0] mgmt_ena[1] mgmt_ena_ro mgmt_in_data[0]
+ mgmt_in_data[10] mgmt_in_data[11] mgmt_in_data[12] mgmt_in_data[13] mgmt_in_data[14]
+ mgmt_in_data[15] mgmt_in_data[16] mgmt_in_data[17] mgmt_in_data[18] mgmt_in_data[19]
+ mgmt_in_data[1] mgmt_in_data[20] mgmt_in_data[21] mgmt_in_data[22] mgmt_in_data[23]
+ mgmt_in_data[24] mgmt_in_data[25] mgmt_in_data[26] mgmt_in_data[27] mgmt_in_data[28]
+ mgmt_in_data[29] mgmt_in_data[2] mgmt_in_data[30] mgmt_in_data[31] mgmt_in_data[32]
+ mgmt_in_data[33] mgmt_in_data[34] mgmt_in_data[35] mgmt_in_data[36] mgmt_in_data[37]
+ mgmt_in_data[3] mgmt_in_data[4] mgmt_in_data[5] mgmt_in_data[6] mgmt_in_data[7]
+ mgmt_in_data[8] mgmt_in_data[9] mgmt_out_data[0] mgmt_out_data[10] mgmt_out_data[11]
+ mgmt_out_data[12] mgmt_out_data[13] mgmt_out_data[14] mgmt_out_data[15] mgmt_out_data[16]
+ mgmt_out_data[17] mgmt_out_data[18] mgmt_out_data[19] mgmt_out_data[1] mgmt_out_data[20]
+ mgmt_out_data[21] mgmt_out_data[22] mgmt_out_data[23] mgmt_out_data[24] mgmt_out_data[25]
+ mgmt_out_data[26] mgmt_out_data[27] mgmt_out_data[28] mgmt_out_data[29] mgmt_out_data[2]
+ mgmt_out_data[30] mgmt_out_data[31] mgmt_out_data[32] mgmt_out_data[33] mgmt_out_data[34]
+ mgmt_out_data[35] mgmt_out_data[36] mgmt_out_data[37] mgmt_out_data[3] mgmt_out_data[4]
+ mgmt_out_data[5] mgmt_out_data[6] mgmt_out_data[7] mgmt_out_data[8] mgmt_out_data[9]
+ mgmt_rdata[0] mgmt_rdata[10] mgmt_rdata[11] mgmt_rdata[12] mgmt_rdata[13] mgmt_rdata[14]
+ mgmt_rdata[15] mgmt_rdata[16] mgmt_rdata[17] mgmt_rdata[18] mgmt_rdata[19] mgmt_rdata[1]
+ mgmt_rdata[20] mgmt_rdata[21] mgmt_rdata[22] mgmt_rdata[23] mgmt_rdata[24] mgmt_rdata[25]
+ mgmt_rdata[26] mgmt_rdata[27] mgmt_rdata[28] mgmt_rdata[29] mgmt_rdata[2] mgmt_rdata[30]
+ mgmt_rdata[31] mgmt_rdata[32] mgmt_rdata[33] mgmt_rdata[34] mgmt_rdata[35] mgmt_rdata[36]
+ mgmt_rdata[37] mgmt_rdata[38] mgmt_rdata[39] mgmt_rdata[3] mgmt_rdata[40] mgmt_rdata[41]
+ mgmt_rdata[42] mgmt_rdata[43] mgmt_rdata[44] mgmt_rdata[45] mgmt_rdata[46] mgmt_rdata[47]
+ mgmt_rdata[48] mgmt_rdata[49] mgmt_rdata[4] mgmt_rdata[50] mgmt_rdata[51] mgmt_rdata[52]
+ mgmt_rdata[53] mgmt_rdata[54] mgmt_rdata[55] mgmt_rdata[56] mgmt_rdata[57] mgmt_rdata[58]
+ mgmt_rdata[59] mgmt_rdata[5] mgmt_rdata[60] mgmt_rdata[61] mgmt_rdata[62] mgmt_rdata[63]
+ mgmt_rdata[6] mgmt_rdata[7] mgmt_rdata[8] mgmt_rdata[9] mgmt_rdata_ro[0] mgmt_rdata_ro[10]
+ mgmt_rdata_ro[11] mgmt_rdata_ro[12] mgmt_rdata_ro[13] mgmt_rdata_ro[14] mgmt_rdata_ro[15]
+ mgmt_rdata_ro[16] mgmt_rdata_ro[17] mgmt_rdata_ro[18] mgmt_rdata_ro[19] mgmt_rdata_ro[1]
+ mgmt_rdata_ro[20] mgmt_rdata_ro[21] mgmt_rdata_ro[22] mgmt_rdata_ro[23] mgmt_rdata_ro[24]
+ mgmt_rdata_ro[25] mgmt_rdata_ro[26] mgmt_rdata_ro[27] mgmt_rdata_ro[28] mgmt_rdata_ro[29]
+ mgmt_rdata_ro[2] mgmt_rdata_ro[30] mgmt_rdata_ro[31] mgmt_rdata_ro[3] mgmt_rdata_ro[4]
+ mgmt_rdata_ro[5] mgmt_rdata_ro[6] mgmt_rdata_ro[7] mgmt_rdata_ro[8] mgmt_rdata_ro[9]
+ mgmt_wdata[0] mgmt_wdata[10] mgmt_wdata[11] mgmt_wdata[12] mgmt_wdata[13] mgmt_wdata[14]
+ mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17] mgmt_wdata[18] mgmt_wdata[19] mgmt_wdata[1]
+ mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23] mgmt_wdata[24] mgmt_wdata[25]
+ mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29] mgmt_wdata[2] mgmt_wdata[30]
+ mgmt_wdata[31] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5] mgmt_wdata[6] mgmt_wdata[7]
+ mgmt_wdata[8] mgmt_wdata[9] mgmt_wen[0] mgmt_wen[1] mgmt_wen_mask[0] mgmt_wen_mask[1]
+ mgmt_wen_mask[2] mgmt_wen_mask[3] mgmt_wen_mask[4] mgmt_wen_mask[5] mgmt_wen_mask[6]
+ mgmt_wen_mask[7] mprj2_vcc_pwrgood mprj2_vdd_pwrgood mprj_ack_i mprj_adr_o[0] mprj_adr_o[10]
+ mprj_adr_o[11] mprj_adr_o[12] mprj_adr_o[13] mprj_adr_o[14] mprj_adr_o[15] mprj_adr_o[16]
+ mprj_adr_o[17] mprj_adr_o[18] mprj_adr_o[19] mprj_adr_o[1] mprj_adr_o[20] mprj_adr_o[21]
+ mprj_adr_o[22] mprj_adr_o[23] mprj_adr_o[24] mprj_adr_o[25] mprj_adr_o[26] mprj_adr_o[27]
+ mprj_adr_o[28] mprj_adr_o[29] mprj_adr_o[2] mprj_adr_o[30] mprj_adr_o[31] mprj_adr_o[3]
+ mprj_adr_o[4] mprj_adr_o[5] mprj_adr_o[6] mprj_adr_o[7] mprj_adr_o[8] mprj_adr_o[9]
+ mprj_cyc_o mprj_dat_i[0] mprj_dat_i[10] mprj_dat_i[11] mprj_dat_i[12] mprj_dat_i[13]
+ mprj_dat_i[14] mprj_dat_i[15] mprj_dat_i[16] mprj_dat_i[17] mprj_dat_i[18] mprj_dat_i[19]
+ mprj_dat_i[1] mprj_dat_i[20] mprj_dat_i[21] mprj_dat_i[22] mprj_dat_i[23] mprj_dat_i[24]
+ mprj_dat_i[25] mprj_dat_i[26] mprj_dat_i[27] mprj_dat_i[28] mprj_dat_i[29] mprj_dat_i[2]
+ mprj_dat_i[30] mprj_dat_i[31] mprj_dat_i[3] mprj_dat_i[4] mprj_dat_i[5] mprj_dat_i[6]
+ mprj_dat_i[7] mprj_dat_i[8] mprj_dat_i[9] mprj_dat_o[0] mprj_dat_o[10] mprj_dat_o[11]
+ mprj_dat_o[12] mprj_dat_o[13] mprj_dat_o[14] mprj_dat_o[15] mprj_dat_o[16] mprj_dat_o[17]
+ mprj_dat_o[18] mprj_dat_o[19] mprj_dat_o[1] mprj_dat_o[20] mprj_dat_o[21] mprj_dat_o[22]
+ mprj_dat_o[23] mprj_dat_o[24] mprj_dat_o[25] mprj_dat_o[26] mprj_dat_o[27] mprj_dat_o[28]
+ mprj_dat_o[29] mprj_dat_o[2] mprj_dat_o[30] mprj_dat_o[31] mprj_dat_o[3] mprj_dat_o[4]
+ mprj_dat_o[5] mprj_dat_o[6] mprj_dat_o[7] mprj_dat_o[8] mprj_dat_o[9] mprj_io_loader_clock
+ mprj_io_loader_data mprj_io_loader_resetn mprj_sel_o[0] mprj_sel_o[1] mprj_sel_o[2]
+ mprj_sel_o[3] mprj_stb_o mprj_vcc_pwrgood mprj_vdd_pwrgood mprj_we_o porb pwr_ctrl_out[0]
+ pwr_ctrl_out[1] pwr_ctrl_out[2] pwr_ctrl_out[3] resetb sdo_out sdo_outenb user_clk
+ VPWR VGND
.ends

* Black-box entry subcircuit for simple_por abstract view
.subckt simple_por vdd3v3 vdd1v8 vss porb_h por_l porb_l
.ends

* Black-box entry subcircuit for user_id_programming abstract view
.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VPWR VGND
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[45] HI[46] HI[47] HI[48] HI[49] HI[4]
+ HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57] HI[58] HI[59] HI[5] HI[60]
+ HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68] HI[69] HI[6] HI[70] HI[71]
+ HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79] HI[7] HI[80] HI[81] HI[82]
+ HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8] HI[90] HI[91] HI[92] HI[93]
+ HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1 vssd1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__decap_8 abstract view
.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__conb_1 abstract view
.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_2 abstract view
.subckt sky130_fd_sc_hvl__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__decap_4 abstract view
.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_1 abstract view
.subckt sky130_fd_sc_hvl__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__lsbufhv2lv_1 abstract view
.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
.ends

.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2
+ vssa2 FILLER_2_300/li_65_797# FILLER_1_260/li_65_797# FILLER_2_115/li_737_n17# FILLER_1_131/li_0_n17#
+ FILLER_1_32/li_161_n17# FILLER_1_8/li_161_n17# FILLER_1_48/li_641_797# FILLER_2_243/li_0_797#
+ FILLER_2_115/li_257_797# FILLER_0_216/li_100_536# FILLER_2_155/li_545_797# FILLER_2_24/li_545_797#
+ FILLER_0_216/li_449_797# mprj2_logic_high_lv/li_514_79# FILLER_1_107/li_353_n17#
+ FILLER_0_264/li_0_797# FILLER_2_227/li_545_n17# mprj2_logic_high_hvl/li_161_797#
+ FILLER_0_32/li_353_797# FILLER_0_176/li_545_797# FILLER_2_187/li_641_n17# mprj2_logic_high_lv/li_161_1611#
+ FILLER_2_16/li_353_n17# FILLER_1_131/li_353_n17# FILLER_1_180/li_161_n17# FILLER_1_24/li_65_n17#
+ FILLER_1_131/li_34_73# FILLER_2_267/li_353_797# FILLER_1_268/li_0_797# FILLER_1_188/li_65_797#
+ FILLER_0_232/li_0_n17# FILLER_0_96/li_65_797# FILLER_2_259/li_161_n17# FILLER_1_156/li_0_797#
+ FILLER_1_268/li_641_n17# FILLER_0_224/li_115_72# FILLER_0_112/li_115_72# FILLER_2_300/li_65_n17#
+ mprj2_logic_high_lv/li_34_216# FILLER_2_171/li_0_797# FILLER_2_32/li_737_797# FILLER_1_48/li_641_n17#
+ FILLER_1_115/li_545_n17# FILLER_2_115/li_257_n17# FILLER_1_260/li_115_72# FILLER_2_243/li_0_n17#
+ FILLER_2_155/li_545_n17# mprj2_logic_high_lv/li_179_1349# FILLER_2_24/li_545_n17#
+ FILLER_1_204/li_100_536# mprj_logic_high_lv/li_545_1611# FILLER_0_264/li_0_n17#
+ FILLER_1_48/li_161_797# mprj2_logic_high_hvl/li_161_n17# FILLER_2_235/li_257_797#
+ FILLER_2_195/li_115_72# FILLER_2_8/li_65_797# FILLER_1_220/li_65_n17# FILLER_0_104/li_641_797#
+ FILLER_2_195/li_353_797# FILLER_0_256/li_257_797# FILLER_1_236/li_545_n17# FILLER_0_160/li_0_n17#
+ FILLER_2_267/li_353_n17# FILLER_1_196/li_641_n17# FILLER_2_187/li_161_n17# FILLER_2_267/li_65_n17#
+ FILLER_2_155/li_65_n17# FILLER_1_16/li_545_n17# FILLER_2_171/li_0_n17# mprj2_logic_high_lv/li_26_452#
+ FILLER_1_188/li_115_72# FILLER_2_32/li_737_n17# mprj_logic_high_lv/m1_0_n23# FILLER_2_219/li_115_72#
+ FILLER_2_107/li_115_72# FILLER_1_268/li_161_n17# FILLER_2_243/li_100_536# FILLER_2_243/li_449_797#
+ FILLER_0_24/li_0_797# FILLER_2_163/li_257_797# FILLER_2_32/li_257_797# FILLER_0_264/li_100_536#
+ FILLER_0_208/li_65_n17# FILLER_1_48/li_161_n17# FILLER_0_264/li_449_797# FILLER_2_235/li_257_n17#
+ FILLER_2_8/li_65_n17# FILLER_0_0/li_545_797# FILLER_1_164/li_545_n17# FILLER_0_184/li_257_797#
+ FILLER_2_195/li_353_n17# FILLER_0_232/li_0_797# FILLER_0_80/li_353_797# mprj2_logic_high_lv/li_1313_1611#
+ FILLER_0_232/li_65_797# FILLER_2_203/li_641_797# FILLER_1_32/li_0_n17# FILLER_0_224/li_641_797#
+ FILLER_0_104/li_161_797# mprj_logic_high_lv/li_1505_797# FILLER_2_195/li_0_797#
+ FILLER_1_62/li_65_797# FILLER_0_88/li_641_797# FILLER_1_196/li_161_n17# FILLER_2_171/li_100_536#
+ FILLER_2_171/li_449_797# FILLER_2_0/li_0_797# FILLER_0_192/li_100_536# FILLER_2_243/li_449_n17#
+ FILLER_2_163/li_257_n17# mprj2_logic_high_lv/li_34_1244# FILLER_0_272/li_115_72#
+ FILLER_0_192/li_449_797# FILLER_0_160/li_115_72# FILLER_1_180/li_0_n17# FILLER_2_32/li_257_n17#
+ FILLER_2_187/li_0_797# FILLER_1_252/li_100_536# FILLER_1_24/li_115_72# FILLER_2_251/li_545_797#
+ FILLER_0_16/li_257_797# FILLER_2_203/li_641_n17# FILLER_0_112/li_353_797# FILLER_1_244/li_257_n17#
+ FILLER_1_32/li_100_536# FILLER_2_8/li_0_797# FILLER_1_8/li_100_536# FILLER_0_104/li_161_n17#
+ FILLER_2_195/li_0_n17# FILLER_1_62/li_65_n17# FILLER_1_204/li_65_797# FILLER_2_115/li_65_797#
+ FILLER_1_24/li_257_n17# FILLER_2_171/li_449_n17# FILLER_0_224/li_161_797# FILLER_0_8/li_353_797#
+ FILLER_0_88/li_161_797# FILLER_2_32/li_0_797# FILLER_2_0/li_0_n17# FILLER_1_140/li_0_797#
+ FILLER_1_220/li_115_72# FILLER_0_24/li_100_536# FILLER_1_180/li_100_536# FILLER_0_208/li_0_797#
+ mprj_logic_high_lv/m1_0_51# FILLER_0_24/li_449_797# FILLER_2_187/li_0_n17# FILLER_2_267/li_115_72#
+ FILLER_0_256/li_65_n17# FILLER_0_96/li_115_72# FILLER_2_259/li_100_536# FILLER_2_155/li_115_72#
+ FILLER_1_62/li_545_797# FILLER_1_172/li_257_n17# FILLER_2_259/li_449_797# FILLER_2_179/li_257_797#
+ FILLER_0_0/li_0_797# FILLER_2_211/li_353_797# FILLER_1_140/li_641_797# FILLER_2_8/li_0_n17#
+ FILLER_1_32/li_449_n17# FILLER_1_196/li_65_n17# FILLER_1_8/li_449_n17# FILLER_2_227/li_65_n17#
+ FILLER_2_203/li_161_n17# FILLER_2_115/li_65_n17# FILLER_0_232/li_353_797# FILLER_1_212/li_641_n17#
+ FILLER_1_0/li_0_n17# FILLER_0_96/li_353_797# FILLER_0_272/li_641_797# FILLER_1_0/li_641_n17#
+ FILLER_2_219/li_641_797# FILLER_2_0/li_257_797# FILLER_1_62/li_0_797# FILLER_2_32/li_0_n17#
+ FILLER_1_140/li_0_n17# mprj_logic_high_lv/li_449_1611# FILLER_2_8/li_115_72# FILLER_2_8/li_545_797#
+ FILLER_0_208/li_0_n17# FILLER_1_16/li_0_n17# FILLER_0_184/li_65_n17# FILLER_2_187/li_100_536#
+ FILLER_2_187/li_449_797# FILLER_1_62/li_545_n17# FILLER_2_259/li_449_n17# FILLER_0_200/li_257_797#
+ mprj_logic_high_lv/li_833_1611# FILLER_2_211/li_353_n17# FILLER_2_179/li_257_n17#
+ FILLER_0_240/li_545_797# FILLER_1_140/li_641_n17# FILLER_2_251/li_641_n17# FILLER_0_160/li_353_797#
+ FILLER_2_107/li_353_797# FILLER_1_268/li_100_536# FILLER_2_16/li_641_797# FILLER_0_272/li_641_n17#
+ FILLER_0_208/li_545_797# FILLER_0_96/li_353_n17# FILLER_2_0/li_257_n17# FILLER_2_219/li_641_n17#
+ FILLER_1_140/li_161_797# mprj2_logic_high_lv/m1_0_51# FILLER_1_48/li_100_536# FILLER_0_168/li_641_797#
+ FILLER_1_48/li_449_797# FILLER_1_212/li_161_n17# mprj2_logic_high_lv/li_1455_797#
+ FILLER_1_32/li_65_n17# FILLER_1_62/li_0_n17# FILLER_0_272/li_161_797# FILLER_1_0/li_161_n17#
+ FILLER_1_220/li_65_797# FILLER_1_164/li_0_797# FILLER_2_8/li_545_n17# FILLER_0_232/li_115_72#
+ FILLER_2_187/li_449_n17# mprj2_logic_high_lv/li_1217_1611# FILLER_1_62/li_115_72#
+ mprj_logic_high_lv/li_34_1244# FILLER_2_115/li_545_797# FILLER_1_196/li_100_536#
+ FILLER_0_224/li_0_797# FILLER_1_107/li_641_n17# mprj_logic_high_lv/li_1121_1611#
+ FILLER_2_107/li_353_n17# FILLER_0_272/li_65_n17# FILLER_0_32/li_641_797# mprj2_logic_high_lv/li_1601_1611#
+ FILLER_2_16/li_641_n17# FILLER_0_16/li_65_797# FILLER_1_188/li_257_n17# mprj_logic_high_lv/li_179_79#
+ FILLER_0_224/li_0_n17# FILLER_1_140/li_161_n17# FILLER_2_251/li_161_n17# FILLER_1_260/li_641_n17#
+ FILLER_2_227/li_353_797# FILLER_1_48/li_449_n17# FILLER_2_267/li_641_797# FILLER_2_16/li_161_797#
+ FILLER_0_248/li_353_797# FILLER_1_228/li_641_n17# FILLER_2_219/li_161_n17# FILLER_2_163/li_65_n17#
+ mprj2_logic_high_lv/li_26_893# FILLER_0_168/li_161_797# FILLER_0_104/li_100_536#
+ FILLER_1_196/li_115_72# FILLER_0_104/li_449_797# FILLER_2_227/li_115_72# FILLER_2_115/li_545_n17#
+ FILLER_2_115/li_115_72# FILLER_0_200/li_65_n17# FILLER_1_268/li_65_n17# mprj2_logic_high_lv/li_384_137#
+ FILLER_1_156/li_65_n17# FILLER_2_235/li_545_797# FILLER_2_155/li_353_797# FILLER_2_24/li_353_797#
+ FILLER_0_216/li_257_797# FILLER_1_107/li_161_n17# FILLER_2_195/li_641_797# FILLER_0_256/li_545_797#
+ FILLER_2_227/li_353_n17# FILLER_0_240/li_65_797# FILLER_0_32/li_161_797# FILLER_1_156/li_641_n17#
+ FILLER_0_176/li_353_797# FILLER_2_267/li_641_n17# FILLER_2_16/li_161_n17# FILLER_1_196/li_0_n17#
+ FILLER_1_268/li_65_797# FILLER_1_228/li_161_n17# FILLER_1_107/li_65_n17# FILLER_2_203/li_100_536#
+ FILLER_2_203/li_449_797# FILLER_2_251/li_0_797# mprj2_logic_high_lv/li_353_1611#
+ FILLER_0_224/li_100_536# FILLER_2_163/li_545_797# FILLER_2_32/li_545_797# FILLER_0_224/li_449_797#
+ FILLER_0_88/li_100_536# FILLER_1_115/li_353_n17# FILLER_0_88/li_449_797# FILLER_2_235/li_545_n17#
+ FILLER_2_155/li_353_n17# FILLER_1_32/li_115_72# FILLER_0_168/li_65_797# FILLER_0_184/li_545_797#
+ FILLER_2_195/li_641_n17# FILLER_2_24/li_353_n17# FILLER_0_80/li_641_797# FILLER_1_260/li_161_n17#
+ FILLER_1_196/li_65_797# FILLER_0_240/li_0_n17# FILLER_1_236/li_0_797# FILLER_1_156/li_161_n17#
+ FILLER_2_267/li_161_n17# mprj_logic_high_lv/li_737_1611# FILLER_2_179/li_0_797#
+ FILLER_1_16/li_353_n17# FILLER_2_203/li_449_n17# FILLER_2_251/li_0_n17# FILLER_0_200/li_0_797#
+ FILLER_2_163/li_545_n17# mprj2_logic_high_hvl/li_43_635# FILLER_2_32/li_545_n17#
+ FILLER_0_216/li_0_797# FILLER_1_212/li_100_536# FILLER_1_0/li_100_536# FILLER_1_260/li_0_797#
+ FILLER_2_243/li_257_797# FILLER_0_16/li_545_797# FILLER_2_163/li_115_72# FILLER_1_300/li_65_n17#
+ FILLER_0_112/li_641_797# FILLER_0_264/li_257_797# FILLER_1_244/li_545_n17# FILLER_0_0/li_353_797#
+ FILLER_0_168/li_0_n17# FILLER_2_195/li_161_n17# mprj2_logic_high_hvl/li_307_57#
+ FILLER_0_80/li_161_797# FILLER_2_235/li_65_n17# FILLER_1_24/li_545_n17# FILLER_1_268/li_115_72#
+ FILLER_0_8/li_641_797# FILLER_1_156/li_115_72# FILLER_2_179/li_0_n17# mprj_logic_high_lv/li_1025_1611#
+ FILLER_0_16/li_115_72# FILLER_1_140/li_100_536# FILLER_0_160/li_0_797# FILLER_2_251/li_100_536#
+ FILLER_1_140/li_449_797# FILLER_1_131/li_257_797# FILLER_1_188/li_0_797# mprj2_logic_high_lv/li_1505_1611#
+ FILLER_0_32/li_0_797# FILLER_2_171/li_257_797# FILLER_0_272/li_100_536# FILLER_1_228/li_65_n17#
+ FILLER_0_216/li_65_n17# FILLER_0_272/li_449_797# FILLER_1_260/li_0_n17# FILLER_2_243/li_257_n17#
+ FILLER_2_219/li_100_536# FILLER_0_192/li_257_797# FILLER_1_0/li_449_n17# FILLER_1_172/li_545_n17#
+ FILLER_2_219/li_449_797# FILLER_2_267/li_0_797# FILLER_2_179/li_545_797# FILLER_2_251/li_353_797#
+ FILLER_2_211/li_641_797# mprj_logic_high_lv/li_384_137# FILLER_0_200/li_65_797#
+ FILLER_1_32/li_737_n17# FILLER_1_107/li_115_72# FILLER_0_232/li_641_797# FILLER_0_112/li_161_797#
+ FILLER_2_16/li_0_797# FILLER_0_96/li_641_797# FILLER_2_0/li_545_797# mprj_logic_high_hvl/li_353_797#
+ FILLER_1_107/li_100_536# FILLER_1_131/li_257_n17# FILLER_1_140/li_449_n17# FILLER_2_251/li_449_n17#
+ FILLER_2_171/li_257_n17# FILLER_0_240/li_115_72# FILLER_0_8/li_161_797# FILLER_1_188/li_0_n17#
+ FILLER_2_16/li_100_536# FILLER_2_16/li_449_797# FILLER_0_272/li_449_n17# FILLER_1_260/li_100_536#
+ FILLER_0_168/li_100_536# FILLER_2_219/li_449_n17# FILLER_0_168/li_449_797# FILLER_2_267/li_0_n17#
+ FILLER_0_200/li_545_797# FILLER_0_24/li_257_797# FILLER_2_179/li_545_n17# FILLER_2_211/li_641_n17#
+ FILLER_1_252/li_257_n17# FILLER_1_228/li_100_536# FILLER_0_160/li_641_797# FILLER_2_107/li_641_797#
+ FILLER_1_62/li_353_797# FILLER_1_268/li_737_797# FILLER_2_259/li_257_797# FILLER_2_16/li_0_n17#
+ FILLER_0_96/li_641_n17# FILLER_0_24/li_65_797# FILLER_1_212/li_65_797# FILLER_2_0/li_545_n17#
+ FILLER_1_32/li_257_n17# mprj_logic_high_hvl/li_353_n17# FILLER_1_8/li_257_n17# FILLER_0_0/li_65_797#
+ mprj_logic_high_lv/li_65_797# mprj2_logic_high_lv/li_257_1611# FILLER_1_48/li_737_797#
+ FILLER_0_232/li_161_797# FILLER_0_168/li_115_72# FILLER_1_48/li_0_797# FILLER_0_96/li_161_797#
+ FILLER_0_112/li_0_n17# FILLER_2_171/li_65_n17# FILLER_0_32/li_100_536# mprj2_logic_high_hvl/li_257_797#
+ FILLER_2_16/li_449_n17# FILLER_0_32/li_449_797# mprj2_logic_high_lv/li_641_1611#
+ FILLER_2_8/li_353_797# FILLER_0_264/li_65_n17# FILLER_2_235/li_115_72# FILLER_1_156/li_100_536#
+ FILLER_1_180/li_257_n17# FILLER_1_204/li_161_n17# FILLER_2_267/li_100_536# FILLER_2_267/li_449_797#
+ FILLER_1_204/li_0_797# FILLER_2_187/li_257_797# mprj_logic_high_hvl/li_43_635# FILLER_0_232/li_65_n17#
+ FILLER_2_107/li_641_n17# FILLER_1_268/li_737_n17# FILLER_1_62/li_353_n17# FILLER_1_164/li_65_n17#
+ FILLER_2_259/li_257_n17# FILLER_1_188/li_545_n17# FILLER_2_211/li_161_n17# FILLER_0_240/li_353_797#
+ FILLER_1_220/li_641_n17# FILLER_0_160/li_161_797# FILLER_2_227/li_641_797# FILLER_2_107/li_161_797#
+ FILLER_1_48/li_737_n17# FILLER_1_228/li_115_72# FILLER_0_208/li_353_797# mprj_logic_high_hvl/li_307_57#
+ FILLER_0_248/li_641_797# FILLER_1_48/li_0_n17# FILLER_1_48/li_257_797# mprj2_logic_high_hvl/li_257_n17#
+ FILLER_2_195/li_100_536# mprj2_logic_high_lv/li_384_1039# FILLER_0_112/li_0_797#
+ FILLER_2_195/li_449_797# FILLER_2_8/li_353_n17# FILLER_1_115/li_65_n17# FILLER_0_160/li_65_n17#
+ FILLER_2_267/li_449_n17# FILLER_1_204/li_0_n17# FILLER_2_187/li_257_n17# FILLER_2_107/li_0_797#
+ FILLER_2_115/li_353_797# mprj_logic_high_lv/li_826_79# FILLER_2_155/li_641_797#
+ FILLER_0_216/li_545_797# FILLER_0_176/li_65_797# FILLER_2_24/li_641_797# FILLER_2_227/li_641_n17#
+ FILLER_2_107/li_161_n17# FILLER_1_268/li_257_n17# FILLER_0_176/li_641_797# mprj2_logic_high_lv/li_1409_1611#
+ FILLER_1_220/li_161_n17# FILLER_1_228/li_65_797# FILLER_1_48/li_257_n17# FILLER_0_200/li_115_72#
+ mprj_logic_high_lv/li_1313_1611# FILLER_0_248/li_161_797# FILLER_0_80/li_100_536#
+ FILLER_2_195/li_449_n17# FILLER_0_80/li_449_797# FILLER_2_107/li_0_n17# FILLER_0_104/li_257_797#
+ FILLER_1_115/li_641_n17# mprj2_logic_high_lv/li_506_1123# FILLER_0_96/li_0_797#
+ FILLER_2_155/li_0_797# FILLER_2_115/li_353_n17# mprj_logic_high_lv/li_514_79# FILLER_2_155/li_641_n17#
+ FILLER_2_24/li_641_n17# FILLER_1_196/li_257_n17# FILLER_2_171/li_115_72# FILLER_2_235/li_353_797#
+ FILLER_1_156/li_65_797# FILLER_2_24/li_161_797# FILLER_0_256/li_353_797# FILLER_1_236/li_641_n17#
+ FILLER_2_243/li_65_n17# FILLER_2_227/li_161_n17# FILLER_0_176/li_161_797# FILLER_2_16/li_65_797#
+ FILLER_0_112/li_100_536# mprj_logic_high_lv/li_34_216# FILLER_1_16/li_641_n17# FILLER_0_112/li_449_797#
+ FILLER_1_164/li_115_72# FILLER_0_24/li_115_72# FILLER_0_0/li_115_72# FILLER_2_155/li_0_n17#
+ FILLER_2_203/li_257_797# mprj2_logic_high_lv/li_0_1611# FILLER_1_236/li_65_n17#
+ FILLER_2_243/li_545_797# FILLER_0_8/li_100_536# FILLER_2_163/li_353_797# FILLER_2_32/li_353_797#
+ FILLER_0_224/li_257_797# FILLER_1_204/li_545_n17# FILLER_0_8/li_449_797# FILLER_1_115/li_161_n17#
+ FILLER_0_264/li_545_797# FILLER_0_88/li_257_797# FILLER_2_235/li_353_n17# FILLER_2_155/li_161_n17#
+ FILLER_1_164/li_641_n17# FILLER_0_184/li_353_797# FILLER_2_24/li_161_n17# FILLER_0_0/li_641_797#
+ FILLER_1_115/li_115_72# mprj2_logic_high_lv/li_545_1611# FILLER_2_16/li_65_n17#
+ FILLER_2_300/li_0_797# FILLER_1_236/li_161_n17# mprj_logic_high_lv/li_26_452# FILLER_2_211/li_100_536#
+ FILLER_2_211/li_449_797# FILLER_1_140/li_737_797# FILLER_0_232/li_100_536# FILLER_2_171/li_545_797#
+ FILLER_1_220/li_0_n17# FILLER_1_16/li_161_n17# FILLER_0_96/li_100_536# FILLER_2_203/li_257_n17#
+ FILLER_0_272/li_737_797# FILLER_0_232/li_449_797# FILLER_0_96/li_449_797# FILLER_2_243/li_545_n17#
+ FILLER_0_248/li_65_797# FILLER_0_192/li_545_797# FILLER_1_8/li_0_n17# FILLER_2_227/li_0_797#
+ FILLER_2_163/li_353_n17# FILLER_2_32/li_353_n17# FILLER_2_251/li_641_797# FILLER_0_16/li_353_797#
+ mprj_logic_high_lv/li_929_1611# mprj2_logic_high_lv/li_756_683# FILLER_0_248/li_0_n17#
+ FILLER_0_32/li_65_797# FILLER_1_164/li_161_n17# FILLER_1_252/li_0_797# FILLER_0_0/li_161_797#
+ FILLER_1_24/li_353_n17# FILLER_0_160/li_100_536# FILLER_0_176/li_115_72# FILLER_2_211/li_449_n17#
+ FILLER_1_140/li_737_n17# FILLER_0_160/li_449_797# FILLER_2_259/li_0_n17# FILLER_2_107/li_100_536#
+ FILLER_2_171/li_545_n17# FILLER_2_107/li_449_797# FILLER_2_24/li_0_797# FILLER_0_272/li_737_n17#
+ FILLER_1_220/li_100_536# FILLER_0_96/li_449_n17# FILLER_2_227/li_0_n17# FILLER_1_140/li_257_797#
+ mprj2_logic_high_lv/li_1505_797# FILLER_0_24/li_545_797# FILLER_2_243/li_115_72#
+ FILLER_1_212/li_257_n17# FILLER_0_272/li_257_797# FILLER_1_252/li_545_n17# FILLER_1_62/li_641_797#
+ FILLER_1_0/li_257_n17# FILLER_0_176/li_0_n17# FILLER_2_219/li_257_797# mprj2_logic_high_hvl/li_0_797#
+ FILLER_1_172/li_65_n17# mprj_logic_high_lv/li_1217_1611# FILLER_2_259/li_545_797#
+ FILLER_2_179/li_353_797# FILLER_2_203/li_65_n17# FILLER_1_252/li_0_n17# FILLER_1_32/li_545_n17#
+ FILLER_0_192/li_0_797# FILLER_1_8/li_545_n17# FILLER_1_236/li_115_72# FILLER_2_0/li_353_797#
+ FILLER_1_115/li_0_n17# FILLER_2_300/li_0_n17# mprj_logic_high_hvl/li_161_797# FILLER_2_107/li_449_n17#
+ mprj_logic_high_lv/li_161_1611# FILLER_0_32/li_737_797# FILLER_2_24/li_0_n17# FILLER_0_224/li_65_n17#
+ FILLER_2_8/li_641_797# FILLER_1_268/li_0_n17# FILLER_1_140/li_257_n17# FILLER_2_251/li_257_n17#
+ FILLER_2_227/li_100_536# FILLER_1_180/li_545_n17# FILLER_2_227/li_449_797# FILLER_2_16/li_115_72#
+ FILLER_2_267/li_737_797# FILLER_2_187/li_545_797# FILLER_2_16/li_257_797# FILLER_0_248/li_100_536#
+ FILLER_2_219/li_257_n17# FILLER_0_248/li_449_797# FILLER_1_236/li_0_n17# FILLER_1_62/li_641_n17#
+ FILLER_0_168/li_257_797# FILLER_2_259/li_545_n17# FILLER_0_200/li_353_797# mprj2_logic_high_hvl/li_0_n17#
+ FILLER_2_179/li_353_n17# FILLER_0_240/li_641_797# FILLER_0_184/li_65_797# FILLER_1_62/li_161_797#
+ mprj_logic_high_lv/li_179_1349# FILLER_1_48/li_65_797# FILLER_0_208/li_641_797#
+ FILLER_2_0/li_353_n17# FILLER_1_115/li_100_536# FILLER_0_80/li_65_797# mprj_logic_high_hvl/li_161_n17#
+ FILLER_2_155/li_100_536# FILLER_1_48/li_545_797# FILLER_2_24/li_100_536# FILLER_2_155/li_449_797#
+ FILLER_2_24/li_449_797# FILLER_2_8/li_641_n17# FILLER_1_107/li_257_n17# FILLER_2_227/li_449_n17#
+ FILLER_2_203/li_0_797# FILLER_0_208/li_65_797# FILLER_1_0/li_65_n17# FILLER_1_164/li_0_n17#
+ FILLER_0_176/li_100_536# FILLER_2_267/li_737_n17# FILLER_2_16/li_257_n17# FILLER_0_32/li_257_797#
+ FILLER_0_176/li_449_797# FILLER_2_187/li_545_n17# FILLER_1_156/li_0_n17# FILLER_2_8/li_161_797#
+ FILLER_1_236/li_100_536# FILLER_2_115/li_641_797# mprj2_logic_high_lv/li_449_1611#
+ FILLER_2_235/li_0_797# FILLER_2_267/li_257_797# FILLER_1_228/li_257_n17# FILLER_1_268/li_545_n17#
+ FILLER_1_16/li_100_536# FILLER_1_48/li_65_n17# FILLER_1_62/li_161_n17# FILLER_0_192/li_0_n17#
+ FILLER_1_180/li_0_797# FILLER_0_240/li_161_797# mprj_logic_high_lv/m1_0_689# mprj_logic_high_lv/li_756_683#
+ mprj2_logic_high_lv/li_833_1611# mprj2_logic_high_hvl/li_65_797# FILLER_0_248/li_115_72#
+ FILLER_1_48/li_545_n17# FILLER_0_80/li_65_n17# FILLER_1_115/li_449_n17# FILLER_2_251/li_65_n17#
+ FILLER_0_208/li_161_797# FILLER_2_155/li_449_n17# FILLER_2_24/li_65_797# FILLER_2_203/li_0_n17#
+ FILLER_2_24/li_449_n17# FILLER_0_88/li_0_797# FILLER_1_172/li_115_72# FILLER_0_32/li_115_72#
+ FILLER_1_164/li_100_536# FILLER_2_203/li_115_72# FILLER_0_104/li_545_797# FILLER_2_195/li_257_797#
+ FILLER_2_8/li_161_n17# FILLER_2_235/li_0_n17# FILLER_2_115/li_641_n17# FILLER_1_244/li_65_n17#
+ FILLER_0_240/li_65_n17# FILLER_1_156/li_257_n17# FILLER_2_267/li_257_n17# FILLER_0_8/li_65_797#
+ FILLER_1_196/li_545_n17# mprj2_logic_high_lv/li_161_797# FILLER_1_16/li_449_n17#
+ FILLER_2_235/li_641_797# FILLER_2_115/li_161_797# FILLER_2_179/li_65_n17# mprj2_logic_high_hvl/li_65_n17#
+ FILLER_0_216/li_353_797# FILLER_0_256/li_641_797# FILLER_2_24/li_65_n17# FILLER_1_300/li_161_n17#
+ mprj_logic_high_lv/li_26_893# FILLER_0_112/li_737_797# FILLER_0_0/li_100_536# FILLER_0_168/li_65_n17#
+ FILLER_0_0/li_449_797# FILLER_2_195/li_257_n17# FILLER_0_80/li_257_797# FILLER_2_203/li_545_797#
+ FILLER_2_163/li_641_797# FILLER_0_256/li_65_797# mprj2_logic_high_lv/li_65_1611#
+ FILLER_2_32/li_641_797# FILLER_0_224/li_545_797# FILLER_0_88/li_545_797# FILLER_2_235/li_641_n17#
+ FILLER_2_115/li_161_n17# FILLER_0_184/li_641_797# mprj_logic_high_lv/li_1505_1611#
+ FILLER_1_260/li_257_n17# FILLER_1_0/li_115_72# FILLER_1_236/li_65_797# FILLER_1_212/li_0_797#
+ FILLER_0_256/li_161_797# FILLER_0_184/li_115_72# FILLER_2_219/li_0_797# FILLER_1_48/li_115_72#
+ FILLER_0_112/li_257_797# FILLER_2_203/li_545_n17# FILLER_0_240/li_0_797# FILLER_0_104/li_0_797#
+ FILLER_2_163/li_641_n17# FILLER_2_32/li_641_n17# FILLER_2_251/li_115_72# FILLER_1_131/li_65_797#
+ FILLER_0_80/li_115_72# mprj2_logic_high_lv/m1_0_689# FILLER_2_243/li_353_797# FILLER_0_16/li_641_797#
+ FILLER_1_164/li_65_797# FILLER_0_8/li_257_797# FILLER_1_180/li_65_n17# FILLER_2_32/li_161_797#
+ FILLER_0_264/li_353_797# FILLER_1_244/li_641_n17# FILLER_0_208/li_115_72# FILLER_2_235/li_161_n17#
+ FILLER_0_184/li_161_797# FILLER_2_211/li_65_n17# FILLER_0_272/li_0_797# mprj_logic_high_lv/li_0_797#
+ mprj_logic_high_hvl/li_65_797# FILLER_1_244/li_115_72# FILLER_1_24/li_641_n17# FILLER_2_219/li_0_n17#
+ FILLER_0_168/li_0_797# FILLER_1_62/li_100_536# FILLER_2_115/li_0_797# FILLER_1_62/li_449_797#
+ FILLER_0_104/li_0_n17# FILLER_1_228/li_0_797# FILLER_2_179/li_115_72# FILLER_2_211/li_257_797#
+ FILLER_1_140/li_545_797# FILLER_1_131/li_65_n17# mprj_logic_high_lv/li_1455_797#
+ FILLER_2_171/li_353_797# FILLER_1_212/li_545_n17# mprj2_logic_high_lv/li_737_1611#
+ FILLER_2_24/li_115_72# FILLER_0_232/li_257_797# FILLER_0_96/li_257_797# FILLER_2_243/li_353_n17#
+ FILLER_0_272/li_545_797# FILLER_0_192/li_353_797# FILLER_1_0/li_545_n17# FILLER_1_172/li_641_n17#
+ FILLER_2_219/li_545_797# FILLER_2_163/li_161_n17# FILLER_2_32/li_161_n17# mprj_logic_high_lv/li_161_797#
+ FILLER_2_179/li_641_797# FILLER_0_192/li_65_797# FILLER_2_251/li_449_797# FILLER_2_8/li_100_536#
+ FILLER_1_300/li_0_n17# FILLER_0_16/li_161_797# FILLER_2_8/li_449_797# FILLER_1_244/li_161_n17#
+ mprj_logic_high_hvl/li_65_n17# FILLER_2_0/li_641_797# FILLER_0_8/li_115_72# FILLER_0_80/li_0_797#
+ FILLER_2_115/li_0_n17# FILLER_1_62/li_449_n17# FILLER_0_240/li_100_536# FILLER_1_228/li_0_n17#
+ FILLER_1_24/li_161_n17# FILLER_2_211/li_257_n17# FILLER_0_240/li_449_797# FILLER_1_140/li_545_n17#
+ FILLER_0_160/li_257_797# FILLER_2_251/li_545_n17# FILLER_2_171/li_353_n17# FILLER_2_107/li_257_797#
+ FILLER_0_216/li_65_797# FILLER_0_208/li_100_536# FILLER_0_104/li_65_797# FILLER_2_211/li_0_797#
+ FILLER_2_16/li_545_797# FILLER_0_272/li_545_n17# FILLER_0_208/li_449_797# FILLER_2_219/li_545_n17#
+ FILLER_0_176/li_0_797# FILLER_0_200/li_641_797# FILLER_0_24/li_353_797# mprj2_logic_high_lv/li_179_79#
+ FILLER_0_168/li_545_797# FILLER_1_252/li_65_797# FILLER_2_179/li_641_n17# mprj_logic_high_lv/li_65_1611#
+ FILLER_1_140/li_65_797# FILLER_0_256/li_0_n17# FILLER_2_8/li_449_n17# FILLER_1_172/li_161_n17#
+ FILLER_2_0/li_65_797# FILLER_2_259/li_353_797# FILLER_1_180/li_65_797# FILLER_0_80/li_0_n17#
+ FILLER_2_0/li_641_n17# FILLER_0_256/li_115_72# FILLER_1_32/li_353_n17# FILLER_1_8/li_353_n17#
+ FILLER_2_115/li_100_536# FILLER_2_115/li_449_797# FILLER_2_32/li_65_797# FILLER_2_163/li_0_797#
+ FILLER_2_0/li_161_797# FILLER_0_112/li_65_n17# FILLER_2_107/li_257_n17# FILLER_1_180/li_115_72#
+ mprj2_logic_high_hvl/li_353_797# FILLER_0_32/li_545_797# FILLER_0_104/li_65_n17#
+ FILLER_0_184/li_0_797# mprj_logic_high_lv/li_1409_1611# FILLER_2_211/li_115_72#
+ FILLER_2_211/li_0_n17# FILLER_2_16/li_545_n17# FILLER_1_220/li_257_n17# FILLER_1_260/li_545_n17#
+ FILLER_1_244/li_0_797# FILLER_0_184/li_0_n17# FILLER_1_204/li_257_n17# FILLER_2_227/li_257_797#
+ FILLER_1_252/li_65_n17# FILLER_1_140/li_65_n17# FILLER_2_267/li_545_797# FILLER_2_187/li_353_797#
+ mprj2_logic_high_lv/li_0_797# FILLER_0_248/li_257_797# FILLER_1_228/li_545_n17#
+ mprj_logic_high_lv/li_353_1611# FILLER_2_259/li_353_n17# FILLER_2_0/li_65_n17# FILLER_0_200/li_161_797#
+ FILLER_1_188/li_641_n17# FILLER_2_179/li_161_n17# FILLER_2_187/li_65_n17# FILLER_1_204/li_115_72#
+ FILLER_1_115/li_737_n17# FILLER_2_115/li_449_n17# FILLER_2_163/li_0_n17# FILLER_2_32/li_65_n17#
+ FILLER_2_300/li_161_797# FILLER_2_0/li_161_n17# FILLER_1_107/li_0_n17# FILLER_2_235/li_100_536#
+ FILLER_1_48/li_353_797# mprj2_logic_high_hvl/li_353_n17# FILLER_2_235/li_449_797#
+ FILLER_1_172/li_0_797# FILLER_2_155/li_257_797# FILLER_2_24/li_257_797# FILLER_0_256/li_100_536#
+ FILLER_2_227/li_257_n17# FILLER_2_195/li_545_797# FILLER_0_256/li_449_797# FILLER_1_244/li_0_n17#
+ FILLER_1_156/li_545_n17# FILLER_2_267/li_545_n17# FILLER_0_176/li_257_797# FILLER_2_187/li_353_n17#
+ FILLER_0_96/li_0_n17# FILLER_0_264/li_65_797# FILLER_1_24/li_0_n17# FILLER_0_216/li_641_797#
+ mprj2_logic_high_lv/li_1121_1611# FILLER_0_272/li_0_n17# FILLER_1_188/li_161_n17#
+ FILLER_2_300/li_161_n17# FILLER_2_163/li_100_536# FILLER_2_32/li_100_536# FILLER_2_163/li_449_797#
+ FILLER_2_32/li_449_797# FILLER_1_48/li_353_n17# FILLER_1_115/li_257_n17# FILLER_0_184/li_100_536#
+ FILLER_0_192/li_115_72# FILLER_2_235/li_449_n17# FILLER_2_155/li_257_n17# FILLER_0_8/li_0_797#
+ FILLER_1_172/li_0_n17# FILLER_0_184/li_449_797# FILLER_2_195/li_545_n17# FILLER_2_24/li_257_n17#
+ FILLER_0_80/li_545_797# FILLER_1_260/li_65_n17# FILLER_1_244/li_100_536# FILLER_0_104/li_353_797#
+ FILLER_1_236/li_257_n17# FILLER_1_24/li_100_536# FILLER_1_16/li_65_n17# FILLER_0_200/li_0_n17#
+ FILLER_0_88/li_65_797# FILLER_1_131/li_50_537# FILLER_0_216/li_115_72# FILLER_1_16/li_257_n17#
+ FILLER_0_104/li_115_72# FILLER_1_8/li_65_n17# FILLER_2_163/li_449_n17# FILLER_0_216/li_161_797#
+ FILLER_2_32/li_449_n17# FILLER_1_252/li_115_72# FILLER_1_140/li_115_72# FILLER_0_16/li_100_536#
+ FILLER_1_172/li_100_536# FILLER_0_16/li_449_797# FILLER_2_0/li_115_72# FILLER_0_112/li_545_797#
+ FILLER_2_187/li_115_72# FILLER_0_248/li_65_n17# FILLER_1_164/li_257_n17# FILLER_1_212/li_65_n17#
+ FILLER_0_0/li_257_797# FILLER_1_24/li_449_n17# FILLER_2_203/li_353_797# FILLER_2_32/li_115_72#
+ FILLER_2_259/li_65_n17# FILLER_2_243/li_641_797# FILLER_1_204/li_641_n17# FILLER_0_224/li_353_797#
+ FILLER_0_8/li_545_797# FILLER_0_88/li_353_797# FILLER_0_264/li_641_797# FILLER_0_176/li_65_n17#
+ FILLER_1_62/li_737_797# FILLER_2_179/li_100_536# FILLER_2_179/li_449_797# mprj_logic_high_lv/li_257_1611#
+ FILLER_2_211/li_545_797# mprj_logic_high_lv/li_0_1611# FILLER_2_171/li_641_797#
+ FILLER_1_212/li_0_n17# FILLER_2_203/li_353_n17# FILLER_0_232/li_545_797# FILLER_0_224/li_65_797#
+ FILLER_0_96/li_545_797# FILLER_0_112/li_65_797# FILLER_2_243/li_641_n17# FILLER_2_0/li_100_536#
+ FILLER_0_256/li_0_797# FILLER_0_192/li_641_797# FILLER_2_0/li_449_797# mprj_logic_high_hvl/li_257_797#
+ FILLER_0_16/li_0_797# mprj_logic_high_lv/li_641_1611# FILLER_2_259/li_0_797# FILLER_1_244/li_65_797#
+ mprj2_logic_high_lv/li_65_797# FILLER_0_264/li_161_797# FILLER_1_196/li_0_797# FILLER_0_264/li_115_72#
+ FILLER_1_62/li_737_n17# FILLER_0_200/li_100_536# FILLER_0_200/li_449_797# FILLER_1_16/li_115_72#
+ FILLER_2_211/li_545_n17# FILLER_2_179/li_449_n17# FILLER_0_248/li_0_797# FILLER_0_160/li_545_797#
+ FILLER_2_171/li_641_n17# FILLER_2_107/li_545_797# FILLER_1_62/li_257_797# FILLER_1_188/li_100_536#
+ FILLER_0_96/li_545_n17# FILLER_1_131/li_161_797# mprj2_logic_high_lv/li_1601_797#
+ FILLER_2_0/li_449_n17# FILLER_1_8/li_115_72# FILLER_1_140/li_353_797# mprj2_logic_high_lv/li_1025_1611#
+ FILLER_0_24/li_641_797# mprj_logic_high_hvl/li_257_n17# mprj_logic_high_lv/li_384_1039#
+ FILLER_1_220/li_0_797# FILLER_1_172/li_65_797# FILLER_0_216/li_0_n17# FILLER_2_107/li_65_797#
+ FILLER_1_252/li_641_n17# FILLER_2_243/li_161_n17# FILLER_0_272/li_353_797# FILLER_1_0/li_353_n17#
+ FILLER_0_192/li_161_797# FILLER_2_219/li_353_797# FILLER_2_259/li_641_797# FILLER_2_195/li_65_n17#
+ FILLER_1_32/li_641_n17# FILLER_2_251/li_257_797# FILLER_1_212/li_115_72# FILLER_1_8/li_641_n17#
+ FILLER_2_8/li_257_797# FILLER_1_204/li_65_n17# FILLER_2_115/li_737_797# mprj2_logic_high_lv/li_929_1611#
+ FILLER_1_131/li_0_797# FILLER_0_88/li_115_72# FILLER_2_259/li_115_72# FILLER_2_107/li_545_n17#
+ FILLER_1_62/li_257_n17# FILLER_0_192/li_65_n17# FILLER_0_240/li_257_797# FILLER_1_220/li_545_n17#
+ mprj2_logic_high_lv/li_826_79# FILLER_1_131/li_161_n17# FILLER_1_140/li_353_n17#
+ FILLER_1_188/li_65_n17# FILLER_2_251/li_353_n17# FILLER_1_180/li_641_n17# FILLER_2_227/li_545_797#
+ FILLER_2_219/li_65_n17# FILLER_2_171/li_161_n17# FILLER_2_107/li_65_n17# FILLER_2_16/li_353_797#
+ FILLER_0_208/li_257_797# FILLER_2_187/li_641_797# FILLER_1_131/li_353_797# FILLER_0_272/li_65_797#
+ FILLER_0_248/li_545_797# FILLER_2_219/li_353_n17# FILLER_0_24/li_161_797# FILLER_0_160/li_65_797#
+ FILLER_0_168/li_353_797# FILLER_2_259/li_641_n17# FILLER_1_252/li_161_n17# mprj_logic_high_lv/li_506_1123#
+ FILLER_2_8/li_257_n17#
XFILLER_2_187 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_24 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_264 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_155 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_232 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_0 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_200 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_180 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_179 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_16 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_256 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_115 vssd vssd FILLER_2_115/VPB FILLER_2_115/VPB sky130_fd_sc_hvl__decap_8
XFILLER_0_224 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_62 vssa2 vssa2 vdda2 vdda2 sky130_fd_sc_hvl__decap_8
Xmprj2_logic_high_hvl vssa2 vssa2 vdda2 vdda2 mprj2_logic_high_lv/A mprj2_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
XFILLER_1_172 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_248 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_216 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_140 vssa1 vssa1 vdda1 vdda1 sky130_fd_sc_hvl__decap_8
XFILLER_2_107 vssd vssd FILLER_2_115/VPB FILLER_2_115/VPB sky130_fd_sc_hvl__decap_8
XFILLER_1_300 vssd vssd vdda1 vdda1 sky130_fd_sc_hvl__fill_2
XFILLER_1_196 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_32 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_164 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_131 vssa1 vssa1 vdda1 vdda1 sky130_fd_sc_hvl__decap_4
XFILLER_1_8 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_208 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_56 vssa2 vssa2 vdda2 vdda2 sky130_fd_sc_hvl__fill_1
XFILLER_1_188 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_156 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
Xmprj_logic_high_hvl vssa1 vssa1 vdda1 vdda1 mprj_logic_high_lv/A mprj_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
XFILLER_1_24 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_251 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_48 vssa2 vssa2 vdda2 vdda2 sky130_fd_sc_hvl__decap_8
XFILLER_1_16 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_243 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_192 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_115 vssd vssd FILLER_2_115/VPB FILLER_2_115/VPB sky130_fd_sc_hvl__decap_8
XFILLER_2_211 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_160 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_267 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_0 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_235 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_184 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_107 vssd vssd FILLER_2_115/VPB FILLER_2_115/VPB sky130_fd_sc_hvl__decap_8
XFILLER_2_203 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_259 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_32 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_0 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_260 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_227 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_176 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_112 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_219 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_168 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_24 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_252 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_220 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_80 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_104 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_8 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_16 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_244 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_212 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_8 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_268 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_171 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_96 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_236 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_1_204 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_195 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_32 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_300 vssd vssd vdda1 vdda1 sky130_fd_sc_hvl__fill_2
Xmprj_logic_high_lv mprj_logic_high_lv/A vccd vssd vssd vdda1 vdda1 mprj_vdd_logic1
+ sky130_fd_sc_hvl__lsbufhv2lv_1
XFILLER_1_228 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_2_163 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_88 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_272 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
XFILLER_0_240 vssd vssd vccd vccd sky130_fd_sc_hvl__decap_8
Xmprj2_logic_high_lv mprj2_logic_high_lv/A vccd vssd vssd vdda2 vdda2 mprj2_vdd_logic1
+ sky130_fd_sc_hvl__lsbufhv2lv_1
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_oen_core[0] la_oen_core[100] la_oen_core[101] la_oen_core[102]
+ la_oen_core[103] la_oen_core[104] la_oen_core[105] la_oen_core[106] la_oen_core[107]
+ la_oen_core[108] la_oen_core[109] la_oen_core[10] la_oen_core[110] la_oen_core[111]
+ la_oen_core[112] la_oen_core[113] la_oen_core[114] la_oen_core[115] la_oen_core[116]
+ la_oen_core[117] la_oen_core[118] la_oen_core[119] la_oen_core[11] la_oen_core[120]
+ la_oen_core[121] la_oen_core[122] la_oen_core[123] la_oen_core[124] la_oen_core[125]
+ la_oen_core[126] la_oen_core[127] la_oen_core[12] la_oen_core[13] la_oen_core[14]
+ la_oen_core[15] la_oen_core[16] la_oen_core[17] la_oen_core[18] la_oen_core[19]
+ la_oen_core[1] la_oen_core[20] la_oen_core[21] la_oen_core[22] la_oen_core[23] la_oen_core[24]
+ la_oen_core[25] la_oen_core[26] la_oen_core[27] la_oen_core[28] la_oen_core[29]
+ la_oen_core[2] la_oen_core[30] la_oen_core[31] la_oen_core[32] la_oen_core[33] la_oen_core[34]
+ la_oen_core[35] la_oen_core[36] la_oen_core[37] la_oen_core[38] la_oen_core[39]
+ la_oen_core[3] la_oen_core[40] la_oen_core[41] la_oen_core[42] la_oen_core[43] la_oen_core[44]
+ la_oen_core[45] la_oen_core[46] la_oen_core[47] la_oen_core[48] la_oen_core[49]
+ la_oen_core[4] la_oen_core[50] la_oen_core[51] la_oen_core[52] la_oen_core[53] la_oen_core[54]
+ la_oen_core[55] la_oen_core[56] la_oen_core[57] la_oen_core[58] la_oen_core[59]
+ la_oen_core[5] la_oen_core[60] la_oen_core[61] la_oen_core[62] la_oen_core[63] la_oen_core[64]
+ la_oen_core[65] la_oen_core[66] la_oen_core[67] la_oen_core[68] la_oen_core[69]
+ la_oen_core[6] la_oen_core[70] la_oen_core[71] la_oen_core[72] la_oen_core[73] la_oen_core[74]
+ la_oen_core[75] la_oen_core[76] la_oen_core[77] la_oen_core[78] la_oen_core[79]
+ la_oen_core[7] la_oen_core[80] la_oen_core[81] la_oen_core[82] la_oen_core[83] la_oen_core[84]
+ la_oen_core[85] la_oen_core[86] la_oen_core[87] la_oen_core[88] la_oen_core[89]
+ la_oen_core[8] la_oen_core[90] la_oen_core[91] la_oen_core[92] la_oen_core[93] la_oen_core[94]
+ la_oen_core[95] la_oen_core[96] la_oen_core[97] la_oen_core[98] la_oen_core[99]
+ la_oen_core[9] la_oen_mprj[0] la_oen_mprj[100] la_oen_mprj[101] la_oen_mprj[102]
+ la_oen_mprj[103] la_oen_mprj[104] la_oen_mprj[105] la_oen_mprj[106] la_oen_mprj[107]
+ la_oen_mprj[108] la_oen_mprj[109] la_oen_mprj[10] la_oen_mprj[110] la_oen_mprj[111]
+ la_oen_mprj[112] la_oen_mprj[113] la_oen_mprj[114] la_oen_mprj[115] la_oen_mprj[116]
+ la_oen_mprj[117] la_oen_mprj[118] la_oen_mprj[119] la_oen_mprj[11] la_oen_mprj[120]
+ la_oen_mprj[121] la_oen_mprj[122] la_oen_mprj[123] la_oen_mprj[124] la_oen_mprj[125]
+ la_oen_mprj[126] la_oen_mprj[127] la_oen_mprj[12] la_oen_mprj[13] la_oen_mprj[14]
+ la_oen_mprj[15] la_oen_mprj[16] la_oen_mprj[17] la_oen_mprj[18] la_oen_mprj[19]
+ la_oen_mprj[1] la_oen_mprj[20] la_oen_mprj[21] la_oen_mprj[22] la_oen_mprj[23] la_oen_mprj[24]
+ la_oen_mprj[25] la_oen_mprj[26] la_oen_mprj[27] la_oen_mprj[28] la_oen_mprj[29]
+ la_oen_mprj[2] la_oen_mprj[30] la_oen_mprj[31] la_oen_mprj[32] la_oen_mprj[33] la_oen_mprj[34]
+ la_oen_mprj[35] la_oen_mprj[36] la_oen_mprj[37] la_oen_mprj[38] la_oen_mprj[39]
+ la_oen_mprj[3] la_oen_mprj[40] la_oen_mprj[41] la_oen_mprj[42] la_oen_mprj[43] la_oen_mprj[44]
+ la_oen_mprj[45] la_oen_mprj[46] la_oen_mprj[47] la_oen_mprj[48] la_oen_mprj[49]
+ la_oen_mprj[4] la_oen_mprj[50] la_oen_mprj[51] la_oen_mprj[52] la_oen_mprj[53] la_oen_mprj[54]
+ la_oen_mprj[55] la_oen_mprj[56] la_oen_mprj[57] la_oen_mprj[58] la_oen_mprj[59]
+ la_oen_mprj[5] la_oen_mprj[60] la_oen_mprj[61] la_oen_mprj[62] la_oen_mprj[63] la_oen_mprj[64]
+ la_oen_mprj[65] la_oen_mprj[66] la_oen_mprj[67] la_oen_mprj[68] la_oen_mprj[69]
+ la_oen_mprj[6] la_oen_mprj[70] la_oen_mprj[71] la_oen_mprj[72] la_oen_mprj[73] la_oen_mprj[74]
+ la_oen_mprj[75] la_oen_mprj[76] la_oen_mprj[77] la_oen_mprj[78] la_oen_mprj[79]
+ la_oen_mprj[7] la_oen_mprj[80] la_oen_mprj[81] la_oen_mprj[82] la_oen_mprj[83] la_oen_mprj[84]
+ la_oen_mprj[85] la_oen_mprj[86] la_oen_mprj[87] la_oen_mprj[88] la_oen_mprj[89]
+ la_oen_mprj[8] la_oen_mprj[90] la_oen_mprj[91] la_oen_mprj[92] la_oen_mprj[93] la_oen_mprj[94]
+ la_oen_mprj[95] la_oen_mprj[96] la_oen_mprj[97] la_oen_mprj[98] la_oen_mprj[99]
+ la_oen_mprj[9] mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12]
+ mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16]
+ mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20]
+ mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24]
+ mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28]
+ mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3]
+ mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8]
+ mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12]
+ mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16]
+ mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20]
+ mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24]
+ mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28]
+ mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3]
+ mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8]
+ mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_o_core[0] mprj_dat_o_core[10]
+ mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14]
+ mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18]
+ mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22]
+ mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26]
+ mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30]
+ mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6]
+ mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10]
+ mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14]
+ mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18]
+ mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22]
+ mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26]
+ mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30]
+ mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6]
+ mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_sel_o_core[0] mprj_sel_o_core[1]
+ mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2]
+ mprj_sel_o_user[3] mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user
+ user1_vcc_powergood user1_vdd_powergood user2_vcc_powergood user2_vdd_powergood
+ user_clock user_clock2 user_reset user_resetn vccd vssd vccd1 vssd1 vccd2 vssd2
+ vdda1 vdda2 FILLER_21_1889/li_0_527# la_buf\[99\]/li_17_51# powergood_check/FILLER_0_112/li_737_797#
+ user_to_mprj_in_gates\[124\]/li_339_n17# PHY_225/li_0_527# FILLER_25_774/li_0_n17#
+ FILLER_27_806/li_155_n17# la_buf\[82\]/li_779_17# PHY_418/li_0_527# user_to_mprj_oen_buffers\[74\]/li_611_17#
+ _470_/li_247_527# la_buf\[95\]/li_1259_527# FILLER_13_1680/li_0_527# user_to_mprj_oen_buffers\[74\]/li_707_n17#
+ PHY_676/li_0_527# user_to_mprj_oen_buffers\[46\]/li_1351_527# PHY_791/li_0_n17#
+ _333_/li_0_n17# user_to_mprj_in_gates\[98\]/li_431_n17# user_to_mprj_in_gates\[54\]/li_18_51#
+ PHY_819/li_0_n17# PHY_692/li_0_527# FILLER_26_1054/li_63_527# FILLER_12_1923/li_155_527#
+ FILLER_11_1627/li_63_n17# user_to_mprj_oen_buffers\[56\]/li_431_n17# user_to_mprj_in_gates\[105\]/li_615_n17#
+ PHY_350/li_0_n17# _614_/li_0_n17# la_buf\[12\]/li_611_17# FILLER_21_1436/li_0_n17#
+ la_buf\[81\]/li_63_527# FILLER_21_471/li_0_527# _546_/li_155_527# la_buf\[15\]/li_0_527#
+ _627_/li_0_n17# _522_/li_0_527# ANTENNA_user_to_mprj_in_gates\[124\]_A/li_63_n17#
+ PHY_797/li_0_n17# FILLER_7_984/li_63_527# _637_/li_0_n17# PHY_772/li_0_n17# user_to_mprj_in_gates\[51\]/li_339_n17#
+ PHY_381/li_0_n17# user_to_mprj_oen_buffers\[10\]/li_207_51# PHY_499/li_0_527# powergood_check/FILLER_1_220/li_115_72#
+ _605_/li_0_527# PHY_321/li_0_n17# la_buf\[24\]/li_891_527# la_buf\[9\]/li_779_17#
+ powergood_check/FILLER_0_168/li_65_n17# mprj_adr_buf\[25\]/li_215_311# PHY_87/li_0_n17#
+ PHY_340/li_0_n17# FILLER_24_1494/li_63_n17# user_to_mprj_in_gates\[88\]/li_63_n17#
+ la_buf\[58\]/li_707_n17# user_to_mprj_in_gates\[77\]/li_431_527# FILLER_11_447/li_0_n17#
+ powergood_check/FILLER_0_24/li_100_536# user_to_mprj_oen_buffers\[36\]/li_17_51#
+ la_buf\[107\]/li_0_527# PHY_652/li_0_n17# _337_/li_155_n17# user_to_mprj_in_gates\[112\]/li_339_n17#
+ user_to_mprj_in_gates\[25\]/li_707_367# _636_/li_0_n17# PHY_820/li_0_n17# user_to_mprj_in_buffers\[45\]/li_51_367#
+ PHY_821/li_0_527# la_buf\[48\]/li_17_51# powergood_check/FILLER_0_96/li_115_72#
+ la_buf\[98\]/li_1259_n17# FILLER_17_231/li_0_527# _641_/li_0_n17# user_to_mprj_in_gates\[30\]/li_339_527#
+ user_to_mprj_oen_buffers\[62\]/li_707_n17# user_to_mprj_in_gates\[33\]/li_523_n17#
+ mprj_dat_buf\[6\]/li_207_51# FILLER_11_996/li_0_n17# FILLER_11_792/li_0_n17# user_to_mprj_in_gates\[86\]/li_431_n17#
+ PHY_269/li_0_527# la_buf\[49\]/li_247_n17# powergood_check/FILLER_0_24/li_449_797#
+ user_to_mprj_in_gates\[90\]/li_63_n17# FILLER_24_1494/li_0_n17# FILLER_11_1004/li_0_527#
+ user_to_mprj_oen_buffers\[44\]/li_431_n17# PHY_721/li_0_n17# _579_/li_0_n17# PHY_600/li_0_n17#
+ user_to_mprj_in_gates\[104\]/li_523_n17# powergood_check/FILLER_2_195/li_257_n17#
+ PHY_413/li_0_527# PHY_289/li_0_527# _463_/li_0_527# PHY_57/li_0_527# user_to_mprj_oen_buffers\[76\]/li_207_51#
+ FILLER_7_921/li_63_527# user_to_mprj_oen_buffers\[42\]/li_431_527# PHY_41/li_0_n17#
+ _454_/li_0_527# FILLER_16_1589/li_63_n17# PHY_707/li_0_527# la_buf\[6\]/li_1535_527#
+ mprj_adr_buf\[2\]/li_1351_527# _464_/li_0_n17# ANTENNA__430__A/li_0_527# mprj_adr_buf\[13\]/li_215_311#
+ PHY_338/li_0_527# la_buf\[106\]/li_1259_n17# PHY_48/li_0_527# mprj_dat_buf\[27\]/li_1167_527#
+ la_buf\[28\]/li_247_527# _348_/li_0_527# PHY_538/li_0_n17# _430_/li_0_n17# user_to_mprj_oen_buffers\[57\]/li_779_17#
+ FILLER_23_1814/li_63_n17# _610_/li_0_527# _538_/li_0_n17# la_buf\[83\]/li_63_527#
+ _475_/li_0_n17# user_to_mprj_in_gates\[100\]/li_339_n17# user_to_mprj_in_gates\[13\]/li_707_367#
+ user_to_mprj_in_gates\[92\]/li_707_n17# PHY_97/li_0_527# PHY_356/li_0_n17# PHY_344/li_0_n17#
+ FILLER_13_1635/li_0_n17# user_to_mprj_in_buffers\[8\]/li_523_n17# _402_/li_0_n17#
+ PHY_600/li_0_527# FILLER_23_1429/li_63_n17# PHY_55/li_0_n17# la_buf\[41\]/li_0_527#
+ PHY_248/li_0_n17# PHY_224/li_0_n17# la_buf\[26\]/li_1075_n17# la_buf\[38\]/li_207_51#
+ powergood_check/FILLER_2_203/li_545_797# user_to_mprj_oen_buffers\[22\]/li_795_379#
+ la_buf\[37\]/li_247_n17# user_to_mprj_in_gates\[74\]/li_431_n17# _477_/li_0_n17#
+ la_buf\[97\]/li_1167_n17# PHY_752/li_0_527# FILLER_13_895/li_63_527# FILLER_25_1768/li_0_n17#
+ user_to_mprj_in_gates\[72\]/li_155_527# PHY_37/li_0_n17# la_buf\[101\]/li_207_51#
+ PHY_443/li_0_n17# ANTENNA__514__A/li_63_n17# user_to_mprj_oen_buffers\[20\]/li_891_n17#
+ PHY_57/li_0_n17# _607_/li_0_527# PHY_62/li_0_527# powergood_check/FILLER_2_267/li_115_72#
+ _483_/li_247_527# user_to_mprj_in_buffers\[127\]/li_404_367# la_buf\[24\]/li_63_n17#
+ _608_/li_0_527# la_buf\[47\]/li_63_527# PHY_664/li_0_527# powergood_check/FILLER_2_8/li_0_n17#
+ FILLER_9_171/li_155_n17# mprj_dat_buf\[14\]/li_523_n17# powergood_check/FILLER_1_62/li_545_797#
+ powergood_check/FILLER_2_155/li_115_72# la_buf\[40\]/li_207_51# PHY_392/li_0_527#
+ user_to_mprj_oen_buffers\[91\]/li_63_n17# mprj_sel_buf\[1\]/li_779_17# _596_/li_247_n17#
+ _494_/li_155_527# powergood_check/FILLER_2_163/li_641_797# FILLER_12_685/li_0_527#
+ _489_/li_0_n17# _432_/li_0_n17# _465_/li_0_n17# PHY_782/li_0_527# la_buf\[114\]/li_63_n17#
+ powergood_check/FILLER_0_224/li_545_797# la_buf\[95\]/li_215_311# user_to_mprj_in_buffers\[69\]/li_339_n17#
+ FILLER_21_1720/li_0_n17# FILLER_23_1413/li_0_527# FILLER_19_530/li_0_n17# FILLER_10_1174/li_63_n17#
+ powergood_check/FILLER_1_8/li_449_n17# FILLER_9_1142/li_0_n17# FILLER_25_1096/li_0_n17#
+ user_to_mprj_oen_buffers\[50\]/li_1535_527# FILLER_16_88/li_0_n17# PHY_53/li_0_527#
+ PHY_394/li_0_527# mprj_adr_buf\[27\]/li_17_51# FILLER_12_890/li_0_527# _510_/li_0_527#
+ FILLER_28_1726/li_63_n17# FILLER_18_40/li_0_527# user_to_mprj_oen_buffers\[20\]/li_431_n17#
+ user_to_mprj_in_gates\[98\]/li_247_527# _607_/li_247_527# _584_/li_155_n17# mprj_adr_buf\[28\]/li_795_379#
+ PHY_691/li_0_527# la_buf\[109\]/li_247_n17# FILLER_18_1899/li_155_527# _648_/li_0_527#
+ user_to_mprj_in_buffers\[115\]/li_404_367# powergood_check/FILLER_2_115/li_161_n17#
+ FILLER_25_974/li_0_n17# user_to_mprj_in_gates\[106\]/li_18_51# user_to_mprj_in_buffers\[49\]/li_339_527#
+ user_to_mprj_in_gates\[123\]/li_431_n17# user_to_mprj_in_buffers\[72\]/li_236_17#
+ PHY_750/li_0_527# PHY_225/li_0_n17# powergood_check/FILLER_2_235/li_641_n17# PHY_900/li_0_527#
+ FILLER_8_1850/li_63_527# user_to_mprj_in_gates\[121\]/li_615_527# la_buf\[79\]/li_707_527#
+ FILLER_23_1510/li_0_527# powergood_check/FILLER_0_184/li_641_797# PHY_23/li_0_n17#
+ FILLER_16_293/li_0_527# _623_/li_247_527# FILLER_14_1986/li_63_527# powergood_check/FILLER_1_32/li_449_n17#
+ powergood_check/FILLER_1_196/li_65_n17# _374_/li_155_527# mprj_dat_buf\[5\]/li_17_51#
+ user_to_mprj_in_gates\[35\]/li_0_n17# FILLER_9_367/li_63_n17# user_to_mprj_in_buffers\[49\]/li_404_17#
+ FILLER_19_48/li_155_527# user_to_mprj_oen_buffers\[105\]/li_247_527# PHY_687/li_0_527#
+ PHY_496/li_0_527# PHY_809/li_0_527# PHY_42/li_0_527# _468_/li_0_527# FILLER_25_1176/li_63_n17#
+ la_buf\[59\]/li_1167_n17# PHY_395/li_0_n17# la_buf\[83\]/li_215_311# PHY_7/li_0_527#
+ FILLER_13_1048/li_63_527# FILLER_25_934/li_155_n17# la_buf\[57\]/li_615_527# powergood_check/FILLER_1_0/li_641_n17#
+ FILLER_13_1199/li_63_527# user_to_mprj_in_gates\[50\]/li_431_n17# PHY_157/li_0_n17#
+ _345_/li_0_527# FILLER_7_984/li_155_527# la_buf\[27\]/li_891_n17# mprj_adr_buf\[10\]/li_611_17#
+ FILLER_13_1199/li_0_527# FILLER_0_58/li_0_527# PHY_701/li_0_n17# user_to_mprj_oen_buffers\[92\]/li_891_527#
+ user_to_mprj_in_buffers\[103\]/li_404_367# powergood_check/FILLER_2_0/li_257_797#
+ user_to_mprj_oen_buffers\[15\]/li_207_51# powergood_check/FILLER_1_260/li_257_n17#
+ FILLER_17_1570/li_0_n17# FILLER_24_1648/li_63_527# mprj_adr_buf\[26\]/li_431_n17#
+ _334_/li_247_n17# PHY_703/li_0_n17# user_to_mprj_in_gates\[111\]/li_431_n17# user_to_mprj_in_gates\[79\]/li_247_527#
+ FILLER_15_1688/li_0_n17# FILLER_12_748/li_155_527# user_to_mprj_oen_buffers\[49\]/li_891_527#
+ powergood_check/FILLER_2_227/li_65_n17# user_to_mprj_oen_buffers\[86\]/li_17_51#
+ mprj_stb_buf/li_1075_n17# la_buf\[47\]/li_0_n17# _425_/li_0_527# user_to_mprj_in_gates\[14\]/li_247_527#
+ FILLER_12_1035/li_63_n17# la_buf\[67\]/li_63_n17# _450_/li_0_n17# _626_/li_0_527#
+ la_buf\[98\]/li_17_51# FILLER_12_1186/li_63_n17# _553_/li_155_527# powergood_check/FILLER_2_115/li_65_n17#
+ FILLER_15_59/li_0_527# PHY_178/li_0_n17# FILLER_22_387/li_0_527# PHY_182/li_0_527#
+ ANTENNA__332__A/li_0_n17# _504_/li_0_n17# FILLER_25_638/li_63_n17# la_buf\[71\]/li_215_311#
+ FILLER_11_798/li_63_n17# FILLER_25_1648/li_63_527# PHY_550/li_0_n17# user_to_mprj_in_gates\[88\]/li_247_n17#
+ PHY_820/li_0_527# powergood_check/FILLER_0_96/li_353_797# la_buf\[44\]/li_1075_527#
+ PHY_718/li_0_n17# la_buf\[45\]/li_615_527# FILLER_0_1346/li_0_527# _422_/li_0_527#
+ user_to_mprj_in_gates\[95\]/li_63_n17# FILLER_21_1405/li_0_n17# PHY_352/li_0_n17#
+ PHY_524/li_0_n17# mprj_dat_buf\[11\]/li_891_n17# mprj_dat_buf\[17\]/li_1351_527#
+ _633_/li_0_n17# user_to_mprj_in_gates\[53\]/li_18_51# mprj_dat_buf\[26\]/li_215_311#
+ FILLER_21_66/li_63_n17# FILLER_16_459/li_63_n17# PHY_864/li_0_527# ANTENNA_user_to_mprj_in_gates\[32\]_A/li_63_527#
+ _344_/li_155_n17# FILLER_16_1927/li_0_n17# powergood_check/FILLER_2_0/li_65_n17#
+ _643_/li_155_n17# mprj_adr_buf\[2\]/li_247_n17# user_to_mprj_oen_buffers\[80\]/li_891_527#
+ PHY_233/li_0_n17# user_to_mprj_oen_buffers\[114\]/li_63_527# user_to_mprj_in_gates\[57\]/li_0_n17#
+ PHY_810/li_0_527# powergood_check/FILLER_1_236/li_65_797# user_to_mprj_in_gates\[69\]/li_523_n17#
+ FILLER_5_617/li_155_527# PHY_676/li_0_n17# powergood_check/FILLER_1_140/li_0_n17#
+ FILLER_12_617/li_0_n17# FILLER_24_1425/li_155_527# PHY_851/li_0_n17# user_to_mprj_oen_buffers\[25\]/li_247_527#
+ user_to_mprj_in_gates\[1\]/li_155_527# la_buf\[120\]/li_0_527# _439_/li_0_n17# FILLER_11_196/li_63_527#
+ FILLER_22_1408/li_0_n17# mprj_adr_buf\[29\]/li_1535_527# la_buf\[98\]/li_795_379#
+ PHY_287/li_0_527# mprj_adr_buf\[12\]/li_207_51# la_buf\[88\]/li_63_527# PHY_896/li_0_n17#
+ user_to_mprj_oen_buffers\[35\]/li_17_51# user_to_mprj_oen_buffers\[8\]/li_1351_527#
+ la_buf\[31\]/li_0_527# PHY_835/li_0_527# _470_/li_0_527# user_to_mprj_oen_buffers\[83\]/li_207_51#
+ user_to_mprj_in_gates\[117\]/li_247_527# PHY_704/li_0_527# user_to_mprj_in_gates\[89\]/li_247_527#
+ PHY_437/li_0_n17# la_buf\[47\]/li_17_51# FILLER_14_1793/li_63_527# PHY_81/li_0_527#
+ FILLER_15_357/li_0_n17# FILLER_16_1601/li_0_527# FILLER_12_978/li_155_n17# _463_/li_247_527#
+ FILLER_23_607/li_0_527# la_buf\[106\]/li_207_51# _346_/li_247_n17# PHY_56/li_0_n17#
+ PHY_816/li_0_n17# PHY_309/li_0_n17# FILLER_9_1234/li_155_527# FILLER_21_1570/li_63_n17#
+ mprj_dat_buf\[14\]/li_215_311# FILLER_12_1552/li_63_n17# FILLER_5_954/li_155_527#
+ la_buf\[18\]/li_215_311# FILLER_26_1247/li_155_527# _559_/li_247_n17# FILLER_11_1606/li_63_n17#
+ PHY_890/li_0_527# FILLER_9_1158/li_0_n17# la_buf\[87\]/li_63_527# _569_/li_0_n17#
+ powergood_check/FILLER_0_256/li_161_797# powergood_check/FILLER_2_8/li_545_797#
+ FILLER_16_1502/li_0_527# _536_/li_0_n17# PHY_502/li_0_527# FILLER_22_2044/li_0_n17#
+ PHY_704/li_0_n17# user_to_mprj_in_gates\[57\]/li_523_n17# user_to_mprj_oen_buffers\[119\]/li_215_311#
+ mprj_dat_buf\[12\]/li_1351_n17# PHY_386/li_0_n17# PHY_352/li_0_527# FILLER_19_1634/li_155_n17#
+ la_buf\[45\]/li_207_51# FILLER_13_733/li_63_527# PHY_505/li_0_527# mprj_dat_buf\[6\]/li_707_527#
+ user_to_mprj_in_buffers\[11\]/li_236_17# user_to_mprj_in_gates\[116\]/li_339_527#
+ PHY_48/li_0_n17# la_buf\[79\]/li_1351_527# la_buf\[86\]/li_795_379# la_buf\[54\]/li_983_527#
+ _345_/li_0_n17# FILLER_7_1035/li_155_527# user_to_mprj_oen_buffers\[90\]/li_1351_n17#
+ user_to_mprj_in_gates\[118\]/li_523_n17# FILLER_9_1099/li_63_527# _612_/li_0_527#
+ user_to_mprj_oen_buffers\[92\]/li_215_311# PHY_364/li_0_n17# user_to_mprj_in_gates\[64\]/li_247_n17#
+ _438_/li_0_527# la_buf\[21\]/li_615_527# FILLER_11_1097/li_0_n17# PHY_743/li_0_n17#
+ _589_/li_155_n17# FILLER_11_716/li_63_n17# PHY_342/li_0_n17# PHY_405/li_0_527# FILLER_11_827/li_63_n17#
+ FILLER_12_593/li_0_527# _612_/li_0_n17# PHY_921/li_0_n17# user_to_mprj_oen_buffers\[85\]/li_1259_n17#
+ FILLER_18_1416/li_63_527# powergood_check/FILLER_2_219/li_0_797# PHY_921/li_0_527#
+ user_to_mprj_in_gates\[125\]/li_247_n17# PHY_477/li_0_n17# PHY_292/li_0_n17# user_to_mprj_in_gates\[45\]/li_523_n17#
+ user_to_mprj_oen_buffers\[91\]/li_1351_527# FILLER_11_838/li_0_n17# PHY_49/li_0_527#
+ user_to_mprj_oen_buffers\[107\]/li_215_311# user_to_mprj_oen_buffers\[20\]/li_611_17#
+ FILLER_14_1808/li_0_527# PHY_742/li_0_527# PHY_63/li_0_527# la_buf\[118\]/li_983_527#
+ PHY_292/li_0_527# FILLER_22_1653/li_155_527# la_buf\[99\]/li_63_527# _492_/li_0_527#
+ _395_/li_0_n17# la_buf\[7\]/li_1075_527# FILLER_19_568/li_0_527# _379_/li_155_527#
+ PHY_550/li_0_527# ANTENNA_user_to_mprj_in_gates\[35\]_B/li_63_n17# user_to_mprj_in_buffers\[82\]/li_404_367#
+ _592_/li_155_n17# la_buf\[60\]/li_0_n17# ANTENNA__365__A/li_63_527# PHY_714/li_0_n17#
+ la_buf\[25\]/li_1167_n17# la_buf\[84\]/li_431_n17# PHY_232/li_0_527# PHY_715/li_0_527#
+ la_buf\[126\]/li_983_527# FILLER_20_2110/li_155_527# user_to_mprj_oen_buffers\[80\]/li_215_311#
+ FILLER_25_303/li_63_527# PHY_682/li_0_527# FILLER_28_55/li_63_527# PHY_720/li_0_n17#
+ la_buf\[6\]/li_983_527# user_to_mprj_oen_buffers\[54\]/li_615_527# FILLER_21_1440/li_63_n17#
+ powergood_check/FILLER_0_112/li_257_797# user_to_mprj_oen_buffers\[65\]/li_63_527#
+ PHY_457/li_0_n17# PHY_79/li_0_n17# FILLER_15_70/li_0_527# user_to_mprj_in_gates\[34\]/li_63_n17#
+ PHY_790/li_0_n17# user_to_mprj_oen_buffers\[39\]/li_215_311# _469_/li_155_n17# la_buf\[51\]/li_983_n17#
+ mprj_adr_buf\[26\]/li_17_51# FILLER_13_1587/li_63_527# powergood_check/FILLER_0_240/li_0_797#
+ _385_/li_0_527# user_to_mprj_oen_buffers\[22\]/li_891_527# FILLER_25_638/li_155_n17#
+ FILLER_13_1021/li_155_527# PHY_841/li_0_527# mprj_adr_buf\[28\]/li_247_n17# user_to_mprj_oen_buffers\[86\]/li_611_17#
+ user_to_mprj_in_gates\[98\]/li_707_367# PHY_530/li_0_n17# user_to_mprj_in_gates\[105\]/li_18_51#
+ PHY_847/li_0_n17# user_to_mprj_oen_buffers\[97\]/li_1535_527# _637_/li_0_527# powergood_check/FILLER_2_203/li_545_n17#
+ user_to_mprj_in_gates\[31\]/li_247_527# PHY_523/li_0_n17# mprj_dat_buf\[18\]/li_431_527#
+ mprj_dat_buf\[7\]/li_63_527# FILLER_12_1610/li_0_527# PHY_424/li_0_n17# PHY_319/li_0_527#
+ powergood_check/mprj_logic_high_lv/m1_0_n23# _597_/li_0_527# FILLER_9_1230/li_155_527#
+ la_buf\[109\]/li_611_17# _419_/li_0_527# PHY_223/li_0_n17# PHY_850/li_0_n17# user_to_mprj_in_buffers\[70\]/li_404_367#
+ powergood_check/mprj2_logic_high_lv/li_0_1611# _558_/li_247_527# mprj_pwrgood/li_19_289#
+ la_buf\[27\]/li_63_527# mprj_dat_buf\[4\]/li_17_51# la_buf\[65\]/li_247_n17# FILLER_20_284/li_0_n17#
+ PHY_32/li_0_n17# PHY_678/li_0_n17# PHY_770/li_0_527# PHY_396/li_0_527# user_to_mprj_oen_buffers\[22\]/li_207_51#
+ PHY_663/li_0_527# powergood_check/FILLER_1_62/li_545_n17# la_buf\[92\]/li_891_527#
+ user_to_mprj_in_gates\[40\]/li_247_n17# user_to_mprj_oen_buffers\[42\]/li_615_527#
+ FILLER_12_693/li_63_527# _651_/li_247_n17# mprj_adr_buf\[3\]/li_523_n17# _460_/li_0_n17#
+ _458_/li_0_527# FILLER_9_1060/li_0_527# FILLER_21_1876/li_0_527# powergood_check/FILLER_2_163/li_641_n17#
+ _571_/li_0_n17# user_to_mprj_in_gates\[60\]/li_707_n17# PHY_786/li_0_527# _349_/li_155_n17#
+ FILLER_2_294/li_0_527# user_to_mprj_oen_buffers\[27\]/li_215_311# _497_/li_0_527#
+ _599_/li_0_527# _646_/li_0_n17# PHY_414/li_0_527# _560_/li_155_527# user_to_mprj_oen_buffers\[44\]/li_1167_527#
+ user_to_mprj_in_gates\[101\]/li_247_n17# user_to_mprj_in_gates\[86\]/li_707_367#
+ FILLER_15_1988/li_155_n17# FILLER_24_512/li_63_n17# PHY_337/li_0_n17# FILLER_25_953/li_63_n17#
+ user_to_mprj_oen_buffers\[88\]/li_1075_n17# mprj_adr_buf\[17\]/li_207_51# mprj_dat_buf\[19\]/li_17_51#
+ la_buf\[50\]/li_611_17# PHY_767/li_0_527# PHY_753/li_0_527# la_buf\[50\]/li_795_379#
+ la_buf\[9\]/li_0_527# user_to_mprj_oen_buffers\[85\]/li_17_51# PHY_330/li_0_527#
+ mprj_sel_buf\[0\]/li_431_n17# _351_/li_155_n17# user_to_mprj_oen_buffers\[88\]/li_207_51#
+ FILLER_18_1805/li_63_527# PHY_769/li_0_n17# FILLER_0_54/li_63_527# PHY_434/li_0_n17#
+ _650_/li_155_n17# FILLER_15_1791/li_0_527# la_buf\[97\]/li_17_51# FILLER_14_359/li_0_527#
+ PHY_346/li_0_n17# FILLER_21_565/li_0_n17# _590_/li_247_527# PHY_415/li_0_527# user_to_mprj_oen_buffers\[29\]/li_0_527#
+ user_to_mprj_in_buffers\[17\]/li_404_367# mprj_adr_buf\[15\]/li_707_527# PHY_299/li_0_n17#
+ FILLER_8_981/li_0_527# _478_/li_0_n17# la_buf\[89\]/li_247_527# PHY_716/li_0_n17#
+ user_to_mprj_oen_buffers\[15\]/li_215_311# PHY_367/li_0_527# user_to_mprj_in_gates\[52\]/li_18_51#
+ PHY_12/li_0_n17# la_buf\[94\]/li_707_527# PHY_182/li_0_n17# user_to_mprj_oen_buffers\[80\]/li_0_527#
+ ANTENNA__350__A/li_63_n17# _537_/li_0_n17# ANTENNA__657__A/li_63_n17# ANTENNA_la_buf\[120\]_A/li_63_n17#
+ user_to_mprj_in_gates\[59\]/li_339_n17# _432_/li_0_527# _440_/li_247_527# _541_/li_247_527#
+ user_to_mprj_oen_buffers\[90\]/li_207_51# user_to_mprj_in_gates\[74\]/li_707_367#
+ PHY_771/li_0_n17# FILLER_12_1021/li_0_527# user_to_mprj_oen_buffers\[59\]/li_1351_n17#
+ PHY_766/li_0_527# la_buf\[84\]/li_1259_n17# FILLER_19_1417/li_155_n17# la_buf\[3\]/li_431_527#
+ PHY_727/li_0_n17# PHY_312/li_0_n17# _353_/li_247_n17# la_buf\[113\]/li_207_51# PHY_713/li_0_527#
+ FILLER_11_996/li_0_527# powergood_check/FILLER_2_243/li_353_797# ANTENNA__575__A/li_63_n17#
+ FILLER_18_1556/li_0_n17# powergood_check/FILLER_2_0/li_257_n17# user_to_mprj_oen_buffers\[34\]/li_17_51#
+ FILLER_24_56/li_155_527# _617_/li_247_527# PHY_857/li_0_527# _560_/li_0_527# la_buf\[46\]/li_17_51#
+ PHY_491/li_0_527# PHY_164/li_0_527# mprj_clk2_buf/li_779_17# la_buf\[52\]/li_207_51#
+ powergood_check/FILLER_1_164/li_65_797# _451_/li_0_527# PHY_484/li_0_527# user_to_mprj_oen_buffers\[60\]/li_983_n17#
+ la_buf\[77\]/li_247_527# _506_/li_0_527# _577_/li_0_n17# ANTENNA_user_to_mprj_in_gates\[71\]_A/li_63_527#
+ FILLER_21_1570/li_0_527# user_to_mprj_oen_buffers\[44\]/li_707_n17# _552_/li_0_527#
+ user_to_mprj_in_gates\[47\]/li_339_n17# FILLER_16_1711/li_0_527# PHY_733/li_0_527#
+ FILLER_11_916/li_155_527# powergood_check/FILLER_0_96/li_353_n17# PHY_411/li_0_527#
+ _430_/li_247_n17# PHY_326/li_0_527# powergood_check/FILLER_1_244/li_641_n17# powergood_check/FILLER_2_16/li_641_797#
+ FILLER_14_1692/li_155_527# FILLER_16_1581/li_63_n17# FILLER_12_1482/li_63_n17# _464_/li_247_527#
+ user_to_mprj_oen_buffers\[71\]/li_795_379# powergood_check/FILLER_0_264/li_353_797#
+ PHY_734/li_0_527# la_buf\[86\]/li_247_n17# _596_/li_155_n17# user_to_mprj_in_gates\[123\]/li_707_367#
+ la_buf\[65\]/li_63_n17# user_to_mprj_in_gates\[28\]/li_615_n17# _335_/li_0_n17#
+ user_to_mprj_oen_buffers\[81\]/li_431_n17# ANTENNA__563__A/li_63_n17# la_buf\[53\]/li_707_527#
+ PHY_407/li_0_n17# powergood_check/FILLER_2_235/li_161_n17# la_buf\[110\]/li_795_379#
+ PHY_401/li_0_n17# mprj_stb_buf/li_63_n17# FILLER_11_1674/li_63_n17# powergood_check/FILLER_0_184/li_161_797#
+ FILLER_9_559/li_155_n17# FILLER_15_1692/li_63_527# user_to_mprj_in_gates\[38\]/li_523_n17#
+ ANTENNA__647__A/li_0_n17# powergood_check/FILLER_1_32/li_65_n17# la_buf\[120\]/li_431_n17#
+ user_to_mprj_oen_buffers\[7\]/li_1443_527# PHY_480/li_0_527# FILLER_12_734/li_0_n17#
+ PHY_719/li_0_527# la_buf\[67\]/li_523_n17# user_to_mprj_oen_buffers\[18\]/li_891_527#
+ mprj_dat_buf\[12\]/li_207_51# _386_/li_155_527# PHY_376/li_0_n17# PHY_416/li_0_527#
+ user_to_mprj_oen_buffers\[37\]/li_707_527# user_to_mprj_in_gates\[32\]/li_0_n17#
+ PHY_220/li_0_n17# powergood_check/FILLER_1_0/li_161_n17# FILLER_9_534/li_63_n17#
+ FILLER_16_1415/li_63_527# powergood_check/FILLER_1_48/li_100_536# PHY_115/li_0_527#
+ PHY_714/li_0_527# PHY_28/li_0_n17# FILLER_12_617/li_0_527# la_buf\[45\]/li_1167_527#
+ PHY_231/li_0_527# PHY_718/li_0_527# FILLER_12_1374/li_63_n17# _598_/li_247_n17#
+ PHY_839/li_0_527# PHY_744/li_0_527# mprj_adr_buf\[22\]/li_611_17# _602_/li_0_527#
+ FILLER_12_748/li_0_527# _476_/li_155_n17# la_buf\[74\]/li_247_n17# powergood_check/FILLER_2_8/li_545_n17#
+ user_to_mprj_in_gates\[88\]/li_707_n17# mprj_adr_buf\[3\]/li_215_311# FILLER_12_1923/li_63_n17#
+ la_buf\[17\]/li_1443_n17# _413_/li_0_527# FILLER_15_543/li_0_527# powergood_check/FILLER_1_48/li_449_797#
+ user_to_mprj_oen_buffers\[27\]/li_207_51# user_to_mprj_in_gates\[104\]/li_0_n17#
+ FILLER_19_1581/li_0_527# PHY_759/li_0_527# FILLER_15_73/li_63_527# FILLER_10_625/li_63_n17#
+ FILLER_9_1273/li_155_527# mprj_dat_buf\[29\]/li_247_n17# user_to_mprj_oen_buffers\[109\]/li_17_51#
+ PHY_423/li_0_n17# PHY_372/li_0_527# user_to_mprj_in_gates\[69\]/li_615_527# FILLER_21_1436/li_63_527#
+ PHY_363/li_0_n17# PHY_788/li_0_527# FILLER_13_1084/li_155_527# la_buf\[88\]/li_0_527#
+ user_to_mprj_in_gates\[90\]/li_431_527# FILLER_10_497/li_0_n17# la_buf\[73\]/li_891_527#
+ mprj_adr_buf\[7\]/li_1351_527# mprj_adr_buf\[25\]/li_17_51# _656_/li_0_527# FILLER_9_1173/li_0_527#
+ FILLER_22_1704/li_0_527# FILLER_19_1754/li_0_n17# FILLER_25_815/li_155_527# user_to_mprj_in_gates\[104\]/li_18_51#
+ user_to_mprj_oen_buffers\[66\]/li_247_527# PHY_358/li_0_527# user_to_mprj_in_gates\[49\]/li_431_527#
+ _402_/li_0_527# FILLER_11_1709/li_63_527# FILLER_16_548/li_0_527# FILLER_20_1983/li_0_527#
+ _654_/li_0_n17# _498_/li_0_527# ANTENNA_user_to_mprj_in_gates\[102\]_B/li_63_n17#
+ _356_/li_155_n17# _409_/li_0_527# powergood_check/FILLER_2_219/li_0_n17# _655_/li_155_n17#
+ user_to_mprj_in_gates\[3\]/li_707_367# FILLER_21_1812/li_0_527# powergood_check/FILLER_0_168/li_0_797#
+ mprj_rstn_buf/li_0_n17# la_buf\[63\]/li_1443_527# mprj_dat_buf\[3\]/li_17_51# user_to_mprj_oen_buffers\[114\]/li_779_17#
+ PHY_38/li_0_527# FILLER_19_1471/li_0_527# FILLER_11_846/li_0_527# mprj_adr_buf\[24\]/li_207_51#
+ _611_/li_0_527# user_to_mprj_oen_buffers\[16\]/li_431_n17# FILLER_13_1048/li_155_527#
+ PHY_302/li_0_n17# powergood_check/FILLER_1_164/li_0_797# _578_/li_0_527# PHY_860/li_0_n17#
+ FILLER_9_386/li_63_n17# la_buf\[41\]/li_247_527# powergood_check/FILLER_0_232/li_115_72#
+ ANTENNA_user_to_mprj_in_gates\[92\]_A/li_63_n17# user_to_mprj_oen_buffers\[95\]/li_207_51#
+ ANTENNA_user_to_mprj_in_gates\[64\]_A/li_63_527# _487_/li_0_527# FILLER_3_759/li_63_527#
+ user_to_mprj_in_gates\[32\]/li_707_n17# PHY_457/li_0_527# PHY_263/li_0_527# PHY_395/li_0_527#
+ mprj_adr_buf\[2\]/li_1075_n17# FILLER_13_1067/li_63_527# FILLER_14_491/li_63_527#
+ FILLER_11_1132/li_63_527# powergood_check/FILLER_2_115/li_0_797# FILLER_25_1099/li_155_n17#
+ PHY_176/li_0_n17# la_buf\[6\]/li_1259_n17# FILLER_21_1741/li_155_n17# FILLER_11_507/li_63_n17#
+ la_buf\[118\]/li_207_51# user_to_mprj_in_gates\[65\]/li_155_n17# FILLER_22_1913/li_0_n17#
+ la_buf\[94\]/li_615_527# mprj_dat_buf\[18\]/li_17_51# PHY_860/li_0_527# user_to_mprj_oen_buffers\[95\]/li_247_n17#
+ PHY_97/li_0_n17# mprj_stb_buf/li_207_51# la_buf\[50\]/li_247_n17# user_to_mprj_oen_buffers\[84\]/li_17_51#
+ powergood_check/FILLER_1_62/li_115_72# _535_/li_155_n17# mprj_stb_buf/li_247_527#
+ la_buf\[79\]/li_215_311# user_to_mprj_oen_buffers\[22\]/li_707_n17# user_to_mprj_in_buffers\[31\]/li_523_n17#
+ la_buf\[96\]/li_17_51# FILLER_0_288/li_63_n17# la_buf\[57\]/li_207_51# PHY_364/li_0_527#
+ _563_/li_247_527# la_buf\[47\]/li_1351_527# FILLER_13_1203/li_63_n17# user_to_mprj_in_buffers\[0\]/li_523_527#
+ mprj_dat_buf\[19\]/li_891_n17# user_to_mprj_in_gates\[44\]/li_155_527# user_to_mprj_oen_buffers\[91\]/li_523_n17#
+ FILLER_12_1931/li_0_527# FILLER_12_978/li_63_527# la_buf\[120\]/li_207_51# PHY_818/li_0_n17#
+ _361_/li_247_527# _479_/li_0_527# user_to_mprj_in_gates\[51\]/li_18_51# PHY_432/li_0_527#
+ FILLER_12_693/li_0_527# ANTENNA__472__A/li_63_527# la_buf\[38\]/li_779_17# powergood_check/FILLER_1_228/li_0_797#
+ la_buf\[113\]/li_247_527# la_buf\[7\]/li_1535_527# FILLER_24_1886/li_63_527# FILLER_21_1383/li_0_527#
+ FILLER_24_1425/li_0_n17# FILLER_19_1756/li_155_n17# FILLER_16_1681/li_0_527# PHY_778/li_0_527#
+ _603_/li_0_527# FILLER_26_876/li_0_527# powergood_check/FILLER_1_140/li_545_797#
+ powergood_check/FILLER_2_211/li_257_797# user_to_mprj_oen_buffers\[83\]/li_247_n17#
+ FILLER_12_1044/li_0_527# FILLER_26_457/li_0_527# _415_/li_155_n17# FILLER_28_1735/li_0_527#
+ FILLER_11_1433/li_0_n17# la_buf\[67\]/li_215_311# user_to_mprj_in_buffers\[39\]/li_615_n17#
+ PHY_450/li_0_n17# user_to_mprj_oen_buffers\[33\]/li_17_51# mprj_pwrgood/li_247_527#
+ mprj_pwrgood/li_607_367# la_buf\[122\]/li_247_n17# FILLER_24_1401/li_0_527# PHY_757/li_0_527#
+ FILLER_25_1047/li_0_n17# PHY_767/li_0_n17# FILLER_13_1207/li_155_527# FILLER_11_1264/li_63_n17#
+ user_to_mprj_in_gates\[34\]/li_431_n17# la_buf\[2\]/li_247_n17# la_buf\[45\]/li_17_51#
+ user_to_mprj_oen_buffers\[4\]/li_215_311# PHY_334/li_0_527# FILLER_15_357/li_63_n17#
+ _512_/li_0_527# la_buf\[31\]/li_1259_527# user_to_mprj_in_gates\[32\]/li_155_527#
+ _655_/li_0_n17# mprj_adr_buf\[28\]/li_707_n17# PHY_318/li_0_527# mprj_dat_buf\[17\]/li_207_51#
+ _441_/li_0_527# la_buf\[72\]/li_63_n17# FILLER_17_1925/li_0_527# user_to_mprj_oen_buffers\[82\]/li_1443_n17#
+ FILLER_12_593/li_63_527# PHY_494/li_0_527# powergood_check/FILLER_2_171/li_353_797#
+ _505_/li_0_n17# PHY_220/li_0_527# _549_/li_0_n17# powergood_check/FILLER_1_212/li_545_n17#
+ FILLER_11_1035/li_63_n17# FILLER_13_925/li_0_527# PHY_331/li_0_527# _452_/li_0_527#
+ PHY_412/li_0_527# user_to_mprj_in_gates\[85\]/li_523_527# powergood_check/FILLER_0_232/li_257_797#
+ PHY_762/li_0_527# PHY_765/li_0_527# mprj_sel_buf\[3\]/li_1259_527# _432_/li_247_n17#
+ mprj_adr_buf\[27\]/li_611_17# FILLER_12_1357/li_155_n17# PHY_271/li_0_n17# FILLER_21_1573/li_63_n17#
+ la_buf\[12\]/li_1259_n17# FILLER_13_911/li_0_527# _393_/li_155_527# _588_/li_0_n17#
+ FILLER_22_1886/li_63_527# user_to_mprj_oen_buffers\[85\]/li_891_n17# FILLER_18_504/li_0_527#
+ user_to_mprj_in_gates\[40\]/li_707_n17# la_buf\[9\]/li_1075_n17# mprj_dat_buf\[3\]/li_891_527#
+ user_to_mprj_in_gates\[19\]/li_18_51# ANTENNA_user_to_mprj_in_gates\[39\]_B/li_63_527#
+ la_buf\[34\]/li_63_527# la_buf\[55\]/li_215_311# mprj_dat_buf\[25\]/li_615_527#
+ FILLER_15_2067/li_63_527# FILLER_17_108/li_0_n17# _528_/li_0_n17# _476_/li_0_n17#
+ FILLER_25_1903/li_63_n17# la_buf\[29\]/li_615_527# FILLER_12_1117/li_63_527# powergood_check/FILLER_0_16/li_65_797#
+ powergood_check/FILLER_0_272/li_545_797# PHY_433/li_0_527# FILLER_18_1459/li_155_n17#
+ FILLER_16_2087/li_0_527# FILLER_13_1203/li_155_527# mprj_logic_high_inst/m1_566_1040#
+ _500_/li_0_527# FILLER_14_1500/li_63_527# _500_/li_247_527# user_to_mprj_in_gates\[92\]/li_247_527#
+ la_buf\[4\]/li_891_n17# _545_/li_0_527# user_to_mprj_in_gates\[101\]/li_707_n17#
+ powergood_check/FILLER_1_172/li_641_n17# powergood_check/FILLER_2_243/li_353_n17#
+ user_to_mprj_oen_buffers\[50\]/li_247_527# powergood_check/mprj2_logic_high_lv/li_1121_1611#
+ mprj2_logic_high_inst/m2_1030_1294# la_buf\[39\]/li_63_527# powergood_check/FILLER_0_192/li_353_797#
+ PHY_229/li_0_n17# FILLER_19_411/li_0_527# FILLER_19_1475/li_155_527# _572_/li_247_527#
+ FILLER_15_1523/li_0_n17# user_to_mprj_oen_buffers\[34\]/li_207_51# FILLER_9_575/li_0_527#
+ la_buf\[102\]/li_63_527# powergood_check/FILLER_2_163/li_161_n17# PHY_26/li_0_527#
+ user_to_mprj_in_gates\[73\]/li_523_527# user_to_mprj_oen_buffers\[2\]/li_611_17#
+ user_to_mprj_oen_buffers\[28\]/li_707_n17# PHY_835/li_0_n17# FILLER_23_1678/li_0_n17#
+ powergood_check/FILLER_2_219/li_545_797# PHY_828/li_0_527# PHY_858/li_0_527# _545_/li_0_n17#
+ FILLER_21_2061/li_63_n17# la_buf\[123\]/li_611_17# user_to_mprj_oen_buffers\[15\]/li_779_17#
+ powergood_check/FILLER_0_32/li_641_797# _572_/li_155_527# PHY_799/li_0_527# user_to_mprj_oen_buffers\[88\]/li_215_311#
+ la_buf\[41\]/li_63_527# mprj_sel_buf\[3\]/li_207_51# la_buf\[43\]/li_215_311# mprj2_logic_high_inst/li_0_527#
+ ANTENNA_user_to_mprj_in_buffers\[18\]_A/li_63_n17# la_buf\[17\]/li_615_527# powergood_check/FILLER_2_16/li_641_n17#
+ FILLER_18_1582/li_0_527# la_buf\[127\]/li_215_311# FILLER_23_493/li_0_n17# la_buf\[50\]/li_0_527#
+ mprj_adr_buf\[29\]/li_207_51# PHY_296/li_0_527# user_to_mprj_oen_buffers\[108\]/li_17_51#
+ PHY_717/li_0_n17# FILLER_9_928/li_155_n17# user_to_mprj_oen_buffers\[40\]/li_523_n17#
+ la_buf\[7\]/li_215_311# FILLER_15_1692/li_0_527# FILLER_13_2020/li_155_n17# user_to_mprj_in_buffers\[109\]/li_155_n17#
+ user_to_mprj_oen_buffers\[63\]/li_707_n17# FILLER_11_409/li_155_527# _363_/li_155_n17#
+ user_to_mprj_oen_buffers\[52\]/li_891_527# FILLER_18_539/li_155_527# PHY_27/li_0_n17#
+ powergood_check/FILLER_2_179/li_641_797# _543_/li_0_n17# user_to_mprj_oen_buffers\[42\]/li_1167_527#
+ mprj_adr_buf\[24\]/li_17_51# user_to_mprj_in_gates\[39\]/li_247_527# PHY_832/li_0_527#
+ user_to_mprj_in_gates\[61\]/li_523_527# user_to_mprj_in_gates\[103\]/li_18_51# PHY_83/li_0_n17#
+ mprj_adr_buf\[31\]/li_207_51# user_to_mprj_in_buffers\[78\]/li_404_367# user_to_mprj_oen_buffers\[91\]/li_615_527#
+ FILLER_25_1204/li_155_n17# FILLER_9_550/li_63_n17# user_to_mprj_oen_buffers\[7\]/li_795_379#
+ FILLER_25_1107/li_63_n17# powergood_check/FILLER_2_251/li_449_797# user_to_mprj_oen_buffers\[76\]/li_215_311#
+ _651_/li_0_527# la_buf\[31\]/li_215_311# user_to_mprj_in_gates\[48\]/li_247_n17#
+ user_to_mprj_oen_buffers\[4\]/li_207_51# PHY_447/li_0_n17# mprj_dat_buf\[2\]/li_17_51#
+ la_buf\[15\]/li_1075_n17# FILLER_26_43/li_0_n17# user_to_mprj_in_buffers\[28\]/li_236_17#
+ PHY_179/li_0_n17# la_buf\[115\]/li_215_311# la_buf\[125\]/li_207_51# PHY_792/li_0_n17#
+ mprj_dat_buf\[22\]/li_611_17# user_to_mprj_in_gates\[109\]/li_247_n17# powergood_check/FILLER_1_48/li_449_n17#
+ _633_/li_0_527# FILLER_6_755/li_0_527# PHY_705/li_0_527# _542_/li_155_n17# la_buf\[11\]/li_63_n17#
+ mprj_dat_buf\[3\]/li_215_311# _477_/li_0_527# user_to_mprj_in_gates\[99\]/li_339_527#
+ user_to_mprj_in_gates\[27\]/li_247_527# FILLER_28_43/li_0_n17# PHY_291/li_0_527#
+ la_buf\[64\]/li_207_51# la_buf\[86\]/li_707_n17# la_buf\[106\]/li_779_17# PHY_628/li_0_527#
+ _400_/li_247_527# FILLER_11_1553/li_63_527# user_to_mprj_in_buffers\[66\]/li_404_367#
+ user_to_mprj_oen_buffers\[4\]/li_1351_527# PHY_760/li_0_527# FILLER_12_1117/li_63_n17#
+ _615_/li_0_527# mprj_dat_buf\[17\]/li_17_51# user_to_mprj_in_gates\[113\]/li_247_527#
+ FILLER_13_1096/li_63_527# _657_/li_0_527# FILLER_11_413/li_63_527# FILLER_9_992/li_155_527#
+ user_to_mprj_oen_buffers\[127\]/li_1351_527# user_to_mprj_oen_buffers\[64\]/li_215_311#
+ user_to_mprj_oen_buffers\[83\]/li_17_51# _633_/li_247_527# powergood_check/FILLER_2_16/li_161_797#
+ powergood_check/FILLER_1_244/li_161_n17# la_buf\[40\]/li_1259_527# la_buf\[74\]/li_1167_n17#
+ la_buf\[14\]/li_983_527# user_to_mprj_in_gates\[110\]/li_523_527# user_to_mprj_in_gates\[36\]/li_247_n17#
+ FILLER_17_245/li_63_527# user_to_mprj_oen_buffers\[37\]/li_611_17# FILLER_13_106/li_63_527#
+ _541_/li_0_n17# la_buf\[95\]/li_17_51# FILLER_9_1036/li_0_527# user_to_mprj_oen_buffers\[120\]/li_215_311#
+ la_buf\[103\]/li_215_311# PHY_481/li_0_527# powergood_check/FILLER_2_300/li_0_797#
+ user_to_mprj_in_buffers\[46\]/li_155_n17# PHY_390/li_0_527# PHY_751/li_0_527# ANTENNA__358__A/li_63_n17#
+ FILLER_12_1044/li_63_n17# powergood_check/FILLER_1_62/li_0_797# user_to_mprj_oen_buffers\[15\]/li_983_n17#
+ FILLER_20_496/li_155_n17# user_to_mprj_in_gates\[90\]/li_431_n17# ANTENNA_user_to_mprj_in_gates\[78\]_A/li_63_n17#
+ user_to_mprj_in_gates\[50\]/li_18_51# la_buf\[109\]/li_523_n17# FILLER_17_56/li_63_527#
+ user_to_mprj_in_gates\[87\]/li_339_527# user_to_mprj_in_buffers\[96\]/li_236_17#
+ FILLER_11_1004/li_63_527# la_buf\[74\]/li_707_n17# user_to_mprj_oen_buffers\[37\]/li_983_n17#
+ FILLER_23_245/li_63_527# PHY_795/li_0_n17# user_to_mprj_in_buffers\[97\]/li_523_n17#
+ ANTENNA__659__A/li_63_527# powergood_check/FILLER_2_163/li_65_n17# FILLER_13_1038/li_63_527#
+ PHY_766/li_0_n17# _449_/li_0_n17# user_to_mprj_in_buffers\[54\]/li_404_367# FILLER_22_387/li_63_n17#
+ FILLER_18_1463/li_63_n17# mprj_dat_buf\[24\]/li_207_51# _475_/li_155_527# PHY_488/li_0_527#
+ user_to_mprj_in_gates\[104\]/li_63_n17# user_to_mprj_in_gates\[69\]/li_18_51# PHY_33/li_0_n17#
+ PHY_353/li_0_527# PHY_724/li_0_527# FILLER_22_520/li_63_527# user_to_mprj_oen_buffers\[52\]/li_215_311#
+ FILLER_20_496/li_0_n17# powergood_check/FILLER_1_8/li_65_n17# FILLER_17_231/li_0_n17#
+ powergood_check/FILLER_2_115/li_0_n17# PHY_332/li_0_n17# _455_/li_0_527# PHY_54/li_0_n17#
+ user_to_mprj_in_gates\[96\]/li_339_n17# PHY_387/li_0_n17# PHY_385/li_0_527# PHY_762/li_0_n17#
+ user_to_mprj_oen_buffers\[32\]/li_17_51# FILLER_19_1609/li_0_527# la_buf\[44\]/li_17_51#
+ PHY_730/li_0_527# FILLER_21_2075/li_0_527# ANTENNA__346__A/li_63_n17# FILLER_22_349/li_63_n17#
+ FILLER_21_527/li_0_n17# user_to_mprj_in_gates\[80\]/li_339_n17# user_to_mprj_oen_buffers\[39\]/li_207_51#
+ _611_/li_247_n17# mprj_adr_buf\[25\]/li_983_n17# FILLER_16_444/li_0_527# user_to_mprj_oen_buffers\[62\]/li_1351_n17#
+ PHY_15/li_0_527# la_buf\[119\]/li_431_527# powergood_check/FILLER_0_240/li_100_536#
+ _542_/li_0_527# la_buf\[6\]/li_0_n17# user_to_mprj_oen_buffers\[7\]/li_611_17# mprj_dat_buf\[30\]/li_795_379#
+ FILLER_14_1399/li_0_527# FILLER_7_1029/li_0_n17# FILLER_16_520/li_63_527# FILLER_23_1896/li_63_n17#
+ user_to_mprj_in_buffers\[49\]/li_523_527# powergood_check/FILLER_1_196/li_115_72#
+ PHY_712/li_0_527# ANTENNA_user_to_mprj_oen_buffers\[108\]_TE/li_63_n17# mprj_dat_buf\[7\]/li_431_527#
+ la_buf\[122\]/li_1351_n17# la_buf\[118\]/li_795_379# _503_/li_0_n17# _577_/li_155_527#
+ la_buf\[46\]/li_63_527# _449_/li_247_527# powergood_check/FILLER_1_228/li_0_n17#
+ _578_/li_0_n17# user_to_mprj_oen_buffers\[40\]/li_215_311# user_to_mprj_in_gates\[18\]/li_18_51#
+ user_to_mprj_oen_buffers\[41\]/li_207_51# powergood_check/FILLER_0_240/li_449_797#
+ la_buf\[95\]/li_891_n17# _339_/li_247_527# user_to_mprj_in_gates\[84\]/li_339_n17#
+ _467_/li_0_n17# la_buf\[67\]/li_611_17# mprj_dat_buf\[6\]/li_795_379# powergood_check/FILLER_1_140/li_545_n17#
+ powergood_check/FILLER_2_211/li_257_n17# FILLER_16_558/li_0_527# FILLER_25_934/li_63_527#
+ _354_/li_0_n17# powergood_check/FILLER_0_160/li_257_797# mprj_adr_buf\[2\]/li_1535_n17#
+ PHY_739/li_0_527# FILLER_17_1457/li_63_527# _368_/li_155_n17# FILLER_10_509/li_0_n17#
+ PHY_715/li_0_n17# PHY_322/li_0_n17# user_to_mprj_in_gates\[65\]/li_615_n17# user_to_mprj_oen_buffers\[93\]/li_1443_527#
+ user_to_mprj_oen_buffers\[66\]/li_0_n17# user_to_mprj_in_gates\[63\]/li_339_527#
+ FILLER_13_855/li_63_527# FILLER_19_1631/li_63_n17# mprj_stb_buf/li_1167_527# _393_/li_0_n17#
+ powergood_check/FILLER_2_251/li_545_n17# user_to_mprj_oen_buffers\[61\]/li_63_527#
+ _638_/li_0_n17# powergood_check/FILLER_2_227/li_115_72# PHY_833/li_0_n17# user_to_mprj_in_gates\[119\]/li_707_367#
+ _617_/li_0_527# PHY_728/li_0_527# la_buf\[101\]/li_707_n17# la_buf\[51\]/li_1259_n17#
+ la_buf\[106\]/li_795_379# la_buf\[32\]/li_431_n17# powergood_check/FILLER_2_115/li_115_72#
+ powergood_check/FILLER_2_107/li_257_797# FILLER_27_798/li_63_n17# ANTENNA_user_to_mprj_in_gates\[106\]_B/li_63_527#
+ powergood_check/FILLER_2_171/li_353_n17# PHY_52/li_0_527# user_to_mprj_oen_buffers\[9\]/li_207_51#
+ powergood_check/FILLER_0_208/li_100_536# ANTENNA__375__A/li_0_n17# la_buf\[116\]/li_431_n17#
+ FILLER_25_324/li_63_n17# FILLER_24_1758/li_0_527# PHY_745/li_0_n17# PHY_800/li_0_n17#
+ user_to_mprj_oen_buffers\[107\]/li_17_51# user_to_mprj_oen_buffers\[44\]/li_1075_n17#
+ user_to_mprj_oen_buffers\[88\]/li_779_17# PHY_259/li_0_527# la_buf\[113\]/li_707_527#
+ _584_/li_0_527# user_to_mprj_in_gates\[120\]/li_615_527# user_to_mprj_oen_buffers\[56\]/li_431_527#
+ PHY_726/li_0_527# FILLER_24_520/li_155_527# la_buf\[14\]/li_63_527# _547_/li_155_n17#
+ powergood_check/FILLER_2_0/li_115_72# user_to_mprj_in_gates\[46\]/li_707_367# FILLER_27_794/li_63_n17#
+ PHY_784/li_0_527# powergood_check/FILLER_0_208/li_449_797# FILLER_20_2087/li_155_n17#
+ PHY_772/li_0_527# powergood_check/FILLER_0_272/li_545_n17# FILLER_25_1422/li_63_n17#
+ mprj_adr_buf\[23\]/li_17_51# la_buf\[69\]/li_207_51# user_to_mprj_oen_buffers\[92\]/li_0_527#
+ user_to_mprj_in_gates\[120\]/li_0_527# FILLER_9_501/li_63_n17# FILLER_9_996/li_0_n17#
+ la_buf\[6\]/li_795_379# user_to_mprj_in_gates\[102\]/li_18_51# PHY_547/li_0_n17#
+ user_to_mprj_in_gates\[107\]/li_707_367# mprj_pwrgood/li_707_527# user_to_mprj_oen_buffers\[90\]/li_779_17#
+ la_buf\[20\]/li_431_n17# la_buf\[34\]/li_1351_n17# _337_/li_155_527# powergood_check/FILLER_1_268/li_65_n17#
+ FILLER_25_1903/li_0_n17# FILLER_26_1195/li_0_527# PHY_756/li_0_527# PHY_360/li_0_n17#
+ user_to_mprj_oen_buffers\[7\]/li_247_n17# user_to_mprj_in_gates\[32\]/li_615_527#
+ _641_/li_0_527# FILLER_24_311/li_0_n17# mprj_cyc_buf/li_1627_n17# powergood_check/FILLER_1_156/li_65_n17#
+ PHY_802/li_0_527# la_buf\[71\]/li_207_51# mprj_dat_buf\[1\]/li_17_51# powergood_check/FILLER_2_219/li_545_n17#
+ FILLER_9_792/li_0_527# user_to_mprj_oen_buffers\[1\]/li_1075_n17# powergood_check/FILLER_0_168/li_545_797#
+ user_to_mprj_in_buffers\[109\]/li_51_17# PHY_366/li_0_n17# user_to_mprj_in_buffers\[3\]/li_404_17#
+ _461_/li_0_527# user_to_mprj_oen_buffers\[23\]/li_63_527# mprj_dat_buf\[30\]/li_707_527#
+ user_to_mprj_oen_buffers\[74\]/li_1259_n17# user_to_mprj_in_gates\[27\]/li_707_n17#
+ user_to_mprj_in_buffers\[14\]/li_404_17# PHY_382/li_0_n17# PHY_486/li_0_527# user_to_mprj_oen_buffers\[80\]/li_1351_527#
+ powergood_check/mprj2_logic_high_hvl/li_0_797# user_to_mprj_oen_buffers\[44\]/li_611_17#
+ powergood_check/FILLER_0_200/li_641_797# _524_/li_0_527# FILLER_14_1533/li_155_527#
+ mprj_adr_buf\[4\]/li_1167_n17# FILLER_16_88/li_63_n17# user_to_mprj_in_gates\[95\]/li_431_n17#
+ mprj_dat_buf\[29\]/li_207_51# FILLER_25_949/li_155_n17# user_to_mprj_in_gates\[109\]/li_63_n17#
+ user_to_mprj_oen_buffers\[56\]/li_0_n17# PHY_324/li_0_n17# la_buf\[84\]/li_63_n17#
+ powergood_check/FILLER_2_179/li_641_n17# powergood_check/mprj_logic_high_lv/li_929_1611#
+ FILLER_26_1066/li_0_527# mprj_dat_buf\[16\]/li_17_51# mprj_adr_buf\[29\]/li_983_527#
+ la_buf\[98\]/li_247_527# PHY_232/li_0_n17# FILLER_15_1998/li_0_527# mprj_adr_buf\[11\]/li_983_n17#
+ user_to_mprj_oen_buffers\[82\]/li_17_51# FILLER_5_954/li_63_527# FILLER_10_463/li_63_527#
+ mprj_dat_buf\[18\]/li_1259_527# PHY_177/li_0_527# PHY_270/li_0_527# FILLER_19_1754/li_0_527#
+ la_buf\[94\]/li_17_51# mprj_adr_buf\[22\]/li_215_311# PHY_843/li_0_527# PHY_371/li_0_527#
+ mprj_dat_buf\[27\]/li_1351_n17# FILLER_7_1774/li_63_n17# mprj_dat_buf\[31\]/li_207_51#
+ powergood_check/FILLER_1_196/li_0_n17# powergood_check/FILLER_2_24/li_353_797# user_to_mprj_in_gates\[111\]/li_63_n17#
+ ANTENNA_user_to_mprj_in_gates\[42\]_A/li_63_n17# powergood_check/FILLER_0_256/li_0_n17#
+ powergood_check/mprj2_logic_high_lv/li_756_683# user_to_mprj_in_gates\[14\]/li_707_367#
+ mprj_clk_buf/li_611_17# la_buf\[0\]/li_207_51# user_to_mprj_in_gates\[22\]/li_707_367#
+ _606_/li_155_n17# FILLER_13_620/li_63_n17# FILLER_15_2039/li_0_527# _518_/li_0_n17#
+ mprj_logic_high_inst/m3_800_851# FILLER_9_989/li_63_527# powergood_check/FILLER_1_172/li_161_n17#
+ PHY_187/li_0_n17# PHY_188/li_0_n17# user_to_mprj_oen_buffers\[91\]/li_63_527# _388_/li_0_527#
+ mprj_dat_buf\[0\]/li_63_527# FILLER_13_1013/li_0_n17# user_to_mprj_in_gates\[60\]/li_63_n17#
+ PHY_764/li_0_n17# PHY_86/li_0_n17# user_to_mprj_in_gates\[81\]/li_155_527# ANTENNA_user_to_mprj_in_gates\[110\]_B/li_63_n17#
+ user_to_mprj_oen_buffers\[57\]/li_63_n17# FILLER_26_676/li_0_527# user_to_mprj_in_gates\[80\]/li_707_n17#
+ user_to_mprj_in_gates\[68\]/li_18_51# PHY_735/li_0_527# user_to_mprj_oen_buffers\[46\]/li_207_51#
+ powergood_check/FILLER_0_240/li_65_797# user_to_mprj_in_buffers\[65\]/li_615_527#
+ PHY_93/li_0_527# user_to_mprj_oen_buffers\[31\]/li_17_51# user_to_mprj_in_buffers\[107\]/li_0_527#
+ la_buf\[27\]/li_523_n17# mprj_dat_buf\[21\]/li_247_527# powergood_check/FILLER_0_32/li_161_797#
+ mprj_adr_buf\[10\]/li_215_311# la_buf\[43\]/li_17_51# PHY_787/li_0_n17# user_to_mprj_oen_buffers\[100\]/li_611_17#
+ _584_/li_155_527# la_buf\[53\]/li_63_527# powergood_check/FILLER_2_16/li_161_n17#
+ FILLER_25_827/li_155_n17# user_to_mprj_in_gates\[3\]/li_0_527# powergood_check/FILLER_2_259/li_353_797#
+ mprj_dat_buf\[29\]/li_0_n17# user_to_mprj_in_gates\[1\]/li_339_n17# FILLER_12_906/li_0_527#
+ mprj_cyc_buf/li_63_527# la_buf\[102\]/li_0_527# user_to_mprj_in_gates\[89\]/li_707_367#
+ FILLER_11_585/li_0_n17# FILLER_1_59/li_63_n17# mprj_adr_buf\[3\]/li_207_51# la_buf\[74\]/li_611_17#
+ user_to_mprj_oen_buffers\[59\]/li_63_n17# FILLER_22_1653/li_155_n17# powergood_check/FILLER_1_180/li_65_797#
+ FILLER_11_1717/li_63_n17# powergood_check/FILLER_1_62/li_0_n17# PHY_99/li_0_527#
+ _375_/li_155_n17# FILLER_17_2088/li_0_n17# user_to_mprj_in_gates\[35\]/li_0_527#
+ FILLER_12_873/li_0_527# la_buf\[110\]/li_1351_527# PHY_799/li_0_n17# _572_/li_0_n17#
+ powergood_check/mprj2_logic_high_lv/li_1455_797# FILLER_9_1234/li_0_527# FILLER_26_1176/li_63_527#
+ FILLER_17_353/li_0_527# FILLER_13_1217/li_0_527# user_to_mprj_in_gates\[17\]/li_18_51#
+ _451_/li_0_n17# FILLER_21_589/li_155_527# user_to_mprj_in_gates\[109\]/li_707_n17#
+ la_buf\[10\]/li_207_51# FILLER_21_62/li_63_n17# PHY_78/li_0_n17# PHY_817/li_0_n17#
+ FILLER_16_88/li_0_527# FILLER_11_2093/li_63_527# FILLER_13_1498/li_0_527# _344_/li_0_n17#
+ PHY_719/li_0_n17# user_to_mprj_oen_buffers\[92\]/li_1259_527# FILLER_25_1502/li_155_527#
+ user_to_mprj_oen_buffers\[50\]/li_891_527# PHY_228/li_0_n17# user_to_mprj_oen_buffers\[114\]/li_247_527#
+ FILLER_25_1922/li_63_n17# PHY_525/li_0_n17# user_to_mprj_oen_buffers\[73\]/li_1351_527#
+ PHY_90/li_0_n17# PHY_343/li_0_n17# mprj_adr_buf\[29\]/li_431_527# FILLER_15_1939/li_155_527#
+ la_buf\[92\]/li_215_311# FILLER_10_2082/li_155_n17# _400_/li_0_527# FILLER_26_1186/li_63_527#
+ FILLER_21_1455/li_63_n17# _334_/li_247_527# _383_/li_0_n17# PHY_231/li_0_n17# la_buf\[66\]/li_63_527#
+ FILLER_22_1771/li_63_n17# user_to_mprj_oen_buffers\[102\]/li_207_51# _598_/li_0_527#
+ PHY_500/li_0_527# PHY_339/li_0_n17# powergood_check/FILLER_2_115/li_100_536# user_to_mprj_in_gates\[36\]/li_707_n17#
+ FILLER_20_1551/li_155_527# la_buf\[47\]/li_0_527# la_buf\[113\]/li_0_n17# ANTENNA_user_to_mprj_in_gates\[17\]_B/li_63_n17#
+ _554_/li_155_n17# user_to_mprj_in_gates\[95\]/li_615_527# _347_/li_0_n17# FILLER_8_793/li_155_n17#
+ user_to_mprj_in_buffers\[112\]/li_404_367# user_to_mprj_in_buffers\[46\]/li_615_n17#
+ ANTENNA__332__A/li_0_527# la_buf\[109\]/li_1259_n17# la_buf\[76\]/li_207_51# FILLER_11_1186/li_63_n17#
+ la_buf\[72\]/li_1075_527# user_to_mprj_in_gates\[16\]/li_155_527# FILLER_11_798/li_0_n17#
+ PHY_855/li_0_n17# user_to_mprj_oen_buffers\[48\]/li_523_n17# la_buf\[50\]/li_891_n17#
+ mprj_stb_buf/li_779_17# powergood_check/FILLER_2_115/li_449_797# user_to_mprj_in_buffers\[8\]/li_404_17#
+ user_to_mprj_oen_buffers\[106\]/li_17_51# FILLER_10_1284/li_155_n17# user_to_mprj_oen_buffers\[38\]/li_1535_n17#
+ _344_/li_155_527# powergood_check/mprj_logic_high_lv/li_179_79# _643_/li_155_527#
+ PHY_490/li_0_527# FILLER_25_815/li_0_n17# user_to_mprj_oen_buffers\[49\]/li_611_17#
+ user_to_mprj_oen_buffers\[116\]/li_891_527# la_buf\[80\]/li_215_311# la_buf\[32\]/li_1351_527#
+ mprj_adr_buf\[22\]/li_17_51# user_to_mprj_in_gates\[25\]/li_155_n17# PHY_303/li_0_527#
+ powergood_check/FILLER_2_163/li_0_797# PHY_851/li_0_527# _521_/li_0_527# FILLER_22_1408/li_0_527#
+ powergood_check/FILLER_0_112/li_65_n17# la_buf\[5\]/li_1259_n17# la_buf\[89\]/li_63_n17#
+ FILLER_13_1431/li_0_527# user_to_mprj_in_gates\[101\]/li_18_51# la_buf\[80\]/li_779_17#
+ user_to_mprj_oen_buffers\[119\]/li_523_n17# FILLER_15_59/li_0_n17# powergood_check/FILLER_1_107/li_65_n17#
+ _414_/li_0_527# la_buf\[39\]/li_215_311# _435_/li_0_n17# user_to_mprj_in_buffers\[7\]/li_236_367#
+ FILLER_14_1724/li_0_n17# user_to_mprj_in_buffers\[100\]/li_404_367# user_to_mprj_in_gates\[78\]/li_523_n17#
+ FILLER_18_1459/li_63_n17# la_buf\[43\]/li_1351_527# user_to_mprj_in_gates\[76\]/li_247_527#
+ PHY_744/li_0_n17# mprj_dat_buf\[0\]/li_17_51# FILLER_11_744/li_155_527# PHY_309/li_0_527#
+ PHY_56/li_0_527# powergood_check/FILLER_2_107/li_257_n17# _576_/li_247_n17# la_buf\[5\]/li_207_51#
+ FILLER_25_1126/li_63_n17# FILLER_5_1209/li_0_527# FILLER_9_420/li_0_n17# FILLER_9_1382/li_63_527#
+ PHY_399/li_0_n17# FILLER_19_1742/li_63_527# FILLER_12_982/li_0_527# powergood_check/FILLER_0_184/li_0_797#
+ ANTENNA__371__A/li_0_n17# mprj_dat_buf\[17\]/li_779_17# user_to_mprj_oen_buffers\[87\]/li_615_527#
+ user_to_mprj_in_gates\[85\]/li_247_n17# FILLER_9_1169/li_63_527# FILLER_23_1728/li_0_527#
+ la_buf\[42\]/li_63_527# _332_/li_0_n17# user_to_mprj_in_gates\[65\]/li_63_n17# ANTENNA_mprj_sel_buf\[2\]_A/li_63_527#
+ user_to_mprj_oen_buffers\[57\]/li_891_n17# la_buf\[12\]/li_891_n17# mprj_dat_buf\[23\]/li_215_311#
+ FILLER_22_1418/li_0_527# PHY_184/li_0_n17# FILLER_19_1417/li_63_527# la_buf\[27\]/li_215_311#
+ _494_/li_247_527# user_to_mprj_in_gates\[118\]/li_523_527# PHY_843/li_0_n17# PHY_449/li_0_527#
+ mprj_dat_buf\[15\]/li_17_51# FILLER_11_1064/li_0_n17# PHY_761/li_0_527# user_to_mprj_in_gates\[66\]/li_523_n17#
+ user_to_mprj_oen_buffers\[81\]/li_17_51# PHY_355/li_0_527# powergood_check/FILLER_1_32/li_115_72#
+ user_to_mprj_in_gates\[64\]/li_247_527# FILLER_19_1446/li_63_n17# ANTENNA_la_buf\[121\]_TE/li_63_n17#
+ user_to_mprj_oen_buffers\[28\]/li_983_527# powergood_check/FILLER_1_220/li_257_n17#
+ la_buf\[93\]/li_17_51# FILLER_19_1742/li_0_527# la_buf\[95\]/li_795_379# FILLER_12_1693/li_0_n17#
+ FILLER_9_829/li_0_527# PHY_442/li_0_527# powergood_check/FILLER_0_88/li_100_536#
+ _407_/li_0_527# user_to_mprj_in_buffers\[7\]/li_339_n17# user_to_mprj_oen_buffers\[53\]/li_207_51#
+ FILLER_18_63/li_0_527# PHY_406/li_0_n17# user_to_mprj_oen_buffers\[53\]/li_0_527#
+ user_to_mprj_in_gates\[33\]/li_0_527# FILLER_12_471/li_0_n17# mprj_dat_buf\[18\]/li_983_527#
+ mprj_adr_buf\[8\]/li_207_51# user_to_mprj_in_gates\[73\]/li_247_n17# powergood_check/FILLER_2_32/li_545_797#
+ ANTENNA__341__A/li_63_527# powergood_check/FILLER_1_260/li_545_n17# la_buf\[30\]/li_615_527#
+ FILLER_22_1522/li_155_n17# _532_/li_0_n17# FILLER_17_507/li_0_527# mprj_dat_buf\[11\]/li_215_311#
+ PHY_492/li_0_527# FILLER_25_1563/li_0_n17# _591_/li_155_527# la_buf\[15\]/li_215_311#
+ user_to_mprj_in_gates\[106\]/li_523_527# la_buf\[126\]/li_1351_527# powergood_check/FILLER_0_88/li_449_797#
+ powergood_check/mprj_logic_high_lv/li_1121_1611# la_buf\[86\]/li_707_527# powergood_check/mprj2_logic_high_hvl/li_0_n17#
+ powergood_check/FILLER_0_184/li_0_n17# powergood_check/FILLER_1_204/li_257_n17#
+ PHY_862/li_0_527# PHY_362/li_0_n17# user_to_mprj_in_gates\[67\]/li_18_51# user_to_mprj_in_gates\[42\]/li_0_n17#
+ mprj_dat_buf\[27\]/li_983_n17# _623_/li_0_527# powergood_check/FILLER_1_244/li_0_797#
+ user_to_mprj_oen_buffers\[116\]/li_215_311# la_buf\[70\]/li_983_n17# user_to_mprj_in_gates\[52\]/li_247_527#
+ la_buf\[15\]/li_207_51# FILLER_25_1422/li_0_n17# FILLER_17_1541/li_0_n17# user_to_mprj_in_gates\[60\]/li_339_n17#
+ user_to_mprj_oen_buffers\[30\]/li_17_51# FILLER_17_2088/li_63_n17# la_buf\[51\]/li_983_527#
+ _382_/li_155_n17# FILLER_10_1188/li_0_n17# FILLER_5_763/li_0_n17# _469_/li_155_527#
+ PHY_356/li_0_527# la_buf\[42\]/li_17_51# powergood_check/FILLER_2_227/li_257_797#
+ PHY_435/li_0_527# user_to_mprj_in_gates\[88\]/li_0_n17# user_to_mprj_oen_buffers\[24\]/li_707_527#
+ user_to_mprj_in_buffers\[90\]/li_51_367# PHY_798/li_0_n17# powergood_check/FILLER_0_168/li_65_797#
+ la_buf\[93\]/li_779_17# mprj_adr_buf\[31\]/li_983_527# mprj_dat_buf\[18\]/li_63_527#
+ mprj_dat_buf\[27\]/li_779_17# user_to_mprj_in_gates\[118\]/li_247_527# PHY_847/li_0_527#
+ PHY_746/li_0_n17# user_to_mprj_in_gates\[33\]/li_523_527# user_to_mprj_oen_buffers\[49\]/li_17_51#
+ user_to_mprj_oen_buffers\[107\]/li_207_51# la_buf\[51\]/li_63_527# _626_/li_0_n17#
+ powergood_check/FILLER_2_24/li_353_n17# _638_/li_0_527# powergood_check/FILLER_2_267/li_545_797#
+ FILLER_23_1978/li_0_527# user_to_mprj_oen_buffers\[48\]/li_215_311# _559_/li_155_n17#
+ FILLER_17_96/li_0_n17# FILLER_14_355/li_0_527# _479_/li_155_527# PHY_247/li_0_n17#
+ PHY_814/li_0_527# powergood_check/FILLER_0_80/li_641_797# FILLER_23_2061/li_155_527#
+ FILLER_7_1774/li_155_n17# user_to_mprj_in_gates\[122\]/li_247_n17# _558_/li_0_n17#
+ mprj_dat_buf\[30\]/li_1167_527# FILLER_23_1774/li_63_527# user_to_mprj_in_gates\[42\]/li_523_n17#
+ mprj_adr_buf\[31\]/li_779_17# FILLER_13_1203/li_0_527# powergood_check/FILLER_2_187/li_353_797#
+ user_to_mprj_oen_buffers\[104\]/li_215_311# FILLER_13_2012/li_0_527# user_to_mprj_in_gates\[16\]/li_18_51#
+ _529_/li_0_527# user_to_mprj_in_gates\[40\]/li_247_527# powergood_check/FILLER_1_228/li_545_n17#
+ _651_/li_247_527# PHY_271/li_0_527# PHY_384/li_0_n17# mprj_dat_buf\[27\]/li_431_527#
+ mprj_dat_buf\[13\]/li_1075_n17# powergood_check/FILLER_0_248/li_257_797# _446_/li_0_n17#
+ _655_/li_247_n17# _593_/li_0_n17# FILLER_9_555/li_155_n17# _349_/li_155_527# _493_/li_0_527#
+ _463_/li_247_n17# user_to_mprj_in_gates\[103\]/li_523_n17# _334_/li_0_n17# user_to_mprj_in_gates\[101\]/li_247_527#
+ FILLER_17_2085/li_63_n17# user_to_mprj_in_gates\[5\]/li_247_527# FILLER_16_2073/li_0_527#
+ PHY_666/li_0_527# la_buf\[83\]/li_207_51# FILLER_9_54/li_155_527# la_buf\[3\]/li_983_527#
+ user_to_mprj_in_buffers\[38\]/li_404_367# _433_/li_0_n17# FILLER_20_1459/li_63_527#
+ PHY_25/li_0_527# _373_/li_0_n17# FILLER_13_1484/li_0_527# FILLER_11_1561/li_63_n17#
+ mprj_adr_buf\[28\]/li_707_527# powergood_check/FILLER_0_200/li_161_797# user_to_mprj_oen_buffers\[36\]/li_215_311#
+ powergood_check/FILLER_1_188/li_641_n17# powergood_check/FILLER_2_259/li_353_n17#
+ _351_/li_155_527# ANTENNA__371__A/li_63_n17# _655_/li_247_527# PHY_741/li_0_n17#
+ FILLER_7_931/li_63_527# user_to_mprj_in_gates\[95\]/li_707_367# user_to_mprj_oen_buffers\[56\]/li_611_17#
+ user_to_mprj_in_gates\[98\]/li_63_n17# FILLER_21_74/li_0_n17# user_to_mprj_in_buffers\[87\]/li_523_n17#
+ powergood_check/FILLER_2_179/li_161_n17# FILLER_21_1989/li_0_527# _424_/li_0_527#
+ FILLER_13_973/li_0_527# la_buf\[19\]/li_431_527# FILLER_10_621/li_0_n17# user_to_mprj_oen_buffers\[105\]/li_17_51#
+ powergood_check/FILLER_0_16/li_0_797# _528_/li_155_527# _441_/li_155_n17# FILLER_20_465/li_63_n17#
+ _467_/li_0_527# user_to_mprj_in_gates\[81\]/li_615_527# user_to_mprj_in_buffers\[69\]/li_523_n17#
+ FILLER_12_978/li_63_n17# user_to_mprj_in_buffers\[26\]/li_404_367# mprj_adr_buf\[21\]/li_17_51#
+ mprj_adr_buf\[9\]/li_1351_527# FILLER_20_1421/li_155_527# user_to_mprj_oen_buffers\[0\]/li_1351_527#
+ FILLER_17_100/li_0_n17# user_to_mprj_in_gates\[123\]/li_63_n17# PHY_805/li_0_527#
+ ANTENNA_user_to_mprj_in_gates\[81\]_B/li_63_527# PHY_347/li_0_n17# user_to_mprj_oen_buffers\[24\]/li_215_311#
+ FILLER_13_1816/li_0_n17# user_to_mprj_in_gates\[100\]/li_18_51# PHY_94/li_0_n17#
+ user_to_mprj_in_gates\[28\]/li_247_527# _530_/li_247_527# PHY_760/li_0_n17# user_to_mprj_in_gates\[83\]/li_707_367#
+ PHY_677/li_0_527# powergood_check/FILLER_1_115/li_737_n17# user_to_mprj_oen_buffers\[24\]/li_1351_527#
+ PHY_737/li_0_n17# la_buf\[110\]/li_983_527# user_to_mprj_oen_buffers\[92\]/li_795_379#
+ user_to_mprj_in_gates\[119\]/li_18_51# user_to_mprj_oen_buffers\[5\]/li_63_527#
+ powergood_check/FILLER_1_236/li_0_797# FILLER_9_1142/li_155_n17# ANTENNA_user_to_mprj_in_gates\[102\]_A/li_63_n17#
+ _408_/li_0_527# _408_/li_155_527# ANTENNA__584__A/li_63_n17# user_to_mprj_oen_buffers\[58\]/li_207_51#
+ _660_/li_0_527# PHY_241/li_0_527# PHY_174/li_0_n17# FILLER_14_532/li_0_527# _559_/li_0_527#
+ PHY_72/li_0_n17# FILLER_25_1004/li_63_n17# powergood_check/mprj_logic_high_hvl/li_161_797#
+ powergood_check/FILLER_2_115/li_449_n17# user_to_mprj_in_buffers\[14\]/li_404_367#
+ PHY_222/li_0_527# powergood_check/mprj2_logic_high_lv/m1_0_51# _447_/li_0_527# FILLER_24_512/li_155_527#
+ PHY_816/li_0_527# user_to_mprj_oen_buffers\[39\]/li_779_17# la_buf\[84\]/li_63_527#
+ _596_/li_155_527# FILLER_25_819/li_0_n17# user_to_mprj_oen_buffers\[12\]/li_215_311#
+ FILLER_16_93/li_63_527# mprj_adr_buf\[28\]/li_1075_n17# _418_/li_0_527# _535_/li_247_n17#
+ user_to_mprj_oen_buffers\[117\]/li_431_n17# user_to_mprj_oen_buffers\[60\]/li_207_51#
+ user_to_mprj_in_gates\[71\]/li_707_367# mprj_dat_buf\[14\]/li_17_51# powergood_check/mprj_logic_high_lv/li_161_1611#
+ mprj_pwrgood/li_155_527# _378_/li_247_n17# powergood_check/FILLER_2_163/li_0_n17#
+ PHY_178/li_0_527# la_buf\[82\]/li_1351_527# la_buf\[86\]/li_611_17# user_to_mprj_oen_buffers\[80\]/li_17_51#
+ user_to_mprj_in_buffers\[102\]/li_615_n17# PHY_448/li_0_n17# user_to_mprj_oen_buffers\[80\]/li_795_379#
+ la_buf\[92\]/li_17_51# FILLER_12_685/li_63_527# _388_/li_0_n17# user_to_mprj_oen_buffers\[41\]/li_779_17#
+ powergood_check/FILLER_2_300/li_161_797# FILLER_20_1893/li_0_n17# ANTENNA__572__A/li_63_n17#
+ user_to_mprj_in_gates\[38\]/li_707_367# _412_/li_0_527# _550_/li_0_527# user_to_mprj_oen_buffers\[99\]/li_17_51#
+ la_buf\[22\]/li_707_n17# FILLER_13_1812/li_63_n17# FILLER_23_332/li_0_n17# mprj_dat_buf\[1\]/li_707_527#
+ PHY_30/li_0_527# powergood_check/FILLER_1_16/li_353_n17# la_buf\[22\]/li_207_51#
+ FILLER_11_1027/li_63_527# FILLER_3_906/li_63_527# powergood_check/FILLER_0_216/li_0_797#
+ PHY_96/li_0_n17# la_buf\[72\]/li_1535_527# PHY_455/li_0_527# la_buf\[50\]/li_1351_n17#
+ user_to_mprj_in_gates\[16\]/li_615_527# FILLER_11_996/li_155_527# PHY_387/li_0_527#
+ FILLER_15_2067/li_0_527# PHY_738/li_0_n17# user_to_mprj_in_gates\[44\]/li_339_n17#
+ mprj_dat_buf\[25\]/li_63_527# PHY_77/li_0_527# user_to_mprj_in_gates\[66\]/li_18_51#
+ user_to_mprj_in_gates\[1\]/li_615_527# FILLER_9_411/li_0_n17# mprj_dat_buf\[29\]/li_247_527#
+ la_buf\[88\]/li_1443_527# mprj_adr_buf\[18\]/li_215_311# user_to_mprj_oen_buffers\[114\]/li_207_51#
+ user_to_mprj_in_gates\[98\]/li_155_n17# powergood_check/FILLER_2_235/li_100_536#
+ user_to_mprj_in_gates\[105\]/li_339_n17# la_buf\[70\]/li_795_379# _566_/li_0_n17#
+ user_to_mprj_in_gates\[120\]/li_707_367# la_buf\[35\]/li_63_n17# FILLER_15_415/li_0_n17#
+ user_to_mprj_in_gates\[25\]/li_615_n17# FILLER_23_1387/li_0_n17# la_buf\[41\]/li_17_51#
+ user_to_mprj_oen_buffers\[64\]/li_1443_n17# FILLER_11_423/li_63_n17# user_to_mprj_in_gates\[23\]/li_339_527#
+ PHY_46/li_0_527# FILLER_27_81/li_0_n17# la_buf\[88\]/li_207_51# FILLER_16_1939/li_63_527#
+ FILLER_13_202/li_63_n17# PHY_852/li_0_n17# PHY_747/li_0_527# user_to_mprj_in_gates\[79\]/li_431_n17#
+ user_to_mprj_oen_buffers\[48\]/li_17_51# powergood_check/FILLER_2_235/li_449_797#
+ powergood_check/FILLER_1_172/li_0_797# user_to_mprj_in_gates\[77\]/li_155_527# user_to_mprj_oen_buffers\[38\]/li_523_n17#
+ PHY_324/li_0_527# powergood_check/FILLER_1_0/li_100_536# PHY_71/li_0_527# mprj_sel_buf\[2\]/li_247_527#
+ FILLER_15_1510/li_0_n17# PHY_482/li_0_527# mprj_dat_buf\[0\]/li_1443_n17# la_buf\[69\]/li_779_17#
+ powergood_check/FILLER_2_155/li_257_797# FILLER_13_1199/li_63_n17# mprj_dat_buf\[19\]/li_523_n17#
+ PHY_398/li_0_527# powergood_check/FILLER_2_32/li_545_n17# la_buf\[90\]/li_207_51#
+ PHY_246/li_0_527# ANTENNA_la_buf\[126\]_A/li_63_527# powergood_check/FILLER_0_256/li_100_536#
+ _548_/li_0_n17# ANTENNA_user_to_mprj_oen_buffers\[45\]_A/li_63_n17# la_buf\[11\]/li_0_527#
+ user_to_mprj_in_gates\[15\]/li_18_51# user_to_mprj_oen_buffers\[17\]/li_1351_527#
+ _535_/li_0_527# user_to_mprj_in_gates\[86\]/li_155_n17# FILLER_13_1931/li_0_n17#
+ FILLER_25_934/li_0_n17# PHY_302/li_0_527# user_to_mprj_oen_buffers\[42\]/li_63_527#
+ PHY_377/li_0_n17# _470_/li_0_n17# PHY_157/li_0_527# _446_/li_155_n17# user_to_mprj_in_gates\[85\]/li_707_n17#
+ powergood_check/FILLER_2_195/li_545_797# _587_/li_0_n17# _600_/li_0_527# mprj_adr_buf\[0\]/li_215_311#
+ la_buf\[113\]/li_615_527# user_to_mprj_in_gates\[119\]/li_431_527# _657_/li_155_n17#
+ powergood_check/FILLER_1_244/li_0_n17# user_to_mprj_oen_buffers\[52\]/li_1075_527#
+ user_to_mprj_oen_buffers\[63\]/li_611_17# FILLER_9_1138/li_0_n17# powergood_check/FILLER_0_256/li_449_797#
+ FILLER_26_1099/li_155_527# la_buf\[6\]/li_1259_527# FILLER_19_1471/li_155_527# FILLER_13_855/li_155_n17#
+ FILLER_17_1713/li_0_n17# mprj_dat_buf\[27\]/li_891_527# powergood_check/FILLER_1_156/li_545_n17#
+ powergood_check/FILLER_2_227/li_257_n17# la_buf\[50\]/li_247_527# powergood_check/FILLER_0_176/li_257_797#
+ la_buf\[95\]/li_983_527# _535_/li_155_527# user_to_mprj_in_gates\[107\]/li_0_527#
+ FILLER_0_288/li_63_527# FILLER_18_2110/li_155_n17# FILLER_16_1331/li_155_527# PHY_504/li_0_527#
+ FILLER_13_752/li_63_527# powergood_check/FILLER_2_267/li_545_n17# FILLER_12_986/li_0_n17#
+ user_to_mprj_in_gates\[74\]/li_155_n17# mprj_adr_buf\[24\]/li_247_527# _342_/li_0_527#
+ PHY_818/li_0_527# FILLER_20_567/li_63_n17# user_to_mprj_in_buffers\[99\]/li_404_17#
+ powergood_check/FILLER_1_32/li_0_n17# powergood_check/FILLER_0_16/li_545_797# PHY_257/li_0_n17#
+ user_to_mprj_in_gates\[73\]/li_707_n17# user_to_mprj_oen_buffers\[104\]/li_17_51#
+ PHY_31/li_0_527# la_buf\[88\]/li_215_311# FILLER_25_1180/li_155_n17# powergood_check/FILLER_2_187/li_353_n17#
+ user_to_mprj_in_gates\[107\]/li_431_527# mprj_dat_buf\[27\]/li_707_527# FILLER_12_1106/li_155_n17#
+ la_buf\[102\]/li_1259_527# user_to_mprj_in_gates\[55\]/li_431_n17# powergood_check/FILLER_2_163/li_115_72#
+ FILLER_26_981/li_0_527# powergood_check/FILLER_1_300/li_65_n17# la_buf\[0\]/li_779_17#
+ user_to_mprj_in_gates\[53\]/li_155_527# user_to_mprj_oen_buffers\[117\]/li_611_17#
+ mprj_adr_buf\[20\]/li_17_51# mprj_sel_buf\[1\]/li_523_n17# user_to_mprj_oen_buffers\[13\]/li_431_n17#
+ powergood_check/FILLER_0_0/li_353_797# user_to_mprj_in_gates\[60\]/li_0_n17# user_to_mprj_oen_buffers\[83\]/li_247_527#
+ user_to_mprj_oen_buffers\[119\]/li_247_n17# powergood_check/FILLER_1_8/li_115_72#
+ _415_/li_155_527# user_to_mprj_in_buffers\[108\]/li_404_367# mprj_adr_buf\[17\]/li_1351_527#
+ user_to_mprj_oen_buffers\[65\]/li_207_51# FILLER_5_743/li_0_527# user_to_mprj_in_gates\[116\]/li_431_n17#
+ FILLER_25_1200/li_155_n17# FILLER_21_1331/li_155_527# PHY_858/li_0_n17# la_buf\[4\]/li_523_n17#
+ PHY_21/li_0_527# FILLER_13_911/li_63_n17# user_to_mprj_in_gates\[10\]/li_615_527#
+ user_to_mprj_in_gates\[118\]/li_18_51# PHY_865/li_0_n17# FILLER_13_883/li_63_n17#
+ _516_/li_0_527# _505_/li_155_n17# la_buf\[76\]/li_215_311# user_to_mprj_in_gates\[9\]/li_18_51#
+ user_to_mprj_in_gates\[123\]/li_155_n17# PHY_780/li_0_n17# PHY_782/li_0_n17# la_buf\[27\]/li_207_51#
+ PHY_728/li_0_n17# user_to_mprj_oen_buffers\[124\]/li_983_n17# PHY_186/li_0_527#
+ la_buf\[109\]/li_17_51# FILLER_19_2061/li_155_527# FILLER_17_530/li_155_527# user_to_mprj_in_gates\[122\]/li_707_n17#
+ powergood_check/mprj_logic_high_lv/li_179_1349# _437_/li_0_527# FILLER_19_1573/li_63_527#
+ FILLER_22_1909/li_155_n17# FILLER_13_1017/li_63_527# FILLER_12_748/li_63_527# FILLER_9_375/li_63_n17#
+ FILLER_17_1957/li_0_n17# la_buf\[109\]/li_0_527# la_buf\[59\]/li_891_n17# PHY_623/li_0_527#
+ user_to_mprj_in_gates\[88\]/li_431_527# mprj_dat_buf\[13\]/li_17_51# FILLER_24_612/li_155_527#
+ FILLER_11_992/li_0_527# powergood_check/FILLER_0_216/li_641_797# user_to_mprj_oen_buffers\[119\]/li_207_51#
+ user_to_mprj_in_gates\[94\]/li_523_527# la_buf\[19\]/li_0_527# _443_/li_0_n17# la_buf\[99\]/li_0_n17#
+ ANTENNA_la_buf\[5\]_TE/li_63_n17# user_to_mprj_in_gates\[50\]/li_155_n17# powergood_check/FILLER_0_80/li_161_797#
+ _507_/li_247_n17# FILLER_5_1196/li_0_527# _483_/li_155_527# la_buf\[91\]/li_17_51#
+ FILLER_19_1587/li_63_527# PHY_434/li_0_527# user_to_mprj_in_gates\[32\]/li_0_527#
+ la_buf\[64\]/li_215_311# powergood_check/mprj_logic_high_lv/li_756_683# la_buf\[10\]/li_779_17#
+ la_buf\[84\]/li_0_n17# user_to_mprj_oen_buffers\[57\]/li_1443_527# user_to_mprj_in_gates\[111\]/li_155_n17#
+ FILLER_19_1475/li_63_527# PHY_332/li_0_527# user_to_mprj_oen_buffers\[98\]/li_17_51#
+ la_buf\[1\]/li_63_527# PHY_803/li_0_n17# la_buf\[57\]/li_1351_527# FILLER_24_602/li_0_527#
+ FILLER_23_1678/li_0_527# user_to_mprj_oen_buffers\[121\]/li_207_51# user_to_mprj_oen_buffers\[1\]/li_215_311#
+ powergood_check/FILLER_0_8/li_641_797# mprj_dat_buf\[19\]/li_215_311# _573_/li_0_527#
+ _561_/li_247_527# powergood_check/FILLER_2_235/li_65_n17# _533_/li_0_527# _573_/li_155_n17#
+ FILLER_11_1030/li_0_n17# PHY_260/li_0_n17# powergood_check/FILLER_1_24/li_545_n17#
+ powergood_check/FILLER_0_272/li_0_n17# PHY_736/li_0_n17# FILLER_12_593/li_155_527#
+ _595_/li_155_527# powergood_check/mprj_logic_high_hvl/li_161_n17# _454_/li_0_n17#
+ la_buf\[95\]/li_207_51# mprj_adr_buf\[2\]/li_779_17# PHY_812/li_0_527# user_to_mprj_in_gates\[65\]/li_18_51#
+ user_to_mprj_oen_buffers\[18\]/li_247_527# la_buf\[58\]/li_707_527# user_to_mprj_in_gates\[82\]/li_523_527#
+ powergood_check/FILLER_1_188/li_161_n17# user_to_mprj_oen_buffers\[47\]/li_63_527#
+ user_to_mprj_in_buffers\[99\]/li_404_367# user_to_mprj_in_gates\[95\]/li_0_n17#
+ PHY_259/li_0_n17# FILLER_7_1131/li_0_527# _363_/li_155_527# user_to_mprj_oen_buffers\[82\]/li_891_n17#
+ PHY_365/li_0_n17# user_to_mprj_oen_buffers\[97\]/li_215_311# la_buf\[40\]/li_17_51#
+ la_buf\[52\]/li_215_311# FILLER_17_1512/li_155_n17# powergood_check/FILLER_0_16/li_115_72#
+ FILLER_0_288/li_155_527# user_to_mprj_in_gates\[69\]/li_247_n17# mprj_dat_buf\[22\]/li_615_527#
+ powergood_check/FILLER_0_160/li_0_797# FILLER_21_66/li_155_527# la_buf\[26\]/li_615_527#
+ FILLER_25_1291/li_0_n17# user_to_mprj_in_gates\[91\]/li_523_n17# PHY_417/li_0_n17#
+ FILLER_21_1402/li_63_527# FILLER_23_2061/li_155_n17# user_to_mprj_oen_buffers\[47\]/li_17_51#
+ _463_/li_0_n17# FILLER_25_953/li_0_n17# mprj_adr_buf\[29\]/li_1259_527# powergood_check/FILLER_2_300/li_161_n17#
+ FILLER_16_1825/li_0_527# FILLER_11_1713/li_0_n17# powergood_check/FILLER_1_268/li_115_72#
+ powergood_check/FILLER_2_163/li_100_536# user_to_mprj_in_buffers\[123\]/li_615_n17#
+ la_buf\[59\]/li_17_51# FILLER_22_1522/li_0_527# FILLER_25_746/li_0_n17# FILLER_17_353/li_63_n17#
+ user_to_mprj_in_buffers\[40\]/li_404_17# FILLER_23_1778/li_0_527# powergood_check/FILLER_1_156/li_115_72#
+ user_to_mprj_oen_buffers\[70\]/li_611_17# FILLER_10_1264/li_155_n17# user_to_mprj_in_gates\[48\]/li_247_527#
+ PHY_96/li_0_527# FILLER_28_43/li_0_527# FILLER_11_933/li_0_527# FILLER_15_365/li_0_527#
+ user_to_mprj_in_gates\[14\]/li_18_51# FILLER_5_1031/li_155_527# PHY_386/li_0_527#
+ powergood_check/FILLER_2_163/li_449_797# user_to_mprj_in_gates\[33\]/li_155_n17#
+ la_buf\[89\]/li_431_n17# user_to_mprj_in_gates\[109\]/li_247_527# powergood_check/FILLER_1_115/li_257_n17#
+ _542_/li_155_527# FILLER_22_1440/li_0_527# la_buf\[11\]/li_63_527# user_to_mprj_oen_buffers\[85\]/li_215_311#
+ FILLER_14_1784/li_0_527# FILLER_0_1326/li_63_527# user_to_mprj_in_buffers\[12\]/li_615_n17#
+ la_buf\[40\]/li_215_311# PHY_824/li_0_527# user_to_mprj_in_gates\[57\]/li_247_n17#
+ la_buf\[14\]/li_615_527# user_to_mprj_oen_buffers\[22\]/li_523_n17# FILLER_12_697/li_0_n17#
+ la_buf\[5\]/li_779_17# la_buf\[124\]/li_215_311# FILLER_13_911/li_0_n17# user_to_mprj_in_gates\[84\]/li_63_n17#
+ FILLER_9_1169/li_155_527# la_buf\[59\]/li_707_n17# powergood_check/FILLER_0_184/li_100_536#
+ la_buf\[4\]/li_215_311# _353_/li_0_n17# PHY_856/li_0_n17# _333_/li_155_n17# user_to_mprj_in_gates\[118\]/li_247_n17#
+ ANTENNA_user_to_mprj_in_gates\[88\]_B/li_63_n17# PHY_161/li_0_527# _634_/li_0_n17#
+ user_to_mprj_in_buffers\[41\]/li_51_367# FILLER_13_703/li_63_527# powergood_check/mprj2_logic_high_lv/li_1025_1611#
+ FILLER_13_1676/li_0_527# PHY_815/li_0_n17# user_to_mprj_in_gates\[36\]/li_247_527#
+ la_buf\[14\]/li_1351_n17# user_to_mprj_oen_buffers\[5\]/li_431_527# PHY_75/li_0_527#
+ powergood_check/FILLER_2_235/li_449_n17# mprj_adr_buf\[23\]/li_1351_527# _392_/li_0_n17#
+ powergood_check/FILLER_1_172/li_0_n17# mprj_dat_buf\[2\]/li_207_51# user_to_mprj_in_buffers\[46\]/li_51_17#
+ la_buf\[67\]/li_795_379# FILLER_14_452/li_63_n17# powergood_check/FILLER_0_184/li_449_797#
+ user_to_mprj_oen_buffers\[124\]/li_611_17# user_to_mprj_in_buffers\[75\]/li_404_367#
+ PHY_823/li_0_n17# la_buf\[77\]/li_63_527# la_buf\[77\]/li_431_n17# FILLER_25_1269/li_155_n17#
+ powergood_check/FILLER_2_155/li_257_n17# FILLER_25_1204/li_155_527# FILLER_19_48/li_63_527#
+ user_to_mprj_oen_buffers\[72\]/li_207_51# user_to_mprj_oen_buffers\[73\]/li_215_311#
+ ANTENNA_user_to_mprj_in_gates\[106\]_A/li_63_527# user_to_mprj_in_gates\[3\]/li_615_527#
+ user_to_mprj_oen_buffers\[103\]/li_17_51# FILLER_25_1749/li_63_527# FILLER_19_407/li_0_n17#
+ powergood_check/mprj2_logic_high_lv/li_353_1611# user_to_mprj_in_gates\[45\]/li_247_n17#
+ FILLER_16_1585/li_0_527# user_to_mprj_oen_buffers\[47\]/li_615_527# la_buf\[98\]/li_611_17#
+ mprj_adr_buf\[8\]/li_523_n17# powergood_check/FILLER_1_0/li_449_n17# PHY_795/li_0_527#
+ la_buf\[112\]/li_215_311# powergood_check/FILLER_0_32/li_0_797# la_buf\[66\]/li_1167_n17#
+ user_to_mprj_oen_buffers\[53\]/li_779_17# _648_/li_0_n17# powergood_check/FILLER_2_195/li_545_n17#
+ FILLER_20_2110/li_63_527# FILLER_17_342/li_0_527# FILLER_23_1896/li_0_n17# user_to_mprj_in_gates\[116\]/li_247_n17#
+ mprj_dat_buf\[0\]/li_215_311# FILLER_13_1115/li_0_n17# powergood_check/FILLER_1_260/li_65_n17#
+ FILLER_28_51/li_155_527# user_to_mprj_in_gates\[24\]/li_247_527# FILLER_22_1929/li_0_527#
+ la_buf\[34\]/li_207_51# _558_/li_247_n17# powergood_check/FILLER_1_228/li_65_n17#
+ PHY_217/li_0_527# powergood_check/FILLER_1_244/li_100_536# ANTENNA__362__A/li_63_527#
+ ANTENNA__626__A/li_63_n17# FILLER_9_563/li_0_n17# la_buf\[65\]/li_431_n17# user_to_mprj_in_gates\[117\]/li_18_51#
+ PHY_284/li_0_527# FILLER_18_1805/li_0_527# user_to_mprj_oen_buffers\[61\]/li_215_311#
+ user_to_mprj_in_gates\[77\]/li_615_527# FILLER_21_66/li_0_n17# ANTENNA__657__A/li_0_527#
+ FILLER_12_693/li_0_n17# _640_/li_0_527# user_to_mprj_in_gates\[8\]/li_18_51# mprj_dat_buf\[6\]/li_1535_527#
+ FILLER_9_1352/li_63_527# FILLER_18_1529/li_155_527# user_to_mprj_oen_buffers\[126\]/li_207_51#
+ la_buf\[100\]/li_215_311# la_buf\[46\]/li_0_527# ANTENNA_user_to_mprj_in_gates\[31\]_B/li_63_527#
+ la_buf\[108\]/li_17_51# _578_/li_155_n17# FILLER_9_534/li_0_n17# la_buf\[50\]/li_0_n17#
+ la_buf\[44\]/li_431_527# _490_/li_155_527# user_to_mprj_in_gates\[79\]/li_707_367#
+ PHY_226/li_0_n17# user_to_mprj_in_gates\[86\]/li_615_n17# FILLER_17_543/li_155_n17#
+ FILLER_25_945/li_155_n17# user_to_mprj_oen_buffers\[107\]/li_779_17# PHY_842/li_0_527#
+ user_to_mprj_in_gates\[12\]/li_247_527# PHY_44/li_0_n17# mprj_dat_buf\[12\]/li_17_51#
+ _480_/li_247_527# _541_/li_0_527# _354_/li_0_527# _368_/li_155_527# powergood_check/FILLER_0_104/li_353_797#
+ PHY_866/li_0_527# _580_/li_155_n17# la_buf\[90\]/li_17_51# PHY_333/li_0_527# PHY_260/li_0_527#
+ la_buf\[7\]/li_795_379# PHY_293/li_0_n17# la_buf\[50\]/li_707_527# FILLER_8_949/li_0_527#
+ user_to_mprj_oen_buffers\[97\]/li_17_51# user_to_mprj_oen_buffers\[54\]/li_63_527#
+ user_to_mprj_oen_buffers\[110\]/li_1167_n17# PHY_833/li_0_527# _570_/li_0_n17# FILLER_19_1916/li_0_527#
+ FILLER_17_1520/li_0_527# powergood_check/FILLER_1_236/li_257_n17# _370_/li_155_527#
+ PHY_410/li_0_527# FILLER_19_109/li_63_n17# la_buf\[32\]/li_431_527# _539_/li_0_527#
+ la_buf\[124\]/li_891_n17# user_to_mprj_in_buffers\[45\]/li_404_17# FILLER_27_868/li_0_n17#
+ la_buf\[83\]/li_779_17# user_to_mprj_in_gates\[67\]/li_707_367# user_to_mprj_oen_buffers\[124\]/li_523_n17#
+ PHY_295/li_0_n17# user_to_mprj_in_gates\[74\]/li_615_n17# mprj_adr_buf\[24\]/li_707_527#
+ FILLER_25_899/li_63_n17# user_to_mprj_in_gates\[72\]/li_339_527# la_buf\[95\]/li_1167_n17#
+ user_to_mprj_in_gates\[82\]/li_0_527# mprj_adr_buf\[16\]/li_1351_527# PHY_800/li_0_527#
+ FILLER_17_2088/li_155_n17# user_to_mprj_in_gates\[64\]/li_18_51# FILLER_11_992/li_0_n17#
+ PHY_341/li_0_527# powergood_check/FILLER_1_32/li_737_n17# powergood_check/FILLER_0_200/li_65_797#
+ user_to_mprj_oen_buffers\[86\]/li_431_n17# mprj_sel_buf\[3\]/li_707_527# PHY_314/li_0_n17#
+ la_buf\[41\]/li_431_n17# FILLER_19_95/li_0_527# _660_/li_247_n17# mprj_clk_buf/li_215_311#
+ FILLER_13_1812/li_0_n17# powergood_check/FILLER_0_200/li_0_n17# user_to_mprj_oen_buffers\[11\]/li_207_51#
+ user_to_mprj_oen_buffers\[59\]/li_1075_n17# FILLER_9_501/li_63_527# la_buf\[37\]/li_779_17#
+ FILLER_25_823/li_155_n17# la_buf\[3\]/li_1443_527# user_to_mprj_in_buffers\[61\]/li_523_527#
+ mprj_dat_buf\[3\]/li_795_379# user_to_mprj_oen_buffers\[56\]/li_891_n17# la_buf\[84\]/li_983_n17#
+ user_to_mprj_oen_buffers\[46\]/li_17_51# _338_/li_155_n17# powergood_check/FILLER_1_107/li_115_72#
+ FILLER_23_1670/li_0_527# PHY_380/li_0_527# FILLER_10_804/li_63_527# _538_/li_247_n17#
+ user_to_mprj_in_gates\[55\]/li_707_367# la_buf\[7\]/li_707_527# la_buf\[58\]/li_17_51#
+ _371_/li_0_527# powergood_check/FILLER_2_0/li_545_797# PHY_340/li_0_527# user_to_mprj_oen_buffers\[7\]/li_247_527#
+ PHY_69/li_0_n17# mprj_stb_buf/li_431_n17# PHY_513/li_0_n17# _573_/li_247_n17# FILLER_12_890/li_155_527#
+ mprj_dat_buf\[7\]/li_207_51# FILLER_21_1570/li_0_n17# user_to_mprj_in_buffers\[96\]/li_51_17#
+ user_to_mprj_in_gates\[31\]/li_0_527# PHY_160/li_0_527# _386_/li_247_527# _357_/li_247_n17#
+ user_to_mprj_in_gates\[91\]/li_63_n17# user_to_mprj_oen_buffers\[24\]/li_63_n17#
+ user_to_mprj_in_gates\[13\]/li_18_51# user_to_mprj_in_gates\[116\]/li_707_367# FILLER_10_1170/li_63_n17#
+ powergood_check/mprj2_logic_high_hvl/li_65_797# user_to_mprj_in_gates\[123\]/li_615_n17#
+ mprj_adr_buf\[8\]/li_215_311# user_to_mprj_oen_buffers\[74\]/li_431_n17# FILLER_11_680/li_0_527#
+ user_to_mprj_oen_buffers\[77\]/li_207_51# PHY_36/li_0_n17# FILLER_13_345/li_63_527#
+ user_to_mprj_in_gates\[121\]/li_431_527# _567_/li_0_n17# FILLER_19_1577/li_155_n17#
+ _395_/li_0_527# powergood_check/FILLER_0_96/li_641_797# FILLER_23_1520/li_63_527#
+ PHY_901/li_0_527# FILLER_15_1437/li_0_527# PHY_335/li_0_527# PHY_908/li_0_n17# PHY_675/li_0_527#
+ _343_/li_0_n17# FILLER_13_1574/li_155_n17# _553_/li_0_n17# FILLER_25_1315/li_0_n17#
+ user_to_mprj_in_gates\[43\]/li_707_367# PHY_693/li_0_527# user_to_mprj_in_gates\[50\]/li_615_n17#
+ PHY_185/li_0_527# PHY_713/li_0_n17# FILLER_11_1682/li_63_n17# FILLER_23_1896/li_63_527#
+ la_buf\[39\]/li_207_51# la_buf\[54\]/li_1075_527# user_to_mprj_oen_buffers\[52\]/li_795_379#
+ FILLER_11_1717/li_0_n17# user_to_mprj_oen_buffers\[7\]/li_1167_527# _382_/li_0_n17#
+ user_to_mprj_in_gates\[104\]/li_707_367# la_buf\[102\]/li_207_51# user_to_mprj_oen_buffers\[45\]/li_1535_527#
+ FILLER_21_467/li_0_527# user_to_mprj_oen_buffers\[60\]/li_779_17# user_to_mprj_in_gates\[111\]/li_615_n17#
+ ANTENNA_user_to_mprj_in_gates\[46\]_A/li_63_527# user_to_mprj_oen_buffers\[62\]/li_431_n17#
+ la_buf\[70\]/li_0_n17# FILLER_13_883/li_63_527# powergood_check/FILLER_0_216/li_161_797#
+ PHY_258/li_0_527# mprj_adr_buf\[21\]/li_63_n17# PHY_300/li_0_n17# la_buf\[120\]/li_247_n17#
+ FILLER_28_40/li_63_n17# user_to_mprj_oen_buffers\[102\]/li_17_51# FILLER_13_206/li_0_527#
+ _536_/li_0_527# la_buf\[41\]/li_207_51# PHY_859/li_0_n17# FILLER_14_1662/li_0_n17#
+ mprj_adr_buf\[31\]/li_215_311# powergood_check/FILLER_2_163/li_449_n17# user_to_mprj_in_gates\[121\]/li_339_n17#
+ FILLER_14_2144/li_63_527# PHY_84/li_0_527# _421_/li_0_527# PHY_793/li_0_527# _652_/li_0_527#
+ PHY_257/li_0_527# user_to_mprj_in_gates\[31\]/li_707_367# ANTENNA_user_to_mprj_in_gates\[99\]_B/li_63_527#
+ powergood_check/FILLER_0_8/li_161_797# FILLER_12_1186/li_155_n17# user_to_mprj_oen_buffers\[52\]/li_247_527#
+ FILLER_22_1444/li_63_527# user_to_mprj_in_gates\[92\]/li_431_n17# user_to_mprj_in_gates\[69\]/li_707_n17#
+ user_to_mprj_in_gates\[90\]/li_155_527# la_buf\[69\]/li_891_n17# _585_/li_155_n17#
+ FILLER_23_1425/li_155_n17# user_to_mprj_oen_buffers\[61\]/li_1167_527# user_to_mprj_in_gates\[116\]/li_18_51#
+ user_to_mprj_in_gates\[1\]/li_339_527# PHY_746/li_0_527# FILLER_9_586/li_63_527#
+ user_to_mprj_oen_buffers\[16\]/li_0_n17# _618_/li_0_n17# PHY_91/li_0_n17# user_to_mprj_oen_buffers\[66\]/li_0_527#
+ user_to_mprj_in_gates\[49\]/li_155_527# user_to_mprj_in_gates\[7\]/li_18_51# FILLER_12_1482/li_155_527#
+ mprj_dat_buf\[30\]/li_247_527# FILLER_24_1656/li_0_527# PHY_826/li_0_n17# la_buf\[89\]/li_1351_527#
+ PHY_404/li_0_n17# user_to_mprj_in_gates\[71\]/li_431_527# FILLER_11_1717/li_63_527#
+ PHY_351/li_0_n17# la_buf\[107\]/li_17_51# ANTENNA__477__A/li_63_527# FILLER_9_1230/li_63_527#
+ powergood_check/FILLER_1_172/li_100_536# _610_/li_247_527# FILLER_16_355/li_0_527#
+ PHY_865/li_0_527# user_to_mprj_oen_buffers\[118\]/li_1351_527# PHY_376/li_0_527#
+ _456_/li_0_527# mprj_dat_buf\[11\]/li_17_51# la_buf\[43\]/li_247_n17# user_to_mprj_in_gates\[57\]/li_707_n17#
+ FILLER_23_1937/li_0_n17# _344_/li_0_527# FILLER_9_394/li_63_n17# user_to_mprj_oen_buffers\[60\]/li_1443_n17#
+ powergood_check/FILLER_0_240/li_115_72# FILLER_5_865/li_0_527# FILLER_25_1827/li_63_527#
+ user_to_mprj_oen_buffers\[16\]/li_207_51# user_to_mprj_oen_buffers\[82\]/li_611_17#
+ user_to_mprj_in_buffers\[65\]/li_615_n17# user_to_mprj_oen_buffers\[91\]/li_1351_n17#
+ user_to_mprj_in_buffers\[61\]/li_339_527# user_to_mprj_oen_buffers\[9\]/li_215_311#
+ powergood_check/FILLER_0_112/li_545_797# user_to_mprj_oen_buffers\[90\]/li_1535_n17#
+ FILLER_21_1558/li_63_n17# user_to_mprj_in_gates\[37\]/li_155_527# powergood_check/FILLER_2_16/li_100_536#
+ user_to_mprj_in_gates\[118\]/li_707_n17# la_buf\[24\]/li_523_n17# _377_/li_247_527#
+ FILLER_9_575/li_0_n17# user_to_mprj_oen_buffers\[96\]/li_17_51# FILLER_21_1506/li_0_527#
+ user_to_mprj_in_gates\[70\]/li_247_527# FILLER_14_495/li_0_527# FILLER_22_2092/li_155_n17#
+ FILLER_19_1778/li_63_n17# _596_/li_247_527# FILLER_26_1835/li_0_527# user_to_mprj_in_buffers\[2\]/li_523_n17#
+ powergood_check/FILLER_2_16/li_449_797# powergood_check/FILLER_0_248/li_65_n17#
+ user_to_mprj_in_gates\[96\]/li_63_n17# PHY_306/li_0_n17# user_to_mprj_in_gates\[63\]/li_18_51#
+ FILLER_0_91/li_63_527# user_to_mprj_in_gates\[45\]/li_707_n17# FILLER_16_1589/li_63_527#
+ _345_/li_155_n17# ANTENNA_user_to_mprj_in_gates\[63\]_A/li_63_n17# _644_/li_155_n17#
+ powergood_check/FILLER_1_164/li_257_n17# FILLER_24_1494/li_155_n17# FILLER_25_815/li_0_527#
+ la_buf\[7\]/li_1259_527# _577_/li_247_n17# FILLER_15_506/li_0_527# user_to_mprj_oen_buffers\[57\]/li_523_n17#
+ la_buf\[9\]/li_891_n17# mprj_adr_buf\[13\]/li_207_51# FILLER_22_1522/li_0_n17# la_buf\[6\]/li_247_527#
+ FILLER_21_1662/li_0_n17# la_buf\[89\]/li_63_527# mprj_rstn_buf/li_1535_527# user_to_mprj_oen_buffers\[45\]/li_17_51#
+ la_buf\[96\]/li_983_527# la_buf\[30\]/li_1443_n17# FILLER_13_620/li_155_n17# user_to_mprj_oen_buffers\[84\]/li_207_51#
+ la_buf\[57\]/li_17_51# powergood_check/FILLER_0_24/li_257_797# FILLER_13_895/li_0_527#
+ FILLER_13_1574/li_63_n17# PHY_837/li_0_527# la_buf\[46\]/li_1351_n17# user_to_mprj_in_gates\[34\]/li_155_n17#
+ PHY_185/li_0_n17# FILLER_13_659/li_63_527# la_buf\[107\]/li_207_51# FILLER_12_1796/li_0_n17#
+ _355_/li_0_n17# _370_/li_0_527# user_to_mprj_oen_buffers\[88\]/li_1351_527# FILLER_12_1547/li_0_n17#
+ FILLER_18_1700/li_0_527# user_to_mprj_in_gates\[12\]/li_18_51# FILLER_11_1706/li_63_n17#
+ la_buf\[48\]/li_215_311# PHY_399/li_0_527# PHY_826/li_0_527# mprj_dat_buf\[18\]/li_615_527#
+ user_to_mprj_oen_buffers\[82\]/li_1167_n17# FILLER_25_945/li_0_n17# PHY_441/li_0_527#
+ la_buf\[46\]/li_207_51# _557_/li_0_n17# user_to_mprj_in_gates\[49\]/li_0_527# la_buf\[121\]/li_1443_527#
+ mprj_dat_buf\[6\]/li_1351_n17# FILLER_14_1529/li_0_527# powergood_check/mprj2_logic_high_lv/li_161_797#
+ la_buf\[84\]/li_983_527# PHY_184/li_0_527# FILLER_13_1096/li_0_527# _596_/li_0_n17#
+ powergood_check/FILLER_2_203/li_353_797# FILLER_13_1025/li_0_n17# la_buf\[27\]/li_779_17#
+ FILLER_13_837/li_0_527# la_buf\[67\]/li_891_527# FILLER_23_1915/li_0_527# powergood_check/FILLER_0_24/li_65_797#
+ user_to_mprj_oen_buffers\[52\]/li_247_n17# _372_/li_0_n17# la_buf\[59\]/li_0_n17#
+ powergood_check/FILLER_2_243/li_641_797# user_to_mprj_oen_buffers\[1\]/li_63_n17#
+ powergood_check/FILLER_2_0/li_545_n17# la_buf\[116\]/li_523_n17# powergood_check/FILLER_1_62/li_353_797#
+ user_to_mprj_oen_buffers\[56\]/li_1351_n17# la_buf\[36\]/li_215_311# FILLER_24_1421/li_63_527#
+ user_to_mprj_oen_buffers\[88\]/li_1259_n17# mprj_adr_buf\[10\]/li_795_379# la_buf\[122\]/li_63_n17#
+ FILLER_16_1711/li_0_n17# FILLER_12_471/li_0_527# PHY_263/li_0_n17# FILLER_14_1500/li_0_527#
+ FILLER_17_1405/li_0_527# user_to_mprj_oen_buffers\[101\]/li_17_51# FILLER_26_939/li_0_527#
+ ANTENNA_mprj_stb_buf_A/li_63_527# powergood_check/FILLER_1_204/li_641_n17# FILLER_13_752/li_155_527#
+ FILLER_24_1522/li_155_527# powergood_check/mprj2_logic_high_hvl/li_65_n17# powergood_check/FILLER_0_224/li_353_797#
+ user_to_mprj_oen_buffers\[45\]/li_891_527# FILLER_20_567/li_0_n17# la_buf\[72\]/li_983_527#
+ mprj_dat_buf\[8\]/li_215_311# user_to_mprj_in_gates\[39\]/li_339_n17# powergood_check/FILLER_1_8/li_257_n17#
+ FILLER_26_685/li_0_527# FILLER_10_1184/li_0_n17# _571_/li_0_527# FILLER_13_2051/li_0_527#
+ FILLER_15_361/li_63_n17# powergood_check/FILLER_0_96/li_641_n17# FILLER_13_1648/li_63_527#
+ FILLER_13_699/li_63_527# user_to_mprj_in_gates\[54\]/li_523_527# PHY_39/li_0_527#
+ FILLER_25_554/li_63_527# user_to_mprj_oen_buffers\[80\]/li_63_527# PHY_265/li_0_n17#
+ FILLER_23_489/li_63_n17# FILLER_12_1543/li_63_n17# PHY_497/li_0_527# powergood_check/FILLER_0_264/li_641_797#
+ user_to_mprj_in_gates\[35\]/li_63_n17# FILLER_7_1031/li_63_n17# mprj_dat_buf\[20\]/li_215_311#
+ user_to_mprj_oen_buffers\[69\]/li_215_311# ANTENNA_user_to_mprj_in_gates\[81\]_A/li_63_527#
+ la_buf\[95\]/li_779_17# la_buf\[24\]/li_215_311# user_to_mprj_oen_buffers\[59\]/li_1535_n17#
+ user_to_mprj_oen_buffers\[42\]/li_891_527# FILLER_14_355/li_0_n17# user_to_mprj_in_gates\[115\]/li_18_51#
+ la_buf\[3\]/li_615_527# powergood_check/FILLER_1_32/li_257_n17# la_buf\[53\]/li_1443_527#
+ la_buf\[108\]/li_215_311# user_to_mprj_oen_buffers\[125\]/li_215_311# user_to_mprj_in_gates\[6\]/li_18_51#
+ FILLER_23_607/li_63_527# user_to_mprj_oen_buffers\[7\]/li_707_527# la_buf\[4\]/li_1351_n17#
+ la_buf\[60\]/li_983_527# _559_/li_155_527# FILLER_15_96/li_0_527# la_buf\[106\]/li_17_51#
+ user_to_mprj_in_gates\[124\]/li_523_n17# user_to_mprj_oen_buffers\[23\]/li_207_51#
+ ANTENNA_mprj_sel_buf\[0\]_TE/li_63_n17# _558_/li_0_527# PHY_264/li_0_527# la_buf\[95\]/li_1443_527#
+ PHY_403/li_0_n17# FILLER_14_456/li_0_n17# la_buf\[99\]/li_1167_527# PHY_373/li_0_n17#
+ mprj_adr_buf\[9\]/li_17_51# _446_/li_0_527# user_to_mprj_in_buffers\[124\]/li_339_527#
+ mprj_dat_buf\[10\]/li_17_51# user_to_mprj_oen_buffers\[57\]/li_215_311# _649_/li_155_n17#
+ _561_/li_155_527# la_buf\[30\]/li_63_527# la_buf\[12\]/li_215_311# FILLER_13_1177/li_63_527#
+ _334_/li_0_527# powergood_check/FILLER_1_48/li_737_797# FILLER_21_1436/li_155_n17#
+ FILLER_6_829/li_0_527# _485_/li_0_527# FILLER_25_1200/li_0_n17# user_to_mprj_in_gates\[51\]/li_523_n17#
+ FILLER_17_1996/li_63_527# user_to_mprj_oen_buffers\[113\]/li_215_311# mprj_dat_buf\[29\]/li_17_51#
+ mprj_adr_buf\[18\]/li_207_51# la_buf\[28\]/li_983_n17# _433_/li_0_527# _373_/li_0_527#
+ la_buf\[51\]/li_611_17# PHY_830/li_0_n17# la_buf\[80\]/li_63_527# user_to_mprj_oen_buffers\[93\]/li_983_527#
+ user_to_mprj_oen_buffers\[95\]/li_17_51# powergood_check/FILLER_0_168/li_115_72#
+ FILLER_11_744/li_0_n17# _352_/li_155_n17# powergood_check/FILLER_0_96/li_161_797#
+ _439_/li_155_527# user_to_mprj_oen_buffers\[89\]/li_207_51# PHY_807/li_0_527# ANTENNA_la_buf\[37\]_TE/li_63_n17#
+ ANTENNA__371__A/li_63_527# _651_/li_155_n17# user_to_mprj_in_buffers\[60\]/li_51_367#
+ user_to_mprj_in_gates\[112\]/li_523_n17# PHY_769/li_0_527# mprj_dat_buf\[31\]/li_1259_n17#
+ PHY_754/li_0_527# FILLER_13_1239/li_0_527# user_to_mprj_in_gates\[110\]/li_247_527#
+ la_buf\[67\]/li_707_n17# la_buf\[14\]/li_707_527# FILLER_21_74/li_0_527# la_buf\[98\]/li_1443_n17#
+ user_to_mprj_in_gates\[30\]/li_523_527# FILLER_12_982/li_63_527# user_to_mprj_in_buffers\[94\]/li_155_527#
+ user_to_mprj_in_buffers\[47\]/li_404_367# la_buf\[86\]/li_779_17# PHY_229/li_0_527#
+ _576_/li_0_n17# mprj_adr_buf\[20\]/li_207_51# user_to_mprj_oen_buffers\[30\]/li_1535_n17#
+ la_buf\[49\]/li_431_n17# PHY_346/li_0_527# FILLER_15_1437/li_155_n17# user_to_mprj_in_gates\[62\]/li_18_51#
+ user_to_mprj_oen_buffers\[45\]/li_215_311# user_to_mprj_in_buffers\[6\]/li_236_17#
+ user_to_mprj_in_gates\[104\]/li_707_n17# user_to_mprj_oen_buffers\[91\]/li_207_51#
+ FILLER_7_942/li_155_527# ANTENNA__380__A/li_63_n17# user_to_mprj_in_gates\[90\]/li_155_n17#
+ FILLER_5_964/li_63_527# user_to_mprj_in_gates\[99\]/li_0_527# powergood_check/mprj_logic_high_lv/li_1025_1611#
+ PHY_17/li_0_527# la_buf\[120\]/li_63_n17# user_to_mprj_oen_buffers\[101\]/li_215_311#
+ PHY_247/li_0_527# FILLER_13_1788/li_63_n17# _354_/li_247_n17# powergood_check/FILLER_2_171/li_65_n17#
+ la_buf\[114\]/li_207_51# ANTENNA__339__A/li_63_n17# ANTENNA_user_to_mprj_oen_buffers\[3\]_A/li_63_n17#
+ la_buf\[29\]/li_0_527# powergood_check/FILLER_0_176/li_65_n17# PHY_452/li_0_n17#
+ FILLER_23_1510/li_0_n17# mprj_dat_buf\[11\]/li_611_17# PHY_223/li_0_527# powergood_check/FILLER_0_32/li_100_536#
+ user_to_mprj_oen_buffers\[44\]/li_17_51# mprj_adr_buf\[15\]/li_523_n17# user_to_mprj_in_gates\[100\]/li_523_n17#
+ FILLER_25_934/li_0_527# la_buf\[70\]/li_1167_527# FILLER_13_1217/li_0_n17# la_buf\[56\]/li_17_51#
+ FILLER_11_2093/li_0_527# FILLER_22_2092/li_63_527# user_to_mprj_in_gates\[90\]/li_615_527#
+ la_buf\[53\]/li_207_51# PHY_842/li_0_n17# FILLER_9_1127/li_63_n17# la_buf\[27\]/li_795_379#
+ FILLER_5_743/li_155_527# powergood_check/FILLER_2_8/li_353_797# la_buf\[37\]/li_431_n17#
+ powergood_check/FILLER_0_32/li_449_797# ANTENNA_user_to_mprj_in_gates\[88\]_A/li_63_527#
+ FILLER_25_957/li_0_n17# user_to_mprj_oen_buffers\[33\]/li_215_311# FILLER_18_1529/li_0_527#
+ user_to_mprj_in_gates\[49\]/li_615_527# user_to_mprj_in_gates\[11\]/li_18_51# powergood_check/FILLER_2_179/li_100_536#
+ _594_/li_0_527# user_to_mprj_oen_buffers\[62\]/li_1075_n17# powergood_check/FILLER_2_16/li_449_n17#
+ PHY_391/li_0_527# user_to_mprj_in_buffers\[15\]/li_236_17# PHY_82/li_0_n17# _597_/li_155_n17#
+ FILLER_13_202/li_155_n17# FILLER_26_819/li_0_527# FILLER_11_548/li_0_n17# PHY_781/li_0_527#
+ PHY_690/li_0_527# powergood_check/FILLER_2_179/li_449_797# _586_/li_0_n17# user_to_mprj_oen_buffers\[88\]/li_707_n17#
+ FILLER_9_1805/li_0_527# FILLER_6_1013/li_63_n17# _378_/li_247_527# la_buf\[3\]/li_247_527#
+ _589_/li_247_n17# user_to_mprj_in_buffers\[23\]/li_404_367# powergood_check/FILLER_2_211/li_545_797#
+ mprj_dat_buf\[13\]/li_207_51# _387_/li_155_527# mprj_adr_buf\[2\]/li_1259_n17# FILLER_12_1796/li_155_527#
+ _362_/li_0_n17# FILLER_11_1135/li_0_527# user_to_mprj_oen_buffers\[21\]/li_215_311#
+ FILLER_11_1449/li_63_n17# PHY_226/li_0_527# ANTENNA__576__A/li_155_n17# user_to_mprj_in_gates\[65\]/li_339_n17#
+ la_buf\[109\]/li_431_n17# user_to_mprj_oen_buffers\[93\]/li_1167_527# _500_/li_155_527#
+ FILLER_16_1939/li_63_n17# FILLER_19_1417/li_0_527# mprj_dat_buf\[19\]/li_1351_527#
+ _464_/li_0_527# la_buf\[74\]/li_0_527# user_to_mprj_oen_buffers\[100\]/li_17_51#
+ user_to_mprj_oen_buffers\[79\]/li_1443_n17# powergood_check/FILLER_2_235/li_115_72#
+ user_to_mprj_oen_buffers\[37\]/li_0_527# user_to_mprj_in_buffers\[117\]/li_51_17#
+ user_to_mprj_in_gates\[42\]/li_63_n17# FILLER_10_325/li_0_n17# PHY_495/li_0_527#
+ PHY_808/li_0_527# user_to_mprj_in_gates\[39\]/li_707_367# user_to_mprj_in_buffers\[64\]/li_404_17#
+ FILLER_9_627/li_0_527# PHY_89/li_0_527# powergood_check/FILLER_2_171/li_641_797#
+ PHY_485/li_0_527# user_to_mprj_oen_buffers\[28\]/li_207_51# ANTENNA__581__A/li_63_n17#
+ user_to_mprj_in_gates\[44\]/li_339_527# PHY_753/li_0_n17# _489_/li_0_527# FILLER_14_1692/li_0_527#
+ user_to_mprj_oen_buffers\[91\]/li_707_n17# _339_/li_247_n17# FILLER_12_1931/li_63_527#
+ user_to_mprj_oen_buffers\[119\]/li_17_51# PHY_790/li_0_527# powergood_check/FILLER_0_232/li_545_797#
+ FILLER_25_544/li_63_527# _595_/li_247_527# PHY_845/li_0_n17# powergood_check/mprj2_logic_high_lv/li_65_1611#
+ PHY_462/li_0_527# FILLER_21_2061/li_63_527# user_to_mprj_oen_buffers\[56\]/li_0_527#
+ powergood_check/FILLER_2_203/li_353_n17# user_to_mprj_in_gates\[120\]/li_339_527#
+ _501_/li_0_527# la_buf\[35\]/li_63_527# _391_/li_155_527# ANTENNA__356__A/li_63_n17#
+ _653_/li_0_n17# user_to_mprj_oen_buffers\[30\]/li_207_51# PHY_852/li_0_527# user_to_mprj_in_gates\[114\]/li_18_51#
+ mprj_adr_buf\[27\]/li_215_311# FILLER_15_1688/li_155_n17# FILLER_23_2085/li_0_n17#
+ powergood_check/FILLER_2_243/li_641_n17# user_to_mprj_oen_buffers\[49\]/li_983_527#
+ user_to_mprj_in_gates\[5\]/li_18_51# _357_/li_155_n17# powergood_check/FILLER_1_62/li_353_n17#
+ powergood_check/FILLER_0_192/li_641_797# FILLER_9_559/li_63_n17# ANTENNA_user_to_mprj_in_gates\[105\]_B/li_63_n17#
+ user_to_mprj_in_gates\[27\]/li_707_367# _656_/li_155_n17# PHY_176/li_0_527# user_to_mprj_in_gates\[76\]/li_339_n17#
+ user_to_mprj_in_gates\[34\]/li_615_n17# ANTENNA_user_to_mprj_in_gates\[49\]_B/li_63_527#
+ la_buf\[105\]/li_17_51# user_to_mprj_in_gates\[32\]/li_339_527# FILLER_12_1552/li_0_n17#
+ mprj_adr_buf\[12\]/li_1351_527# powergood_check/FILLER_1_164/li_65_n17# _548_/li_0_527#
+ user_to_mprj_in_buffers\[42\]/li_523_n17# ANTENNA_user_to_mprj_oen_buffers\[73\]_A/li_63_n17#
+ user_to_mprj_in_gates\[88\]/li_431_n17# mprj_adr_buf\[25\]/li_207_51# FILLER_11_1666/li_0_n17#
+ FILLER_26_986/li_155_527# FILLER_12_1527/li_0_n17# la_buf\[84\]/li_523_n17# mprj_adr_buf\[8\]/li_17_51#
+ FILLER_21_1405/li_63_n17# PHY_377/li_0_527# FILLER_13_1279/li_63_527# FILLER_25_520/li_155_n17#
+ PHY_40/li_0_n17# _446_/li_155_527# user_to_mprj_oen_buffers\[96\]/li_207_51# _587_/li_0_527#
+ ANTENNA_user_to_mprj_in_gates\[95\]_A/li_63_n17# PHY_837/li_0_n17# user_to_mprj_in_gates\[41\]/li_339_n17#
+ FILLER_14_1533/li_63_527# powergood_check/FILLER_2_8/li_65_797# mprj_adr_buf\[2\]/li_431_n17#
+ FILLER_20_1625/li_0_527# mprj_adr_buf\[15\]/li_215_311# la_buf\[39\]/li_1351_527#
+ la_buf\[9\]/li_1259_n17# la_buf\[119\]/li_207_51# _359_/li_247_n17# la_buf\[80\]/li_0_527#
+ user_to_mprj_in_gates\[95\]/li_155_n17# mprj_dat_buf\[28\]/li_17_51# FILLER_25_1502/li_0_527#
+ FILLER_25_1071/li_63_n17# PHY_735/li_0_n17# _363_/li_0_527# _567_/li_0_527# FILLER_18_1994/li_0_n17#
+ PHY_374/li_0_527# user_to_mprj_in_gates\[15\]/li_707_367# la_buf\[80\]/li_247_n17#
+ user_to_mprj_oen_buffers\[94\]/li_17_51# la_buf\[38\]/li_891_n17# FILLER_16_2087/li_155_527#
+ user_to_mprj_oen_buffers\[121\]/li_1351_527# mprj_adr_buf\[11\]/li_707_n17# la_buf\[58\]/li_207_51#
+ _369_/li_0_527# user_to_mprj_oen_buffers\[0\]/li_207_51# PHY_764/li_0_527# ANTENNA__339__A/li_0_n17#
+ FILLER_12_1338/li_63_527# FILLER_10_621/li_155_n17# _336_/li_247_n17# FILLER_26_978/li_63_527#
+ _361_/li_247_n17# la_buf\[121\]/li_207_51# mprj_dat_buf\[27\]/li_1075_n17# _574_/li_247_n17#
+ _397_/li_247_527# powergood_check/FILLER_2_259/li_0_797# user_to_mprj_in_gates\[61\]/li_18_51#
+ la_buf\[94\]/li_1535_527# _625_/li_0_527# FILLER_5_861/li_0_527# FILLER_17_1405/li_63_527#
+ PHY_430/li_0_527# la_buf\[60\]/li_207_51# PHY_773/li_0_527# FILLER_12_1106/li_63_527#
+ powergood_check/FILLER_1_244/li_65_797# user_to_mprj_in_buffers\[113\]/li_236_17#
+ PHY_849/li_0_n17# user_to_mprj_in_gates\[83\]/li_155_n17# FILLER_9_888/li_0_527#
+ powergood_check/FILLER_1_48/li_737_n17# FILLER_25_1204/li_0_n17# user_to_mprj_in_buffers\[107\]/li_155_n17#
+ FILLER_23_493/li_155_n17# FILLER_3_759/li_155_527# la_buf\[97\]/li_215_311# la_buf\[41\]/li_779_17#
+ user_to_mprj_oen_buffers\[43\]/li_17_51# user_to_mprj_oen_buffers\[40\]/li_707_n17#
+ la_buf\[50\]/li_1075_527# mprj_adr_buf\[21\]/li_0_n17# FILLER_10_1382/li_63_n17#
+ powergood_check/FILLER_1_228/li_115_72# la_buf\[55\]/li_17_51# FILLER_15_1928/li_63_527#
+ mprj_dat_buf\[18\]/li_207_51# user_to_mprj_oen_buffers\[42\]/li_1351_527# la_buf\[73\]/li_63_n17#
+ FILLER_19_1587/li_0_527# FILLER_17_1883/li_0_527# user_to_mprj_in_buffers\[117\]/li_404_367#
+ user_to_mprj_oen_buffers\[85\]/li_1443_n17# powergood_check/mprj_logic_high_hvl/li_65_797#
+ user_to_mprj_in_gates\[10\]/li_18_51# mprj_adr_buf\[7\]/li_1443_527# FILLER_10_481/li_63_n17#
+ user_to_mprj_in_buffers\[45\]/li_523_527# FILLER_26_93/li_63_527# powergood_check/FILLER_0_264/li_161_797#
+ _649_/li_0_n17# user_to_mprj_in_buffers\[92\]/li_236_17# FILLER_26_1233/li_63_527#
+ FILLER_26_1054/li_0_527# FILLER_12_1482/li_0_n17# user_to_mprj_in_gates\[47\]/li_63_n17#
+ mprj_adr_buf\[28\]/li_611_17# mprj_dat_buf\[20\]/li_207_51# la_buf\[118\]/li_1167_527#
+ _394_/li_155_527# user_to_mprj_in_gates\[100\]/li_63_n17# FILLER_21_70/li_63_n17#
+ user_to_mprj_in_buffers\[69\]/li_404_17# user_to_mprj_in_gates\[29\]/li_18_51# FILLER_11_1210/li_155_527#
+ PHY_836/li_0_527# la_buf\[85\]/li_215_311# PHY_863/li_0_n17# PHY_456/li_0_n17# user_to_mprj_oen_buffers\[38\]/li_1351_527#
+ _403_/li_0_527# FILLER_14_1500/li_155_n17# FILLER_12_1588/li_0_n17# FILLER_26_841/li_63_527#
+ FILLER_14_2096/li_0_n17# user_to_mprj_oen_buffers\[82\]/li_523_n17# FILLER_13_1013/li_155_527#
+ FILLER_22_1444/li_0_527# mprj_adr_buf\[11\]/li_1443_n17# _391_/li_0_n17# user_to_mprj_in_buffers\[71\]/li_404_17#
+ FILLER_11_794/li_155_n17# ANTENNA__392__A/li_0_527# user_to_mprj_oen_buffers\[35\]/li_207_51#
+ mprj2_pwrgood/li_155_527# FILLER_21_1812/li_63_527# mprj_adr_buf\[28\]/li_431_n17#
+ FILLER_13_345/li_0_527# powergood_check/FILLER_0_200/li_100_536# la_buf\[2\]/li_63_n17#
+ FILLER_21_1451/li_155_n17# la_buf\[111\]/li_0_527# powergood_check/FILLER_2_8/li_353_n17#
+ FILLER_25_1265/li_155_n17# FILLER_22_1886/li_0_527# PHY_829/li_0_527# FILLER_15_1506/li_0_n17#
+ FILLER_16_1839/li_63_527# user_to_mprj_in_gates\[31\]/li_431_527# FILLER_8_1020/li_155_527#
+ powergood_check/FILLER_1_48/li_257_797# la_buf\[14\]/li_1167_527# FILLER_13_1071/li_0_527#
+ FILLER_9_1246/li_0_527# mprj_rstn_buf/li_215_311# FILLER_13_727/li_0_527# la_buf\[65\]/li_523_n17#
+ user_to_mprj_oen_buffers\[114\]/li_1535_527# la_buf\[73\]/li_215_311# powergood_check/FILLER_0_200/li_449_797#
+ user_to_mprj_in_buffers\[46\]/li_339_n17# user_to_mprj_in_buffers\[77\]/li_51_17#
+ la_buf\[109\]/li_983_n17# user_to_mprj_oen_buffers\[118\]/li_17_51# FILLER_21_1444/li_0_n17#
+ la_buf\[96\]/li_1351_527# user_to_mprj_in_gates\[40\]/li_431_n17# FILLER_21_1440/li_155_n17#
+ PHY_785/li_0_527# mprj_dat_buf\[13\]/li_891_n17# mprj_dat_buf\[28\]/li_215_311#
+ la_buf\[109\]/li_707_n17# PHY_29/li_0_n17# powergood_check/FILLER_2_179/li_449_n17#
+ _379_/li_155_n17# user_to_mprj_oen_buffers\[38\]/li_1259_n17# FILLER_11_1274/li_0_n17#
+ powergood_check/FILLER_0_248/li_0_797# user_to_mprj_in_buffers\[28\]/li_339_n17#
+ PHY_74/li_0_527# PHY_872/li_0_527# PHY_777/li_0_527# user_to_mprj_in_gates\[101\]/li_431_n17#
+ powergood_check/FILLER_2_211/li_545_n17# user_to_mprj_in_gates\[113\]/li_18_51#
+ FILLER_21_523/li_0_527# FILLER_13_1025/li_0_527# powergood_check/FILLER_0_160/li_545_797#
+ user_to_mprj_in_gates\[127\]/li_707_n17# user_to_mprj_oen_buffers\[108\]/li_1351_n17#
+ FILLER_12_1186/li_0_n17# user_to_mprj_in_gates\[4\]/li_18_51# FILLER_11_1713/li_0_527#
+ powergood_check/FILLER_1_115/li_65_n17# _453_/li_155_527# ANTENNA_la_buf\[37\]_A/li_63_n17#
+ PHY_311/li_0_n17# mprj_sel_buf\[1\]/li_215_311# user_to_mprj_oen_buffers\[5\]/li_207_51#
+ la_buf\[61\]/li_215_311# FILLER_12_772/li_63_n17# la_buf\[104\]/li_17_51# user_to_mprj_in_gates\[78\]/li_247_n17#
+ la_buf\[57\]/li_707_527# FILLER_19_1916/li_0_n17# user_to_mprj_in_buffers\[63\]/li_0_527#
+ la_buf\[126\]/li_207_51# mprj_adr_buf\[15\]/li_891_527# FILLER_11_996/li_63_n17#
+ mprj_adr_buf\[22\]/li_707_n17# mprj_dat_buf\[16\]/li_215_311# FILLER_26_1544/li_63_527#
+ FILLER_25_554/li_0_527# user_to_mprj_oen_buffers\[62\]/li_1535_n17# FILLER_9_375/li_155_n17#
+ powergood_check/FILLER_2_107/li_545_797# mprj_adr_buf\[7\]/li_17_51# FILLER_11_1569/li_0_n17#
+ powergood_check/FILLER_2_171/li_641_n17# _426_/li_0_527# la_buf\[89\]/li_431_527#
+ FILLER_9_1138/li_63_527# la_buf\[11\]/li_0_n17# FILLER_12_1693/li_63_n17# powergood_check/FILLER_2_107/li_0_797#
+ user_to_mprj_oen_buffers\[90\]/li_1167_n17# powergood_check/FILLER_1_188/li_100_536#
+ user_to_mprj_in_gates\[59\]/li_523_n17# FILLER_11_1287/li_0_527# powergood_check/mprj_logic_high_lv/li_65_797#
+ la_buf\[65\]/li_207_51# mprj_dat_buf\[7\]/li_615_527# la_buf\[122\]/li_1535_n17#
+ FILLER_13_655/li_155_527# la_buf\[90\]/li_891_n17# FILLER_12_1044/li_0_n17# _465_/li_0_527#
+ mprj_dat_buf\[3\]/li_1075_527# _340_/li_0_527# user_to_mprj_oen_buffers\[29\]/li_891_527#
+ _448_/li_0_527# FILLER_11_1338/li_155_527# user_to_mprj_in_gates\[54\]/li_0_527#
+ PHY_305/li_0_n17# powergood_check/FILLER_1_140/li_0_797# FILLER_19_109/li_0_527#
+ mprj_dat_buf\[27\]/li_17_51# la_buf\[61\]/li_1259_n17# ANTENNA_user_to_mprj_oen_buffers\[7\]_A/li_63_527#
+ _353_/li_0_527# PHY_856/li_0_527# la_buf\[98\]/li_431_n17# _333_/li_155_527# FILLER_22_1698/li_0_527#
+ PHY_665/li_0_527# user_to_mprj_oen_buffers\[93\]/li_17_51# FILLER_12_886/li_63_527#
+ user_to_mprj_oen_buffers\[94\]/li_215_311# FILLER_18_1541/li_0_527# FILLER_22_1408/li_63_n17#
+ user_to_mprj_oen_buffers\[38\]/li_611_17# FILLER_13_1084/li_63_527# user_to_mprj_in_gates\[66\]/li_247_n17#
+ FILLER_17_1921/li_63_527# _335_/li_0_527# user_to_mprj_oen_buffers\[24\]/li_247_n17#
+ ANTENNA__654__A/li_63_n17# powergood_check/FILLER_1_131/li_161_797# user_to_mprj_in_buffers\[76\]/li_155_n17#
+ FILLER_10_2077/li_0_n17# PHY_823/li_0_527# mprj_stb_buf/li_1259_527# la_buf\[67\]/li_0_527#
+ FILLER_22_1418/li_63_n17# FILLER_15_226/li_0_527# user_to_mprj_in_gates\[60\]/li_18_51#
+ ANTENNA_user_to_mprj_in_gates\[109\]_A/li_63_n17# user_to_mprj_oen_buffers\[7\]/li_63_n17#
+ FILLER_10_463/li_63_n17# FILLER_5_613/li_0_527# user_to_mprj_in_gates\[47\]/li_523_n17#
+ user_to_mprj_in_buffers\[97\]/li_236_17# user_to_mprj_oen_buffers\[109\]/li_215_311#
+ powergood_check/FILLER_1_140/li_353_797# user_to_mprj_in_gates\[45\]/li_247_527#
+ user_to_mprj_oen_buffers\[40\]/li_611_17# _468_/li_0_n17# user_to_mprj_in_gates\[49\]/li_615_n17#
+ mprj_adr_buf\[10\]/li_63_527# la_buf\[78\]/li_1351_527# la_buf\[44\]/li_983_527#
+ mprj_dat_buf\[25\]/li_207_51# user_to_mprj_in_gates\[105\]/li_63_n17# FILLER_10_505/li_63_n17#
+ ANTENNA__647__A/li_63_n17# user_to_mprj_in_gates\[79\]/li_18_51# la_buf\[100\]/li_0_527#
+ la_buf\[80\]/li_63_n17# FILLER_8_1008/li_0_527# FILLER_23_1451/li_63_n17# FILLER_17_342/li_0_n17#
+ user_to_mprj_in_gates\[106\]/li_247_527# powergood_check/FILLER_2_8/li_65_n17# _512_/li_155_527#
+ la_buf\[53\]/li_891_527# user_to_mprj_oen_buffers\[82\]/li_215_311# user_to_mprj_oen_buffers\[42\]/li_17_51#
+ user_to_mprj_oen_buffers\[107\]/li_1351_527# FILLER_18_1439/li_0_527# user_to_mprj_in_gates\[56\]/li_339_n17#
+ FILLER_21_1634/li_155_527# la_buf\[54\]/li_17_51# la_buf\[121\]/li_215_311# user_to_mprj_in_gates\[54\]/li_63_n17#
+ FILLER_7_1080/li_63_527# powergood_check/FILLER_1_172/li_65_797# user_to_mprj_in_buffers\[0\]/li_51_367#
+ la_buf\[1\]/li_215_311# powergood_check/FILLER_0_216/li_0_n17# user_to_mprj_in_buffers\[76\]/li_404_17#
+ FILLER_15_1517/li_0_527# FILLER_12_1017/li_155_527# user_to_mprj_in_buffers\[92\]/li_51_17#
+ FILLER_18_539/li_0_527# FILLER_9_563/li_0_527# _379_/li_0_527# user_to_mprj_in_gates\[115\]/li_247_n17#
+ powergood_check/FILLER_0_176/li_65_797# _595_/li_0_527# _561_/li_0_527# user_to_mprj_in_gates\[35\]/li_523_n17#
+ PHY_1/li_0_n17# user_to_mprj_oen_buffers\[37\]/li_1351_527# FILLER_10_471/li_63_n17#
+ user_to_mprj_in_gates\[33\]/li_247_527# _639_/li_0_n17# FILLER_0_201/li_155_527#
+ FILLER_13_620/li_0_n17# la_buf\[95\]/li_891_527# user_to_mprj_oen_buffers\[77\]/li_983_527#
+ powergood_check/FILLER_2_24/li_641_797# _472_/li_0_527# user_to_mprj_in_buffers\[72\]/li_404_367#
+ powergood_check/FILLER_1_252/li_641_n17# _527_/li_0_n17# user_to_mprj_in_gates\[46\]/li_0_527#
+ powergood_check/FILLER_0_272/li_353_797# la_buf\[74\]/li_431_n17# powergood_check/mprj_logic_high_lv/li_161_797#
+ user_to_mprj_in_gates\[28\]/li_18_51# PHY_431/li_0_527# PHY_26/li_0_n17# user_to_mprj_oen_buffers\[42\]/li_207_51#
+ FILLER_13_1207/li_63_n17# _415_/li_0_n17# user_to_mprj_oen_buffers\[70\]/li_215_311#
+ la_buf\[110\]/li_63_527# la_buf\[45\]/li_779_17# powergood_check/FILLER_2_243/li_161_n17#
+ mprj_dat_buf\[30\]/li_891_527# user_to_mprj_in_gates\[42\]/li_247_n17# mprj_dat_buf\[29\]/li_431_n17#
+ powergood_check/FILLER_0_192/li_161_797# user_to_mprj_in_buffers\[94\]/li_523_527#
+ FILLER_25_1208/li_0_n17# mprj_dat_buf\[14\]/li_0_n17# FILLER_17_1921/li_0_527# la_buf\[119\]/li_0_527#
+ la_buf\[41\]/li_983_n17# la_buf\[3\]/li_779_17# user_to_mprj_oen_buffers\[29\]/li_215_311#
+ _575_/li_0_527# la_buf\[105\]/li_0_527# FILLER_13_911/li_155_527# _386_/li_247_n17#
+ la_buf\[73\]/li_983_527# FILLER_15_1951/li_0_527# _580_/li_155_527# user_to_mprj_in_gates\[103\]/li_247_n17#
+ user_to_mprj_in_gates\[88\]/li_707_367# _342_/li_0_n17# FILLER_11_897/li_63_n17#
+ powergood_check/FILLER_2_219/li_353_797# user_to_mprj_in_gates\[95\]/li_615_n17#
+ la_buf\[122\]/li_523_n17# FILLER_24_56/li_63_527# PHY_787/li_0_527# user_to_mprj_in_gates\[21\]/li_247_527#
+ FILLER_11_1429/li_63_n17# FILLER_12_1069/li_63_527# FILLER_9_782/li_0_527# PHY_323/li_0_n17#
+ FILLER_7_1148/li_155_n17# la_buf\[70\]/li_611_17# PHY_747/li_0_n17# la_buf\[0\]/li_1351_n17#
+ _570_/li_0_527# FILLER_25_1922/li_0_n17# _371_/li_155_n17# FILLER_11_1468/li_63_n17#
+ ANTENNA__589__A/li_63_n17# mprj_stb_buf/li_983_n17# powergood_check/mprj_logic_high_hvl/li_65_n17#
+ powergood_check/FILLER_2_259/li_641_797# FILLER_20_449/li_0_527# mprj_dat_buf\[27\]/li_1535_n17#
+ _390_/li_247_n17# user_to_mprj_in_gates\[30\]/li_247_n17# user_to_mprj_in_buffers\[19\]/li_404_367#
+ powergood_check/mprj2_logic_high_lv/li_257_1611# FILLER_9_992/li_0_527# user_to_mprj_oen_buffers\[117\]/li_17_51#
+ FILLER_13_669/li_63_527# user_to_mprj_oen_buffers\[74\]/li_983_n17# FILLER_9_516/li_155_n17#
+ mprj_dat_buf\[28\]/li_611_17# user_to_mprj_oen_buffers\[17\]/li_215_311# ANTENNA__352__A/li_63_n17#
+ _624_/li_0_527# _548_/li_155_n17# FILLER_13_202/li_0_527# user_to_mprj_in_gates\[76\]/li_707_367#
+ ANTENNA_user_to_mprj_in_gates\[127\]_B/li_63_527# PHY_76/li_0_527# ANTENNA_user_to_mprj_in_gates\[99\]_A/li_63_527#
+ FILLER_13_1013/li_155_n17# user_to_mprj_in_gates\[81\]/li_339_527# user_to_mprj_in_gates\[38\]/li_247_n17#
+ user_to_mprj_oen_buffers\[119\]/li_707_527# user_to_mprj_oen_buffers\[63\]/li_1351_n17#
+ la_buf\[6\]/li_1443_n17# user_to_mprj_oen_buffers\[87\]/li_0_527# PHY_830/li_0_527#
+ powergood_check/FILLER_2_251/li_257_797# la_buf\[99\]/li_1351_n17# PHY_230/li_0_n17#
+ user_to_mprj_in_gates\[112\]/li_18_51# FILLER_13_1017/li_0_527# mprj_cyc_buf/li_207_51#
+ user_to_mprj_oen_buffers\[91\]/li_779_17# ANTENNA__331__A/li_63_527# la_buf\[116\]/li_983_n17#
+ user_to_mprj_oen_buffers\[95\]/li_431_n17# la_buf\[44\]/li_0_527# user_to_mprj_in_gates\[3\]/li_18_51#
+ la_buf\[47\]/li_611_17# FILLER_13_2091/li_63_n17# _550_/li_155_n17# la_buf\[27\]/li_707_n17#
+ mprj_stb_buf/li_431_527# FILLER_11_322/li_63_n17# la_buf\[4\]/li_795_379# la_buf\[15\]/li_0_n17#
+ la_buf\[114\]/li_779_17# la_buf\[72\]/li_207_51# user_to_mprj_oen_buffers\[92\]/li_707_527#
+ la_buf\[103\]/li_17_51# powergood_check/FILLER_1_48/li_257_n17# user_to_mprj_in_buffers\[6\]/li_155_n17#
+ FILLER_10_471/li_155_n17# user_to_mprj_oen_buffers\[24\]/li_63_527# la_buf\[79\]/li_247_527#
+ user_to_mprj_oen_buffers\[62\]/li_983_n17# ANTENNA__361__A/li_0_527# FILLER_13_1574/li_0_n17#
+ mprj_adr_buf\[6\]/li_17_51# user_to_mprj_in_buffers\[15\]/li_404_17# powergood_check/FILLER_1_204/li_65_n17#
+ user_to_mprj_oen_buffers\[111\]/li_63_n17# user_to_mprj_in_gates\[64\]/li_707_367#
+ user_to_mprj_oen_buffers\[45\]/li_611_17# mprj_clk_buf/li_17_51# FILLER_12_693/li_155_527#
+ user_to_mprj_oen_buffers\[83\]/li_1351_527# la_buf\[113\]/li_431_527# mprj_cyc_buf/li_431_527#
+ mprj_dat_buf\[3\]/li_983_n17# powergood_check/FILLER_0_200/li_115_72# powergood_check/FILLER_2_115/li_737_797#
+ la_buf\[110\]/li_1535_527# ANTENNA_user_to_mprj_in_gates\[52\]_B/li_63_527# user_to_mprj_in_gates\[80\]/li_155_n17#
+ mprj_adr_buf\[2\]/li_891_n17# la_buf\[85\]/li_63_n17# _401_/li_0_n17# user_to_mprj_oen_buffers\[83\]/li_431_n17#
+ mprj_dat_buf\[26\]/li_17_51# FILLER_21_593/li_0_527# _430_/li_155_n17# _343_/li_0_527#
+ FILLER_25_1071/li_155_n17# FILLER_25_1051/li_63_n17# FILLER_9_1138/li_63_n17# FILLER_17_2033/li_0_527#
+ la_buf\[13\]/li_1167_527# la_buf\[15\]/li_707_n17# powergood_check/FILLER_0_80/li_100_536#
+ user_to_mprj_oen_buffers\[92\]/li_17_51# _494_/li_0_527# FILLER_13_1199/li_155_527#
+ FILLER_7_2083/li_0_527# FILLER_25_1506/li_0_n17# la_buf\[122\]/li_431_n17# FILLER_12_1683/li_0_527#
+ powergood_check/mprj2_logic_high_hvl/li_257_797# user_to_mprj_oen_buffers\[80\]/li_707_527#
+ PHY_80/li_0_527# la_buf\[29\]/li_1075_527# FILLER_11_1717/li_0_527# user_to_mprj_in_gates\[59\]/li_63_n17#
+ FILLER_23_1998/li_0_n17# _589_/li_247_527# la_buf\[2\]/li_431_n17# FILLER_13_1816/li_155_527#
+ la_buf\[82\]/li_983_n17# powergood_check/mprj2_logic_high_lv/li_1313_1611# la_buf\[77\]/li_891_527#
+ user_to_mprj_in_gates\[112\]/li_63_n17# la_buf\[1\]/li_207_51# user_to_mprj_in_gates\[111\]/li_615_527#
+ FILLER_25_849/li_63_n17# user_to_mprj_oen_buffers\[48\]/li_1535_n17# mprj_adr_buf\[29\]/li_615_527#
+ FILLER_27_798/li_155_n17# powergood_check/FILLER_0_80/li_449_797# user_to_mprj_in_gates\[52\]/li_707_367#
+ FILLER_25_1200/li_0_527# mprj_adr_buf\[21\]/li_63_527# FILLER_12_581/li_63_527#
+ _580_/li_0_527# mprj_dat_buf\[13\]/li_779_17# la_buf\[30\]/li_0_527# user_to_mprj_in_buffers\[4\]/li_404_367#
+ user_to_mprj_oen_buffers\[61\]/li_795_379# powergood_check/FILLER_2_107/li_545_n17#
+ mprj_sel_buf\[3\]/li_1443_527# user_to_mprj_in_gates\[113\]/li_707_367# FILLER_25_558/li_0_527#
+ la_buf\[109\]/li_1443_n17# powergood_check/mprj2_logic_high_lv/li_641_1611# mprj_adr_buf\[5\]/li_215_311#
+ powergood_check/FILLER_2_107/li_0_n17# la_buf\[72\]/li_1259_527# user_to_mprj_oen_buffers\[71\]/li_431_n17#
+ la_buf\[12\]/li_1443_n17# user_to_mprj_in_gates\[16\]/li_339_527# user_to_mprj_in_gates\[78\]/li_18_51#
+ FILLER_21_1448/li_63_n17# la_buf\[50\]/li_1075_n17# user_to_mprj_oen_buffers\[47\]/li_207_51#
+ FILLER_13_699/li_0_n17# FILLER_11_669/li_63_n17# user_to_mprj_oen_buffers\[41\]/li_17_51#
+ FILLER_20_465/li_0_527# la_buf\[28\]/li_1351_n17# user_to_mprj_oen_buffers\[6\]/li_1443_527#
+ la_buf\[53\]/li_17_51# FILLER_19_1658/li_0_n17# la_buf\[75\]/li_983_n17# user_to_mprj_oen_buffers\[50\]/li_431_527#
+ la_buf\[54\]/li_63_527# powergood_check/FILLER_0_192/li_65_n17# user_to_mprj_in_gates\[25\]/li_339_n17#
+ powergood_check/mprj_logic_high_lv/li_1455_797# user_to_mprj_in_buffers\[91\]/li_51_17#
+ mprj_dat_buf\[15\]/li_1351_527# powergood_check/FILLER_2_155/li_0_797# mprj_adr_buf\[4\]/li_207_51#
+ FILLER_25_303/li_0_n17# la_buf\[75\]/li_779_17# user_to_mprj_in_gates\[79\]/li_155_n17#
+ FILLER_22_1677/li_0_527# powergood_check/FILLER_1_131/li_161_n17# powergood_check/FILLER_1_220/li_545_n17#
+ powergood_check/FILLER_0_240/li_257_797# _376_/li_155_n17# mprj_rstn_buf/li_207_51#
+ user_to_mprj_in_gates\[101\]/li_707_367# user_to_mprj_in_gates\[78\]/li_707_n17#
+ mprj_adr_buf\[23\]/li_1351_n17# FILLER_15_1437/li_63_n17# PHY_278/li_0_527# powergood_check/FILLER_1_140/li_353_n17#
+ user_to_mprj_in_gates\[119\]/li_707_n17# user_to_mprj_in_gates\[27\]/li_18_51# user_to_mprj_in_buffers\[18\]/li_615_n17#
+ FILLER_26_990/li_0_527# mprj_dat_buf\[25\]/li_983_n17# _556_/li_0_n17# la_buf\[11\]/li_207_51#
+ FILLER_15_226/li_63_527# FILLER_13_1714/li_155_n17# user_to_mprj_oen_buffers\[62\]/li_63_n17#
+ _535_/li_0_n17# powergood_check/FILLER_0_96/li_0_797# _436_/li_0_527# user_to_mprj_oen_buffers\[47\]/li_707_527#
+ powergood_check/FILLER_2_251/li_353_n17# la_buf\[55\]/li_707_527# user_to_mprj_oen_buffers\[63\]/li_891_n17#
+ powergood_check/FILLER_1_180/li_641_n17# _595_/li_0_n17# FILLER_17_583/li_0_527#
+ user_to_mprj_in_gates\[119\]/li_155_527# la_buf\[7\]/li_779_17# mprj_adr_buf\[25\]/li_779_17#
+ user_to_mprj_in_buffers\[40\]/li_51_17# powergood_check/mprj2_logic_high_lv/li_179_79#
+ la_buf\[7\]/li_247_527# user_to_mprj_in_gates\[39\]/li_431_527# PHY_227/li_0_n17#
+ _483_/li_0_n17# powergood_check/FILLER_2_171/li_161_n17# PHY_429/li_0_527# user_to_mprj_oen_buffers\[103\]/li_207_51#
+ PHY_266/li_0_n17# _374_/li_0_527# _371_/li_0_n17# powergood_check/FILLER_2_227/li_545_797#
+ ANTENNA_user_to_mprj_in_gates\[73\]_B/li_63_n17# user_to_mprj_in_gates\[66\]/li_707_n17#
+ _555_/li_155_n17# la_buf\[4\]/li_611_17# mprj_cyc_buf/li_247_527# user_to_mprj_oen_buffers\[24\]/li_707_n17#
+ la_buf\[26\]/li_983_527# user_to_mprj_in_buffers\[111\]/li_155_527# user_to_mprj_in_buffers\[76\]/li_615_n17#
+ la_buf\[77\]/li_207_51# PHY_390/li_0_n17# user_to_mprj_in_gates\[46\]/li_155_527#
+ powergood_check/FILLER_2_24/li_641_n17# la_buf\[116\]/li_247_n17# FILLER_11_992/li_155_527#
+ _380_/li_247_n17# FILLER_13_1574/li_155_527# user_to_mprj_oen_buffers\[116\]/li_17_51#
+ powergood_check/FILLER_0_208/li_257_797# FILLER_17_176/li_0_527# FILLER_19_1417/li_63_n17#
+ ANTENNA_user_to_mprj_in_gates\[91\]_A/li_63_n17# ANTENNA_user_to_mprj_in_gates\[63\]_B/li_63_527#
+ PHY_729/li_0_n17# powergood_check/mprj_logic_high_lv/li_65_1611# la_buf\[58\]/li_779_17#
+ FILLER_15_1569/li_0_527# user_to_mprj_in_gates\[48\]/li_615_n17# user_to_mprj_in_gates\[109\]/li_431_n17#
+ user_to_mprj_in_gates\[107\]/li_155_527# powergood_check/FILLER_2_187/li_641_797#
+ mprj_dat_buf\[3\]/li_431_527# _577_/li_247_527# la_buf\[60\]/li_1075_n17# user_to_mprj_in_gates\[99\]/li_523_527#
+ user_to_mprj_in_gates\[27\]/li_431_527# FILLER_13_1704/li_0_n17# ANTENNA_user_to_mprj_in_buffers\[2\]_A/li_63_n17#
+ _554_/li_247_n17# user_to_mprj_in_gates\[55\]/li_155_n17# PHY_824/li_0_n17# la_buf\[126\]/li_1535_527#
+ powergood_check/FILLER_0_248/li_545_797# powergood_check/FILLER_2_171/li_115_72#
+ _557_/li_247_n17# FILLER_24_1522/li_0_527# user_to_mprj_in_gates\[111\]/li_18_51#
+ PHY_616/li_0_527# _435_/li_155_n17# powergood_check/FILLER_2_219/li_353_n17# user_to_mprj_in_buffers\[104\]/li_0_n17#
+ la_buf\[69\]/li_215_311# PHY_327/li_0_n17# user_to_mprj_in_gates\[60\]/li_523_n17#
+ user_to_mprj_in_gates\[2\]/li_18_51# powergood_check/FILLER_0_168/li_353_797# PHY_385/li_0_n17#
+ user_to_mprj_oen_buffers\[52\]/li_611_17# user_to_mprj_in_gates\[116\]/li_155_n17#
+ _540_/li_0_527# FILLER_11_1402/li_0_n17# FILLER_25_222/li_0_n17# mprj_vdd_pwrgood/li_19_289#
+ _557_/li_0_527# user_to_mprj_in_gates\[36\]/li_431_n17# _482_/li_247_n17# la_buf\[46\]/li_1351_527#
+ FILLER_10_1931/li_63_n17# user_to_mprj_oen_buffers\[6\]/li_215_311# FILLER_26_685/li_63_527#
+ la_buf\[102\]/li_17_51# user_to_mprj_in_gates\[115\]/li_707_n17# FILLER_10_1170/li_155_527#
+ user_to_mprj_in_gates\[118\]/li_431_527# la_buf\[6\]/li_207_51# powergood_check/FILLER_2_259/li_641_n17#
+ _524_/li_155_527# user_to_mprj_oen_buffers\[22\]/li_1351_n17# mprj_adr_buf\[29\]/li_63_527#
+ FILLER_12_1660/li_63_527# user_to_mprj_in_buffers\[111\]/li_404_17# user_to_mprj_oen_buffers\[57\]/li_1167_n17#
+ mprj_adr_buf\[5\]/li_17_51# FILLER_9_456/li_63_n17# FILLER_14_1447/li_155_527# user_to_mprj_in_gates\[87\]/li_523_527#
+ FILLER_25_1265/li_63_n17# PHY_95/li_0_n17# PHY_689/li_0_527# FILLER_17_1684/li_0_527#
+ la_buf\[14\]/li_611_17# user_to_mprj_oen_buffers\[124\]/li_707_n17# user_to_mprj_in_gates\[66\]/li_63_n17#
+ la_buf\[72\]/li_615_527# user_to_mprj_in_buffers\[88\]/li_404_17# user_to_mprj_in_gates\[42\]/li_707_n17#
+ mprj_dat_buf\[6\]/li_983_527# FILLER_18_154/li_63_527# mprj2_logic_high_inst/m3_800_806#
+ _596_/li_0_527# la_buf\[57\]/li_215_311# FILLER_19_1778/li_0_n17# FILLER_21_2061/li_155_527#
+ mprj_dat_buf\[25\]/li_17_51# FILLER_12_1923/li_155_n17# mprj_dat_buf\[27\]/li_615_527#
+ mprj_dat_buf\[13\]/li_1259_n17# FILLER_13_1207/li_0_527# _333_/li_0_527# FILLER_24_612/li_0_527#
+ powergood_check/FILLER_2_16/li_65_797# user_to_mprj_oen_buffers\[91\]/li_17_51#
+ powergood_check/FILLER_2_24/li_161_797# user_to_mprj_in_gates\[96\]/li_523_n17#
+ powergood_check/FILLER_1_252/li_161_n17# user_to_mprj_in_gates\[94\]/li_247_527#
+ w_144678_3514# la_buf\[6\]/li_891_n17# mprj_adr_buf\[18\]/li_707_n17# user_to_mprj_in_gates\[103\]/li_707_n17#
+ user_to_mprj_oen_buffers\[90\]/li_891_n17# _372_/li_0_527# FILLER_11_1196/li_0_527#
+ la_buf\[21\]/li_891_527# user_to_mprj_oen_buffers\[81\]/li_1443_n17# FILLER_25_839/li_63_n17#
+ PHY_370/li_0_n17# user_to_mprj_oen_buffers\[54\]/li_207_51# mprj_adr_buf\[9\]/li_207_51#
+ PHY_506/li_0_527# mprj_adr_buf\[28\]/li_891_527# la_buf\[63\]/li_891_527# la_buf\[113\]/li_1443_527#
+ _579_/li_0_527# FILLER_12_689/li_0_527# powergood_check/mprj_logic_high_lv/li_826_79#
+ powergood_check/FILLER_2_243/li_65_n17# FILLER_8_1020/li_63_527# _597_/li_155_527#
+ la_buf\[61\]/li_63_527# la_buf\[45\]/li_215_311# FILLER_21_1989/li_63_527# user_to_mprj_in_gates\[77\]/li_18_51#
+ FILLER_21_123/li_63_n17# FILLER_9_1142/li_0_527# FILLER_16_56/li_0_527# powergood_check/FILLER_2_115/li_737_n17#
+ user_to_mprj_in_gates\[82\]/li_0_n17# la_buf\[16\]/li_207_51# la_buf\[82\]/li_611_17#
+ user_to_mprj_in_gates\[82\]/li_247_527# user_to_mprj_oen_buffers\[40\]/li_17_51#
+ la_buf\[58\]/li_431_527# FILLER_14_1543/li_63_527# la_buf\[25\]/li_0_n17# powergood_check/FILLER_1_260/li_65_797#
+ la_buf\[9\]/li_215_311# FILLER_11_1351/li_63_n17# _383_/li_155_n17# la_buf\[52\]/li_17_51#
+ FILLER_9_928/li_0_n17# ANTENNA_user_to_mprj_in_gates\[112\]_A/li_63_n17# FILLER_25_693/li_63_n17#
+ PHY_337/li_0_527# powergood_check/mprj2_logic_high_hvl/li_257_n17# FILLER_16_536/li_0_527#
+ powergood_check/FILLER_0_24/li_115_72# mprj_adr_buf\[20\]/li_707_527# FILLER_15_502/li_63_527#
+ user_to_mprj_oen_buffers\[59\]/li_17_51# FILLER_25_891/li_63_527# la_buf\[81\]/li_1351_527#
+ FILLER_13_1816/li_155_n17# FILLER_24_2076/li_0_527# la_buf\[99\]/li_523_n17# user_to_mprj_oen_buffers\[108\]/li_207_51#
+ user_to_mprj_in_gates\[91\]/li_247_n17# user_to_mprj_oen_buffers\[93\]/li_615_527#
+ FILLER_11_451/li_63_n17# PHY_727/li_0_527# FILLER_17_60/li_0_527# la_buf\[9\]/li_611_17#
+ la_buf\[29\]/li_63_n17# _472_/li_155_527# user_to_mprj_oen_buffers\[78\]/li_215_311#
+ FILLER_13_1115/li_0_527# _507_/li_0_n17# powergood_check/FILLER_2_32/li_0_797# user_to_mprj_in_buffers\[6\]/li_615_n17#
+ la_buf\[51\]/li_1443_n17# user_to_mprj_oen_buffers\[114\]/li_1167_527# user_to_mprj_in_gates\[44\]/li_0_527#
+ la_buf\[33\]/li_215_311# PHY_34/li_0_527# FILLER_1_1985/li_155_527# FILLER_17_350/li_63_n17#
+ _591_/li_247_527# powergood_check/mprj2_logic_high_lv/li_384_1039# FILLER_20_457/li_0_n17#
+ FILLER_12_471/li_63_527# powergood_check/FILLER_1_16/li_641_n17# ANTENNA_user_to_mprj_in_buffers\[17\]_A/li_63_n17#
+ user_to_mprj_in_gates\[26\]/li_18_51# mprj_dat_buf\[21\]/li_63_527# powergood_check/FILLER_1_164/li_115_72#
+ FILLER_27_873/li_0_n17# la_buf\[117\]/li_215_311# la_buf\[67\]/li_1351_n17# _509_/li_0_527#
+ user_to_mprj_oen_buffers\[110\]/li_207_51# user_to_mprj_in_gates\[125\]/li_615_n17#
+ _546_/li_0_n17# FILLER_12_1664/li_0_527# FILLER_25_1008/li_0_n17# _562_/li_0_n17#
+ FILLER_20_500/li_0_n17# la_buf\[77\]/li_523_n17# mprj_dat_buf\[5\]/li_215_311# ANTENNA__392__A/li_63_527#
+ _585_/li_0_n17# PHY_478/li_0_527# la_buf\[84\]/li_207_51# _473_/li_0_n17# FILLER_15_1569/li_63_527#
+ user_to_mprj_in_buffers\[68\]/li_404_367# FILLER_21_2105/li_63_n17# FILLER_17_1428/li_0_n17#
+ FILLER_16_40/li_63_n17# _361_/li_0_n17# _352_/li_155_527# user_to_mprj_oen_buffers\[66\]/li_215_311#
+ powergood_check/FILLER_2_155/li_0_n17# PHY_862/li_0_n17# _651_/li_155_527# FILLER_26_1195/li_155_527#
+ la_buf\[21\]/li_215_311# powergood_check/FILLER_2_115/li_257_797# user_to_mprj_oen_buffers\[57\]/li_611_17#
+ user_to_mprj_oen_buffers\[7\]/li_431_n17# FILLER_23_56/li_0_n17# la_buf\[105\]/li_215_311#
+ PHY_408/li_0_527# PHY_838/li_0_527# PHY_382/li_0_527# user_to_mprj_oen_buffers\[122\]/li_215_311#
+ _343_/li_247_n17# ANTENNA_la_buf\[121\]_A/li_63_527# powergood_check/FILLER_0_216/li_100_536#
+ powergood_check/FILLER_2_243/li_0_797# mprj_dat_buf\[16\]/li_523_n17# la_buf\[97\]/li_0_n17#
+ FILLER_24_56/li_0_527# FILLER_14_359/li_63_n17# user_to_mprj_oen_buffers\[115\]/li_17_51#
+ FILLER_17_104/li_0_527# FILLER_26_1236/li_0_527# powergood_check/FILLER_2_155/li_545_797#
+ user_to_mprj_oen_buffers\[74\]/li_1443_n17# FILLER_11_1030/li_0_527# FILLER_12_927/li_63_n17#
+ powergood_check/FILLER_1_107/li_353_n17# powergood_check/FILLER_0_216/li_449_797#
+ mprj_adr_buf\[8\]/li_247_n17# la_buf\[50\]/li_63_527# user_to_mprj_oen_buffers\[114\]/li_707_527#
+ mprj_adr_buf\[31\]/li_17_51# _478_/li_155_n17# powergood_check/FILLER_0_8/li_100_536#
+ FILLER_5_861/li_155_527# la_buf\[43\]/li_63_527# _354_/li_247_527# user_to_mprj_in_gates\[124\]/li_63_n17#
+ FILLER_16_289/li_0_n17# user_to_mprj_in_gates\[110\]/li_18_51# FILLER_12_628/li_0_527#
+ user_to_mprj_oen_buffers\[54\]/li_215_311# _378_/li_0_527# _531_/li_155_527# user_to_mprj_in_gates\[28\]/li_339_n17#
+ la_buf\[98\]/li_431_527# user_to_mprj_in_gates\[98\]/li_339_n17# FILLER_24_1401/li_63_527#
+ FILLER_15_70/li_63_527# powergood_check/FILLER_0_264/li_0_797# user_to_mprj_in_gates\[1\]/li_18_51#
+ FILLER_5_909/li_63_527# mprj_dat_buf\[25\]/li_779_17# PHY_717/li_0_527# user_to_mprj_oen_buffers\[110\]/li_215_311#
+ mprj_dat_buf\[18\]/li_1443_527# user_to_mprj_oen_buffers\[27\]/li_1075_527# powergood_check/FILLER_0_8/li_449_797#
+ powergood_check/FILLER_1_236/li_65_n17# FILLER_11_716/li_155_n17# user_to_mprj_in_gates\[73\]/li_63_n17#
+ la_buf\[21\]/li_611_17# powergood_check/FILLER_2_227/li_545_n17# la_buf\[119\]/li_891_527#
+ la_buf\[101\]/li_17_51# FILLER_9_407/li_63_n17# FILLER_19_52/li_155_527# FILLER_12_1106/li_0_527#
+ powergood_check/FILLER_0_176/li_545_797# FILLER_11_1196/li_0_n17# user_to_mprj_oen_buffers\[52\]/li_523_n17#
+ FILLER_28_91/li_0_n17# _409_/li_155_527# ANTENNA_user_to_mprj_in_gates\[105\]_A/li_63_n17#
+ user_to_mprj_in_gates\[79\]/li_615_n17# user_to_mprj_oen_buffers\[59\]/li_207_51#
+ PHY_256/li_0_527# PHY_379/li_0_n17# ANTENNA_user_to_mprj_in_gates\[49\]_A/li_63_527#
+ _659_/li_0_527# user_to_mprj_in_gates\[77\]/li_339_527# FILLER_13_472/li_0_n17#
+ FILLER_13_1239/li_63_527# mprj_adr_buf\[4\]/li_17_51# _370_/li_0_n17# mprj_dat_buf\[6\]/li_1259_527#
+ _590_/li_0_527# la_buf\[72\]/li_0_n17# _553_/li_0_527# user_to_mprj_in_gates\[45\]/li_0_n17#
+ FILLER_12_849/li_0_527# FILLER_7_810/li_0_527# FILLER_9_334/li_63_n17# user_to_mprj_in_gates\[44\]/li_0_n17#
+ user_to_mprj_oen_buffers\[1\]/li_707_n17# mprj_dat_buf\[19\]/li_707_n17# la_buf\[41\]/li_707_527#
+ PHY_221/li_0_n17# FILLER_14_1696/li_63_527# user_to_mprj_oen_buffers\[42\]/li_215_311#
+ powergood_check/FILLER_2_187/li_641_n17# ANTENNA__593__A/li_63_527# user_to_mprj_oen_buffers\[61\]/li_207_51#
+ _586_/li_0_527# FILLER_11_1338/li_0_n17# user_to_mprj_in_gates\[86\]/li_339_n17#
+ la_buf\[22\]/li_0_n17# user_to_mprj_in_gates\[5\]/li_707_n17# mprj_dat_buf\[24\]/li_17_51#
+ FILLER_5_763/li_63_527# FILLER_25_1337/li_155_527# FILLER_7_931/li_0_527# user_to_mprj_oen_buffers\[90\]/li_17_51#
+ mprj_dat_buf\[8\]/li_891_527# _474_/li_0_527# powergood_check/FILLER_0_0/li_641_797#
+ mprj_dat_buf\[21\]/li_431_527# user_to_mprj_in_gates\[119\]/li_615_527# FILLER_10_463/li_0_n17#
+ FILLER_8_1071/li_0_527# powergood_check/FILLER_2_32/li_353_797# user_to_mprj_oen_buffers\[93\]/li_707_527#
+ mprj_dat_buf\[20\]/li_795_379# la_buf\[23\]/li_207_51# FILLER_17_1829/li_63_527#
+ PHY_14/li_0_527# user_to_mprj_oen_buffers\[37\]/li_983_527# la_buf\[24\]/li_795_379#
+ _387_/li_0_527# user_to_mprj_oen_buffers\[74\]/li_63_n17# powergood_check/FILLER_0_88/li_257_797#
+ ANTENNA_la_buf\[7\]_A/li_63_527# powergood_check/FILLER_1_180/li_161_n17# PHY_45/li_0_n17#
+ FILLER_10_430/li_0_n17# user_to_mprj_oen_buffers\[110\]/li_891_n17# FILLER_22_1663/li_0_n17#
+ FILLER_24_1553/li_0_527# _477_/li_155_527# _546_/li_247_n17# _390_/li_155_n17# FILLER_11_1225/li_63_527#
+ user_to_mprj_in_gates\[94\]/li_0_527# user_to_mprj_oen_buffers\[30\]/li_215_311#
+ PHY_731/li_0_n17# user_to_mprj_in_gates\[74\]/li_339_n17# PHY_402/li_0_n17# mprj_adr_buf\[24\]/li_431_527#
+ user_to_mprj_in_gates\[76\]/li_18_51# user_to_mprj_oen_buffers\[115\]/li_207_51#
+ _606_/li_0_n17# PHY_765/li_0_n17# user_to_mprj_in_gates\[107\]/li_615_527# ANTENNA__609__A/li_63_n17#
+ FILLER_12_685/li_155_527# _567_/li_155_n17# la_buf\[51\]/li_17_51# user_to_mprj_in_gates\[55\]/li_615_n17#
+ ANTENNA_mprj_cyc_buf_A/li_63_n17# mprj_clk2_buf/li_1351_527# ANTENNA__366__A/li_155_527#
+ ANTENNA__590__A/li_63_n17# FILLER_23_1520/li_0_n17# user_to_mprj_oen_buffers\[50\]/li_1075_527#
+ FILLER_22_520/li_63_n17# powergood_check/FILLER_2_16/li_65_n17# user_to_mprj_oen_buffers\[114\]/li_431_527#
+ user_to_mprj_in_gates\[53\]/li_339_527# la_buf\[89\]/li_207_51# powergood_check/FILLER_2_24/li_161_n17#
+ mprj_dat_buf\[3\]/li_707_527# powergood_check/FILLER_2_267/li_353_797# user_to_mprj_oen_buffers\[57\]/li_891_527#
+ user_to_mprj_oen_buffers\[58\]/li_17_51# _482_/li_155_527# FILLER_20_75/li_0_527#
+ FILLER_24_2040/li_63_527# FILLER_15_558/li_0_n17# user_to_mprj_in_buffers\[20\]/li_404_367#
+ user_to_mprj_in_gates\[116\]/li_615_n17# powergood_check/FILLER_1_115/li_115_72#
+ powergood_check/FILLER_1_188/li_65_797# ANTENNA_user_to_mprj_in_gates\[120\]_B/li_63_527#
+ FILLER_21_1335/li_0_527# la_buf\[4\]/li_707_n17# powergood_check/FILLER_0_232/li_0_n17#
+ user_to_mprj_in_buffers\[89\]/li_236_367# user_to_mprj_in_gates\[62\]/li_339_n17#
+ la_buf\[91\]/li_207_51# user_to_mprj_in_buffers\[49\]/li_615_527# user_to_mprj_in_gates\[25\]/li_18_51#
+ ANTENNA__336__A/li_0_527# FILLER_19_1403/li_0_527# ANTENNA__528__A/li_63_527# la_buf\[95\]/li_707_n17#
+ powergood_check/mprj_logic_high_lv/li_514_79# user_to_mprj_in_gates\[123\]/li_339_n17#
+ FILLER_10_1077/li_63_n17# powergood_check/FILLER_1_268/li_641_n17# FILLER_15_1386/li_63_n17#
+ user_to_mprj_oen_buffers\[3\]/li_1443_527# FILLER_10_501/li_0_n17# user_to_mprj_in_gates\[5\]/li_0_527#
+ ANTENNA__337__A/li_63_n17# user_to_mprj_oen_buffers\[83\]/li_1075_n17# _575_/li_0_n17#
+ user_to_mprj_oen_buffers\[45\]/li_795_379# FILLER_25_693/li_155_n17# powergood_check/FILLER_2_259/li_161_n17#
+ la_buf\[67\]/li_1351_527# FILLER_25_891/li_0_n17# FILLER_13_925/li_63_527# _359_/li_247_527#
+ PHY_88/li_0_527# mprj2_pwrgood/li_707_n17# la_buf\[5\]/li_1351_n17# user_to_mprj_in_gates\[88\]/li_615_527#
+ la_buf\[19\]/li_17_51# FILLER_25_1261/li_155_n17# user_to_mprj_in_buffers\[123\]/li_404_17#
+ _351_/li_0_n17# FILLER_13_1820/li_0_527# user_to_mprj_in_gates\[50\]/li_339_n17#
+ user_to_mprj_oen_buffers\[52\]/li_707_527# FILLER_18_1416/li_0_527# _336_/li_247_527#
+ mprj_adr_buf\[24\]/li_215_311# FILLER_11_838/li_63_n17# user_to_mprj_in_gates\[78\]/li_63_n17#
+ user_to_mprj_in_gates\[76\]/li_431_527# _390_/li_0_n17# powergood_check/FILLER_2_32/li_0_n17#
+ FILLER_24_1648/li_0_527# user_to_mprj_oen_buffers\[114\]/li_17_51# user_to_mprj_in_gates\[111\]/li_339_n17#
+ PHY_902/li_0_527# user_to_mprj_in_buffers\[35\]/li_51_367# FILLER_12_1927/li_63_n17#
+ PHY_483/li_0_527# _547_/li_0_n17# user_to_mprj_in_gates\[85\]/li_431_n17# FILLER_13_1021/li_0_n17#
+ mprj_adr_buf\[30\]/li_17_51# FILLER_10_983/li_63_n17# powergood_check/FILLER_2_171/li_0_797#
+ PHY_465/li_0_527# FILLER_23_621/li_155_n17# FILLER_10_1170/li_0_n17# user_to_mprj_in_gates\[83\]/li_155_527#
+ _332_/li_155_n17# powergood_check/FILLER_1_115/li_545_n17# powergood_check/mprj_logic_high_lv/li_1313_1611#
+ powergood_check/FILLER_2_8/li_115_72# FILLER_26_1115/li_0_527# user_to_mprj_oen_buffers\[66\]/li_207_51#
+ FILLER_9_1230/li_0_527# la_buf\[58\]/li_891_527# FILLER_12_1635/li_0_527# PHY_773/li_0_n17#
+ user_to_mprj_in_buffers\[65\]/li_236_367# FILLER_11_2022/li_155_527# user_to_mprj_in_gates\[0\]/li_18_51#
+ mprj_dat_buf\[23\]/li_247_527# FILLER_26_1180/li_0_527# user_to_mprj_in_gates\[64\]/li_431_527#
+ mprj_adr_buf\[12\]/li_215_311# FILLER_22_1408/li_63_527# user_to_mprj_in_gates\[92\]/li_155_n17#
+ user_to_mprj_oen_buffers\[22\]/li_431_527# la_buf\[100\]/li_17_51# la_buf\[53\]/li_0_527#
+ FILLER_21_70/li_0_527# _506_/li_155_n17# powergood_check/FILLER_2_115/li_257_n17#
+ FILLER_21_2101/li_155_n17# user_to_mprj_in_gates\[91\]/li_707_n17# user_to_mprj_in_buffers\[7\]/li_523_n17#
+ powergood_check/FILLER_2_243/li_0_n17# la_buf\[28\]/li_207_51# mprj_adr_buf\[3\]/li_17_51#
+ FILLER_17_1428/li_155_527# FILLER_22_1653/li_0_n17# user_to_mprj_in_gates\[73\]/li_431_n17#
+ la_buf\[119\]/li_17_51# FILLER_11_1717/li_155_n17# PHY_489/li_0_527# _537_/li_0_527#
+ user_to_mprj_in_gates\[71\]/li_155_527# _331_/li_247_n17# powergood_check/FILLER_1_16/li_0_n17#
+ FILLER_25_1035/li_0_n17# PHY_831/li_0_n17# powergood_check/FILLER_2_155/li_545_n17#
+ user_to_mprj_in_buffers\[8\]/li_51_17# PHY_280/li_0_n17# FILLER_22_515/li_0_527#
+ FILLER_15_502/li_0_527# FILLER_8_1896/li_63_527# la_buf\[86\]/li_1351_527# FILLER_15_62/li_155_n17#
+ mprj_dat_buf\[23\]/li_17_51# powergood_check/FILLER_1_8/li_0_n17# FILLER_18_1556/li_0_527#
+ la_buf\[30\]/li_207_51# PHY_359/li_0_527# user_to_mprj_oen_buffers\[81\]/li_63_n17#
+ user_to_mprj_in_gates\[52\]/li_431_527# FILLER_14_528/li_63_527# FILLER_14_1537/li_0_527#
+ mprj2_vdd_pwrgood/li_19_289# FILLER_14_1647/li_63_n17# FILLER_16_113/li_0_527# powergood_check/FILLER_1_204/li_100_536#
+ powergood_check/FILLER_1_16/li_161_n17# user_to_mprj_oen_buffers\[60\]/li_1167_n17#
+ FILLER_19_2061/li_63_527# user_to_mprj_in_buffers\[109\]/li_615_n17# powergood_check/FILLER_0_264/li_0_n17#
+ FILLER_24_307/li_0_n17# la_buf\[11\]/li_779_17# mprj_adr_buf\[28\]/li_431_527# la_buf\[94\]/li_215_311#
+ FILLER_25_819/li_63_n17# powergood_check/FILLER_0_96/li_100_536# user_to_mprj_oen_buffers\[91\]/li_1075_n17#
+ la_buf\[58\]/li_0_527# FILLER_25_1265/li_155_527# user_to_mprj_oen_buffers\[122\]/li_207_51#
+ FILLER_14_1510/li_0_527# _391_/li_0_527# mprj_clk2_buf/li_0_527# la_buf\[24\]/li_247_n17#
+ _574_/li_155_n17# user_to_mprj_oen_buffers\[5\]/li_615_527# PHY_813/li_0_527# la_buf\[43\]/li_63_n17#
+ FILLER_18_1782/li_0_n17# PHY_708/li_0_527# powergood_check/mprj2_logic_high_lv/li_506_1123#
+ FILLER_25_1004/li_0_n17# powergood_check/FILLER_0_96/li_449_797# user_to_mprj_in_buffers\[41\]/li_236_367#
+ FILLER_25_746/li_63_n17# la_buf\[96\]/li_207_51# FILLER_25_1107/li_155_n17# user_to_mprj_in_gates\[122\]/li_431_n17#
+ la_buf\[70\]/li_247_527# FILLER_12_1103/li_63_527# user_to_mprj_in_gates\[75\]/li_18_51#
+ user_to_mprj_in_gates\[120\]/li_155_527# FILLER_13_777/li_155_527# user_to_mprj_oen_buffers\[48\]/li_247_527#
+ user_to_mprj_oen_buffers\[48\]/li_63_527# _336_/li_0_527# FILLER_16_1585/li_155_527#
+ user_to_mprj_in_buffers\[39\]/li_404_17# la_buf\[77\]/li_779_17# mprj_adr_buf\[8\]/li_707_n17#
+ la_buf\[50\]/li_17_51# powergood_check/FILLER_2_235/li_257_797# FILLER_21_1558/li_155_n17#
+ _366_/li_0_527# la_buf\[82\]/li_215_311# powergood_check/FILLER_0_248/li_65_797#
+ FILLER_9_611/li_63_527# PHY_341/li_0_n17# la_buf\[56\]/li_615_527# user_to_mprj_oen_buffers\[41\]/li_611_17#
+ user_to_mprj_oen_buffers\[57\]/li_17_51# user_to_mprj_oen_buffers\[50\]/li_63_527#
+ powergood_check/FILLER_0_104/li_641_797# FILLER_18_528/li_63_527# la_buf\[98\]/li_983_n17#
+ _399_/li_0_n17# la_buf\[69\]/li_17_51# powergood_check/FILLER_2_32/li_353_n17# FILLER_28_55/li_0_527#
+ _569_/li_0_527# user_to_mprj_in_buffers\[9\]/li_236_367# mprj_adr_buf\[15\]/li_795_379#
+ powergood_check/mprj_logic_high_lv/li_34_216# FILLER_16_1581/li_155_527# PHY_311/li_0_527#
+ user_to_mprj_in_buffers\[102\]/li_404_367# user_to_mprj_in_gates\[69\]/li_0_n17#
+ user_to_mprj_in_gates\[78\]/li_247_527# PHY_75/li_0_n17# FILLER_18_1439/li_0_n17#
+ FILLER_11_728/li_155_527# powergood_check/FILLER_2_195/li_353_797# user_to_mprj_in_gates\[24\]/li_18_51#
+ powergood_check/FILLER_1_236/li_545_n17# FILLER_12_1543/li_0_527# _568_/li_0_527#
+ ANTENNA_user_to_mprj_in_gates\[34\]_A/li_63_n17# FILLER_15_1928/li_0_527# powergood_check/FILLER_0_256/li_257_797#
+ FILLER_9_1234/li_63_527# _543_/li_155_527# FILLER_9_563/li_155_n17# FILLER_19_44/li_0_527#
+ PHY_834/li_0_527# la_buf\[70\]/li_215_311# la_buf\[31\]/li_1351_527# ANTENNA__359__A/li_63_n17#
+ powergood_check/FILLER_0_160/li_0_n17# la_buf\[13\]/li_0_527# FILLER_12_1039/li_0_n17#
+ _565_/li_0_n17# la_buf\[6\]/li_779_17# la_buf\[44\]/li_615_527# user_to_mprj_in_gates\[85\]/li_63_n17#
+ user_to_mprj_oen_buffers\[59\]/li_891_n17# FILLER_17_547/li_0_n17# _393_/li_247_n17#
+ la_buf\[2\]/li_1443_n17# mprj_dat_buf\[25\]/li_215_311# FILLER_18_1961/li_63_527#
+ FILLER_13_1177/li_0_527# la_buf\[29\]/li_215_311# _334_/li_155_n17# FILLER_22_1559/li_63_527#
+ user_to_mprj_in_buffers\[42\]/li_51_367# la_buf\[18\]/li_17_51# _469_/li_247_n17#
+ ANTENNA__348__A/li_0_n17# la_buf\[45\]/li_1535_527# powergood_check/FILLER_2_267/li_353_n17#
+ _341_/li_0_n17# powergood_check/FILLER_1_196/li_641_n17# powergood_check/mprj_logic_high_lv/li_353_1611#
+ la_buf\[42\]/li_1351_527# user_to_mprj_in_gates\[66\]/li_247_527# PHY_493/li_0_527#
+ mprj_dat_buf\[3\]/li_207_51# powergood_check/FILLER_0_16/li_353_797# user_to_mprj_oen_buffers\[24\]/li_247_527#
+ FILLER_16_593/li_155_527# powergood_check/FILLER_0_32/li_65_797# PHY_783/li_0_n17#
+ user_to_mprj_oen_buffers\[20\]/li_63_n17# powergood_check/FILLER_2_187/li_161_n17#
+ la_buf\[78\]/li_63_527# FILLER_18_1945/li_155_527# FILLER_11_1569/li_63_n17# PHY_720/li_0_527#
+ user_to_mprj_oen_buffers\[56\]/li_1075_n17# _423_/li_155_527# user_to_mprj_in_gates\[127\]/li_247_527#
+ user_to_mprj_oen_buffers\[73\]/li_207_51# la_buf\[106\]/li_0_n17# user_to_mprj_oen_buffers\[113\]/li_17_51#
+ user_to_mprj_oen_buffers\[3\]/li_1075_527# FILLER_13_699/li_0_527# FILLER_9_512/li_155_n17#
+ FILLER_22_1771/li_0_n17# powergood_check/FILLER_0_0/li_161_797# la_buf\[99\]/li_611_17#
+ user_to_mprj_in_gates\[75\]/li_247_n17# FILLER_13_106/li_0_527# powergood_check/FILLER_1_252/li_0_797#
+ FILLER_25_1896/li_63_n17# mprj_dat_buf\[13\]/li_215_311# FILLER_10_505/li_0_n17#
+ la_buf\[17\]/li_215_311# ANTENNA__397__A/li_63_n17# FILLER_21_1451/li_63_527# FILLER_14_1696/li_155_527#
+ la_buf\[86\]/li_431_527# FILLER_11_1394/li_63_n17# FILLER_21_1985/li_155_n17# FILLER_11_992/li_155_n17#
+ la_buf\[76\]/li_1443_n17# FILLER_25_895/li_0_n17# user_to_mprj_oen_buffers\[118\]/li_215_311#
+ user_to_mprj_in_gates\[56\]/li_523_n17# la_buf\[35\]/li_207_51# user_to_mprj_in_gates\[54\]/li_247_527#
+ user_to_mprj_oen_buffers\[86\]/li_63_n17# mprj_sel_buf\[3\]/li_795_379# FILLER_9_171/li_63_n17#
+ FILLER_9_600/li_63_n17# FILLER_9_888/li_63_527# FILLER_24_616/li_0_527# PHY_446/li_0_527#
+ la_buf\[85\]/li_63_527# user_to_mprj_in_buffers\[93\]/li_404_367# _380_/li_247_527#
+ user_to_mprj_in_gates\[127\]/li_18_51# user_to_mprj_oen_buffers\[59\]/li_1259_n17#
+ la_buf\[109\]/li_63_n17# FILLER_4_905/li_0_527# user_to_mprj_in_buffers\[115\]/li_51_17#
+ user_to_mprj_oen_buffers\[91\]/li_215_311# FILLER_11_744/li_63_527# PHY_59/li_0_527#
+ la_buf\[7\]/li_63_527# FILLER_21_1436/li_155_527# FILLER_23_1670/li_155_527# mprj_dat_buf\[1\]/li_891_527#
+ user_to_mprj_oen_buffers\[127\]/li_207_51# mprj_adr_buf\[2\]/li_17_51# la_buf\[118\]/li_17_51#
+ PHY_35/li_0_527# FILLER_12_890/li_0_n17# FILLER_12_839/li_63_n17# PHY_296/li_0_n17#
+ FILLER_5_967/li_63_527# _579_/li_155_n17# la_buf\[48\]/li_63_n17# _491_/li_155_527#
+ FILLER_15_1802/li_0_527# PHY_5/li_0_n17# user_to_mprj_in_gates\[124\]/li_247_n17#
+ FILLER_0_87/li_155_527# _415_/li_0_527# user_to_mprj_in_buffers\[7\]/li_51_17# PHY_326/li_0_n17#
+ FILLER_27_806/li_63_n17# FILLER_3_893/li_0_n17# user_to_mprj_oen_buffers\[106\]/li_215_311#
+ FILLER_13_2020/li_63_n17# FILLER_8_1221/li_0_527# PHY_779/li_0_527# la_buf\[95\]/li_1167_527#
+ mprj_dat_buf\[29\]/li_431_527# mprj_dat_buf\[22\]/li_17_51# FILLER_5_743/li_63_527#
+ FILLER_14_1571/li_63_527# powergood_check/FILLER_2_171/li_0_n17# FILLER_25_1208/li_0_527#
+ FILLER_15_1441/li_0_n17# _369_/li_155_527# la_buf\[25\]/li_0_527# FILLER_26_450/li_0_527#
+ FILLER_12_1923/li_63_527# ANTENNA__644__A/li_63_n17# ANTENNA_user_to_mprj_in_gates\[52\]_A/li_63_527#
+ _581_/li_155_n17# user_to_mprj_oen_buffers\[23\]/li_0_527# user_to_mprj_in_gates\[105\]/li_523_n17#
+ la_buf\[50\]/li_63_n17# user_to_mprj_in_gates\[31\]/li_615_n17# user_to_mprj_in_gates\[103\]/li_247_527#
+ user_to_mprj_oen_buffers\[40\]/li_1075_n17# FILLER_12_1357/li_63_n17# FILLER_23_625/li_63_527#
+ _475_/li_0_527# user_to_mprj_oen_buffers\[110\]/li_779_17# FILLER_11_1186/li_0_n17#
+ user_to_mprj_in_gates\[51\]/li_247_n17# FILLER_15_1437/li_63_527# PHY_732/li_0_527#
+ PHY_323/li_0_527# FILLER_7_1148/li_155_527# _591_/li_0_527# powergood_check/FILLER_1_24/li_353_n17#
+ powergood_check/FILLER_1_268/li_161_n17# FILLER_19_1634/li_63_n17# PHY_317/li_0_n17#
+ _381_/li_0_527# user_to_mprj_in_gates\[24\]/li_63_n17# ANTENNA_user_to_mprj_oen_buffers\[7\]_TE/li_63_527#
+ mprj_sel_buf\[2\]/li_431_527# user_to_mprj_oen_buffers\[38\]/li_215_311# FILLER_17_1925/li_155_527#
+ powergood_check/FILLER_0_176/li_115_72# ANTENNA__589__A/li_63_527# la_buf\[75\]/li_63_527#
+ user_to_mprj_in_gates\[110\]/li_0_527# user_to_mprj_in_buffers\[46\]/li_404_17#
+ la_buf\[84\]/li_779_17# PHY_831/li_0_527# FILLER_20_2087/li_0_n17# FILLER_14_1673/li_63_527#
+ FILLER_13_1931/li_63_n17# user_to_mprj_in_gates\[112\]/li_247_n17# user_to_mprj_in_gates\[97\]/li_707_367#
+ user_to_mprj_in_buffers\[24\]/li_339_n17# PHY_774/li_0_n17# la_buf\[98\]/li_1167_n17#
+ la_buf\[35\]/li_1351_527# user_to_mprj_in_gates\[30\]/li_247_527# PHY_175/li_0_n17#
+ user_to_mprj_in_gates\[74\]/li_18_51# FILLER_18_63/li_63_527# _393_/li_0_527# FILLER_9_825/li_63_527#
+ la_buf\[72\]/li_431_527# ANTENNA__333__A/li_63_527# FILLER_10_578/li_0_n17# powergood_check/FILLER_2_243/li_100_536#
+ _548_/li_155_527# la_buf\[17\]/li_63_527# PHY_781/li_0_n17# _632_/li_0_n17# PHY_706/li_0_n17#
+ FILLER_9_390/li_0_n17# PHY_394/li_0_n17# FILLER_26_969/li_0_527# user_to_mprj_in_gates\[104\]/li_431_n17#
+ PHY_43/li_0_527# user_to_mprj_oen_buffers\[12\]/li_207_51# la_buf\[113\]/li_795_379#
+ user_to_mprj_oen_buffers\[87\]/li_1075_527# PHY_159/li_0_n17# mprj_adr_buf\[2\]/li_523_n17#
+ la_buf\[6\]/li_1443_527# FILLER_9_1038/li_63_527# _634_/li_247_527# FILLER_19_1573/li_155_n17#
+ user_to_mprj_oen_buffers\[56\]/li_17_51# powergood_check/FILLER_2_243/li_449_797#
+ mprj_dat_buf\[27\]/li_1075_527# _339_/li_155_n17# user_to_mprj_oen_buffers\[26\]/li_215_311#
+ _638_/li_155_n17# la_buf\[68\]/li_17_51# user_to_mprj_oen_buffers\[109\]/li_63_527#
+ mprj_dat_buf\[23\]/li_707_527# la_buf\[50\]/li_431_527# PHY_739/li_0_n17# user_to_mprj_in_gates\[100\]/li_247_n17#
+ FILLER_21_1989/li_0_n17# FILLER_11_996/li_63_527# FILLER_14_491/li_63_n17# user_to_mprj_in_gates\[92\]/li_615_n17#
+ mprj_dat_buf\[8\]/li_207_51# powergood_check/FILLER_2_163/li_257_797# user_to_mprj_in_gates\[90\]/li_339_527#
+ FILLER_17_530/li_0_527# powergood_check/FILLER_0_208/li_65_n17# user_to_mprj_in_gates\[92\]/li_63_n17#
+ PHY_261/li_0_527# powergood_check/FILLER_0_264/li_100_536# user_to_mprj_in_gates\[23\]/li_18_51#
+ user_to_mprj_in_buffers\[18\]/li_0_527# FILLER_18_2110/li_155_527# FILLER_14_1571/li_155_527#
+ _341_/li_155_n17# FILLER_15_2107/li_63_527# user_to_mprj_oen_buffers\[78\]/li_207_51#
+ user_to_mprj_in_gates\[49\]/li_339_527# powergood_check/FILLER_0_96/li_449_n17#
+ _641_/li_155_n17# FILLER_18_1463/li_155_n17# user_to_mprj_in_gates\[71\]/li_615_527#
+ powergood_check/FILLER_2_24/li_0_797# FILLER_20_200/li_0_n17# FILLER_19_2000/li_155_n17#
+ powergood_check/FILLER_0_264/li_449_797# _555_/li_0_n17# FILLER_11_728/li_0_527#
+ user_to_mprj_oen_buffers\[109\]/li_795_379# user_to_mprj_oen_buffers\[59\]/li_779_17#
+ la_buf\[88\]/li_247_527# la_buf\[89\]/li_0_n17# user_to_mprj_oen_buffers\[122\]/li_1351_527#
+ mprj_sel_buf\[1\]/li_707_n17# user_to_mprj_oen_buffers\[14\]/li_215_311# FILLER_17_1570/li_0_527#
+ powergood_check/FILLER_2_235/li_257_n17# powergood_check/FILLER_1_164/li_545_n17#
+ user_to_mprj_oen_buffers\[119\]/li_431_n17# la_buf\[68\]/li_0_527# user_to_mprj_oen_buffers\[80\]/li_207_51#
+ powergood_check/FILLER_0_184/li_257_797# _594_/li_0_n17# la_buf\[17\]/li_17_51#
+ FILLER_3_763/li_0_527# FILLER_7_810/li_63_527# _659_/li_0_n17# FILLER_12_1374/li_155_527#
+ _482_/li_0_n17# FILLER_12_1796/li_63_527# user_to_mprj_in_buffers\[104\]/li_615_n17#
+ la_buf\[103\]/li_207_51# ANTENNA_user_to_mprj_in_gates\[73\]_A/li_63_n17# user_to_mprj_oen_buffers\[91\]/li_1535_n17#
+ powergood_check/FILLER_1_0/li_257_n17# ANTENNA__574__A/li_63_n17# FILLER_11_728/li_63_527#
+ _607_/li_155_527# user_to_mprj_oen_buffers\[69\]/li_707_n17# powergood_check/FILLER_0_24/li_545_797#
+ la_buf\[24\]/li_707_n17# FILLER_25_1158/li_0_n17# FILLER_18_1899/li_63_527# user_to_mprj_oen_buffers\[112\]/li_17_51#
+ PHY_290/li_0_n17# powergood_check/FILLER_2_195/li_353_n17# la_buf\[42\]/li_207_51#
+ _342_/li_247_n17# mprj_we_buf/li_17_51# user_to_mprj_in_buffers\[3\]/li_155_n17#
+ FILLER_11_413/li_155_527# la_buf\[91\]/li_0_527# user_to_mprj_in_gates\[16\]/li_0_527#
+ FILLER_13_507/li_63_527# powergood_check/FILLER_2_243/li_115_72# FILLER_9_407/li_0_n17#
+ FILLER_23_1629/li_0_527# FILLER_19_1577/li_0_527# user_to_mprj_in_gates\[61\]/li_707_367#
+ la_buf\[116\]/li_63_n17# _635_/li_0_527# FILLER_9_670/li_0_527# user_to_mprj_oen_buffers\[22\]/li_779_17#
+ powergood_check/mprj_logic_high_lv/li_26_452# la_buf\[59\]/li_1075_n17# user_to_mprj_oen_buffers\[18\]/li_983_n17#
+ FILLER_13_2020/li_63_527# FILLER_9_440/li_155_n17# FILLER_25_1502/li_0_n17# FILLER_6_711/li_0_527#
+ PHY_417/li_0_527# la_buf\[85\]/li_779_17# _586_/li_155_n17# FILLER_21_1695/li_63_527#
+ powergood_check/FILLER_2_203/li_641_797# user_to_mprj_in_gates\[122\]/li_707_367#
+ PHY_310/li_0_527# ANTENNA__562__A/li_63_n17# _443_/li_247_527# user_to_mprj_oen_buffers\[57\]/li_707_n17#
+ la_buf\[49\]/li_1535_n17# user_to_mprj_in_gates\[126\]/li_18_51# la_buf\[12\]/li_707_n17#
+ user_to_mprj_oen_buffers\[29\]/li_795_379# _597_/li_0_n17# FILLER_25_303/li_0_527#
+ _630_/li_0_527# FILLER_20_1421/li_155_n17# FILLER_15_335/li_0_527# user_to_mprj_oen_buffers\[103\]/li_1167_n17#
+ mprj_adr_buf\[1\]/li_17_51# FILLER_11_1817/li_63_527# FILLER_9_416/li_63_n17# la_buf\[117\]/li_17_51#
+ powergood_check/FILLER_1_62/li_641_797# la_buf\[89\]/li_779_17# FILLER_19_249/li_63_n17#
+ PHY_736/li_0_527# user_to_mprj_in_gates\[34\]/li_339_n17# FILLER_11_1196/li_63_527#
+ powergood_check/FILLER_0_192/li_0_797# FILLER_12_689/li_63_n17# _405_/li_0_527#
+ user_to_mprj_in_buffers\[6\]/li_51_17# FILLER_19_1742/li_155_527# powergood_check/FILLER_0_104/li_161_797#
+ powergood_check/FILLER_1_252/li_0_n17# powergood_check/FILLER_1_172/li_65_n17# _556_/li_0_527#
+ user_to_mprj_in_gates\[88\]/li_155_n17# FILLER_5_609/li_155_527# PHY_361/li_0_n17#
+ mprj_dat_buf\[21\]/li_17_51# FILLER_12_1527/li_0_527# powergood_check/FILLER_0_224/li_641_797#
+ FILLER_9_1273/li_0_527# FILLER_26_43/li_63_n17# FILLER_25_1219/li_0_n17# user_to_mprj_in_gates\[31\]/li_63_n17#
+ powergood_check/FILLER_1_8/li_545_n17# FILLER_25_899/li_0_n17# FILLER_13_1502/li_0_527#
+ user_to_mprj_in_gates\[110\]/li_707_367# mprj_adr_buf\[2\]/li_215_311# FILLER_13_585/li_0_527#
+ FILLER_17_1925/li_63_n17# user_to_mprj_oen_buffers\[17\]/li_207_51# user_to_mprj_oen_buffers\[83\]/li_611_17#
+ PHY_751/li_0_n17# _332_/li_0_527# FILLER_11_1196/li_155_n17# PHY_840/li_0_n17# user_to_mprj_in_gates\[69\]/li_431_n17#
+ user_to_mprj_in_buffers\[90\]/li_236_367# _483_/li_0_527# PHY_227/li_0_527# FILLER_23_324/li_0_527#
+ mprj_adr_buf\[29\]/li_1443_527# FILLER_23_1915/li_63_527# user_to_mprj_in_gates\[52\]/li_339_n17#
+ _555_/li_155_527# la_buf\[24\]/li_63_527# powergood_check/mprj2_logic_high_lv/li_1217_1611#
+ user_to_mprj_in_buffers\[49\]/li_236_367# FILLER_18_170/li_63_527# powergood_check/FILLER_1_32/li_545_n17#
+ powergood_check/FILLER_2_203/li_65_n17# user_to_mprj_oen_buffers\[5\]/li_1167_527#
+ la_buf\[101\]/li_707_527# FILLER_16_1449/li_0_n17# FILLER_16_508/li_63_n17# PHY_9/li_0_n17#
+ user_to_mprj_in_gates\[73\]/li_18_51# FILLER_23_324/li_63_527# FILLER_16_2069/li_0_527#
+ powergood_check/FILLER_1_196/li_161_n17# _346_/li_155_n17# FILLER_18_1416/li_155_527#
+ _645_/li_155_n17# user_to_mprj_in_gates\[2\]/li_707_367# ANTENNA_user_to_mprj_in_gates\[39\]_A/li_63_527#
+ FILLER_26_1247/li_63_527# powergood_check/mprj2_logic_high_lv/li_545_1611# FILLER_23_625/li_0_n17#
+ PHY_291/li_0_n17# FILLER_10_2082/li_63_n17# PHY_375/li_0_527# user_to_mprj_in_gates\[57\]/li_431_n17#
+ mprj_adr_buf\[14\]/li_207_51# powergood_check/FILLER_2_0/li_353_797# user_to_mprj_oen_buffers\[22\]/li_611_17#
+ FILLER_21_1638/li_0_527# user_to_mprj_oen_buffers\[55\]/li_17_51# FILLER_11_196/li_0_527#
+ user_to_mprj_oen_buffers\[85\]/li_207_51# FILLER_10_55/li_155_527# ANTENNA_la_buf\[110\]_TE/li_63_n17#
+ powergood_check/FILLER_2_171/li_100_536# la_buf\[67\]/li_17_51# PHY_327/li_0_527#
+ la_buf\[1\]/li_611_17# FILLER_18_335/li_0_527# FILLER_13_1067/li_0_527# la_buf\[4\]/li_247_527#
+ powergood_check/FILLER_1_236/li_115_72# FILLER_16_1601/li_63_n17# mprj_dat_buf\[23\]/li_1075_527#
+ la_buf\[108\]/li_207_51# user_to_mprj_oen_buffers\[42\]/li_1075_527# user_to_mprj_in_gates\[22\]/li_18_51#
+ mprj_sel_buf\[3\]/li_17_51# _357_/li_0_527# powergood_check/FILLER_2_171/li_449_797#
+ user_to_mprj_in_buffers\[2\]/li_236_17# la_buf\[78\]/li_215_311# user_to_mprj_oen_buffers\[85\]/li_1167_n17#
+ PHY_365/li_0_527# la_buf\[47\]/li_207_51# FILLER_25_1265/li_63_527# user_to_mprj_in_gates\[45\]/li_431_n17#
+ user_to_mprj_in_gates\[48\]/li_707_n17# user_to_mprj_in_buffers\[13\]/li_236_17#
+ user_to_mprj_in_gates\[124\]/li_707_n17# la_buf\[110\]/li_207_51# la_buf\[118\]/li_891_527#
+ FILLER_22_1653/li_63_527# powergood_check/FILLER_0_192/li_100_536# FILLER_20_567/li_0_527#
+ la_buf\[114\]/li_523_n17# la_buf\[28\]/li_779_17# la_buf\[21\]/li_1075_527# FILLER_13_1013/li_0_527#
+ _584_/li_0_n17# la_buf\[99\]/li_1075_527# la_buf\[16\]/li_17_51# FILLER_23_2106/li_155_527#
+ FILLER_25_1075/li_0_n17# la_buf\[6\]/li_891_527# _335_/li_247_527# FILLER_21_1440/li_0_n17#
+ powergood_check/FILLER_1_180/li_0_n17# powergood_check/FILLER_2_243/li_449_n17#
+ FILLER_13_1812/li_0_527# user_to_mprj_oen_buffers\[82\]/li_247_n17# powergood_check/FILLER_0_192/li_449_797#
+ user_to_mprj_in_gates\[51\]/li_707_n17# FILLER_15_554/li_0_527# la_buf\[51\]/li_891_n17#
+ _360_/li_0_n17# la_buf\[66\]/li_215_311# la_buf\[123\]/li_63_n17# FILLER_13_973/li_63_527#
+ powergood_check/FILLER_2_163/li_257_n17# powergood_check/mprj2_logic_high_lv/li_1601_1611#
+ FILLER_25_1019/li_0_n17# user_to_mprj_oen_buffers\[111\]/li_17_51# FILLER_23_1678/li_63_527#
+ powergood_check/FILLER_2_8/li_641_797# user_to_mprj_oen_buffers\[3\]/li_215_311#
+ user_to_mprj_in_gates\[31\]/li_155_527# user_to_mprj_in_gates\[112\]/li_707_n17#
+ FILLER_13_1279/li_0_527# user_to_mprj_oen_buffers\[67\]/li_983_527# la_buf\[14\]/li_891_527#
+ powergood_check/FILLER_0_32/li_737_797# FILLER_9_615/li_0_527# powergood_check/FILLER_2_24/li_0_n17#
+ FILLER_26_389/li_63_527# FILLER_0_58/li_155_527# la_buf\[92\]/li_795_379# user_to_mprj_in_gates\[40\]/li_155_n17#
+ user_to_mprj_in_gates\[36\]/li_63_n17# PHY_839/li_0_n17# FILLER_23_1919/li_0_527#
+ FILLER_5_964/li_0_527# FILLER_9_1352/li_0_527# powergood_check/FILLER_2_187/li_0_797#
+ powergood_check/FILLER_1_252/li_100_536# user_to_mprj_oen_buffers\[99\]/li_215_311#
+ FILLER_5_1775/li_155_527# user_to_mprj_oen_buffers\[88\]/li_611_17# ANTENNA_user_to_mprj_in_gates\[72\]_B/li_63_n17#
+ la_buf\[54\]/li_215_311# powergood_check/FILLER_2_16/li_115_72# ANTENNA__359__A/li_0_n17#
+ FILLER_28_55/li_63_n17# user_to_mprj_in_gates\[125\]/li_18_51# user_to_mprj_in_gates\[101\]/li_155_n17#
+ FILLER_24_512/li_0_n17# FILLER_21_1573/li_63_527# FILLER_12_1440/li_0_n17# powergood_check/FILLER_2_0/li_0_797#
+ _469_/li_0_n17# PHY_811/li_0_527# PHY_461/li_0_527# user_to_mprj_in_gates\[91\]/li_247_527#
+ FILLER_5_1196/li_63_527# user_to_mprj_in_gates\[100\]/li_707_n17# mprj_adr_buf\[0\]/li_17_51#
+ _473_/li_155_n17# la_buf\[29\]/li_63_527# powergood_check/FILLER_2_251/li_545_797#
+ la_buf\[89\]/li_0_527# PHY_294/li_0_n17# FILLER_12_1623/li_63_n17# la_buf\[116\]/li_17_51#
+ _507_/li_0_527# user_to_mprj_in_buffers\[6\]/li_615_527# la_buf\[26\]/li_1443_n17#
+ user_to_mprj_oen_buffers\[90\]/li_611_17# user_to_mprj_oen_buffers\[24\]/li_207_51#
+ mprj_dat_buf\[23\]/li_779_17# FILLER_15_1609/li_0_n17# la_buf\[102\]/li_891_527#
+ FILLER_11_581/li_63_n17# FILLER_25_1103/li_63_n17# user_to_mprj_in_gates\[55\]/li_0_527#
+ PHY_794/li_0_n17# la_buf\[95\]/li_1351_n17# FILLER_25_953/li_155_n17# FILLER_9_596/li_63_n17#
+ mprj_dat_buf\[20\]/li_17_51# FILLER_14_518/li_0_n17# user_to_mprj_oen_buffers\[62\]/li_1259_n17#
+ la_buf\[101\]/li_0_527# _562_/li_155_527# FILLER_9_600/li_0_n17# user_to_mprj_oen_buffers\[87\]/li_215_311#
+ la_buf\[31\]/li_63_527# powergood_check/FILLER_0_112/li_353_797# la_buf\[34\]/li_0_527#
+ la_buf\[42\]/li_215_311# ANTENNA__657__A/li_0_n17# user_to_mprj_in_gates\[59\]/li_247_n17#
+ la_buf\[122\]/li_1259_n17# PHY_815/li_0_527# mprj_adr_buf\[19\]/li_207_51# la_buf\[126\]/li_215_311#
+ user_to_mprj_oen_buffers\[37\]/li_0_n17# user_to_mprj_in_buffers\[67\]/li_155_n17#
+ FILLER_9_407/li_155_n17# FILLER_16_1425/li_0_527# la_buf\[6\]/li_215_311# powergood_check/FILLER_2_203/li_641_n17#
+ la_buf\[84\]/li_1167_n17# FILLER_13_1052/li_0_527# _353_/li_155_n17# user_to_mprj_oen_buffers\[54\]/li_0_527#
+ _361_/li_0_527# _592_/li_0_n17# _652_/li_155_n17# user_to_mprj_in_buffers\[60\]/li_0_527#
+ powergood_check/FILLER_2_16/li_257_797# user_to_mprj_oen_buffers\[123\]/li_63_527#
+ PHY_498/li_0_527# powergood_check/FILLER_1_244/li_257_n17# FILLER_16_508/li_0_n17#
+ user_to_mprj_in_gates\[38\]/li_247_527# user_to_mprj_oen_buffers\[7\]/li_431_527#
+ la_buf\[10\]/li_0_n17# _343_/li_247_527# ANTENNA_la_buf\[123\]_A/li_63_n17# FILLER_10_804/li_155_527#
+ mprj_adr_buf\[21\]/li_207_51# user_to_mprj_in_buffers\[77\]/li_404_367# powergood_check/FILLER_1_62/li_641_n17#
+ FILLER_24_56/li_0_n17# FILLER_17_108/li_63_527# user_to_mprj_in_gates\[30\]/li_707_n17#
+ user_to_mprj_in_gates\[72\]/li_18_51# user_to_mprj_oen_buffers\[60\]/li_891_n17#
+ user_to_mprj_in_gates\[98\]/li_431_527# user_to_mprj_in_buffers\[7\]/li_236_17#
+ _440_/li_0_527# user_to_mprj_oen_buffers\[92\]/li_207_51# user_to_mprj_oen_buffers\[75\]/li_215_311#
+ user_to_mprj_in_buffers\[3\]/li_615_n17# la_buf\[30\]/li_215_311# powergood_check/FILLER_0_104/li_161_n17#
+ FILLER_5_609/li_63_527# user_to_mprj_in_gates\[47\]/li_247_n17# user_to_mprj_oen_buffers\[37\]/li_63_527#
+ user_to_mprj_in_buffers\[18\]/li_236_17# la_buf\[114\]/li_215_311# FILLER_21_1889/li_63_527#
+ _382_/li_247_n17# user_to_mprj_oen_buffers\[9\]/li_17_51# FILLER_16_1927/li_63_n17#
+ la_buf\[115\]/li_207_51# _363_/li_0_n17# FILLER_22_1559/li_63_n17# FILLER_14_1692/li_63_527#
+ user_to_mprj_oen_buffers\[54\]/li_17_51# user_to_mprj_in_gates\[87\]/li_707_n17#
+ FILLER_16_548/li_0_n17# FILLER_12_597/li_0_527# mprj_dat_buf\[30\]/li_1535_527#
+ user_to_mprj_in_gates\[28\]/li_523_n17# mprj_dat_buf\[2\]/li_215_311# user_to_mprj_in_gates\[98\]/li_339_527#
+ user_to_mprj_in_gates\[26\]/li_247_527# la_buf\[66\]/li_17_51# la_buf\[54\]/li_207_51#
+ FILLER_14_2009/li_0_527# mprj_adr_buf\[22\]/li_1535_527# la_buf\[57\]/li_795_379#
+ user_to_mprj_in_buffers\[63\]/li_51_367# powergood_check/FILLER_1_48/li_65_797#
+ FILLER_25_1261/li_0_n17# user_to_mprj_oen_buffers\[7\]/li_1351_527# FILLER_8_1265/li_63_n17#
+ la_buf\[67\]/li_431_n17# FILLER_13_1603/li_0_n17# la_buf\[109\]/li_983_527# mprj_sel_buf\[2\]/li_17_51#
+ ANTENNA_user_to_mprj_in_gates\[120\]_A/li_63_527# user_to_mprj_oen_buffers\[63\]/li_215_311#
+ user_to_mprj_in_gates\[21\]/li_18_51# PHY_487/li_0_527# la_buf\[35\]/li_779_17#
+ FILLER_15_1692/li_0_n17# powergood_check/FILLER_0_184/li_65_797# user_to_mprj_oen_buffers\[37\]/li_615_527#
+ user_to_mprj_in_gates\[39\]/li_707_n17# FILLER_16_1415/li_0_527# _647_/li_0_n17#
+ user_to_mprj_in_buffers\[87\]/li_523_527# la_buf\[77\]/li_1351_n17# la_buf\[102\]/li_215_311#
+ powergood_check/FILLER_1_204/li_65_797# FILLER_10_1188/li_63_n17# ANTENNA__607__A/li_63_527#
+ ANTENNA__357__A/li_63_n17# PHY_469/li_0_n17# user_to_mprj_in_gates\[9\]/li_707_n17#
+ user_to_mprj_in_gates\[88\]/li_615_n17# _620_/li_0_527# PHY_732/li_0_n17# FILLER_11_996/li_155_n17#
+ FILLER_20_2087/li_63_527# _574_/li_0_n17# la_buf\[15\]/li_17_51# powergood_check/FILLER_2_0/li_353_n17#
+ user_to_mprj_in_buffers\[99\]/li_615_n17# la_buf\[45\]/li_795_379# user_to_mprj_in_buffers\[111\]/li_615_527#
+ powergood_check/FILLER_1_62/li_161_797# FILLER_16_88/li_63_527# user_to_mprj_in_buffers\[53\]/li_404_367#
+ mprj_dat_buf\[14\]/li_207_51# FILLER_20_1625/li_155_527# user_to_mprj_in_buffers\[53\]/li_51_17#
+ mprj_dat_buf\[4\]/li_63_527# user_to_mprj_oen_buffers\[51\]/li_215_311# _350_/li_0_n17#
+ user_to_mprj_in_gates\[95\]/li_339_n17# FILLER_25_1502/li_63_527# user_to_mprj_in_gates\[1\]/li_523_527#
+ powergood_check/FILLER_0_224/li_161_797# user_to_mprj_oen_buffers\[110\]/li_17_51#
+ FILLER_13_760/li_0_527# PHY_47/li_0_527# _535_/li_247_527# mprj_dat_buf\[30\]/li_431_527#
+ FILLER_10_2082/li_0_n17# FILLER_24_1656/li_63_527# _546_/li_247_527# _390_/li_155_527#
+ powergood_check/FILLER_2_171/li_449_n17# user_to_mprj_in_gates\[69\]/li_707_367#
+ la_buf\[3\]/li_1535_n17# user_to_mprj_oen_buffers\[29\]/li_207_51# _611_/li_0_n17#
+ FILLER_19_1631/li_0_n17# powergood_check/FILLER_0_80/li_65_797# la_buf\[118\]/li_431_527#
+ la_buf\[63\]/li_1351_527# mprj_dat_buf\[27\]/li_1259_n17# _652_/li_247_n17# FILLER_5_763/li_0_527#
+ user_to_mprj_oen_buffers\[88\]/li_431_n17# la_buf\[43\]/li_431_n17# _567_/li_155_527#
+ mprj_stb_buf/li_611_17# mprj_cyc_buf/li_795_379# PHY_342/li_0_527# user_to_mprj_oen_buffers\[31\]/li_207_51#
+ user_to_mprj_in_gates\[116\]/li_615_527# user_to_mprj_in_gates\[83\]/li_339_n17#
+ user_to_mprj_in_gates\[124\]/li_18_51# mprj_dat_buf\[6\]/li_891_527# PHY_117/li_0_n17#
+ la_buf\[6\]/li_1167_n17# la_buf\[10\]/li_983_n17# FILLER_21_1741/li_63_n17# _358_/li_155_n17#
+ user_to_mprj_in_gates\[60\]/li_615_n17# la_buf\[115\]/li_17_51# mprj_sel_buf\[0\]/li_207_51#
+ ANTENNA__365__A/li_0_n17# powergood_check/FILLER_1_180/li_100_536# FILLER_26_1835/li_63_527#
+ la_buf\[94\]/li_1167_n17# la_buf\[126\]/li_795_379# FILLER_11_914/li_0_527# powergood_check/FILLER_2_8/li_641_n17#
+ user_to_mprj_in_buffers\[9\]/li_404_367# mprj_adr_buf\[15\]/li_1535_527# user_to_mprj_oen_buffers\[66\]/li_795_379#
+ FILLER_22_134/li_0_527# mprj_adr_buf\[26\]/li_207_51# ANTENNA__343__A/li_0_n17#
+ FILLER_10_467/li_155_n17# user_to_mprj_oen_buffers\[44\]/li_63_n17# ANTENNA_la_buf\[97\]_TE/li_63_n17#
+ powergood_check/FILLER_1_48/li_545_797# FILLER_9_386/li_155_n17# ANTENNA_la_buf\[6\]_TE/li_63_527#
+ FILLER_11_1943/li_0_527# user_to_mprj_in_gates\[118\]/li_707_367# FILLER_9_586/li_63_n17#
+ FILLER_19_1475/li_0_527# _360_/li_155_n17# _447_/li_155_527# user_to_mprj_oen_buffers\[97\]/li_207_51#
+ PHY_161/li_0_n17# powergood_check/FILLER_0_208/li_0_797# FILLER_5_1087/li_63_527#
+ FILLER_25_544/li_0_527# la_buf\[7\]/li_1443_527# FILLER_25_891/li_0_527# ANTENNA__361__A/li_63_n17#
+ powergood_check/FILLER_2_187/li_0_n17# powergood_check/FILLER_2_24/li_100_536# FILLER_22_1415/li_63_527#
+ FILLER_19_1756/li_63_n17# ANTENNA__537__A/li_63_527# la_buf\[6\]/li_431_527# FILLER_25_1261/li_155_527#
+ FILLER_25_670/li_0_n17# _351_/li_0_527# powergood_check/FILLER_2_0/li_0_n17# la_buf\[59\]/li_207_51#
+ user_to_mprj_oen_buffers\[82\]/li_707_n17# user_to_mprj_oen_buffers\[1\]/li_207_51#
+ FILLER_13_1103/li_63_n17# FILLER_19_1471/li_63_527# PHY_298/li_0_n17# la_buf\[122\]/li_207_51#
+ user_to_mprj_in_gates\[106\]/li_707_367# powergood_check/FILLER_0_256/li_65_n17#
+ powergood_check/FILLER_2_24/li_449_797# _390_/li_0_527# FILLER_11_322/li_155_n17#
+ FILLER_25_1103/li_155_n17# user_to_mprj_in_gates\[71\]/li_18_51# FILLER_26_1186/li_0_527#
+ FILLER_21_1455/li_0_n17# FILLER_18_1907/li_0_527# FILLER_26_1241/li_0_527# PHY_803/li_0_527#
+ user_to_mprj_in_gates\[31\]/li_615_527# user_to_mprj_oen_buffers\[82\]/li_1351_n17#
+ powergood_check/FILLER_1_156/li_0_n17# powergood_check/mprj2_logic_high_lv/li_1505_797#
+ user_to_mprj_oen_buffers\[61\]/li_707_527# FILLER_13_1454/li_0_n17# powergood_check/FILLER_1_172/li_257_n17#
+ la_buf\[61\]/li_207_51# FILLER_17_1428/li_155_n17# user_to_mprj_oen_buffers\[8\]/li_17_51#
+ FILLER_19_249/li_0_527# mprj_dat_buf\[4\]/li_983_527# FILLER_14_1529/li_155_527#
+ powergood_check/FILLER_0_208/li_65_797# la_buf\[109\]/li_1167_n17# FILLER_19_568/li_155_527#
+ la_buf\[11\]/li_983_n17# user_to_mprj_in_gates\[33\]/li_707_367# powergood_check/FILLER_2_259/li_100_536#
+ la_buf\[96\]/li_1535_527# user_to_mprj_in_gates\[40\]/li_615_n17# FILLER_16_1585/li_63_n17#
+ user_to_mprj_oen_buffers\[53\]/li_17_51# la_buf\[42\]/li_779_17# powergood_check/FILLER_2_8/li_161_797#
+ user_to_mprj_oen_buffers\[34\]/li_611_17# PHY_378/li_0_527# powergood_check/FILLER_0_32/li_257_797#
+ la_buf\[65\]/li_17_51# la_buf\[28\]/li_1075_n17# user_to_mprj_oen_buffers\[42\]/li_795_379#
+ FILLER_12_1117/li_0_527# mprj_dat_buf\[19\]/li_207_51# mprj_dat_buf\[26\]/li_1351_527#
+ FILLER_25_849/li_155_n17# FILLER_13_96/li_0_527# FILLER_26_1038/li_155_527# user_to_mprj_in_gates\[101\]/li_615_n17#
+ la_buf\[74\]/li_63_n17# user_to_mprj_oen_buffers\[52\]/li_431_n17# powergood_check/FILLER_2_16/li_257_n17#
+ FILLER_17_1935/li_0_527# FILLER_10_430/li_63_n17# powergood_check/FILLER_2_259/li_449_797#
+ _506_/li_155_527# user_to_mprj_in_gates\[3\]/li_339_527# user_to_mprj_in_gates\[20\]/li_18_51#
+ mprj_sel_buf\[1\]/li_17_51# powergood_check/FILLER_2_235/li_0_797# FILLER_24_1652/li_63_527#
+ user_to_mprj_oen_buffers\[20\]/li_1259_n17# powergood_check/FILLER_2_179/li_257_797#
+ mprj_adr_buf\[21\]/li_215_311# user_to_mprj_in_gates\[61\]/li_247_527# FILLER_26_939/li_155_527#
+ mprj_dat_buf\[27\]/li_611_17# FILLER_11_1717/li_155_527# user_to_mprj_in_gates\[48\]/li_63_n17#
+ mprj_dat_buf\[21\]/li_207_51# _397_/li_247_n17# user_to_mprj_in_gates\[101\]/li_63_n17#
+ user_to_mprj_in_gates\[39\]/li_18_51# _658_/li_247_n17# FILLER_22_1913/li_63_n17#
+ FILLER_11_1713/li_63_n17# powergood_check/FILLER_1_140/li_641_797# powergood_check/FILLER_2_211/li_353_797#
+ mprj_dat_buf\[16\]/li_1535_527# user_to_mprj_in_buffers\[86\]/li_339_n17# PHY_822/li_0_527#
+ ANTENNA__653__A/li_0_n17# FILLER_19_407/li_0_527# user_to_mprj_oen_buffers\[29\]/li_63_527#
+ FILLER_11_1601/li_63_n17# _564_/li_0_n17# _396_/li_0_n17# la_buf\[14\]/li_17_51#
+ FILLER_17_1883/li_63_527# user_to_mprj_in_gates\[50\]/li_63_n17# user_to_mprj_in_gates\[59\]/li_707_n17#
+ user_to_mprj_in_gates\[80\]/li_155_527# user_to_mprj_oen_buffers\[40\]/li_431_n17#
+ PHY_336/li_0_n17# la_buf\[36\]/li_63_527# _644_/li_0_527# FILLER_5_1205/li_155_527#
+ user_to_mprj_in_buffers\[72\]/li_404_17# la_buf\[9\]/li_17_51# user_to_mprj_oen_buffers\[36\]/li_207_51#
+ user_to_mprj_in_buffers\[60\]/li_0_n17# PHY_438/li_0_527# la_buf\[104\]/li_63_527#
+ FILLER_26_819/li_63_527# la_buf\[7\]/li_611_17# la_buf\[3\]/li_63_n17# _340_/li_0_n17#
+ user_to_mprj_in_gates\[39\]/li_155_527# user_to_mprj_in_gates\[87\]/li_339_n17#
+ PHY_316/li_0_527# powergood_check/FILLER_1_48/li_65_n17# la_buf\[0\]/li_891_527#
+ PHY_303/li_0_n17# PHY_50/li_0_n17# FILLER_13_756/li_0_527# powergood_check/FILLER_1_212/li_641_n17#
+ _510_/li_247_527# la_buf\[44\]/li_1535_n17# powergood_check/FILLER_0_232/li_353_797#
+ PHY_408/li_0_n17# PHY_380/li_0_n17# ANTENNA__578__A/li_63_n17# user_to_mprj_in_buffers\[76\]/li_339_n17#
+ powergood_check/FILLER_2_203/li_161_n17# la_buf\[99\]/li_0_527# la_buf\[99\]/li_1351_527#
+ user_to_mprj_in_gates\[47\]/li_707_n17# la_buf\[50\]/li_707_n17# _365_/li_155_n17#
+ powergood_check/FILLER_0_272/li_641_797# FILLER_16_1419/li_0_n17# FILLER_24_528/li_63_n17#
+ user_to_mprj_in_gates\[109\]/li_155_n17# powergood_check/mprj_logic_high_lv/li_1217_1611#
+ user_to_mprj_in_gates\[99\]/li_247_527# powergood_check/FILLER_1_62/li_161_n17#
+ user_to_mprj_in_gates\[27\]/li_155_527# user_to_mprj_in_gates\[123\]/li_18_51# user_to_mprj_oen_buffers\[59\]/li_523_n17#
+ powergood_check/FILLER_1_16/li_100_536# la_buf\[2\]/li_1075_n17# PHY_845/li_0_527#
+ la_buf\[106\]/li_983_527# user_to_mprj_oen_buffers\[51\]/li_63_n17# powergood_check/FILLER_0_0/li_0_797#
+ FILLER_9_456/li_155_n17# PHY_402/li_0_527# powergood_check/mprj2_logic_high_lv/li_65_797#
+ FILLER_22_1886/li_0_n17# ANTENNA_user_to_mprj_in_gates\[16\]_B/li_63_527# la_buf\[107\]/li_1351_527#
+ powergood_check/FILLER_2_219/li_641_797# user_to_mprj_oen_buffers\[6\]/li_207_51#
+ la_buf\[114\]/li_17_51# la_buf\[91\]/li_215_311# user_to_mprj_oen_buffers\[12\]/li_1351_527#
+ user_to_mprj_in_gates\[110\]/li_431_527# user_to_mprj_in_gates\[36\]/li_155_n17#
+ FILLER_24_215/li_63_n17# _576_/li_0_527# la_buf\[127\]/li_207_51# _367_/li_247_n17#
+ user_to_mprj_oen_buffers\[85\]/li_779_17# FILLER_20_129/li_0_n17# user_to_mprj_in_buffers\[3\]/li_51_17#
+ user_to_mprj_in_gates\[35\]/li_707_n17# FILLER_24_1425/li_0_527# la_buf\[35\]/li_891_n17#
+ powergood_check/FILLER_0_80/li_65_n17# FILLER_9_563/li_155_527# user_to_mprj_oen_buffers\[15\]/li_891_n17#
+ la_buf\[66\]/li_207_51# user_to_mprj_in_gates\[90\]/li_339_n17# la_buf\[49\]/li_0_n17#
+ FILLER_15_550/li_63_527# user_to_mprj_in_gates\[87\]/li_247_527# _656_/li_247_n17#
+ PHY_451/li_0_n17# user_to_mprj_oen_buffers\[18\]/li_63_527# ANTENNA__659__A/li_0_527#
+ powergood_check/FILLER_1_180/li_0_797# _453_/li_0_527# _334_/li_155_527# FILLER_1_892/li_155_527#
+ FILLER_20_496/li_63_n17# ANTENNA_user_to_mprj_in_gates\[119\]_B/li_63_527# FILLER_12_1687/li_0_n17#
+ powergood_check/FILLER_0_248/li_115_72# user_to_mprj_oen_buffers\[40\]/li_63_n17#
+ FILLER_13_850/li_0_527# FILLER_25_934/li_155_527# FILLER_22_515/li_155_n17# la_buf\[45\]/li_1351_n17#
+ powergood_check/FILLER_1_0/li_0_n17# user_to_mprj_in_gates\[96\]/li_247_n17# powergood_check/FILLER_2_24/li_65_797#
+ FILLER_17_1921/li_155_527# la_buf\[53\]/li_615_527# FILLER_25_1099/li_63_n17# mprj_dat_buf\[29\]/li_891_n17#
+ FILLER_25_899/li_155_n17# FILLER_18_2110/li_63_n17# user_to_mprj_oen_buffers\[12\]/li_1259_n17#
+ la_buf\[122\]/li_707_n17# _380_/li_0_527# la_buf\[95\]/li_983_n17# FILLER_12_1569/li_63_527#
+ la_buf\[38\]/li_215_311# FILLER_9_334/li_155_n17# mprj_adr_buf\[7\]/li_1535_527#
+ user_to_mprj_in_gates\[70\]/li_18_51# user_to_mprj_oen_buffers\[107\]/li_611_17#
+ FILLER_14_2009/li_63_527# mprj_adr_buf\[25\]/li_891_n17# user_to_mprj_in_gates\[75\]/li_247_527#
+ powergood_check/FILLER_1_48/li_545_n17# FILLER_15_1487/li_63_n17# FILLER_12_1378/li_63_527#
+ mprj_dat_buf\[26\]/li_207_51# PHY_780/li_0_527# FILLER_13_1021/li_0_527# user_to_mprj_oen_buffers\[7\]/li_17_51#
+ user_to_mprj_in_gates\[116\]/li_63_n17# la_buf\[60\]/li_1535_527# user_to_mprj_in_gates\[89\]/li_18_51#
+ powergood_check/FILLER_2_251/li_65_n17# powergood_check/FILLER_0_184/li_65_n17#
+ _566_/li_0_527# la_buf\[108\]/li_1259_n17# powergood_check/FILLER_0_208/li_0_n17#
+ PHY_284/li_0_n17# _513_/li_155_527# FILLER_26_895/li_0_527# user_to_mprj_oen_buffers\[52\]/li_17_51#
+ user_to_mprj_in_gates\[84\]/li_247_n17# mprj_dat_buf\[9\]/li_891_527# powergood_check/FILLER_2_300/li_0_n17#
+ la_buf\[64\]/li_17_51# la_buf\[41\]/li_615_527# user_to_mprj_in_gates\[55\]/li_63_n17#
+ FILLER_15_1666/li_155_527# mprj_dat_buf\[22\]/li_215_311# la_buf\[83\]/li_983_n17#
+ mprj_adr_buf\[2\]/li_1443_n17# la_buf\[26\]/li_215_311# _331_/li_0_527# FILLER_25_91/li_0_n17#
+ PHY_393/li_0_527# FILLER_25_730/li_0_n17# FILLER_21_467/li_0_n17# mprj_sel_buf\[0\]/li_17_51#
+ powergood_check/FILLER_2_187/li_100_536# user_to_mprj_in_gates\[65\]/li_523_n17#
+ user_to_mprj_oen_buffers\[93\]/li_1351_527# user_to_mprj_oen_buffers\[127\]/li_215_311#
+ powergood_check/FILLER_0_32/li_115_72# user_to_mprj_oen_buffers\[68\]/li_1351_n17#
+ mprj_sel_buf\[1\]/li_1259_n17# powergood_check/FILLER_2_24/li_449_n17# FILLER_17_1424/li_0_527#
+ FILLER_21_1989/li_155_527# la_buf\[94\]/li_795_379# PHY_165/li_0_527# mprj_stb_buf/li_615_527#
+ FILLER_12_839/li_63_527# user_to_mprj_oen_buffers\[104\]/li_1351_527# user_to_mprj_in_gates\[62\]/li_247_527#
+ _579_/li_155_527# la_buf\[48\]/li_63_527# powergood_check/FILLER_0_88/li_0_797#
+ user_to_mprj_in_gates\[38\]/li_18_51# user_to_mprj_in_buffers\[6\]/li_339_n17# la_buf\[51\]/li_1167_n17#
+ user_to_mprj_oen_buffers\[43\]/li_207_51# user_to_mprj_in_gates\[124\]/li_247_527#
+ FILLER_13_669/li_0_527# la_buf\[111\]/li_63_527# powergood_check/FILLER_2_187/li_449_797#
+ user_to_mprj_in_gates\[42\]/li_0_527# la_buf\[69\]/li_611_17# ANTENNA_user_to_mprj_oen_buffers\[33\]_A/li_63_n17#
+ powergood_check/FILLER_1_172/li_115_72# FILLER_25_324/li_0_n17# user_to_mprj_in_gates\[125\]/li_431_n17#
+ FILLER_15_1441/li_0_527# _554_/li_0_n17# la_buf\[13\]/li_17_51# FILLER_12_697/li_0_527#
+ mprj_dat_buf\[10\]/li_215_311# FILLER_11_1742/li_63_n17# FILLER_17_1580/li_63_527#
+ user_to_mprj_oen_buffers\[59\]/li_215_311# FILLER_7_984/li_0_527# _581_/li_155_527#
+ FILLER_25_681/li_0_n17# la_buf\[14\]/li_215_311# powergood_check/FILLER_2_8/li_161_n17#
+ FILLER_24_520/li_63_527# la_buf\[8\]/li_17_51# la_buf\[53\]/li_1351_527# user_to_mprj_oen_buffers\[115\]/li_215_311#
+ user_to_mprj_in_gates\[51\]/li_247_527# mprj_adr_buf\[0\]/li_207_51# _330_/li_0_n17#
+ powergood_check/mprj_logic_high_lv/li_257_1611# _365_/li_0_n17# powergood_check/FILLER_0_200/li_257_797#
+ _372_/li_155_n17# powergood_check/FILLER_2_259/li_449_n17# la_buf\[50\]/li_983_527#
+ user_to_mprj_in_buffers\[90\]/li_404_367# FILLER_25_1071/li_0_n17# ANTENNA__653__A/li_63_n17#
+ ANTENNA_la_buf\[51\]_A/li_63_n17# powergood_check/FILLER_2_235/li_0_n17# user_to_mprj_in_gates\[112\]/li_247_527#
+ mprj_adr_buf\[27\]/li_247_527# FILLER_11_733/li_155_n17# la_buf\[69\]/li_707_n17#
+ FILLER_11_507/li_0_n17# powergood_check/FILLER_2_203/li_115_72# user_to_mprj_in_gates\[32\]/li_523_527#
+ powergood_check/FILLER_2_179/li_257_n17# user_to_mprj_in_gates\[60\]/li_247_n17#
+ _589_/li_0_527# user_to_mprj_in_buffers\[49\]/li_404_367# FILLER_28_55/li_0_n17#
+ user_to_mprj_oen_buffers\[127\]/li_17_51# powergood_check/FILLER_0_240/li_545_797#
+ FILLER_9_526/li_155_n17# FILLER_18_2110/li_0_n17# user_to_mprj_oen_buffers\[47\]/li_215_311#
+ _549_/li_155_n17# la_buf\[101\]/li_615_527# ANTENNA__382__A/li_63_n17# powergood_check/FILLER_1_140/li_641_n17#
+ powergood_check/FILLER_2_211/li_353_n17# user_to_mprj_oen_buffers\[74\]/li_1167_n17#
+ user_to_mprj_in_gates\[27\]/li_615_n17# FILLER_16_2069/li_63_527# FILLER_14_1872/li_63_527#
+ PHY_262/li_0_527# FILLER_14_1396/li_63_n17# powergood_check/FILLER_0_160/li_353_797#
+ FILLER_16_1589/li_155_n17# FILLER_21_1937/li_0_527# PHY_314/li_0_527# user_to_mprj_oen_buffers\[103\]/li_215_311#
+ FILLER_20_56/li_0_n17# user_to_mprj_in_gates\[122\]/li_18_51# mprj_rstn_buf/li_0_527#
+ _339_/li_155_527# powergood_check/FILLER_2_251/li_641_n17# _551_/li_155_n17# la_buf\[0\]/li_611_17#
+ FILLER_25_1269/li_0_n17# la_buf\[80\]/li_431_n17# mprj_dat_buf\[16\]/li_795_379#
+ powergood_check/FILLER_1_268/li_100_536# user_to_mprj_in_gates\[100\]/li_247_527#
+ mprj_adr_buf\[29\]/li_891_527# mprj_dat_buf\[21\]/li_0_527# user_to_mprj_in_gates\[20\]/li_523_527#
+ la_buf\[73\]/li_207_51# la_buf\[29\]/li_795_379# user_to_mprj_in_gates\[51\]/li_0_n17#
+ la_buf\[113\]/li_17_51# powergood_check/FILLER_2_107/li_353_797# mprj_adr_buf\[11\]/li_891_n17#
+ la_buf\[7\]/li_983_527# mprj_dat_buf\[18\]/li_1167_527# user_to_mprj_oen_buffers\[50\]/li_615_527#
+ FILLER_23_1915/li_0_n17# powergood_check/FILLER_1_244/li_65_n17# user_to_mprj_oen_buffers\[25\]/li_63_527#
+ user_to_mprj_in_buffers\[2\]/li_51_17# user_to_mprj_oen_buffers\[35\]/li_215_311#
+ PHY_748/li_0_n17# _341_/li_155_527# user_to_mprj_in_gates\[79\]/li_339_n17# _640_/li_155_527#
+ user_to_mprj_in_gates\[94\]/li_707_367# FILLER_9_303/li_63_n17# user_to_mprj_oen_buffers\[46\]/li_611_17#
+ powergood_check/mprj_logic_high_hvl/li_257_797# la_buf\[33\]/li_0_527# _404_/li_0_527#
+ powergood_check/FILLER_0_208/li_545_797# _555_/li_0_527# powergood_check/FILLER_0_272/li_641_n17#
+ la_buf\[86\]/li_63_n17# FILLER_14_1808/li_63_527# user_to_mprj_oen_buffers\[110\]/li_707_n17#
+ _463_/li_155_n17# _518_/li_247_527# _443_/li_0_527# ANTENNA__595__A/li_63_n17# FILLER_22_1444/li_155_527#
+ user_to_mprj_oen_buffers\[54\]/li_983_527# la_buf\[17\]/li_795_379# _330_/li_0_527#
+ user_to_mprj_in_buffers\[25\]/li_404_367# FILLER_14_1500/li_0_n17# user_to_mprj_in_buffers\[6\]/li_51_367#
+ la_buf\[27\]/li_431_n17# FILLER_12_581/li_155_527# user_to_mprj_in_gates\[119\]/li_339_527#
+ powergood_check/mprj_logic_high_lv/li_641_1611# la_buf\[9\]/li_707_n17# FILLER_22_1771/li_155_n17#
+ la_buf\[2\]/li_207_51# powergood_check/FILLER_1_140/li_161_797# user_to_mprj_oen_buffers\[23\]/li_215_311#
+ FILLER_25_949/li_63_n17# powergood_check/FILLER_2_219/li_641_n17# user_to_mprj_in_gates\[39\]/li_615_527#
+ user_to_mprj_oen_buffers\[92\]/li_431_527# _608_/li_155_n17# ANTENNA__595__A/li_63_527#
+ FILLER_9_1082/li_63_527# powergood_check/FILLER_0_168/li_641_797# FILLER_13_855/li_63_n17#
+ user_to_mprj_in_gates\[82\]/li_707_367# powergood_check/FILLER_1_16/li_449_n17#
+ mprj_adr_buf\[26\]/li_891_n17# PHY_290/li_0_527# la_buf\[73\]/li_1351_n17# user_to_mprj_in_gates\[19\]/li_0_n17#
+ FILLER_9_1778/li_0_527# FILLER_7_1214/li_63_527# la_buf\[10\]/li_611_17# FILLER_16_1581/li_63_527#
+ FILLER_25_823/li_0_n17# _649_/li_247_n17# user_to_mprj_oen_buffers\[6\]/li_17_51#
+ user_to_mprj_in_gates\[88\]/li_18_51# mprj_adr_buf\[27\]/li_1075_527# user_to_mprj_oen_buffers\[48\]/li_207_51#
+ la_buf\[15\]/li_1443_n17# user_to_mprj_in_gates\[46\]/li_339_527# FILLER_17_156/li_63_527#
+ FILLER_26_859/li_0_527# user_to_mprj_oen_buffers\[51\]/li_17_51# la_buf\[56\]/li_1351_527#
+ powergood_check/FILLER_1_212/li_161_n17# user_to_mprj_in_gates\[109\]/li_615_n17#
+ la_buf\[63\]/li_17_51# mprj_adr_buf\[2\]/li_611_17# powergood_check/FILLER_2_179/li_65_n17#
+ user_to_mprj_in_gates\[107\]/li_339_527# _609_/li_247_n17# PHY_301/li_0_527# _586_/li_155_527#
+ _520_/li_0_527# user_to_mprj_in_gates\[27\]/li_615_527# user_to_mprj_oen_buffers\[11\]/li_215_311#
+ user_to_mprj_oen_buffers\[84\]/li_983_527# PHY_85/li_0_527# user_to_mprj_in_gates\[55\]/li_339_n17#
+ user_to_mprj_oen_buffers\[92\]/li_1167_527# user_to_mprj_oen_buffers\[50\]/li_207_51#
+ user_to_mprj_in_gates\[70\]/li_707_367# powergood_check/FILLER_2_24/li_65_n17# mprj_adr_buf\[5\]/li_207_51#
+ user_to_mprj_in_buffers\[35\]/li_523_527# mprj_adr_buf\[29\]/li_215_311# powergood_check/FILLER_0_272/li_161_797#
+ FILLER_25_1337/li_63_527# FILLER_24_2037/li_63_527# _571_/li_247_527# FILLER_16_88/li_155_n17#
+ _380_/li_155_n17# user_to_mprj_in_gates\[29\]/li_707_367# user_to_mprj_in_gates\[116\]/li_339_n17#
+ la_buf\[70\]/li_707_n17# user_to_mprj_in_gates\[36\]/li_615_n17# FILLER_17_249/li_63_527#
+ FILLER_23_2106/li_63_527# ANTENNA__571__A/li_63_n17# mprj_dat_buf\[22\]/li_523_n17#
+ user_to_mprj_in_gates\[37\]/li_18_51# FILLER_12_1357/li_0_527# _656_/li_0_n17# la_buf\[12\]/li_207_51#
+ _464_/li_155_527# user_to_mprj_oen_buffers\[63\]/li_63_n17# user_to_mprj_oen_buffers\[22\]/li_1535_n17#
+ FILLER_21_1444/li_155_n17# _396_/li_0_527# powergood_check/FILLER_1_220/li_65_797#
+ mprj_sel_buf\[1\]/li_63_n17# la_buf\[12\]/li_17_51# user_to_mprj_oen_buffers\[38\]/li_1443_n17#
+ user_to_mprj_oen_buffers\[45\]/li_707_527# FILLER_21_1985/li_0_527# mprj_adr_buf\[26\]/li_779_17#
+ la_buf\[7\]/li_17_51# user_to_mprj_oen_buffers\[19\]/li_17_51# mprj_adr_buf\[17\]/li_215_311#
+ _583_/li_0_n17# user_to_mprj_oen_buffers\[104\]/li_207_51# user_to_mprj_in_gates\[97\]/li_155_n17#
+ FILLER_9_1795/li_0_n17# la_buf\[70\]/li_0_527# _351_/li_247_n17# _556_/li_155_n17#
+ user_to_mprj_in_gates\[96\]/li_707_n17# user_to_mprj_in_buffers\[69\]/li_51_17#
+ FILLER_20_1778/li_0_527# FILLER_19_530/li_0_527# la_buf\[78\]/li_207_51# mprj_adr_buf\[11\]/li_1351_527#
+ user_to_mprj_in_gates\[78\]/li_431_n17# PHY_180/li_0_n17# FILLER_16_1581/li_0_n17#
+ user_to_mprj_in_gates\[76\]/li_155_527# FILLER_11_1597/li_63_n17# PHY_9/li_0_527#
+ _468_/li_247_527# user_to_mprj_oen_buffers\[126\]/li_17_51# FILLER_22_234/li_0_527#
+ powergood_check/FILLER_0_0/li_100_536# la_buf\[63\]/li_523_n17# mprj_sel_buf\[1\]/li_247_527#
+ _588_/li_0_527# la_buf\[72\]/li_0_527# la_buf\[59\]/li_779_17# FILLER_15_2039/li_63_527#
+ _645_/li_247_527# FILLER_13_1203/li_0_n17# powergood_check/FILLER_2_187/li_449_n17#
+ PHY_456/li_0_527# user_to_mprj_in_gates\[48\]/li_339_n17# PHY_47/li_0_n17# la_buf\[80\]/li_207_51#
+ FILLER_15_1928/li_155_527# mprj_sel_buf\[2\]/li_0_527# la_buf\[45\]/li_1259_527#
+ ANTENNA_user_to_mprj_in_buffers\[5\]_A/li_63_n17# powergood_check/FILLER_0_0/li_449_797#
+ user_to_mprj_in_gates\[85\]/li_155_n17# user_to_mprj_in_gates\[121\]/li_18_51# FILLER_12_1357/li_155_527#
+ PHY_855/li_0_527# FILLER_17_56/li_0_527# FILLER_5_954/li_0_527# la_buf\[70\]/li_247_n17#
+ la_buf\[90\]/li_983_n17# user_to_mprj_in_gates\[84\]/li_707_n17# user_to_mprj_oen_buffers\[120\]/li_1075_527#
+ PHY_442/li_0_n17# la_buf\[99\]/li_215_311# la_buf\[58\]/li_615_527# user_to_mprj_in_buffers\[56\]/li_155_527#
+ user_to_mprj_oen_buffers\[53\]/li_611_17# mprj_adr_buf\[8\]/li_611_17# user_to_mprj_in_gates\[66\]/li_431_n17#
+ la_buf\[112\]/li_17_51# la_buf\[29\]/li_247_n17# user_to_mprj_in_gates\[64\]/li_155_527#
+ mprj_sel_buf\[1\]/li_63_527# FILLER_19_1446/li_0_n17# PHY_234/li_0_n17# FILLER_13_1177/li_63_n17#
+ la_buf\[7\]/li_207_51# la_buf\[51\]/li_523_n17# mprj_sel_buf\[3\]/li_891_527# user_to_mprj_in_buffers\[119\]/li_404_367#
+ FILLER_11_1210/li_0_527# mprj_adr_buf\[27\]/li_63_527# powergood_check/FILLER_2_115/li_545_797#
+ user_to_mprj_in_buffers\[46\]/li_236_367# _539_/li_247_527# FILLER_26_1670/li_0_527#
+ mprj_dat_buf\[19\]/li_779_17# user_to_mprj_in_gates\[125\]/li_155_527# powergood_check/FILLER_1_196/li_100_536#
+ la_buf\[121\]/li_0_527# mprj_dat_buf\[18\]/li_891_527# FILLER_16_1421/li_155_527#
+ la_buf\[15\]/li_611_17# PHY_230/li_0_527# user_to_mprj_in_gates\[67\]/li_63_n17#
+ FILLER_13_202/li_0_n17# PHY_857/li_0_n17# user_to_mprj_in_gates\[73\]/li_155_n17#
+ mprj_dat_buf\[9\]/li_1443_527# FILLER_19_1756/li_155_527# la_buf\[6\]/li_0_527#
+ _506_/li_0_n17# FILLER_25_1103/li_0_n17# user_to_mprj_oen_buffers\[109\]/li_247_527#
+ la_buf\[92\]/li_1535_527# FILLER_27_873/li_155_n17# la_buf\[87\]/li_215_311# powergood_check/mprj2_logic_high_lv/li_826_79#
+ powergood_check/FILLER_1_107/li_641_n17# FILLER_15_1437/li_0_n17# user_to_mprj_in_gates\[106\]/li_431_527#
+ FILLER_13_1013/li_63_527# powergood_check/FILLER_0_224/li_0_797# FILLER_25_1180/li_0_n17#
+ FILLER_23_1382/li_0_n17# mprj_dat_buf\[27\]/li_891_n17# powergood_check/FILLER_0_80/li_257_797#
+ user_to_mprj_in_gates\[52\]/li_155_527# FILLER_25_1180/li_63_n17# FILLER_26_640/li_0_527#
+ PHY_233/li_0_527# FILLER_16_93/li_63_n17# FILLER_7_1148/li_0_527# FILLER_10_2105/li_63_n17#
+ _442_/li_0_527# FILLER_10_1264/li_63_527# user_to_mprj_oen_buffers\[55\]/li_207_51#
+ FILLER_12_1701/li_0_n17# la_buf\[123\]/li_523_n17# powergood_check/FILLER_2_107/li_353_n17#
+ FILLER_25_827/li_63_n17# user_to_mprj_in_gates\[33\]/li_431_527# FILLER_21_70/li_63_527#
+ user_to_mprj_oen_buffers\[91\]/li_247_n17# FILLER_23_56/li_155_n17# user_to_mprj_in_gates\[122\]/li_247_527#
+ PHY_443/li_0_527# ANTENNA_user_to_mprj_in_gates\[94\]_B/li_63_527# mprj_sel_buf\[1\]/li_247_n17#
+ powergood_check/FILLER_0_272/li_65_n17# user_to_mprj_oen_buffers\[5\]/li_17_51#
+ la_buf\[27\]/li_891_527# FILLER_1_929/li_155_527# user_to_mprj_in_gates\[87\]/li_18_51#
+ la_buf\[75\]/li_215_311# powergood_check/mprj_logic_high_hvl/li_257_n17# user_to_mprj_oen_buffers\[1\]/li_1443_n17#
+ FILLER_27_864/li_0_n17# la_buf\[17\]/li_207_51# powergood_check/mprj2_logic_high_lv/li_449_1611#
+ _649_/li_0_527# powergood_check/FILLER_1_188/li_257_n17# mprj_dat_buf\[30\]/li_1075_527#
+ user_to_mprj_in_gates\[42\]/li_431_n17# user_to_mprj_oen_buffers\[50\]/li_17_51#
+ ANTENNA_user_to_mprj_oen_buffers\[37\]_A/li_63_527# FILLER_26_797/li_155_527# FILLER_11_1646/li_0_n17#
+ user_to_mprj_in_gates\[31\]/li_247_n17# user_to_mprj_oen_buffers\[72\]/li_523_n17#
+ FILLER_13_925/li_155_527# la_buf\[62\]/li_17_51# FILLER_16_1415/li_155_n17# user_to_mprj_in_gates\[65\]/li_0_n17#
+ powergood_check/mprj_logic_high_lv/li_384_1039# FILLER_23_1774/li_0_527# powergood_check/FILLER_0_224/li_0_n17#
+ _482_/li_247_527# FILLER_10_625/li_155_n17# user_to_mprj_in_gates\[103\]/li_431_n17#
+ user_to_mprj_oen_buffers\[69\]/li_17_51# FILLER_13_1520/li_63_n17# powergood_check/FILLER_0_256/li_65_797#
+ user_to_mprj_oen_buffers\[109\]/li_207_51# user_to_mprj_oen_buffers\[30\]/li_983_527#
+ _371_/li_247_n17# user_to_mprj_in_gates\[93\]/li_523_527# FILLER_11_413/li_0_527#
+ FILLER_10_551/li_63_n17# user_to_mprj_oen_buffers\[115\]/li_1351_n17# FILLER_10_1109/li_63_n17#
+ user_to_mprj_oen_buffers\[85\]/li_707_527# la_buf\[3\]/li_891_527# powergood_check/FILLER_1_140/li_161_n17#
+ FILLER_17_1921/li_0_n17# FILLER_5_1151/li_0_527# FILLER_6_1037/li_0_527# powergood_check/FILLER_2_32/li_641_797#
+ powergood_check/FILLER_1_260/li_641_n17# mprj_sel_buf\[3\]/li_215_311# FILLER_11_744/li_0_527#
+ user_to_mprj_oen_buffers\[7\]/li_983_527# la_buf\[63\]/li_215_311# FILLER_14_2092/li_63_527#
+ user_to_mprj_in_buffers\[49\]/li_236_17# user_to_mprj_in_gates\[36\]/li_18_51# FILLER_15_428/li_63_527#
+ FILLER_25_827/li_0_n17# FILLER_12_748/li_155_n17# la_buf\[58\]/li_523_n17# powergood_check/FILLER_0_88/li_545_797#
+ powergood_check/FILLER_2_251/li_161_n17# user_to_mprj_oen_buffers\[111\]/li_207_51#
+ user_to_mprj_oen_buffers\[0\]/li_215_311# mprj_dat_buf\[18\]/li_215_311# FILLER_9_596/li_63_527#
+ user_to_mprj_oen_buffers\[60\]/li_523_n17# FILLER_9_575/li_155_n17# FILLER_12_1539/li_63_527#
+ _563_/li_155_n17# la_buf\[32\]/li_63_n17# _534_/li_0_n17# la_buf\[11\]/li_17_51#
+ user_to_mprj_oen_buffers\[43\]/li_1351_527# _586_/li_247_n17# user_to_mprj_in_gates\[59\]/li_247_527#
+ PHY_267/li_0_527# la_buf\[85\]/li_207_51# powergood_check/FILLER_2_227/li_353_797#
+ FILLER_11_1610/li_63_n17# PHY_235/li_0_527# la_buf\[6\]/li_17_51# user_to_mprj_in_gates\[81\]/li_523_527#
+ _573_/li_0_n17# user_to_mprj_oen_buffers\[18\]/li_17_51# user_to_mprj_in_buffers\[98\]/li_404_367#
+ FILLER_19_1425/li_0_n17# FILLER_24_1425/li_63_527# _353_/li_155_527# FILLER_11_1394/li_155_n17#
+ user_to_mprj_oen_buffers\[124\]/li_63_n17# user_to_mprj_oen_buffers\[96\]/li_215_311#
+ la_buf\[51\]/li_215_311# FILLER_11_1548/li_63_n17# FILLER_9_928/li_63_n17# powergood_check/FILLER_2_267/li_641_797#
+ mprj_dat_buf\[21\]/li_615_527# FILLER_11_716/li_0_n17# FILLER_12_685/li_155_n17#
+ FILLER_5_1173/li_63_527# powergood_check/mprj2_logic_high_lv/li_1505_1611# la_buf\[67\]/li_983_n17#
+ la_buf\[110\]/li_891_527# FILLER_13_850/li_63_527# la_buf\[70\]/li_891_n17# user_to_mprj_oen_buffers\[125\]/li_17_51#
+ powergood_check/FILLER_2_16/li_0_797# FILLER_15_361/li_0_527# ANTENNA_mprj_rstn_buf_A/li_63_n17#
+ powergood_check/FILLER_1_228/li_641_n17# FILLER_12_748/li_0_n17# FILLER_5_1775/li_0_527#
+ powergood_check/FILLER_0_248/li_353_797# user_to_mprj_in_gates\[47\]/li_247_527#
+ user_to_mprj_oen_buffers\[60\]/li_611_17# FILLER_22_532/li_0_527# _482_/li_0_527#
+ powergood_check/FILLER_2_219/li_161_n17# user_to_mprj_in_buffers\[86\]/li_404_367#
+ user_to_mprj_in_gates\[125\]/li_63_n17# powergood_check/FILLER_0_168/li_161_797#
+ powergood_check/mprj2_logic_high_lv/li_833_1611# FILLER_24_512/li_63_527# FILLER_13_883/li_0_n17#
+ user_to_mprj_in_gates\[120\]/li_18_51# user_to_mprj_in_gates\[115\]/li_247_527#
+ PHY_755/li_0_527# FILLER_12_689/li_63_527# user_to_mprj_oen_buffers\[84\]/li_215_311#
+ _412_/li_247_527# FILLER_0_232/li_155_527# user_to_mprj_in_gates\[56\]/li_247_n17#
+ FILLER_11_562/li_0_n17# la_buf\[123\]/li_215_311# user_to_mprj_in_gates\[74\]/li_63_n17#
+ la_buf\[22\]/li_611_17# FILLER_14_452/li_63_527# FILLER_15_1666/li_0_527# la_buf\[111\]/li_17_51#
+ user_to_mprj_oen_buffers\[7\]/li_63_527# user_to_mprj_oen_buffers\[114\]/li_615_527#
+ la_buf\[3\]/li_215_311# user_to_mprj_in_buffers\[96\]/li_404_17# FILLER_9_1082/li_63_n17#
+ la_buf\[77\]/li_983_527# mprj_stb_buf/li_17_51# FILLER_17_108/li_0_527# la_buf\[4\]/li_431_527#
+ FILLER_13_1714/li_0_n17# user_to_mprj_in_gates\[37\]/li_523_n17# FILLER_25_1204/li_63_n17#
+ FILLER_25_1200/li_155_527# mprj_dat_buf\[1\]/li_615_527# powergood_check/FILLER_1_212/li_0_797#
+ user_to_mprj_in_buffers\[74\]/li_404_367# FILLER_14_491/li_155_n17# FILLER_13_590/li_0_n17#
+ powergood_check/FILLER_0_104/li_100_536# _546_/li_0_527# la_buf\[67\]/li_63_527#
+ FILLER_9_803/li_0_527# FILLER_25_1261/li_0_527# FILLER_13_1115/li_63_527# user_to_mprj_oen_buffers\[72\]/li_215_311#
+ user_to_mprj_oen_buffers\[62\]/li_207_51# FILLER_22_294/li_63_527# mprj_logic_high_inst/li_1380_1071#
+ user_to_mprj_in_gates\[16\]/li_523_527# FILLER_11_846/li_63_527# la_buf\[50\]/li_1259_n17#
+ la_buf\[22\]/li_0_527# user_to_mprj_oen_buffers\[106\]/li_1351_527# _423_/li_0_527#
+ FILLER_27_802/li_155_n17# _574_/li_0_527# PHY_859/li_0_527# la_buf\[88\]/li_1351_527#
+ la_buf\[111\]/li_215_311# user_to_mprj_oen_buffers\[88\]/li_983_n17# user_to_mprj_in_gates\[106\]/li_0_527#
+ powergood_check/FILLER_0_104/li_449_797# _389_/li_155_n17# PHY_367/li_0_n17# ANTENNA__356__A/li_0_n17#
+ _462_/li_0_527# FILLER_19_1577/li_63_n17# _657_/li_247_n17# _520_/li_247_527# user_to_mprj_in_gates\[105\]/li_247_n17#
+ user_to_mprj_in_gates\[9\]/li_247_n17# user_to_mprj_in_gates\[97\]/li_615_n17# user_to_mprj_in_gates\[25\]/li_523_n17#
+ FILLER_12_1557/li_155_n17# FILLER_11_409/li_63_527# la_buf\[24\]/li_207_51# powergood_check/FILLER_1_48/li_115_72#
+ PHY_403/li_0_527# PHY_441/li_0_n17# FILLER_26_797/li_0_n17# FILLER_20_1663/li_0_n17#
+ _478_/li_247_527# _391_/li_155_n17# FILLER_13_1017/li_155_n17# powergood_check/FILLER_2_115/li_545_n17#
+ powergood_check/FILLER_0_184/li_115_72# user_to_mprj_oen_buffers\[0\]/li_1259_n17#
+ user_to_mprj_oen_buffers\[4\]/li_17_51# user_to_mprj_in_gates\[76\]/li_615_527#
+ user_to_mprj_oen_buffers\[60\]/li_215_311# FILLER_23_2061/li_63_527# user_to_mprj_in_gates\[86\]/li_18_51#
+ powergood_check/mprj_logic_high_lv/m1_0_51# user_to_mprj_in_gates\[35\]/li_615_n17#
+ mprj_dat_buf\[19\]/li_431_n17# FILLER_13_1199/li_0_n17# user_to_mprj_oen_buffers\[116\]/li_207_51#
+ FILLER_25_1107/li_0_n17# user_to_mprj_oen_buffers\[91\]/li_983_n17# FILLER_25_895/li_63_n17#
+ user_to_mprj_in_buffers\[40\]/li_155_n17# user_to_mprj_oen_buffers\[19\]/li_215_311#
+ mprj_adr_buf\[4\]/li_1535_n17# ANTENNA__346__A/li_0_n17# ANTENNA_user_to_mprj_in_gates\[51\]_A/li_63_n17#
+ FILLER_19_1707/li_0_527# _572_/li_155_n17# la_buf\[37\]/li_63_n17# _480_/li_155_527#
+ la_buf\[61\]/li_17_51# powergood_check/FILLER_0_200/li_65_n17# FILLER_25_520/li_63_n17#
+ powergood_check/mprj2_logic_high_lv/li_514_79# FILLER_25_1047/li_155_n17# FILLER_11_1011/li_0_527#
+ PHY_222/li_0_n17# user_to_mprj_oen_buffers\[68\]/li_17_51# FILLER_12_1788/li_63_527#
+ FILLER_22_1653/li_0_527# la_buf\[7\]/li_431_527# la_buf\[6\]/li_1167_527# PHY_702/li_0_527#
+ _358_/li_155_527# FILLER_11_428/li_63_n17# _657_/li_155_527# _570_/li_155_n17# user_to_mprj_in_gates\[53\]/li_0_527#
+ user_to_mprj_in_gates\[64\]/li_615_527# ANTENNA__365__A/li_0_527# la_buf\[92\]/li_207_51#
+ user_to_mprj_oen_buffers\[22\]/li_615_527# user_to_mprj_in_gates\[92\]/li_339_n17#
+ FILLER_10_1138/li_63_n17# user_to_mprj_in_gates\[35\]/li_18_51# user_to_mprj_in_buffers\[8\]/li_155_n17#
+ la_buf\[71\]/li_0_n17# user_to_mprj_oen_buffers\[76\]/li_1535_527# ANTENNA__345__A/li_63_n17#
+ _563_/li_0_n17# PHY_729/li_0_527# FILLER_13_1578/li_0_527# la_buf\[67\]/li_0_n17#
+ powergood_check/FILLER_0_80/li_115_72# la_buf\[31\]/li_431_527# _360_/li_155_527#
+ user_to_mprj_in_gates\[66\]/li_707_367# la_buf\[73\]/li_779_17# mprj_dat_buf\[21\]/li_1351_527#
+ user_to_mprj_oen_buffers\[20\]/li_523_n17# PHY_359/li_0_n17# user_to_mprj_in_gates\[73\]/li_615_n17#
+ la_buf\[10\]/li_17_51# powergood_check/FILLER_0_104/li_0_797# user_to_mprj_in_gates\[71\]/li_339_527#
+ _341_/li_0_527# ANTENNA_user_to_mprj_oen_buffers\[71\]_A/li_63_n17# la_buf\[44\]/li_63_527#
+ la_buf\[5\]/li_17_51# FILLER_14_359/li_155_527# user_to_mprj_oen_buffers\[17\]/li_17_51#
+ user_to_mprj_in_gates\[127\]/li_707_367# powergood_check/mprj_logic_high_lv/li_26_893#
+ FILLER_13_1239/li_155_527# ANTENNA__567__A/li_63_n17# user_to_mprj_oen_buffers\[85\]/li_431_n17#
+ mprj_sel_buf\[1\]/li_431_n17# ANTENNA__336__A/li_0_n17# la_buf\[29\]/li_17_51# _537_/li_155_527#
+ PHY_73/li_0_n17# powergood_check/FILLER_2_235/li_545_797# user_to_mprj_in_gates\[52\]/li_615_527#
+ FILLER_3_889/li_155_n17# _363_/li_247_527# user_to_mprj_oen_buffers\[118\]/li_707_n17#
+ user_to_mprj_in_gates\[79\]/li_63_n17# FILLER_21_493/li_63_n17# la_buf\[27\]/li_611_17#
+ PHY_357/li_0_527# user_to_mprj_in_buffers\[61\]/li_615_527# la_buf\[4\]/li_431_n17#
+ powergood_check/FILLER_2_155/li_353_797# powergood_check/FILLER_2_32/li_641_n17#
+ _389_/li_0_n17# mprj_adr_buf\[28\]/li_615_527# powergood_check/FILLER_1_107/li_161_n17#
+ user_to_mprj_oen_buffers\[91\]/li_1259_n17# user_to_mprj_in_gates\[118\]/li_615_527#
+ powergood_check/FILLER_0_216/li_257_797# user_to_mprj_oen_buffers\[124\]/li_17_51#
+ user_to_mprj_in_gates\[54\]/li_707_367# PHY_793/li_0_n17# PHY_688/li_0_527# FILLER_22_1665/li_63_n17#
+ ANTENNA__368__A/li_63_527# powergood_check/FILLER_1_131/li_65_797# PHY_265/li_0_527#
+ powergood_check/FILLER_2_195/li_641_797# user_to_mprj_in_buffers\[6\]/li_404_367#
+ mprj_adr_buf\[7\]/li_1351_n17# la_buf\[2\]/li_779_17# user_to_mprj_oen_buffers\[119\]/li_611_17#
+ user_to_mprj_in_gates\[81\]/li_63_n17# _559_/li_0_n17# mprj_adr_buf\[27\]/li_0_527#
+ user_to_mprj_in_gates\[115\]/li_707_367# user_to_mprj_oen_buffers\[124\]/li_891_n17#
+ powergood_check/FILLER_0_256/li_545_797# powergood_check/FILLER_2_251/li_115_72#
+ mprj_adr_buf\[7\]/li_215_311# la_buf\[70\]/li_431_527# user_to_mprj_in_gates\[122\]/li_615_n17#
+ la_buf\[102\]/li_795_379# _330_/li_155_n17# FILLER_9_1286/li_0_527# user_to_mprj_oen_buffers\[67\]/li_207_51#
+ powergood_check/FILLER_0_8/li_257_797# user_to_mprj_in_gates\[44\]/li_247_527# powergood_check/FILLER_1_156/li_641_n17#
+ powergood_check/FILLER_2_227/li_353_n17# mprj_dat_buf\[13\]/li_1443_n17# FILLER_11_1721/li_0_n17#
+ powergood_check/FILLER_0_176/li_353_797# user_to_mprj_oen_buffers\[90\]/li_983_n17#
+ FILLER_12_772/li_155_n17# user_to_mprj_oen_buffers\[40\]/li_983_n17# _563_/li_247_n17#
+ la_buf\[57\]/li_247_527# user_to_mprj_in_gates\[94\]/li_431_527# la_buf\[110\]/li_17_51#
+ user_to_mprj_oen_buffers\[52\]/li_431_527# ANTENNA_user_to_mprj_in_gates\[44\]_A/li_63_n17#
+ ANTENNA_user_to_mprj_in_gates\[16\]_A/li_63_527# user_to_mprj_oen_buffers\[29\]/li_707_527#
+ _507_/li_155_n17# powergood_check/FILLER_2_267/li_641_n17# FILLER_22_1440/li_63_527#
+ la_buf\[41\]/li_1351_527# mprj_clk2_buf/li_891_n17# la_buf\[29\]/li_207_51# powergood_check/FILLER_0_16/li_641_797#
+ _653_/li_247_n17# user_to_mprj_oen_buffers\[51\]/li_795_379# powergood_check/FILLER_2_16/li_0_n17#
+ _396_/li_155_n17# FILLER_13_1217/li_63_527# FILLER_23_1429/li_155_n17# user_to_mprj_in_gates\[7\]/li_707_367#
+ la_buf\[46\]/li_1259_n17# FILLER_9_575/li_63_n17# FILLER_16_508/li_155_n17# _658_/li_247_527#
+ FILLER_11_1713/li_63_527# la_buf\[52\]/li_1351_527# mprj_dat_buf\[19\]/li_1535_n17#
+ FILLER_12_697/li_63_n17# powergood_check/FILLER_0_272/li_0_797# _518_/li_0_527#
+ la_buf\[31\]/li_207_51# FILLER_9_1238/li_0_527# user_to_mprj_oen_buffers\[82\]/li_63_n17#
+ powergood_check/FILLER_1_180/li_65_n17# powergood_check/FILLER_2_32/li_161_797#
+ mprj_adr_buf\[30\]/li_215_311# powergood_check/FILLER_0_208/li_115_72# user_to_mprj_in_gates\[82\]/li_431_527#
+ la_buf\[45\]/li_247_527# FILLER_12_701/li_0_n17# PHY_336/li_0_527# _485_/li_155_527#
+ FILLER_9_416/li_0_n17# user_to_mprj_in_gates\[30\]/li_707_367# powergood_check/mprj_logic_high_lv/li_506_1123#
+ mprj_dat_buf\[14\]/li_1351_527# FILLER_25_895/li_155_n17# FILLER_17_1921/li_155_n17#
+ ANTENNA_user_to_mprj_in_gates\[119\]_A/li_63_527# FILLER_13_1084/li_0_527# FILLER_10_1815/li_0_n17#
+ la_buf\[9\]/li_247_527# FILLER_13_1788/li_155_n17# user_to_mprj_in_buffers\[95\]/li_339_n17#
+ user_to_mprj_in_gates\[69\]/li_155_n17# user_to_mprj_oen_buffers\[123\]/li_207_51#
+ la_buf\[98\]/li_615_527# FILLER_15_242/li_0_n17# la_buf\[123\]/li_1167_n17# user_to_mprj_in_gates\[91\]/li_431_n17#
+ FILLER_13_1071/li_63_527# FILLER_23_2061/li_63_n17# _575_/li_155_n17# la_buf\[44\]/li_0_n17#
+ mprj_adr_buf\[29\]/li_1167_527# FILLER_19_1451/li_63_527# powergood_check/FILLER_0_0/li_65_797#
+ FILLER_10_1264/li_155_527# la_buf\[97\]/li_207_51# FILLER_17_353/li_0_n17# user_to_mprj_oen_buffers\[3\]/li_17_51#
+ user_to_mprj_oen_buffers\[88\]/li_523_n17# user_to_mprj_in_gates\[85\]/li_18_51#
+ powergood_check/mprj2_logic_high_lv/li_34_216# powergood_check/FILLER_2_211/li_65_n17#
+ FILLER_23_1915/li_63_n17# FILLER_17_2059/li_0_n17# _487_/li_247_527# la_buf\[35\]/li_523_n17#
+ la_buf\[109\]/li_891_n17# _365_/li_155_527# powergood_check/FILLER_1_268/li_65_797#
+ FILLER_12_1069/li_63_n17# ANTENNA__510__A/li_63_527# la_buf\[60\]/li_17_51# FILLER_13_1048/li_0_527#
+ user_to_mprj_in_gates\[57\]/li_155_n17# _623_/li_247_n17# user_to_mprj_oen_buffers\[67\]/li_17_51#
+ powergood_check/FILLER_1_228/li_161_n17# user_to_mprj_oen_buffers\[51\]/li_63_527#
+ FILLER_20_1785/li_0_527# mprj_dat_buf\[5\]/li_0_527# mprj_adr_buf\[28\]/li_1443_n17#
+ la_buf\[79\]/li_17_51# mprj_clk_buf/li_431_n17# user_to_mprj_in_gates\[56\]/li_707_n17#
+ la_buf\[38\]/li_0_527# powergood_check/FILLER_1_48/li_0_797# FILLER_11_798/li_155_n17#
+ powergood_check/mprj_logic_high_lv/m1_0_689# FILLER_25_1051/li_0_n17# user_to_mprj_in_gates\[100\]/li_0_n17#
+ user_to_mprj_oen_buffers\[72\]/li_611_17# FILLER_13_1177/li_155_n17# user_to_mprj_in_gates\[52\]/li_0_527#
+ user_to_mprj_oen_buffers\[48\]/li_707_527# user_to_mprj_oen_buffers\[8\]/li_215_311#
+ la_buf\[57\]/li_0_527# FILLER_26_737/li_155_527# FILLER_18_1459/li_0_n17# powergood_check/FILLER_1_24/li_641_n17#
+ FILLER_17_1512/li_63_n17# powergood_check/FILLER_1_244/li_115_72# user_to_mprj_in_gates\[34\]/li_18_51#
+ FILLER_15_1998/li_0_n17# FILLER_13_1570/li_63_n17# la_buf\[21\]/li_247_527# powergood_check/FILLER_2_203/li_100_536#
+ mprj_pwrgood/li_339_527# user_to_mprj_in_buffers\[6\]/li_523_527# FILLER_18_1899/li_0_527#
+ FILLER_10_1167/li_63_n17# mprj_adr_buf\[22\]/li_983_n17# FILLER_22_1665/li_155_n17#
+ FILLER_23_1629/li_63_527# user_to_mprj_in_gates\[45\]/li_155_n17# PHY_444/li_0_n17#
+ user_to_mprj_in_gates\[86\]/li_63_n17# FILLER_12_982/li_155_n17# mprj_rstn_buf/li_17_51#
+ mprj_adr_buf\[8\]/li_431_n17# FILLER_10_481/li_155_n17# user_to_mprj_oen_buffers\[16\]/li_17_51#
+ la_buf\[4\]/li_17_51# user_to_mprj_in_gates\[44\]/li_707_n17# FILLER_24_1907/li_0_527#
+ user_to_mprj_oen_buffers\[89\]/li_891_n17# powergood_check/FILLER_2_203/li_449_797#
+ _335_/li_155_n17# powergood_check/FILLER_1_62/li_100_536# la_buf\[95\]/li_1351_527#
+ la_buf\[59\]/li_215_311# _634_/li_155_n17# FILLER_20_2110/li_0_527# la_buf\[28\]/li_17_51#
+ user_to_mprj_oen_buffers\[105\]/li_63_527# la_buf\[114\]/li_247_n17# user_to_mprj_in_buffers\[120\]/li_404_367#
+ _441_/li_0_n17# user_to_mprj_in_gates\[98\]/li_523_n17# mprj_dat_buf\[4\]/li_207_51#
+ user_to_mprj_in_gates\[96\]/li_247_527# user_to_mprj_in_gates\[105\]/li_707_n17#
+ FILLER_26_1099/li_63_527# user_to_mprj_oen_buffers\[54\]/li_247_527# ANTENNA_mprj_adr_buf\[29\]_A/li_63_527#
+ user_to_mprj_in_buffers\[104\]/li_339_527# FILLER_21_1436/li_63_n17# FILLER_19_1421/li_63_n17#
+ FILLER_18_2110/li_63_527# powergood_check/FILLER_0_224/li_100_536# powergood_check/FILLER_2_251/li_0_797#
+ la_buf\[79\]/li_63_527# FILLER_10_501/li_155_n17# FILLER_21_367/li_63_527# powergood_check/FILLER_1_62/li_449_797#
+ _432_/li_247_527# user_to_mprj_oen_buffers\[52\]/li_707_n17# user_to_mprj_oen_buffers\[74\]/li_207_51#
+ ANTENNA__564__A/li_155_n17# user_to_mprj_oen_buffers\[123\]/li_17_51# la_buf\[24\]/li_983_527#
+ mprj_stb_buf/li_1535_527# powergood_check/FILLER_2_163/li_545_797# user_to_mprj_in_gates\[77\]/li_523_527#
+ FILLER_23_1896/li_0_527# powergood_check/FILLER_1_115/li_353_n17# mprj_dat_buf\[6\]/li_1443_527#
+ powergood_check/FILLER_0_224/li_449_797# user_to_mprj_oen_buffers\[35\]/li_779_17#
+ FILLER_21_1878/li_63_527# la_buf\[38\]/li_707_n17# _655_/li_0_527# FILLER_17_231/li_63_527#
+ FILLER_19_568/li_63_527# la_buf\[47\]/li_215_311# powergood_check/FILLER_0_104/li_0_n17#
+ FILLER_25_1524/li_0_n17# PHY_439/li_0_527# _645_/li_0_n17# user_to_mprj_in_gates\[86\]/li_523_n17#
+ FILLER_17_543/li_63_n17# la_buf\[36\]/li_207_51# FILLER_15_554/li_155_527# la_buf\[41\]/li_0_n17#
+ FILLER_22_557/li_63_527# FILLER_10_611/li_63_n17# powergood_check/FILLER_2_179/li_115_72#
+ user_to_mprj_oen_buffers\[42\]/li_247_527# FILLER_21_1993/li_0_n17# powergood_check/FILLER_2_235/li_545_n17#
+ powergood_check/FILLER_0_184/li_545_797# mprj_adr_buf\[2\]/li_707_n17# _603_/li_155_527#
+ FILLER_26_91/li_0_527# FILLER_9_1042/li_0_527# la_buf\[91\]/li_983_n17# powergood_check/FILLER_2_24/li_115_72#
+ FILLER_28_63/li_63_n17# user_to_mprj_in_gates\[72\]/li_247_527# mprj_dat_buf\[27\]/li_1259_527#
+ powergood_check/FILLER_2_155/li_353_n17# PHY_183/li_0_n17# FILLER_9_526/li_63_n17#
+ la_buf\[50\]/li_615_527# user_to_mprj_oen_buffers\[51\]/li_247_n17# _627_/li_0_527#
+ FILLER_21_1812/li_155_527# la_buf\[49\]/li_63_n17# _492_/li_155_527# mprj_dat_buf\[31\]/li_215_311#
+ user_to_mprj_oen_buffers\[110\]/li_1075_n17# FILLER_13_1207/li_63_527# powergood_check/FILLER_1_0/li_545_n17#
+ user_to_mprj_in_buffers\[8\]/li_615_n17# la_buf\[35\]/li_215_311# user_to_mprj_in_buffers\[9\]/li_339_527#
+ powergood_check/FILLER_1_131/li_65_n17# FILLER_19_109/li_0_n17# powergood_check/FILLER_2_195/li_641_n17#
+ user_to_mprj_in_buffers\[68\]/li_236_17# user_to_mprj_in_gates\[74\]/li_523_n17#
+ user_to_mprj_oen_buffers\[11\]/li_611_17# la_buf\[119\]/li_215_311# mprj_adr_buf\[24\]/li_615_527#
+ la_buf\[95\]/li_1075_n17# FILLER_12_1357/li_0_n17# powergood_check/FILLER_1_260/li_161_n17#
+ FILLER_15_1437/li_155_527# FILLER_12_581/li_155_n17# FILLER_12_927/li_0_527# FILLER_11_1742/li_63_527#
+ FILLER_19_2000/li_63_527# FILLER_12_685/li_0_n17# _582_/li_155_n17# _394_/li_247_527#
+ la_buf\[51\]/li_63_n17# mprj_dat_buf\[7\]/li_215_311# ANTENNA__394__A/li_63_527#
+ FILLER_11_1725/li_0_n17# _660_/li_155_n17# FILLER_20_465/li_0_n17# PHY_453/li_0_527#
+ mprj_sel_buf\[1\]/li_891_n17# mprj_dat_buf\[7\]/li_611_17# user_to_mprj_in_gates\[84\]/li_0_n17#
+ FILLER_17_1570/li_63_527# user_to_mprj_oen_buffers\[56\]/li_63_527# FILLER_18_63/li_155_527#
+ user_to_mprj_in_gates\[25\]/li_63_n17# la_buf\[3\]/li_1351_527# FILLER_16_2087/li_0_n17#
+ FILLER_12_1921/li_0_527# _365_/li_0_527# powergood_check/FILLER_0_96/li_257_797#
+ la_buf\[84\]/li_891_n17# user_to_mprj_oen_buffers\[68\]/li_215_311# la_buf\[23\]/li_215_311#
+ FILLER_15_498/li_0_527# la_buf\[7\]/li_615_527# mprj2_pwrgood/li_19_289# la_buf\[107\]/li_215_311#
+ user_to_mprj_oen_buffers\[2\]/li_17_51# FILLER_25_303/li_63_n17# user_to_mprj_oen_buffers\[124\]/li_215_311#
+ la_buf\[45\]/li_707_527# PHY_280/li_0_527# FILLER_9_348/li_155_n17# user_to_mprj_in_gates\[84\]/li_18_51#
+ FILLER_12_890/li_63_527# _464_/li_247_n17# _549_/li_155_527# user_to_mprj_in_gates\[123\]/li_523_n17#
+ user_to_mprj_in_buffers\[3\]/li_339_n17# FILLER_16_1396/li_63_527# user_to_mprj_oen_buffers\[13\]/li_207_51#
+ mprj_dat_buf\[11\]/li_63_n17# FILLER_18_1439/li_63_n17# user_to_mprj_in_gates\[5\]/li_155_527#
+ PHY_445/li_0_n17# powergood_check/FILLER_2_32/li_161_n17# la_buf\[18\]/li_983_527#
+ FILLER_19_1577/li_63_527# user_to_mprj_in_buffers\[58\]/li_404_367# powergood_check/FILLER_2_8/li_100_536#
+ _645_/li_247_n17# user_to_mprj_oen_buffers\[66\]/li_17_51# FILLER_24_1482/li_155_n17#
+ powergood_check/mprj_logic_high_lv/li_1505_1611# user_to_mprj_oen_buffers\[56\]/li_215_311#
+ _639_/li_155_n17# la_buf\[78\]/li_17_51# la_buf\[59\]/li_1259_n17# la_buf\[20\]/li_63_527#
+ la_buf\[11\]/li_215_311# FILLER_25_1096/li_0_527# powergood_check/FILLER_1_196/li_65_797#
+ FILLER_25_1269/li_0_527# user_to_mprj_in_gates\[28\]/li_247_n17# powergood_check/FILLER_0_240/li_0_n17#
+ user_to_mprj_in_gates\[50\]/li_523_n17# mprj_dat_buf\[9\]/li_207_51# FILLER_26_721/li_0_527#
+ user_to_mprj_oen_buffers\[112\]/li_215_311# powergood_check/FILLER_2_8/li_449_797#
+ user_to_mprj_in_gates\[38\]/li_155_n17# la_buf\[41\]/li_611_17# FILLER_16_2069/li_155_527#
+ FILLER_10_551/li_155_n17# PHY_796/li_0_n17# user_to_mprj_oen_buffers\[7\]/li_1075_527#
+ user_to_mprj_in_gates\[33\]/li_18_51# user_to_mprj_oen_buffers\[92\]/li_983_527#
+ FILLER_21_1745/li_0_n17# FILLER_13_1989/li_0_527# powergood_check/FILLER_1_156/li_161_n17#
+ _342_/li_155_n17# user_to_mprj_oen_buffers\[79\]/li_207_51# PHY_384/li_0_527# FILLER_24_1648/li_155_527#
+ PHY_748/li_0_527# user_to_mprj_in_gates\[111\]/li_523_n17# mprj_adr_buf\[26\]/li_523_n17#
+ FILLER_15_1644/li_155_527# powergood_check/FILLER_0_192/li_65_797# la_buf\[45\]/li_63_527#
+ mprj_stb_buf/li_1167_n17# mprj_adr_buf\[10\]/li_207_51# powergood_check/FILLER_2_267/li_161_n17#
+ user_to_mprj_oen_buffers\[2\]/li_1351_527# la_buf\[84\]/li_0_527# PHY_351/li_0_527#
+ FILLER_16_186/li_63_n17# ANTENNA_user_to_mprj_in_gates\[83\]_B/li_63_527# user_to_mprj_oen_buffers\[15\]/li_17_51#
+ FILLER_25_141/li_63_n17# la_buf\[3\]/li_17_51# user_to_mprj_oen_buffers\[44\]/li_215_311#
+ powergood_check/FILLER_0_16/li_161_797# user_to_mprj_oen_buffers\[81\]/li_207_51#
+ user_to_mprj_in_gates\[88\]/li_339_n17# FILLER_4_1896/li_63_527# la_buf\[44\]/li_1167_527#
+ la_buf\[27\]/li_17_51# FILLER_13_1177/li_0_n17# PHY_716/li_0_527# mprj_dat_buf\[11\]/li_983_n17#
+ user_to_mprj_oen_buffers\[100\]/li_215_311# la_buf\[103\]/li_891_527# _582_/li_0_n17#
+ la_buf\[15\]/li_983_n17# powergood_check/FILLER_2_0/li_641_797# mprj_dat_buf\[23\]/li_431_527#
+ la_buf\[104\]/li_207_51# ANTENNA__338__A/li_63_n17# powergood_check/mprj2_logic_high_lv/li_26_452#
+ powergood_check/FILLER_1_48/li_0_n17# user_to_mprj_oen_buffers\[62\]/li_779_17#
+ user_to_mprj_oen_buffers\[80\]/li_983_527# FILLER_7_848/li_63_527# user_to_mprj_in_gates\[69\]/li_615_n17#
+ FILLER_11_1437/li_0_n17# user_to_mprj_in_gates\[76\]/li_707_n17# mprj_adr_buf\[7\]/li_983_527#
+ FILLER_22_1522/li_155_527# user_to_mprj_oen_buffers\[122\]/li_17_51# mprj_adr_buf\[30\]/li_891_n17#
+ FILLER_23_625/li_155_527# la_buf\[43\]/li_207_51# FILLER_12_1106/li_0_n17# FILLER_18_2110/li_0_527#
+ la_buf\[26\]/li_795_379# user_to_mprj_in_buffers\[34\]/li_404_367# user_to_mprj_oen_buffers\[53\]/li_0_n17#
+ powergood_check/mprj2_logic_high_lv/m1_0_689# FILLER_26_823/li_0_527# _497_/li_155_527#
+ la_buf\[89\]/li_707_527# user_to_mprj_in_gates\[41\]/li_247_527# user_to_mprj_oen_buffers\[32\]/li_215_311#
+ powergood_check/FILLER_2_179/li_0_797# _469_/li_0_527# la_buf\[117\]/li_0_n17# _610_/li_155_527#
+ la_buf\[24\]/li_779_17# user_to_mprj_oen_buffers\[16\]/li_611_17# user_to_mprj_in_buffers\[56\]/li_523_527#
+ la_buf\[86\]/li_1535_527# FILLER_21_1451/li_63_n17# user_to_mprj_in_gates\[109\]/li_615_527#
+ powergood_check/FILLER_2_203/li_449_n17# FILLER_13_703/li_155_527# user_to_mprj_in_buffers\[14\]/li_51_17#
+ _587_/li_155_n17# PHY_301/li_0_n17# user_to_mprj_in_gates\[57\]/li_615_n17# mprj_clk2_buf/li_891_527#
+ _401_/li_155_n17# user_to_mprj_oen_buffers\[60\]/li_1351_n17# user_to_mprj_oen_buffers\[95\]/li_1167_n17#
+ user_to_mprj_oen_buffers\[117\]/li_63_n17# FILLER_12_1491/li_63_527# la_buf\[14\]/li_795_379#
+ FILLER_7_1031/li_155_n17# la_buf\[1\]/li_1351_527# user_to_mprj_in_buffers\[22\]/li_404_367#
+ powergood_check/FILLER_2_251/li_0_n17# powergood_check/FILLER_1_62/li_449_n17# FILLER_9_516/li_63_n17#
+ user_to_mprj_oen_buffers\[90\]/li_1443_n17# powergood_check/FILLER_0_200/li_0_797#
+ FILLER_20_276/li_63_n17# _377_/li_155_527# la_buf\[127\]/li_17_51# la_buf\[24\]/li_431_n17#
+ la_buf\[1\]/li_779_17# mprj2_pwrgood/li_607_17# user_to_mprj_oen_buffers\[20\]/li_215_311#
+ powergood_check/FILLER_2_163/li_545_n17# FILLER_25_1126/li_0_n17# FILLER_12_890/li_63_n17#
+ FILLER_18_1782/li_155_n17# FILLER_9_555/li_63_n17# la_buf\[21\]/li_707_527# la_buf\[112\]/li_1351_527#
+ mprj_dat_buf\[31\]/li_17_51# FILLER_19_1446/li_0_527# user_to_mprj_in_gates\[32\]/li_63_n17#
+ la_buf\[98\]/li_1259_527# user_to_mprj_in_buffers\[54\]/li_404_17# PHY_241/li_0_n17#
+ powergood_check/FILLER_1_212/li_100_536# user_to_mprj_in_gates\[45\]/li_615_n17#
+ FILLER_16_1589/li_0_527# la_buf\[92\]/li_779_17# la_buf\[116\]/li_1351_n17# user_to_mprj_oen_buffers\[18\]/li_207_51#
+ FILLER_11_810/li_0_527# powergood_check/FILLER_1_24/li_161_n17# user_to_mprj_oen_buffers\[47\]/li_795_379#
+ user_to_mprj_in_buffers\[53\]/li_523_n17# FILLER_25_1291/li_63_n17# _583_/li_0_527#
+ la_buf\[7\]/li_1167_527# FILLER_22_2065/li_0_527# user_to_mprj_in_buffers\[10\]/li_404_367#
+ la_buf\[114\]/li_707_n17# FILLER_21_1380/li_63_527# _351_/li_247_527# la_buf\[99\]/li_1259_527#
+ la_buf\[82\]/li_247_527# _556_/li_155_527# ANTENNA_user_to_mprj_in_gates\[76\]_B/li_63_527#
+ FILLER_28_55/li_155_527# la_buf\[96\]/li_891_527# powergood_check/mprj_logic_high_lv/li_545_1611#
+ FILLER_9_966/li_0_527# user_to_mprj_oen_buffers\[20\]/li_207_51# FILLER_6_739/li_63_527#
+ user_to_mprj_oen_buffers\[72\]/li_1443_527# FILLER_19_1451/li_63_n17# mprj_adr_buf\[26\]/li_215_311#
+ user_to_mprj_oen_buffers\[19\]/li_1351_527# user_to_mprj_oen_buffers\[1\]/li_17_51#
+ PHY_180/li_0_527# FILLER_21_1436/li_0_527# FILLER_11_1597/li_63_527# user_to_mprj_in_gates\[83\]/li_18_51#
+ _347_/li_155_n17# powergood_check/FILLER_2_211/li_0_797# powergood_check/FILLER_1_260/li_0_797#
+ PHY_375/li_0_n17# ANTENNA_user_to_mprj_in_gates\[94\]_A/li_63_527# FILLER_26_1321/li_0_527#
+ ANTENNA_user_to_mprj_in_gates\[69\]_A/li_63_n17# powergood_check/FILLER_0_176/li_0_797#
+ user_to_mprj_in_gates\[31\]/li_339_527# user_to_mprj_oen_buffers\[82\]/li_1075_n17#
+ PHY_768/li_0_n17# powergood_check/FILLER_1_236/li_0_n17# powergood_check/FILLER_2_243/li_257_797#
+ la_buf\[66\]/li_1351_527# PHY_345/li_0_n17# mprj_adr_buf\[15\]/li_207_51# FILLER_18_1681/li_63_n17#
+ user_to_mprj_in_gates\[85\]/li_155_527# la_buf\[124\]/li_0_527# user_to_mprj_oen_buffers\[65\]/li_17_51#
+ powergood_check/FILLER_0_216/li_65_797# user_to_mprj_oen_buffers\[86\]/li_207_51#
+ powergood_check/FILLER_0_112/li_641_797# la_buf\[84\]/li_891_527# la_buf\[77\]/li_17_51#
+ la_buf\[92\]/li_983_527# FILLER_17_184/li_63_527# FILLER_1_892/li_63_527# user_to_mprj_in_gates\[40\]/li_339_n17#
+ FILLER_25_1265/li_0_n17# PHY_275/li_0_n17# mprj_dat_buf\[27\]/li_523_n17# powergood_check/FILLER_0_104/li_65_797#
+ FILLER_16_1711/li_63_n17# mprj_dat_buf\[25\]/li_247_527# PHY_699/li_0_527# mprj_adr_buf\[14\]/li_215_311#
+ FILLER_26_716/li_0_527# FILLER_11_897/li_0_n17# la_buf\[109\]/li_207_51# la_buf\[29\]/li_247_527#
+ FILLER_17_1428/li_63_527# user_to_mprj_oen_buffers\[24\]/li_431_527# user_to_mprj_in_gates\[32\]/li_18_51#
+ FILLER_11_436/li_63_527# user_to_mprj_in_gates\[101\]/li_339_n17# powergood_check/FILLER_2_16/li_545_797#
+ powergood_check/FILLER_1_244/li_545_n17# mprj_adr_buf\[28\]/li_63_n17# user_to_mprj_in_buffers\[3\]/li_236_17#
+ powergood_check/FILLER_0_264/li_257_797# user_to_mprj_oen_buffers\[56\]/li_1259_n17#
+ PHY_547/li_0_527# user_to_mprj_oen_buffers\[88\]/li_1167_n17# la_buf\[48\]/li_207_51#
+ FILLER_13_1115/li_155_527# user_to_mprj_in_buffers\[14\]/li_236_17# la_buf\[38\]/li_247_n17#
+ powergood_check/FILLER_0_168/li_0_n17# la_buf\[111\]/li_207_51# FILLER_18_1805/li_155_527#
+ FILLER_21_565/li_63_n17# FILLER_16_1415/li_63_n17# la_buf\[72\]/li_891_527# la_buf\[2\]/li_17_51#
+ mprj_adr_buf\[19\]/li_1351_527# user_to_mprj_oen_buffers\[14\]/li_17_51# _615_/li_155_527#
+ la_buf\[90\]/li_1075_n17# FILLER_11_1721/li_63_n17# FILLER_28_55/li_155_n17# la_buf\[26\]/li_17_51#
+ FILLER_8_981/li_63_527# la_buf\[50\]/li_207_51# FILLER_23_1382/li_0_527# la_buf\[17\]/li_247_527#
+ user_to_mprj_in_gates\[54\]/li_431_527# la_buf\[105\]/li_1351_527# FILLER_10_880/li_0_n17#
+ powergood_check/FILLER_0_24/li_353_797# FILLER_12_1543/li_0_n17# FILLER_9_892/li_0_527#
+ ANTENNA_user_to_mprj_in_gates\[40\]_A/li_63_n17# FILLER_15_1688/li_0_527# powergood_check/FILLER_2_195/li_161_n17#
+ user_to_mprj_in_buffers\[41\]/li_339_527# la_buf\[96\]/li_215_311# _359_/li_0_n17#
+ user_to_mprj_oen_buffers\[59\]/li_1443_n17# FILLER_3_893/li_63_n17# _601_/li_247_n17#
+ powergood_check/FILLER_2_8/li_449_n17# user_to_mprj_oen_buffers\[121\]/li_17_51#
+ la_buf\[84\]/li_1351_n17# mprj_dat_buf\[23\]/li_983_n17# la_buf\[70\]/li_63_527#
+ user_to_mprj_in_gates\[61\]/li_155_527# FILLER_11_2107/li_63_n17# user_to_mprj_oen_buffers\[7\]/li_615_527#
+ powergood_check/FILLER_1_252/li_65_797# _594_/li_155_n17# la_buf\[20\]/li_707_527#
+ user_to_mprj_oen_buffers\[91\]/li_247_527# user_to_mprj_in_buffers\[116\]/li_404_367#
+ la_buf\[60\]/li_891_527# user_to_mprj_in_buffers\[43\]/li_236_367# powergood_check/FILLER_1_140/li_65_797#
+ user_to_mprj_in_gates\[124\]/li_431_n17# user_to_mprj_in_gates\[80\]/li_523_n17#
+ ANTENNA__639__A/li_0_n17# FILLER_26_864/li_0_527# user_to_mprj_oen_buffers\[65\]/li_1351_527#
+ FILLER_15_1506/li_155_527# FILLER_17_1996/li_63_n17# _353_/li_247_527# mprj_dat_buf\[10\]/li_207_51#
+ FILLER_22_1634/li_63_527# user_to_mprj_in_buffers\[13\]/li_51_17# FILLER_11_332/li_0_n17#
+ mprj_dat_buf\[10\]/li_1351_527# ANTENNA_user_to_mprj_in_gates\[87\]_A/li_63_527#
+ la_buf\[84\]/li_215_311# FILLER_8_1221/li_63_n17# powergood_check/FILLER_2_0/li_641_n17#
+ user_to_mprj_oen_buffers\[59\]/li_247_n17# FILLER_28_43/li_63_n17# user_to_mprj_in_gates\[51\]/li_431_n17#
+ user_to_mprj_in_gates\[28\]/li_707_n17# FILLER_13_883/li_0_527# _595_/li_247_n17#
+ la_buf\[28\]/li_891_n17# user_to_mprj_oen_buffers\[81\]/li_523_n17# _441_/li_247_n17#
+ user_to_mprj_oen_buffers\[93\]/li_891_527# la_buf\[126\]/li_17_51# FILLER_25_1315/li_63_n17#
+ user_to_mprj_in_gates\[38\]/li_615_n17# user_to_mprj_in_buffers\[111\]/li_0_527#
+ user_to_mprj_oen_buffers\[25\]/li_207_51# la_buf\[75\]/li_247_527# user_to_mprj_oen_buffers\[91\]/li_611_17#
+ FILLER_20_2087/li_63_n17# user_to_mprj_in_gates\[112\]/li_431_n17# FILLER_23_2085/li_63_n17#
+ user_to_mprj_oen_buffers\[7\]/li_1535_527# user_to_mprj_in_gates\[110\]/li_155_527#
+ powergood_check/FILLER_1_8/li_353_n17# la_buf\[52\]/li_63_527# FILLER_13_1404/li_63_527#
+ la_buf\[98\]/li_1351_n17# user_to_mprj_in_gates\[30\]/li_431_527# _646_/li_0_527#
+ mprj_dat_buf\[30\]/li_17_51# la_buf\[114\]/li_611_17# powergood_check/FILLER_2_179/li_0_n17#
+ la_buf\[66\]/li_0_n17# FILLER_16_1415/li_155_527# la_buf\[32\]/li_63_527# _534_/li_0_527#
+ FILLER_12_617/li_63_527# la_buf\[72\]/li_215_311# user_to_mprj_in_gates\[104\]/li_615_n17#
+ FILLER_9_586/li_0_n17# FILLER_18_1961/li_0_527# FILLER_12_1610/li_63_527# mprj_dat_buf\[27\]/li_215_311#
+ powergood_check/FILLER_1_32/li_353_n17# _354_/li_155_n17# FILLER_15_548/li_0_n17#
+ _653_/li_155_n17# FILLER_9_1082/li_0_n17# mprj_stb_buf/li_795_379# FILLER_13_850/li_0_n17#
+ FILLER_12_772/li_63_527# powergood_check/FILLER_0_256/li_115_72# FILLER_21_1989/li_155_n17#
+ powergood_check/FILLER_1_140/li_100_536# user_to_mprj_in_gates\[100\]/li_431_n17#
+ la_buf\[70\]/li_1075_527# FILLER_20_1421/li_63_527# powergood_check/FILLER_2_32/li_65_797#
+ user_to_mprj_in_gates\[90\]/li_523_527# mprj_adr_buf\[22\]/li_207_51# _399_/li_0_527#
+ la_buf\[126\]/li_1351_n17# powergood_check/FILLER_1_131/li_257_797# user_to_mprj_oen_buffers\[0\]/li_17_51#
+ la_buf\[98\]/li_63_527# user_to_mprj_in_gates\[82\]/li_18_51# user_to_mprj_in_buffers\[8\]/li_236_17#
+ _443_/li_155_527# user_to_mprj_oen_buffers\[93\]/li_207_51# mprj_sel_buf\[0\]/li_215_311#
+ powergood_check/FILLER_2_251/li_100_536# FILLER_14_1399/li_0_n17# user_to_mprj_in_gates\[49\]/li_523_527#
+ powergood_check/FILLER_2_0/li_161_797# powergood_check/FILLER_1_140/li_449_797#
+ PHY_470/li_0_527# la_buf\[60\]/li_215_311# mprj_dat_buf\[30\]/li_615_527# user_to_mprj_oen_buffers\[79\]/li_615_527#
+ la_buf\[121\]/li_1535_527# la_buf\[116\]/li_207_51# mprj_dat_buf\[15\]/li_215_311#
+ user_to_mprj_oen_buffers\[74\]/li_779_17# la_buf\[118\]/li_615_527# la_buf\[63\]/li_1535_527#
+ la_buf\[19\]/li_215_311# mprj_dat_buf\[13\]/li_611_17# user_to_mprj_in_buffers\[115\]/li_404_17#
+ user_to_mprj_oen_buffers\[64\]/li_17_51# powergood_check/FILLER_1_188/li_0_797#
+ FILLER_10_1284/li_0_527# FILLER_10_501/li_63_n17# la_buf\[76\]/li_17_51# _338_/li_0_527#
+ la_buf\[55\]/li_207_51# user_to_mprj_oen_buffers\[16\]/li_523_n17# user_to_mprj_oen_buffers\[58\]/li_1351_527#
+ powergood_check/FILLER_2_171/li_257_797# user_to_mprj_in_gates\[61\]/li_431_527#
+ user_to_mprj_in_buffers\[95\]/li_404_367# ANTENNA__361__A/li_0_n17# powergood_check/FILLER_0_216/li_65_n17#
+ FILLER_25_1176/li_0_n17# FILLER_15_230/li_0_527# powergood_check/FILLER_0_272/li_100_536#
+ mprj_adr_buf\[2\]/li_1167_n17# user_to_mprj_in_gates\[31\]/li_18_51# FILLER_13_1714/li_0_527#
+ user_to_mprj_oen_buffers\[93\]/li_215_311# user_to_mprj_in_gates\[37\]/li_523_527#
+ FILLER_22_1400/li_155_n17# user_to_mprj_oen_buffers\[89\]/li_0_n17# FILLER_25_1204/li_63_527#
+ user_to_mprj_in_gates\[65\]/li_247_n17# FILLER_25_226/li_0_527# user_to_mprj_oen_buffers\[93\]/li_1075_527#
+ PHY_817/li_0_527# user_to_mprj_in_gates\[68\]/li_0_527# mprj_dat_buf\[1\]/li_1351_527#
+ la_buf\[22\]/li_615_527# ANTENNA_user_to_mprj_oen_buffers\[75\]_TE/li_63_n17# FILLER_19_1577/li_155_527#
+ powergood_check/FILLER_1_260/li_0_n17# powergood_check/FILLER_2_211/li_0_n17# PHY_19/li_0_n17#
+ user_to_mprj_oen_buffers\[123\]/li_615_527# la_buf\[126\]/li_891_527# powergood_check/FILLER_0_272/li_449_797#
+ _635_/li_0_n17# user_to_mprj_in_buffers\[117\]/li_0_n17# powergood_check/FILLER_2_219/li_100_536#
+ FILLER_13_1203/li_155_n17# user_to_mprj_oen_buffers\[13\]/li_17_51# FILLER_10_625/li_0_527#
+ PHY_453/li_0_n17# la_buf\[1\]/li_17_51# powergood_check/FILLER_1_172/li_545_n17#
+ powergood_check/FILLER_2_243/li_257_n17# user_to_mprj_oen_buffers\[108\]/li_215_311#
+ user_to_mprj_in_gates\[125\]/li_707_n17# user_to_mprj_oen_buffers\[108\]/li_983_n17#
+ FILLER_10_481/li_0_n17# powergood_check/FILLER_0_192/li_257_797# _575_/li_247_n17#
+ la_buf\[25\]/li_17_51# mprj_adr_buf\[21\]/li_0_527# powergood_check/FILLER_1_180/li_115_72#
+ mprj_dat_buf\[15\]/li_207_51# user_to_mprj_in_buffers\[83\]/li_404_367# la_buf\[70\]/li_63_n17#
+ FILLER_17_1577/li_63_527# ANTENNA__366__A/li_63_527# la_buf\[116\]/li_891_n17# powergood_check/FILLER_2_219/li_449_797#
+ user_to_mprj_in_gates\[120\]/li_247_527# _507_/li_247_527# user_to_mprj_oen_buffers\[81\]/li_215_311#
+ powergood_check/FILLER_0_104/li_65_n17# _349_/li_0_n17# powergood_check/FILLER_0_32/li_545_797#
+ user_to_mprj_oen_buffers\[122\]/li_1259_n17# user_to_mprj_oen_buffers\[120\]/li_17_51#
+ la_buf\[6\]/li_615_527# user_to_mprj_oen_buffers\[51\]/li_1167_n17# FILLER_11_1572/li_0_527#
+ la_buf\[120\]/li_215_311# FILLER_27_802/li_0_n17# mprj_adr_buf\[25\]/li_611_17#
+ FILLER_9_1099/li_155_527# FILLER_15_1688/li_63_n17# ANTENNA_user_to_mprj_in_gates\[33\]_B/li_63_527#
+ powergood_check/FILLER_2_16/li_545_n17# FILLER_11_981/li_0_527# la_buf\[0\]/li_215_311#
+ ANTENNA__375__A/li_63_n17# powergood_check/mprj2_logic_high_lv/li_1409_1611# powergood_check/FILLER_2_267/li_0_797#
+ mprj_dat_buf\[27\]/li_247_n17# user_to_mprj_in_gates\[99\]/li_707_367# mprj_dat_buf\[28\]/li_63_n17#
+ user_to_mprj_in_gates\[34\]/li_523_n17# user_to_mprj_in_gates\[32\]/li_247_527#
+ powergood_check/FILLER_2_211/li_115_72# FILLER_18_1439/li_155_n17# FILLER_11_1200/li_0_527#
+ powergood_check/FILLER_2_179/li_545_797# la_buf\[63\]/li_795_379# FILLER_26_895/li_63_527#
+ FILLER_13_777/li_63_527# mprj_rstn_buf/li_431_n17# user_to_mprj_oen_buffers\[82\]/li_1535_n17#
+ powergood_check/mprj2_logic_high_lv/li_737_1611# powergood_check/FILLER_2_211/li_641_797#
+ mprj_dat_buf\[18\]/li_795_379# FILLER_18_1459/li_63_527# user_to_mprj_oen_buffers\[32\]/li_207_51#
+ mprj_adr_buf\[30\]/li_523_n17# FILLER_26_389/li_0_527# la_buf\[58\]/li_611_17# FILLER_14_1533/li_0_527#
+ powergood_check/FILLER_2_251/li_353_797# FILLER_22_2092/li_63_n17# la_buf\[70\]/li_707_527#
+ FILLER_13_1502/li_63_527# user_to_mprj_in_gates\[48\]/li_431_n17# _393_/li_247_527#
+ FILLER_17_1829/li_0_527# la_buf\[9\]/li_1167_n17# mprj_dat_buf\[3\]/li_983_527#
+ user_to_mprj_oen_buffers\[85\]/li_983_n17# PHY_297/li_0_527# _359_/li_155_n17# user_to_mprj_oen_buffers\[28\]/li_215_311#
+ FILLER_15_543/li_0_n17# _658_/li_155_n17# user_to_mprj_in_gates\[122\]/li_155_n17#
+ mprj_dat_buf\[25\]/li_707_527# _570_/li_155_527# FILLER_17_108/li_63_n17# FILLER_12_982/li_63_n17#
+ la_buf\[29\]/li_707_527# user_to_mprj_in_gates\[87\]/li_707_367# mprj_sel_buf\[1\]/li_207_51#
+ la_buf\[125\]/li_17_51# FILLER_16_2087/li_63_527# mprj_adr_buf\[11\]/li_611_17#
+ FILLER_10_459/li_63_527# mprj_adr_buf\[27\]/li_207_51# mprj_adr_buf\[18\]/li_1351_527#
+ powergood_check/FILLER_0_112/li_161_797# FILLER_22_1634/li_63_n17# powergood_check/FILLER_1_252/li_65_n17#
+ _563_/li_0_527# _361_/li_155_n17# user_to_mprj_oen_buffers\[98\]/li_207_51# powergood_check/FILLER_0_232/li_641_797#
+ ANTENNA__588__A/li_63_n17# FILLER_15_73/li_0_527# mprj_adr_buf\[24\]/li_523_n17#
+ powergood_check/FILLER_1_140/li_65_n17# FILLER_9_596/li_0_527# FILLER_21_2061/li_155_n17#
+ _639_/li_247_n17# FILLER_25_1019/li_63_n17# la_buf\[98\]/li_1351_527# FILLER_25_891/li_155_n17#
+ FILLER_13_703/li_0_527# FILLER_9_416/li_155_n17# user_to_mprj_oen_buffers\[16\]/li_215_311#
+ FILLER_20_2079/li_0_527# _538_/li_155_n17# _450_/li_155_527# la_buf\[17\]/li_707_527#
+ powergood_check/mprj_logic_high_lv/li_1505_797# FILLER_23_493/li_63_n17# user_to_mprj_oen_buffers\[2\]/li_207_51#
+ mprj_adr_buf\[10\]/li_779_17# mprj_dat_buf\[17\]/li_1167_n17# user_to_mprj_oen_buffers\[84\]/li_891_527#
+ la_buf\[123\]/li_207_51# FILLER_13_1792/li_0_n17# _363_/li_247_n17# user_to_mprj_oen_buffers\[52\]/li_983_527#
+ _490_/li_0_527# FILLER_20_453/li_0_n17# _389_/li_0_527# mprj_pwrgood/li_523_527#
+ user_to_mprj_oen_buffers\[42\]/li_1259_527# user_to_mprj_in_gates\[81\]/li_18_51#
+ ANTENNA__576__A/li_63_n17# user_to_mprj_in_gates\[39\]/li_339_527# FILLER_12_617/li_155_n17#
+ _627_/li_155_527# user_to_mprj_in_buffers\[53\]/li_404_17# la_buf\[3\]/li_795_379#
+ user_to_mprj_oen_buffers\[85\]/li_1351_n17# la_buf\[62\]/li_207_51# la_buf\[67\]/li_247_n17#
+ FILLER_16_1581/li_0_527# user_to_mprj_in_buffers\[115\]/li_236_17# FILLER_11_581/li_155_n17#
+ FILLER_0_58/li_63_527# FILLER_25_733/li_63_n17# FILLER_13_1376/li_0_527# PHY_455/li_0_n17#
+ la_buf\[118\]/li_1075_527# _330_/li_155_527# la_buf\[9\]/li_1535_n17# user_to_mprj_in_gates\[63\]/li_707_367#
+ FILLER_21_70/li_0_n17# user_to_mprj_oen_buffers\[63\]/li_17_51# FILLER_12_1610/li_0_n17#
+ la_buf\[99\]/li_1535_527# la_buf\[75\]/li_17_51# PHY_740/li_0_n17# FILLER_15_2107/li_0_527#
+ user_to_mprj_oen_buffers\[7\]/li_523_n17# _376_/li_0_n17# user_to_mprj_in_gates\[109\]/li_339_n17#
+ powergood_check/FILLER_2_187/li_65_n17# ANTENNA_user_to_mprj_in_gates\[100\]_A/li_63_n17#
+ user_to_mprj_oen_buffers\[82\]/li_431_n17# ANTENNA__564__A/li_63_n17# FILLER_13_1812/li_155_527#
+ user_to_mprj_in_gates\[27\]/li_339_527# user_to_mprj_oen_buffers\[59\]/li_707_n17#
+ powergood_check/FILLER_1_204/li_115_72# la_buf\[2\]/li_1259_n17# user_to_mprj_in_gates\[30\]/li_18_51#
+ FILLER_22_1421/li_63_n17# FILLER_12_1186/li_155_527# powergood_check/FILLER_2_32/li_65_n17#
+ la_buf\[16\]/li_1351_527# powergood_check/FILLER_1_107/li_100_536# powergood_check/FILLER_1_131/li_257_n17#
+ PHY_261/li_0_n17# FILLER_16_1839/li_0_527# mprj_dat_buf\[22\]/li_207_51# FILLER_13_699/li_63_n17#
+ user_to_mprj_oen_buffers\[61\]/li_431_527# la_buf\[14\]/li_1075_527# user_to_mprj_in_gates\[110\]/li_615_527#
+ user_to_mprj_in_gates\[49\]/li_18_51# la_buf\[74\]/li_1259_n17# FILLER_12_734/li_0_527#
+ user_to_mprj_in_gates\[36\]/li_339_n17# la_buf\[46\]/li_1259_527# powergood_check/FILLER_1_140/li_449_n17#
+ powergood_check/FILLER_2_0/li_161_n17# FILLER_22_1418/li_0_n17# mprj_adr_buf\[11\]/li_63_527#
+ user_to_mprj_in_gates\[95\]/li_339_527# user_to_mprj_oen_buffers\[12\]/li_17_51#
+ la_buf\[0\]/li_17_51# FILLER_17_1829/li_155_527# FILLER_18_1968/li_0_527# la_buf\[24\]/li_17_51#
+ FILLER_20_1907/li_0_n17# user_to_mprj_oen_buffers\[22\]/li_1259_n17# user_to_mprj_in_gates\[51\]/li_63_n17#
+ user_to_mprj_in_gates\[90\]/li_523_n17# powergood_check/FILLER_2_251/li_449_n17#
+ mprj_adr_buf\[4\]/li_215_311# powergood_check/FILLER_1_107/li_0_n17# powergood_check/FILLER_1_188/li_0_n17#
+ _552_/li_0_n17# FILLER_15_1506/li_63_527# user_to_mprj_in_gates\[15\]/li_339_527#
+ user_to_mprj_oen_buffers\[37\]/li_207_51# user_to_mprj_oen_buffers\[38\]/li_1167_n17#
+ FILLER_26_895/li_155_527# FILLER_23_426/li_0_527# FILLER_13_1177/li_155_527# _339_/li_0_n17#
+ powergood_check/FILLER_2_171/li_257_n17# powergood_check/mprj2_logic_high_lv/li_34_1244#
+ FILLER_11_1274/li_63_n17# FILLER_12_1017/li_0_527# la_buf\[70\]/li_1535_527# la_buf\[68\]/li_983_527#
+ FILLER_17_231/li_63_n17# powergood_check/mprj_logic_high_lv/li_0_797# _378_/li_0_n17#
+ FILLER_9_1809/li_63_527# user_to_mprj_in_buffers\[79\]/li_155_527# PHY_266/li_0_527#
+ _610_/li_0_n17# FILLER_16_1581/li_155_n17# la_buf\[65\]/li_611_17# user_to_mprj_in_gates\[78\]/li_155_n17#
+ powergood_check/FILLER_0_272/li_449_n17# FILLER_21_434/li_0_n17# _366_/li_155_n17#
+ user_to_mprj_oen_buffers\[20\]/li_779_17# user_to_mprj_oen_buffers\[62\]/li_1443_n17#
+ FILLER_15_550/li_155_527# powergood_check/FILLER_0_168/li_100_536# FILLER_13_655/li_63_527#
+ powergood_check/FILLER_1_260/li_100_536# user_to_mprj_in_buffers\[11\]/li_51_17#
+ user_to_mprj_in_buffers\[15\]/li_615_n17# PHY_806/li_0_527# FILLER_8_1005/li_63_527#
+ user_to_mprj_in_gates\[59\]/li_431_n17# la_buf\[122\]/li_1443_n17# user_to_mprj_oen_buffers\[52\]/li_63_n17#
+ user_to_mprj_oen_buffers\[87\]/li_247_527# powergood_check/FILLER_2_219/li_449_n17#
+ user_to_mprj_in_gates\[19\]/li_247_527# powergood_check/FILLER_0_168/li_449_797#
+ powergood_check/FILLER_1_48/li_353_797# user_to_mprj_oen_buffers\[7\]/li_207_51#
+ user_to_mprj_in_gates\[118\]/li_155_527# la_buf\[124\]/li_17_51# FILLER_26_1062/li_0_527#
+ PHY_397/li_0_n17# mprj_clk2_buf/li_215_311# user_to_mprj_in_gates\[66\]/li_155_n17#
+ FILLER_18_1459/li_0_527# _368_/li_247_n17# user_to_mprj_oen_buffers\[86\]/li_779_17#
+ powergood_check/FILLER_0_200/li_545_797# powergood_check/FILLER_2_267/li_0_n17#
+ mprj_dat_buf\[19\]/li_0_n17# la_buf\[51\]/li_247_n17# user_to_mprj_in_gates\[65\]/li_707_n17#
+ user_to_mprj_oen_buffers\[71\]/li_0_527# la_buf\[98\]/li_891_527# powergood_check/FILLER_0_0/li_115_72#
+ la_buf\[67\]/li_207_51# la_buf\[109\]/li_779_17# _514_/li_0_527# powergood_check/FILLER_2_179/li_545_n17#
+ la_buf\[62\]/li_1351_527# user_to_mprj_in_gates\[47\]/li_431_n17# la_buf\[4\]/li_1259_527#
+ ANTENNA__591__A/li_63_527# FILLER_26_784/li_155_527# mprj_dat_buf\[3\]/li_63_527#
+ FILLER_20_518/li_0_n17# la_buf\[32\]/li_523_n17# PHY_381/li_0_527# FILLER_25_1261/li_63_n17#
+ FILLER_26_1087/li_0_527# _335_/li_155_527# FILLER_22_198/li_0_527# powergood_check/FILLER_2_211/li_641_n17#
+ la_buf\[29\]/li_523_n17# la_buf\[67\]/li_1259_n17# ANTENNA_la_buf\[125\]_TE/li_63_n17#
+ _634_/li_155_527# mprj2_vdd_pwrgood/li_155_527# user_to_mprj_in_gates\[119\]/li_0_527#
+ powergood_check/FILLER_0_160/li_641_797# powergood_check/FILLER_1_228/li_100_536#
+ user_to_mprj_in_gates\[106\]/li_155_527# powergood_check/FILLER_2_24/li_257_797#
+ powergood_check/FILLER_1_252/li_257_n17# mprj_dat_buf\[0\]/li_891_527# FILLER_13_1021/li_63_527#
+ user_to_mprj_in_gates\[98\]/li_523_527# FILLER_12_986/li_0_527# user_to_mprj_in_buffers\[117\]/li_523_n17#
+ user_to_mprj_oen_buffers\[21\]/li_63_527# FILLER_15_1709/li_0_n17# _480_/li_0_527#
+ FILLER_27_794/li_155_n17# ANTENNA__463__A/li_63_n17# la_buf\[68\]/li_215_311# user_to_mprj_in_gates\[80\]/li_18_51#
+ user_to_mprj_in_buffers\[12\]/li_404_17# la_buf\[50\]/li_779_17# user_to_mprj_in_buffers\[99\]/li_236_17#
+ la_buf\[123\]/li_247_n17# FILLER_21_1331/li_155_n17# powergood_check/FILLER_2_107/li_641_797#
+ la_buf\[3\]/li_247_n17# user_to_mprj_oen_buffers\[5\]/li_215_311# user_to_mprj_in_gates\[33\]/li_155_527#
+ mprj_dat_buf\[27\]/li_207_51# FILLER_13_895/li_155_527# user_to_mprj_in_gates\[107\]/li_63_n17#
+ FILLER_17_1520/li_63_527# user_to_mprj_in_gates\[99\]/li_18_51# PHY_179/li_0_527#
+ powergood_check/FILLER_1_268/li_737_797# _514_/li_155_527# la_buf\[102\]/li_247_527#
+ _644_/li_247_n17# FILLER_0_87/li_63_527# user_to_mprj_oen_buffers\[62\]/li_17_51#
+ FILLER_13_1207/li_0_n17# FILLER_11_744/li_63_n17# FILLER_21_2075/li_0_n17# FILLER_12_1588/li_63_n17#
+ la_buf\[101\]/li_1351_527# la_buf\[74\]/li_17_51# user_to_mprj_oen_buffers\[87\]/li_63_527#
+ la_buf\[107\]/li_1167_n17# powergood_check/FILLER_2_259/li_257_797# PHY_435/li_0_n17#
+ user_to_mprj_in_gates\[42\]/li_155_n17# user_to_mprj_in_gates\[54\]/li_0_n17# FILLER_21_1993/li_0_527#
+ user_to_mprj_oen_buffers\[72\]/li_247_n17# user_to_mprj_oen_buffers\[86\]/li_891_n17#
+ FILLER_15_206/li_0_n17# la_buf\[56\]/li_215_311# FILLER_9_611/li_155_527# user_to_mprj_in_gates\[103\]/li_155_n17#
+ FILLER_25_59/li_0_n17# la_buf\[9\]/li_0_n17# la_buf\[101\]/li_0_n17# user_to_mprj_in_gates\[95\]/li_523_n17#
+ powergood_check/FILLER_0_264/li_65_797# FILLER_13_837/li_155_527# user_to_mprj_oen_buffers\[51\]/li_247_527#
+ powergood_check/FILLER_1_212/li_65_797# la_buf\[21\]/li_523_n17# FILLER_13_1071/li_63_n17#
+ FILLER_10_463/li_155_527# mprj_dat_buf\[11\]/li_1535_n17# user_to_mprj_in_gates\[48\]/li_18_51#
+ user_to_mprj_oen_buffers\[44\]/li_207_51# FILLER_5_1896/li_63_n17# FILLER_5_1209/li_63_527#
+ mprj_stb_buf/li_891_n17# powergood_check/FILLER_1_24/li_0_n17# FILLER_25_373/li_0_527#
+ FILLER_17_2047/li_0_n17# mprj_dat_buf\[27\]/li_1443_n17# user_to_mprj_oen_buffers\[11\]/li_17_51#
+ _593_/li_0_527# FILLER_12_886/li_155_n17# la_buf\[23\]/li_17_51# user_to_mprj_oen_buffers\[60\]/li_247_n17#
+ FILLER_15_324/li_63_527# user_to_mprj_oen_buffers\[74\]/li_891_n17# user_to_mprj_in_buffers\[79\]/li_51_367#
+ la_buf\[115\]/li_0_527# _582_/li_155_527# user_to_mprj_oen_buffers\[89\]/li_215_311#
+ la_buf\[44\]/li_215_311# _542_/li_0_n17# _379_/li_0_n17# mprj_adr_buf\[1\]/li_207_51#
+ FILLER_13_1013/li_63_n17# la_buf\[72\]/li_611_17# PHY_731/li_0_527# la_buf\[55\]/li_1351_527#
+ powergood_check/FILLER_0_232/li_161_797# FILLER_9_1138/li_155_527# user_to_mprj_in_gates\[81\]/li_247_527#
+ _581_/li_0_n17# FILLER_18_1700/li_155_527# la_buf\[8\]/li_215_311# mprj_clk_buf/li_207_51#
+ la_buf\[6\]/li_1351_n17# _373_/li_155_n17# FILLER_23_621/li_155_527# la_buf\[27\]/li_0_527#
+ _368_/li_0_n17# mprj2_logic_high_inst/m1_0_496# PHY_228/li_0_527# FILLER_25_1164/li_63_n17#
+ _598_/li_0_n17# user_to_mprj_oen_buffers\[92\]/li_615_527# user_to_mprj_in_gates\[90\]/li_247_n17#
+ FILLER_9_966/li_63_527# FILLER_23_1362/li_0_527# user_to_mprj_oen_buffers\[62\]/li_891_n17#
+ _462_/li_155_527# user_to_mprj_oen_buffers\[77\]/li_215_311# user_to_mprj_in_gates\[5\]/li_707_367#
+ la_buf\[32\]/li_215_311# powergood_check/FILLER_0_112/li_0_n17# FILLER_14_355/li_63_n17#
+ mprj_adr_buf\[22\]/li_779_17# FILLER_10_459/li_63_n17# user_to_mprj_in_buffers\[38\]/li_236_17#
+ PHY_445/li_0_527# la_buf\[116\]/li_215_311# FILLER_19_52/li_63_527# _385_/li_0_n17#
+ user_to_mprj_oen_buffers\[100\]/li_207_51# la_buf\[113\]/li_523_n17# user_to_mprj_oen_buffers\[93\]/li_779_17#
+ user_to_mprj_oen_buffers\[42\]/li_707_527# la_buf\[110\]/li_1443_527# FILLER_23_1693/li_0_n17#
+ FILLER_22_515/li_63_n17# _552_/li_155_n17# la_buf\[21\]/li_63_n17# FILLER_17_353/li_63_527#
+ mprj_dat_buf\[4\]/li_215_311# la_buf\[38\]/li_0_n17# FILLER_16_88/li_155_527# la_buf\[74\]/li_207_51#
+ la_buf\[116\]/li_779_17# la_buf\[123\]/li_17_51# FILLER_11_1721/li_155_n17# FILLER_11_2093/li_155_527#
+ PHY_297/li_0_n17# user_to_mprj_in_buffers\[40\]/li_236_17# ANTENNA_la_buf\[122\]_A/li_63_n17#
+ user_to_mprj_in_buffers\[6\]/li_404_17# user_to_mprj_oen_buffers\[80\]/li_615_527#
+ user_to_mprj_in_buffers\[67\]/li_404_367# FILLER_21_1570/li_63_527# FILLER_9_54/li_63_527#
+ PHY_437/li_0_527# FILLER_12_1044/li_155_n17# powergood_check/FILLER_1_300/li_0_n17#
+ la_buf\[82\]/li_891_n17# FILLER_9_394/li_155_n17# user_to_mprj_oen_buffers\[50\]/li_891_n17#
+ _342_/li_155_527# user_to_mprj_oen_buffers\[65\]/li_215_311# _641_/li_155_527# la_buf\[20\]/li_215_311#
+ FILLER_21_1455/li_155_n17# FILLER_28_91/li_63_n17# FILLER_26_1186/li_155_527# FILLER_13_1515/li_63_n17#
+ la_buf\[104\]/li_215_311# user_to_mprj_oen_buffers\[121\]/li_215_311# powergood_check/mprj2_logic_high_lv/li_0_797#
+ mprj_dat_buf\[29\]/li_523_n17# FILLER_13_1498/li_63_527# la_buf\[48\]/li_431_527#
+ mprj_sel_buf\[3\]/li_1351_527# _543_/li_0_527# powergood_check/FILLER_2_32/li_100_536#
+ la_buf\[109\]/li_1351_n17# la_buf\[72\]/li_1167_527# la_buf\[12\]/li_1351_n17# user_to_mprj_in_gates\[16\]/li_247_527#
+ la_buf\[50\]/li_983_n17# user_to_mprj_in_gates\[118\]/li_0_527# ANTENNA__368__A/li_63_n17#
+ user_to_mprj_oen_buffers\[54\]/li_1351_527# powergood_check/FILLER_0_8/li_0_797#
+ la_buf\[88\]/li_1075_527# FILLER_15_1506/li_0_527# user_to_mprj_in_gates\[1\]/li_247_527#
+ PHY_725/li_0_n17# PHY_459/li_0_n17# FILLER_12_1117/li_155_527# la_buf\[3\]/li_207_51#
+ powergood_check/FILLER_2_32/li_449_797# PHY_511/li_0_n17# _609_/li_155_n17# powergood_check/FILLER_1_48/li_353_n17#
+ powergood_check/FILLER_0_264/li_65_n17# user_to_mprj_in_buffers\[6\]/li_339_527#
+ user_to_mprj_oen_buffers\[53\]/li_215_311# FILLER_19_2059/li_0_527# user_to_mprj_in_gates\[25\]/li_247_n17#
+ _339_/li_0_527# user_to_mprj_in_gates\[3\]/li_523_527# PHY_274/li_0_n17# powergood_check/FILLER_1_156/li_100_536#
+ FILLER_5_967/li_0_527# powergood_check/FILLER_1_180/li_257_n17# powergood_check/FILLER_1_204/li_161_n17#
+ la_buf\[12\]/li_779_17# FILLER_15_59/li_63_n17# FILLER_14_452/li_155_n17# FILLER_13_855/li_155_527#
+ user_to_mprj_in_buffers\[85\]/li_404_17# FILLER_21_467/li_63_n17# user_to_mprj_in_gates\[98\]/li_18_51#
+ user_to_mprj_oen_buffers\[49\]/li_207_51# user_to_mprj_in_buffers\[107\]/li_51_367#
+ _564_/li_247_n17# user_to_mprj_in_gates\[78\]/li_615_n17# FILLER_26_528/li_0_527#
+ powergood_check/FILLER_0_192/li_115_72# user_to_mprj_in_gates\[76\]/li_339_527#
+ user_to_mprj_oen_buffers\[108\]/li_431_n17# FILLER_14_2028/li_0_527# powergood_check/FILLER_2_267/li_100_536#
+ mprj_dat_buf\[31\]/li_795_379# user_to_mprj_oen_buffers\[61\]/li_17_51# la_buf\[73\]/li_17_51#
+ user_to_mprj_in_gates\[48\]/li_523_n17# mprj_dat_buf\[1\]/li_0_527# la_buf\[119\]/li_795_379#
+ la_buf\[56\]/li_63_527# powergood_check/mprj2_logic_high_hvl/li_353_797# user_to_mprj_oen_buffers\[41\]/li_215_311#
+ FILLER_9_992/li_63_527# user_to_mprj_in_gates\[63\]/li_247_527# powergood_check/FILLER_2_24/li_257_n17#
+ powergood_check/mprj_logic_high_lv/li_1409_1611# _401_/li_155_527# user_to_mprj_oen_buffers\[51\]/li_207_51#
+ user_to_mprj_in_gates\[85\]/li_339_n17# powergood_check/FILLER_2_267/li_449_797#
+ user_to_mprj_oen_buffers\[87\]/li_707_527# la_buf\[126\]/li_0_527# powergood_check/FILLER_1_204/li_0_797#
+ mprj_adr_buf\[6\]/li_207_51# la_buf\[77\]/li_611_17# user_to_mprj_in_buffers\[65\]/li_523_527#
+ mprj_dat_buf\[7\]/li_795_379# la_buf\[9\]/li_431_n17# user_to_mprj_oen_buffers\[57\]/li_983_n17#
+ powergood_check/FILLER_0_80/li_545_797# user_to_mprj_oen_buffers\[93\]/li_0_527#
+ _378_/li_155_n17# powergood_check/FILLER_2_187/li_257_797# la_buf\[0\]/li_983_527#
+ FILLER_9_996/li_0_527# FILLER_9_667/li_63_527# user_to_mprj_in_gates\[59\]/li_707_367#
+ la_buf\[6\]/li_707_527# powergood_check/FILLER_0_232/li_65_n17# user_to_mprj_in_gates\[66\]/li_615_n17#
+ FILLER_23_1449/li_0_n17# user_to_mprj_in_gates\[47\]/li_18_51# user_to_mprj_in_gates\[64\]/li_339_527#
+ PHY_274/li_0_527# powergood_check/FILLER_2_107/li_641_n17# la_buf\[51\]/li_707_n17#
+ user_to_mprj_oen_buffers\[68\]/li_795_379# FILLER_17_462/li_0_n17# la_buf\[13\]/li_207_51#
+ la_buf\[79\]/li_0_n17# ANTENNA__660__A/li_0_n17# user_to_mprj_oen_buffers\[10\]/li_17_51#
+ user_to_mprj_in_buffers\[31\]/li_404_367# _644_/li_0_n17# FILLER_28_51/li_155_n17#
+ powergood_check/FILLER_1_268/li_737_n17# mprj_stb_buf/li_1443_527# la_buf\[22\]/li_17_51#
+ user_to_mprj_in_gates\[125\]/li_431_527# user_to_mprj_in_gates\[53\]/li_247_527#
+ FILLER_25_1008/li_155_n17# user_to_mprj_in_gates\[73\]/li_339_n17# PHY_814/li_0_n17#
+ FILLER_18_1945/li_0_527# user_to_mprj_oen_buffers\[29\]/li_17_51# powergood_check/FILLER_1_188/li_545_n17#
+ powergood_check/FILLER_2_259/li_257_n17# user_to_mprj_in_buffers\[45\]/li_0_527#
+ user_to_mprj_in_gates\[99\]/li_431_527# user_to_mprj_oen_buffers\[105\]/li_207_51#
+ FILLER_12_1701/li_63_n17# ANTENNA_user_to_mprj_oen_buffers\[4\]_TE/li_63_n17# user_to_mprj_oen_buffers\[45\]/li_63_527#
+ PHY_829/li_0_n17# user_to_mprj_in_gates\[106\]/li_615_527# la_buf\[126\]/li_1443_527#
+ FILLER_15_62/li_63_n17# _557_/li_155_n17# user_to_mprj_in_gates\[47\]/li_707_367#
+ la_buf\[6\]/li_611_17# FILLER_21_1947/li_155_527# powergood_check/FILLER_1_220/li_641_n17#
+ powergood_check/FILLER_1_16/li_65_n17# la_buf\[79\]/li_207_51# user_to_mprj_in_gates\[52\]/li_339_527#
+ powergood_check/FILLER_0_240/li_353_797# _358_/li_0_n17# mprj_adr_buf\[14\]/li_1351_527#
+ FILLER_18_1439/li_155_527# user_to_mprj_oen_buffers\[75\]/li_1351_n17# powergood_check/FILLER_2_211/li_161_n17#
+ user_to_mprj_in_gates\[108\]/li_707_367# la_buf\[123\]/li_707_n17# powergood_check/FILLER_0_160/li_161_797#
+ _397_/li_0_n17# la_buf\[21\]/li_431_n17# _355_/li_0_527# FILLER_12_693/li_155_n17#
+ _646_/li_155_527# user_to_mprj_in_gates\[33\]/li_615_527# powergood_check/FILLER_0_88/li_65_797#
+ _391_/li_247_n17# la_buf\[81\]/li_207_51# la_buf\[123\]/li_779_17# PHY_768/li_0_527#
+ _368_/li_247_527# user_to_mprj_oen_buffers\[57\]/li_1075_n17# FILLER_14_1447/li_63_527#
+ PHY_92/li_0_527# user_to_mprj_in_gates\[87\]/li_431_527# FILLER_23_1774/li_0_n17#
+ FILLER_10_1935/li_0_n17# FILLER_14_355/li_63_527# FILLER_12_1378/li_0_527# powergood_check/FILLER_1_24/li_100_536#
+ la_buf\[26\]/li_891_527# user_to_mprj_in_gates\[122\]/li_339_n17# user_to_mprj_in_gates\[35\]/li_707_367#
+ powergood_check/FILLER_2_107/li_161_797# FILLER_10_625/li_0_n17# FILLER_23_2106/li_0_527#
+ user_to_mprj_in_gates\[42\]/li_615_n17# FILLER_22_1440/li_155_527# user_to_mprj_in_buffers\[28\]/li_51_17#
+ user_to_mprj_oen_buffers\[72\]/li_707_n17# powergood_check/FILLER_2_227/li_641_797#
+ FILLER_25_1265/li_0_527# mprj_dat_buf\[13\]/li_1167_n17# la_buf\[122\]/li_17_51#
+ mprj_sel_buf\[2\]/li_63_527# user_to_mprj_in_gates\[96\]/li_431_n17# la_buf\[56\]/li_611_17#
+ user_to_mprj_in_gates\[94\]/li_155_527# PHY_268/li_0_n17# la_buf\[8\]/li_207_51#
+ user_to_mprj_in_gates\[103\]/li_615_n17# mprj_adr_buf\[28\]/li_63_527# _606_/li_0_527#
+ FILLER_17_1577/li_63_n17# powergood_check/FILLER_0_208/li_353_797# user_to_mprj_in_buffers\[9\]/li_523_527#
+ FILLER_20_1459/li_155_527# user_to_mprj_oen_buffers\[110\]/li_431_n17# mprj_adr_buf\[3\]/li_1351_527#
+ PHY_164/li_0_n17# FILLER_20_1663/li_0_527# mprj_adr_buf\[23\]/li_215_311# _345_/li_247_n17#
+ powergood_check/FILLER_1_131/li_50_537# user_to_mprj_in_gates\[22\]/li_247_527#
+ _645_/li_0_527# FILLER_14_1396/li_0_n17# FILLER_16_520/li_155_527# user_to_mprj_in_gates\[23\]/li_707_367#
+ powergood_check/FILLER_0_248/li_641_797# FILLER_25_1241/li_63_n17# FILLER_11_1027/li_63_n17#
+ user_to_mprj_oen_buffers\[60\]/li_707_n17# FILLER_19_1756/li_63_527# FILLER_5_861/li_63_527#
+ mprj_dat_buf\[22\]/li_779_17# user_to_mprj_in_gates\[84\]/li_431_n17# powergood_check/FILLER_0_216/li_115_72#
+ _572_/li_0_527# user_to_mprj_in_gates\[82\]/li_155_527# _528_/li_247_527# powergood_check/FILLER_1_16/li_257_n17#
+ FILLER_26_925/li_0_527# user_to_mprj_in_buffers\[92\]/li_404_17# user_to_mprj_oen_buffers\[56\]/li_207_51#
+ powergood_check/FILLER_0_104/li_115_72# FILLER_14_456/li_0_527# _359_/li_0_527#
+ la_buf\[12\]/li_1535_527# powergood_check/mprj_logic_high_lv/li_449_1611# _488_/li_0_527#
+ FILLER_9_1169/li_0_527# la_buf\[28\]/li_523_n17# FILLER_14_2096/li_0_527# ANTENNA__349__A/li_0_n17#
+ mprj_adr_buf\[11\]/li_215_311# FILLER_17_100/li_0_527# FILLER_13_1816/li_63_n17#
+ user_to_mprj_in_gates\[91\]/li_155_n17# FILLER_25_815/li_63_n17# user_to_mprj_oen_buffers\[110\]/li_611_17#
+ FILLER_17_1424/li_155_527# user_to_mprj_oen_buffers\[37\]/li_779_17# mprj_adr_buf\[25\]/li_1535_n17#
+ user_to_mprj_in_gates\[97\]/li_247_527# la_buf\[113\]/li_983_527# user_to_mprj_in_gates\[97\]/li_18_51#
+ user_to_mprj_in_buffers\[6\]/li_523_n17# la_buf\[51\]/li_1351_n17# powergood_check/FILLER_0_96/li_0_n17#
+ la_buf\[18\]/li_207_51# la_buf\[79\]/li_615_527# la_buf\[84\]/li_611_17# user_to_mprj_oen_buffers\[60\]/li_17_51#
+ user_to_mprj_in_gates\[72\]/li_431_n17# la_buf\[35\]/li_247_n17# FILLER_15_73/li_155_n17#
+ FILLER_11_629/li_155_527# la_buf\[72\]/li_17_51# _385_/li_155_n17# user_to_mprj_in_gates\[125\]/li_523_n17#
+ FILLER_25_1770/li_155_n17# FILLER_12_1035/li_0_n17# user_to_mprj_in_buffers\[125\]/li_404_367#
+ user_to_mprj_oen_buffers\[79\]/li_17_51# la_buf\[20\]/li_207_51# powergood_check/FILLER_2_195/li_100_536#
+ FILLER_24_1886/li_0_527# FILLER_12_1486/li_0_527# mprj_dat_buf\[7\]/li_247_n17#
+ mprj_adr_buf\[24\]/li_63_527# _528_/li_0_527# powergood_check/FILLER_0_112/li_0_797#
+ la_buf\[14\]/li_247_527# powergood_check/FILLER_2_32/li_449_n17# la_buf\[28\]/li_0_527#
+ FILLER_21_2105/li_0_n17# user_to_mprj_oen_buffers\[117\]/li_523_n17# _474_/li_155_527#
+ user_to_mprj_in_gates\[64\]/li_0_527# mprj_adr_buf\[27\]/li_431_527# la_buf\[93\]/li_215_311#
+ mprj_dat_buf\[23\]/li_63_527# user_to_mprj_in_gates\[46\]/li_18_51# FILLER_26_1195/li_63_527#
+ powergood_check/FILLER_2_195/li_449_797# la_buf\[67\]/li_615_527# la_buf\[67\]/li_1259_527#
+ user_to_mprj_oen_buffers\[112\]/li_207_51# powergood_check/FILLER_1_252/li_115_72#
+ FILLER_11_1557/li_0_n17# _564_/li_155_n17# FILLER_25_1204/li_0_527# mprj_adr_buf\[29\]/li_795_379#
+ la_buf\[21\]/li_17_51# user_to_mprj_oen_buffers\[121\]/li_779_17# powergood_check/FILLER_1_140/li_115_72#
+ la_buf\[113\]/li_0_527# FILLER_0_54/li_155_527# FILLER_13_2020/li_0_527# powergood_check/FILLER_0_160/li_65_n17#
+ la_buf\[86\]/li_207_51# user_to_mprj_oen_buffers\[74\]/li_1351_n17# user_to_mprj_in_gates\[31\]/li_0_n17#
+ user_to_mprj_in_gates\[3\]/li_247_527# FILLER_17_1402/li_63_n17# powergood_check/FILLER_0_16/li_100_536#
+ user_to_mprj_oen_buffers\[28\]/li_17_51# _555_/li_247_n17# user_to_mprj_oen_buffers\[60\]/li_983_527#
+ PHY_306/li_0_527# FILLER_21_297/li_0_527# powergood_check/mprj2_logic_high_hvl/li_353_n17#
+ la_buf\[80\]/li_0_n17# powergood_check/mprj_logic_high_lv/li_34_1244# _354_/li_155_527#
+ la_buf\[67\]/li_779_17# FILLER_18_1778/li_155_n17# FILLER_13_1676/li_63_527# powergood_check/FILLER_2_267/li_449_n17#
+ powergood_check/FILLER_1_204/li_0_n17# FILLER_13_911/li_63_527# user_to_mprj_oen_buffers\[59\]/li_611_17#
+ FILLER_15_1666/li_63_527# la_buf\[81\]/li_215_311# FILLER_26_1066/li_63_527# mprj_dat_buf\[16\]/li_983_527#
+ _348_/li_0_n17# user_to_mprj_in_gates\[98\]/li_247_n17# powergood_check/FILLER_0_16/li_449_797#
+ _574_/li_247_527# la_buf\[55\]/li_615_527# powergood_check/FILLER_2_187/li_257_n17#
+ powergood_check/mprj_logic_high_lv/li_833_1611# mprj_dat_buf\[18\]/li_1351_527#
+ FILLER_19_1425/li_0_527# la_buf\[99\]/li_63_n17# la_buf\[12\]/li_523_n17# user_to_mprj_in_gates\[25\]/li_707_n17#
+ ANTENNA_user_to_mprj_in_gates\[33\]_A/li_63_527# FILLER_10_459/li_155_527# user_to_mprj_in_gates\[55\]/li_0_n17#
+ powergood_check/FILLER_0_0/li_257_797# PHY_436/li_0_527# user_to_mprj_in_gates\[79\]/li_523_n17#
+ la_buf\[24\]/li_707_527# user_to_mprj_in_gates\[77\]/li_247_527# FILLER_19_1451/li_155_527#
+ mprj_dat_buf\[6\]/li_1167_527# FILLER_22_1400/li_63_n17# user_to_mprj_in_buffers\[90\]/li_155_527#
+ mprj_adr_buf\[15\]/li_1075_n17# FILLER_18_1744/li_63_n17# _533_/li_155_527# FILLER_5_1217/li_63_n17#
+ FILLER_14_1696/li_0_527# FILLER_15_1692/li_63_n17# user_to_mprj_in_buffers\[40\]/li_339_n17#
+ FILLER_23_1376/li_0_527# user_to_mprj_in_gates\[86\]/li_247_n17# user_to_mprj_in_gates\[5\]/li_615_n17#
+ user_to_mprj_oen_buffers\[44\]/li_247_n17# user_to_mprj_in_gates\[75\]/li_63_n17#
+ la_buf\[121\]/li_17_51# powergood_check/FILLER_2_115/li_353_797# powergood_check/FILLER_2_187/li_115_72#
+ mprj_dat_buf\[24\]/li_215_311# user_to_mprj_in_buffers\[97\]/li_404_17# FILLER_26_1176/li_0_527#
+ la_buf\[28\]/li_215_311# user_to_mprj_in_gates\[119\]/li_523_527# user_to_mprj_oen_buffers\[48\]/li_0_527#
+ _623_/li_155_n17# FILLER_16_1589/li_0_n17# FILLER_25_1481/li_63_527# user_to_mprj_in_gates\[67\]/li_523_n17#
+ powergood_check/FILLER_1_212/li_65_n17# powergood_check/FILLER_2_32/li_115_72# mprj_dat_buf\[27\]/li_983_527#
+ FILLER_12_617/li_63_n17# powergood_check/FILLER_2_155/li_641_797# user_to_mprj_oen_buffers\[23\]/li_247_527#
+ FILLER_15_1609/li_63_n17# user_to_mprj_oen_buffers\[37\]/li_891_527# la_buf\[96\]/li_795_379#
+ la_buf\[64\]/li_983_527# la_buf\[68\]/li_63_527# powergood_check/FILLER_0_216/li_545_797#
+ user_to_mprj_in_buffers\[111\]/li_523_527# FILLER_22_1415/li_0_527# _413_/li_155_527#
+ user_to_mprj_in_buffers\[8\]/li_339_n17# user_to_mprj_in_gates\[126\]/li_247_527#
+ user_to_mprj_oen_buffers\[63\]/li_207_51# PHY_454/li_0_n17# FILLER_13_752/li_0_527#
+ FILLER_25_815/li_63_527# la_buf\[89\]/li_611_17# user_to_mprj_oen_buffers\[109\]/li_1351_527#
+ user_to_mprj_in_gates\[74\]/li_247_n17# FILLER_13_1103/li_63_527# mprj_adr_buf\[19\]/li_17_51#
+ la_buf\[31\]/li_615_527# user_to_mprj_in_gates\[104\]/li_155_n17# mprj_dat_buf\[12\]/li_215_311#
+ user_to_mprj_in_gates\[80\]/li_431_n17# _562_/li_0_527# FILLER_16_1415/li_0_n17#
+ powergood_check/FILLER_2_107/li_161_n17# la_buf\[16\]/li_215_311# FILLER_17_1909/li_63_n17#
+ FILLER_21_467/li_63_527# user_to_mprj_in_gates\[107\]/li_523_527# FILLER_5_1217/li_155_n17#
+ powergood_check/FILLER_0_8/li_545_797# powergood_check/FILLER_2_227/li_641_n17#
+ user_to_mprj_oen_buffers\[83\]/li_0_n17# user_to_mprj_in_gates\[55\]/li_523_n17#
+ FILLER_16_1663/li_0_527# user_to_mprj_oen_buffers\[67\]/li_1351_n17# _349_/li_0_527#
+ powergood_check/FILLER_0_176/li_641_797# user_to_mprj_oen_buffers\[117\]/li_215_311#
+ user_to_mprj_oen_buffers\[50\]/li_983_527# la_buf\[25\]/li_207_51# mprj_sel_buf\[1\]/li_611_17#
+ powergood_check/FILLER_1_268/li_257_n17# mprj_dat_buf\[3\]/li_615_527# powergood_check/FILLER_1_24/li_449_n17#
+ FILLER_12_1044/li_63_527# la_buf\[86\]/li_983_527# FILLER_13_1680/li_0_n17# FILLER_24_2040/li_0_527#
+ la_buf\[3\]/li_1075_527# _392_/li_155_n17# user_to_mprj_in_buffers\[92\]/li_404_367#
+ FILLER_25_1096/li_63_n17# ANTENNA__655__A/li_63_n17# user_to_mprj_in_gates\[116\]/li_523_n17#
+ FILLER_11_2107/li_0_n17# user_to_mprj_in_gates\[96\]/li_18_51# user_to_mprj_oen_buffers\[90\]/li_215_311#
+ PHY_783/li_0_527# mprj_dat_buf\[22\]/li_707_n17# mprj_clk_buf/li_779_17# FILLER_13_911/li_155_n17#
+ PHY_360/li_0_527# FILLER_12_1186/li_0_527# user_to_mprj_oen_buffers\[117\]/li_207_51#
+ user_to_mprj_oen_buffers\[20\]/li_247_n17# FILLER_17_2033/li_0_n17# powergood_check/FILLER_1_220/li_161_n17#
+ la_buf\[119\]/li_1351_527# user_to_mprj_oen_buffers\[49\]/li_215_311# la_buf\[38\]/li_63_n17#
+ la_buf\[71\]/li_17_51# powergood_check/FILLER_2_259/li_65_n17# PHY_316/li_0_n17#
+ FILLER_13_1714/li_63_n17# user_to_mprj_in_gates\[123\]/li_247_n17# mprj_dat_buf\[30\]/li_63_527#
+ user_to_mprj_oen_buffers\[124\]/li_1075_n17# user_to_mprj_oen_buffers\[105\]/li_215_311#
+ user_to_mprj_oen_buffers\[78\]/li_17_51# la_buf\[72\]/li_795_379# _359_/li_155_527#
+ user_to_mprj_in_buffers\[80\]/li_404_367# _658_/li_155_527# _571_/li_155_n17# la_buf\[59\]/li_983_n17#
+ powergood_check/FILLER_0_88/li_353_797# powergood_check/mprj2_logic_high_lv/li_26_893#
+ user_to_mprj_in_gates\[6\]/li_247_527# mprj_dat_buf\[27\]/li_795_379# user_to_mprj_in_gates\[94\]/li_615_527#
+ la_buf\[93\]/li_207_51# FILLER_16_1601/li_0_n17# user_to_mprj_in_gates\[50\]/li_247_n17#
+ user_to_mprj_in_gates\[45\]/li_18_51# user_to_mprj_oen_buffers\[52\]/li_615_527#
+ user_to_mprj_in_buffers\[41\]/li_155_527# user_to_mprj_oen_buffers\[65\]/li_707_527#
+ user_to_mprj_oen_buffers\[22\]/li_891_n17# user_to_mprj_in_gates\[5\]/li_523_n17#
+ FILLER_21_1503/li_63_527# user_to_mprj_oen_buffers\[37\]/li_215_311# _392_/li_0_527#
+ powergood_check/FILLER_1_228/li_65_797# user_to_mprj_in_gates\[38\]/li_431_n17#
+ PHY_460/li_0_527# la_buf\[74\]/li_779_17# _660_/li_155_527# user_to_mprj_oen_buffers\[57\]/li_1535_527#
+ mprj_adr_buf\[31\]/li_983_n17# user_to_mprj_in_gates\[111\]/li_247_n17# user_to_mprj_in_gates\[96\]/li_707_367#
+ la_buf\[20\]/li_17_51# mprj_we_buf/li_215_311# FILLER_16_2031/li_63_n17# la_buf\[120\]/li_0_n17#
+ PHY_239/li_0_n17# user_to_mprj_oen_buffers\[27\]/li_17_51# la_buf\[60\]/li_795_379#
+ FILLER_5_1205/li_63_527# FILLER_25_891/li_155_527# FILLER_9_1127/li_0_527# FILLER_23_1778/li_63_527#
+ la_buf\[39\]/li_17_51# FILLER_17_1817/li_63_527# _597_/li_247_n17# _551_/li_0_n17#
+ FILLER_20_510/li_0_n17# PHY_345/li_0_527# mprj_dat_buf\[15\]/li_795_379# la_buf\[50\]/li_523_n17#
+ user_to_mprj_in_gates\[82\]/li_615_527# FILLER_21_493/li_63_527# la_buf\[58\]/li_795_379#
+ FILLER_10_1931/li_155_n17# FILLER_24_1482/li_63_n17# la_buf\[28\]/li_611_17# FILLER_11_2022/li_63_527#
+ _338_/li_0_n17# FILLER_25_733/li_155_n17# _590_/li_0_n17# FILLER_12_1791/li_0_527#
+ user_to_mprj_in_buffers\[90\]/li_523_527# la_buf\[29\]/li_431_n17# powergood_check/FILLER_0_248/li_161_797#
+ user_to_mprj_oen_buffers\[82\]/li_983_n17# FILLER_16_1585/li_0_n17# user_to_mprj_oen_buffers\[25\]/li_215_311#
+ ANTENNA__610__A/li_63_527# user_to_mprj_oen_buffers\[5\]/li_707_527# user_to_mprj_in_gates\[69\]/li_339_n17#
+ _540_/li_155_527# user_to_mprj_in_gates\[84\]/li_707_367# _380_/li_0_n17# FILLER_21_2101/li_63_n17#
+ user_to_mprj_in_gates\[3\]/li_247_n17# user_to_mprj_in_gates\[91\]/li_615_n17# powergood_check/FILLER_2_195/li_449_n17#
+ mprj_adr_buf\[22\]/li_1535_n17# user_to_mprj_oen_buffers\[93\]/li_795_379# user_to_mprj_in_gates\[82\]/li_63_n17#
+ user_to_mprj_oen_buffers\[15\]/li_63_n17# FILLER_22_1522/li_63_527# FILLER_16_355/li_0_n17#
+ ANTENNA_user_to_mprj_in_gates\[82\]_B/li_63_n17# ANTENNA_user_to_mprj_in_gates\[54\]_B/li_63_527#
+ _331_/li_155_n17# FILLER_11_484/li_0_n17# _450_/li_0_527# user_to_mprj_oen_buffers\[68\]/li_207_51#
+ FILLER_10_1249/li_63_527# FILLER_13_1704/li_0_527# la_buf\[35\]/li_707_n17# ANTENNA_user_to_mprj_oen_buffers\[50\]_A/li_63_527#
+ user_to_mprj_oen_buffers\[58\]/li_611_17# mprj_clk2_buf/li_17_51# la_buf\[86\]/li_1259_527#
+ user_to_mprj_in_buffers\[15\]/li_404_367# mprj_dat_buf\[0\]/li_207_51# mprj_dat_buf\[13\]/li_431_n17#
+ FILLER_21_406/li_0_n17# FILLER_11_744/li_155_n17# FILLER_25_1770/li_63_n17# FILLER_26_1247/li_0_527#
+ FILLER_17_1405/li_63_n17# ANTENNA__371__A/li_0_527# FILLER_11_1601/li_0_n17# FILLER_7_1148/li_63_n17#
+ la_buf\[120\]/li_17_51# _549_/li_0_527# user_to_mprj_oen_buffers\[13\]/li_215_311#
+ user_to_mprj_in_gates\[57\]/li_339_n17# _659_/li_247_527# user_to_mprj_in_gates\[19\]/li_707_367#
+ user_to_mprj_oen_buffers\[70\]/li_207_51# user_to_mprj_in_gates\[72\]/li_707_367#
+ user_to_mprj_oen_buffers\[60\]/li_1075_n17# FILLER_16_334/li_0_527# ANTENNA__649__A/li_63_n17#
+ user_to_mprj_oen_buffers\[94\]/li_983_527# PHY_740/li_0_527# _397_/li_155_n17# user_to_mprj_in_gates\[107\]/li_0_n17#
+ powergood_check/FILLER_1_62/li_737_797# user_to_mprj_oen_buffers\[51\]/li_779_17#
+ user_to_mprj_in_gates\[4\]/li_431_n17# la_buf\[72\]/li_523_n17# FILLER_22_1886/li_63_n17#
+ FILLER_23_60/li_0_n17# PHY_777/li_0_n17# user_to_mprj_oen_buffers\[91\]/li_431_n17#
+ ANTENNA__573__A/li_63_n17# user_to_mprj_oen_buffers\[68\]/li_707_n17# FILLER_11_1813/li_63_527#
+ powergood_check/FILLER_0_104/li_257_797# user_to_mprj_in_buffers\[46\]/li_523_n17#
+ FILLER_9_1809/li_155_527# FILLER_9_563/li_63_n17# _513_/li_0_527# la_buf\[32\]/li_207_51#
+ powergood_check/FILLER_1_115/li_641_n17# user_to_mprj_oen_buffers\[83\]/li_63_n17#
+ user_to_mprj_in_buffers\[2\]/li_155_n17# mprj_adr_buf\[18\]/li_17_51# FILLER_12_685/li_63_n17#
+ _401_/li_0_527# powergood_check/FILLER_1_212/li_0_n17# FILLER_25_1008/li_63_n17#
+ la_buf\[101\]/li_611_17# user_to_mprj_in_gates\[45\]/li_339_n17# FILLER_16_1585/li_63_527#
+ FILLER_9_338/li_0_n17# user_to_mprj_oen_buffers\[90\]/li_707_n17# FILLER_9_1001/li_63_527#
+ PHY_452/li_0_527# mprj_adr_buf\[19\]/li_215_311# la_buf\[4\]/li_63_527# FILLER_25_1047/li_63_n17#
+ user_to_mprj_oen_buffers\[124\]/li_207_51# powergood_check/FILLER_2_115/li_353_n17#
+ user_to_mprj_oen_buffers\[29\]/li_431_527# user_to_mprj_oen_buffers\[97\]/li_983_527#
+ la_buf\[84\]/li_247_n17# _576_/li_155_n17# FILLER_13_1115/li_63_n17# la_buf\[98\]/li_891_n17#
+ FILLER_18_295/li_0_527# mprj_rstn_buf/li_1167_527# la_buf\[98\]/li_207_51# ANTENNA__357__A/li_0_n17#
+ _636_/li_0_527# user_to_mprj_in_gates\[95\]/li_18_51# powergood_check/FILLER_2_155/li_641_n17#
+ FILLER_26_995/li_155_527# user_to_mprj_oen_buffers\[52\]/li_891_n17# powergood_check/FILLER_2_0/li_100_536#
+ user_to_mprj_in_gates\[19\]/li_63_n17# powergood_check/FILLER_1_196/li_257_n17#
+ PHY_458/li_0_n17# la_buf\[60\]/li_0_527# _366_/li_155_527# ANTENNA__657__A/li_63_527#
+ la_buf\[70\]/li_17_51# user_to_mprj_oen_buffers\[119\]/li_63_527# _586_/li_247_527#
+ FILLER_16_1927/li_0_527# FILLER_13_1704/li_63_n17# FILLER_13_1217/li_63_n17# powergood_check/FILLER_0_256/li_0_797#
+ user_to_mprj_in_buffers\[90\]/li_615_527# mprj_dat_buf\[18\]/li_247_527# user_to_mprj_oen_buffers\[77\]/li_17_51#
+ powergood_check/FILLER_2_0/li_449_797# FILLER_20_1778/li_63_527# FILLER_10_621/li_155_527#
+ PHY_295/li_0_527# _490_/li_247_527# la_buf\[89\]/li_17_51# FILLER_12_1017/li_63_527#
+ PHY_67/li_0_527# la_buf\[72\]/li_247_n17# FILLER_12_1927/li_0_527# FILLER_25_1422/li_155_n17#
+ user_to_mprj_in_gates\[86\]/li_707_n17# mprj_adr_buf\[1\]/li_215_311# user_to_mprj_in_gates\[14\]/li_615_n17#
+ powergood_check/FILLER_0_224/li_65_797# FILLER_10_1174/li_0_n17# la_buf\[4\]/li_1167_527#
+ FILLER_13_1631/li_63_n17# PHY_183/li_0_527# FILLER_9_1038/li_63_n17# PHY_397/li_0_527#
+ powergood_check/FILLER_0_112/li_65_797# FILLER_21_1335/li_0_n17# user_to_mprj_in_gates\[44\]/li_18_51#
+ FILLER_26_917/li_63_527# powergood_check/FILLER_0_96/li_545_797# FILLER_18_1945/li_63_527#
+ user_to_mprj_oen_buffers\[56\]/li_983_n17# user_to_mprj_in_gates\[127\]/li_155_527#
+ la_buf\[89\]/li_891_527# user_to_mprj_oen_buffers\[110\]/li_1259_n17# la_buf\[35\]/li_611_17#
+ FILLER_13_472/li_63_n17# powergood_check/FILLER_2_235/li_353_797# FILLER_12_1796/li_63_n17#
+ user_to_mprj_oen_buffers\[26\]/li_17_51# _336_/li_155_n17# FILLER_25_1261/li_63_527#
+ user_to_mprj_in_gates\[74\]/li_707_n17# mprj_dat_buf\[23\]/li_0_527# _635_/li_155_n17#
+ PHY_412/li_0_n17# user_to_mprj_in_gates\[1\]/li_707_367# user_to_mprj_in_buffers\[44\]/li_51_367#
+ FILLER_19_1728/li_0_527# la_buf\[95\]/li_1259_n17# la_buf\[89\]/li_215_311# la_buf\[38\]/li_17_51#
+ _362_/li_0_527# powergood_check/FILLER_1_156/li_65_797# FILLER_11_992/li_63_n17#
+ mprj_clk_buf/li_707_n17# FILLER_10_463/li_155_n17# _590_/li_247_n17# mprj_dat_buf\[5\]/li_207_51#
+ user_to_mprj_in_buffers\[76\]/li_51_17# user_to_mprj_in_gates\[56\]/li_431_n17#
+ FILLER_8_978/li_63_527# FILLER_13_309/li_63_n17# FILLER_25_544/li_155_527# FILLER_14_45/li_0_n17#
+ user_to_mprj_in_gates\[54\]/li_155_527# user_to_mprj_oen_buffers\[86\]/li_523_n17#
+ la_buf\[41\]/li_523_n17# _580_/li_0_n17# FILLER_19_1609/li_63_527# FILLER_12_1539/li_63_n17#
+ FILLER_23_1520/li_0_527# user_to_mprj_oen_buffers\[75\]/li_207_51# la_buf\[12\]/li_1167_527#
+ PHY_343/li_0_527# FILLER_22_1965/li_0_527# la_buf\[4\]/li_707_527# _367_/li_0_n17#
+ user_to_mprj_oen_buffers\[59\]/li_1167_n17# powergood_check/FILLER_1_236/li_641_n17#
+ FILLER_19_1331/li_155_527# powergood_check/FILLER_0_256/li_353_797# la_buf\[84\]/li_1075_n17#
+ mprj_adr_buf\[29\]/li_707_527# mprj_dat_buf\[1\]/li_795_379# user_to_mprj_oen_buffers\[56\]/li_779_17#
+ powergood_check/FILLER_2_227/li_161_n17# la_buf\[82\]/li_63_527# mprj_stb_buf/li_523_n17#
+ user_to_mprj_in_gates\[71\]/li_155_n17# powergood_check/FILLER_0_176/li_161_797#
+ la_buf\[45\]/li_891_527# FILLER_13_756/li_63_527# la_buf\[77\]/li_215_311# FILLER_14_1521/li_63_n17#
+ user_to_mprj_in_gates\[124\]/li_155_n17# la_buf\[37\]/li_207_51# FILLER_13_1587/li_155_527#
+ FILLER_27_806/li_0_n17# FILLER_13_2020/li_0_n17# FILLER_16_44/li_0_n17# FILLER_5_1087/li_155_527#
+ user_to_mprj_in_gates\[44\]/li_615_527# user_to_mprj_in_gates\[123\]/li_707_n17#
+ user_to_mprj_oen_buffers\[74\]/li_523_n17# FILLER_10_459/li_155_n17# la_buf\[100\]/li_207_51#
+ FILLER_15_1390/li_63_n17# _340_/li_247_n17# PHY_471/li_0_n17# FILLER_14_2096/li_63_n17#
+ user_to_mprj_oen_buffers\[83\]/li_1443_n17# FILLER_12_1697/li_0_n17# user_to_mprj_in_gates\[105\]/li_431_n17#
+ la_buf\[9\]/li_63_527# user_to_mprj_in_gates\[7\]/li_155_527# FILLER_14_1521/li_0_527#
+ PHY_392/li_0_n17# PHY_808/li_0_n17# user_to_mprj_in_gates\[51\]/li_155_n17# user_to_mprj_oen_buffers\[81\]/li_707_527#
+ FILLER_25_853/li_0_n17# FILLER_28_51/li_63_n17# user_to_mprj_oen_buffers\[81\]/li_247_n17#
+ FILLER_12_748/li_63_n17# FILLER_9_825/li_155_527# user_to_mprj_in_gates\[50\]/li_707_n17#
+ powergood_check/FILLER_0_112/li_100_536# la_buf\[65\]/li_215_311# user_to_mprj_in_gates\[38\]/li_339_n17#
+ FILLER_14_509/li_0_n17# la_buf\[75\]/li_0_527# user_to_mprj_in_buffers\[69\]/li_236_17#
+ user_to_mprj_in_gates\[112\]/li_155_n17# user_to_mprj_oen_buffers\[7\]/li_1259_527#
+ user_to_mprj_in_gates\[60\]/li_431_n17# user_to_mprj_oen_buffers\[2\]/li_215_311#
+ la_buf\[98\]/li_1075_n17# user_to_mprj_in_gates\[30\]/li_155_527# FILLER_24_1652/li_0_527#
+ mprj_adr_buf\[26\]/li_707_n17# user_to_mprj_oen_buffers\[62\]/li_523_n17# user_to_mprj_in_gates\[111\]/li_707_n17#
+ _654_/li_0_527# mprj_adr_buf\[17\]/li_17_51# FILLER_20_1419/li_0_527# FILLER_12_1503/li_63_527#
+ FILLER_23_1503/li_63_n17# _583_/li_155_n17# FILLER_25_1341/li_0_527# powergood_check/FILLER_0_112/li_449_797#
+ FILLER_22_520/li_155_n17# user_to_mprj_in_gates\[104\]/li_339_n17# la_buf\[113\]/li_891_527#
+ user_to_mprj_in_buffers\[71\]/li_236_17# la_buf\[83\]/li_1351_527# FILLER_23_1629/li_155_527#
+ _581_/li_0_527# user_to_mprj_in_gates\[26\]/li_63_n17# FILLER_7_1148/li_63_527#
+ la_buf\[6\]/li_1351_527# _373_/li_155_527# FILLER_19_1573/li_63_n17# user_to_mprj_oen_buffers\[98\]/li_215_311#
+ powergood_check/FILLER_1_196/li_0_797# la_buf\[53\]/li_215_311# _368_/li_0_527#
+ powergood_check/FILLER_1_16/li_115_72# mprj_dat_buf\[23\]/li_615_527# powergood_check/FILLER_0_264/li_115_72#
+ user_to_mprj_in_gates\[100\]/li_155_n17# FILLER_25_1126/li_155_n17# user_to_mprj_in_gates\[92\]/li_523_n17#
+ user_to_mprj_in_gates\[94\]/li_18_51# user_to_mprj_in_gates\[90\]/li_247_527# la_buf\[69\]/li_983_n17#
+ powergood_check/FILLER_1_62/li_737_n17# user_to_mprj_oen_buffers\[50\]/li_523_n17#
+ FILLER_13_1071/li_155_527# la_buf\[19\]/li_63_527# FILLER_18_170/li_0_527# FILLER_21_70/li_155_527#
+ user_to_mprj_oen_buffers\[114\]/li_63_n17# user_to_mprj_oen_buffers\[14\]/li_207_51#
+ user_to_mprj_oen_buffers\[66\]/li_63_527# user_to_mprj_in_gates\[49\]/li_247_527#
+ user_to_mprj_oen_buffers\[20\]/li_707_n17# user_to_mprj_in_gates\[71\]/li_523_527#
+ mprj_cyc_buf/li_1167_n17# FILLER_11_733/li_63_n17# user_to_mprj_in_buffers\[88\]/li_404_367#
+ user_to_mprj_oen_buffers\[76\]/li_17_51# mprj_cyc_buf/li_17_51# FILLER_10_621/li_63_n17#
+ la_buf\[88\]/li_17_51# _552_/li_155_527# la_buf\[21\]/li_63_527# la_buf\[79\]/li_0_527#
+ FILLER_13_655/li_0_527# user_to_mprj_oen_buffers\[86\]/li_215_311# la_buf\[41\]/li_215_311#
+ user_to_mprj_oen_buffers\[16\]/li_247_n17# FILLER_9_627/li_63_527# la_buf\[125\]/li_215_311#
+ la_buf\[42\]/li_611_17# FILLER_7_1128/li_63_527# user_to_mprj_in_buffers\[69\]/li_155_n17#
+ user_to_mprj_oen_buffers\[60\]/li_1535_n17# FILLER_12_1796/li_0_527# FILLER_12_1374/li_63_527#
+ user_to_mprj_in_gates\[43\]/li_18_51# la_buf\[5\]/li_215_311# FILLER_9_1138/li_155_n17#
+ FILLER_13_1660/li_63_n17# _343_/li_155_n17# FILLER_9_394/li_155_527# PHY_467/li_0_n17#
+ powergood_check/FILLER_1_0/li_65_n17# _643_/li_0_n17# user_to_mprj_oen_buffers\[91\]/li_1443_n17#
+ FILLER_9_582/li_155_n17# PHY_460/li_0_n17# ANTENNA__655__A/li_0_n17# mprj_stb_buf/li_215_311#
+ powergood_check/mprj2_logic_high_lv/li_384_137# powergood_check/FILLER_2_203/li_257_797#
+ la_buf\[58\]/li_63_527# _337_/li_0_527# mprj_adr_buf\[11\]/li_207_51# ANTENNA__639__A/li_63_n17#
+ FILLER_25_1004/li_155_n17# FILLER_25_1506/li_0_527# user_to_mprj_oen_buffers\[25\]/li_17_51#
+ user_to_mprj_oen_buffers\[5\]/li_795_379# user_to_mprj_in_gates\[114\]/li_247_527#
+ user_to_mprj_oen_buffers\[82\]/li_207_51# user_to_mprj_oen_buffers\[74\]/li_215_311#
+ la_buf\[70\]/li_615_527# FILLER_10_1184/li_63_n17# user_to_mprj_in_buffers\[2\]/li_615_n17#
+ la_buf\[37\]/li_17_51# user_to_mprj_in_gates\[120\]/li_523_527# FILLER_10_621/li_63_527#
+ FILLER_19_1446/li_155_527# powergood_check/FILLER_2_243/li_545_797# powergood_check/FILLER_2_0/li_449_n17#
+ powergood_check/FILLER_1_62/li_257_797# FILLER_14_1662/li_63_527# la_buf\[113\]/li_215_311#
+ FILLER_12_1927/li_63_527# mprj_dat_buf\[8\]/li_983_527# FILLER_16_1589/li_155_527#
+ FILLER_11_1274/li_155_n17# la_buf\[105\]/li_207_51# user_to_mprj_oen_buffers\[63\]/li_779_17#
+ powergood_check/FILLER_2_163/li_353_797# FILLER_25_222/li_0_527# user_to_mprj_oen_buffers\[23\]/li_1167_n17#
+ user_to_mprj_in_gates\[118\]/li_615_n17# powergood_check/FILLER_1_115/li_161_n17#
+ powergood_check/FILLER_1_204/li_545_n17# mprj_dat_buf\[1\]/li_215_311# user_to_mprj_in_gates\[107\]/li_707_n17#
+ powergood_check/FILLER_0_224/li_257_797# user_to_mprj_in_gates\[25\]/li_247_527#
+ la_buf\[9\]/li_983_n17# _478_/li_247_n17# la_buf\[44\]/li_207_51# _357_/li_0_n17#
+ user_to_mprj_oen_buffers\[95\]/li_63_n17# la_buf\[76\]/li_1351_527# FILLER_17_350/li_0_527#
+ powergood_check/FILLER_0_96/li_545_n17# FILLER_0_232/li_63_527# FILLER_11_1433/li_63_n17#
+ powergood_check/FILLER_0_264/li_545_797# FILLER_14_456/li_63_n17# FILLER_11_1584/li_63_n17#
+ user_to_mprj_oen_buffers\[62\]/li_215_311# FILLER_19_249/li_0_n17# user_to_mprj_in_gates\[34\]/li_247_n17#
+ FILLER_0_1326/li_155_527# powergood_check/FILLER_2_235/li_353_n17# FILLER_11_1472/li_63_n17#
+ powergood_check/FILLER_1_164/li_641_n17# FILLER_9_1001/li_0_527# la_buf\[87\]/li_1351_527#
+ la_buf\[101\]/li_215_311# PHY_454/li_0_527# FILLER_14_1662/li_63_n17# user_to_mprj_in_buffers\[42\]/li_155_n17#
+ powergood_check/FILLER_0_184/li_353_797# _588_/li_155_n17# user_to_mprj_oen_buffers\[82\]/li_1259_n17#
+ mprj_dat_buf\[18\]/li_707_527# la_buf\[45\]/li_431_527# powergood_check/FILLER_2_155/li_161_n17#
+ FILLER_9_559/li_0_n17# _402_/li_155_n17# PHY_370/li_0_527# user_to_mprj_oen_buffers\[117\]/li_779_17#
+ FILLER_11_992/li_63_527# user_to_mprj_in_buffers\[76\]/li_236_17# FILLER_17_1925/li_0_n17#
+ powergood_check/FILLER_1_0/li_353_n17# FILLER_11_1196/li_63_n17# la_buf\[44\]/li_795_379#
+ mprj_we_buf/li_63_527# powergood_check/FILLER_0_24/li_641_797# FILLER_5_617/li_0_527#
+ FILLER_19_109/li_63_527# _378_/li_155_527# FILLER_14_1510/li_63_527# mprj_dat_buf\[27\]/li_707_n17#
+ _588_/li_247_n17# _590_/li_155_n17# FILLER_12_1035/li_0_527# la_buf\[67\]/li_983_527#
+ user_to_mprj_oen_buffers\[50\]/li_215_311# mprj_adr_buf\[29\]/li_1351_527# FILLER_24_56/li_63_n17#
+ user_to_mprj_oen_buffers\[24\]/li_615_527# FILLER_25_1176/li_155_n17# FILLER_12_1503/li_63_n17#
+ FILLER_11_916/li_63_527# FILLER_14_1543/li_155_527# powergood_check/FILLER_1_220/li_0_797#
+ user_to_mprj_oen_buffers\[56\]/li_1443_n17# FILLER_12_689/li_155_n17# FILLER_24_1421/li_155_527#
+ ANTENNA_user_to_mprj_in_gates\[50\]_A/li_63_n17# mprj_adr_buf\[16\]/li_17_51# _380_/li_155_527#
+ FILLER_17_1457/li_0_527# user_to_mprj_in_gates\[73\]/li_155_527# powergood_check/FILLER_2_107/li_65_797#
+ user_to_mprj_oen_buffers\[19\]/li_207_51# user_to_mprj_oen_buffers\[85\]/li_611_17#
+ FILLER_17_56/li_0_n17# FILLER_13_2012/li_0_n17# FILLER_9_582/li_63_n17# FILLER_26_939/li_63_527#
+ user_to_mprj_oen_buffers\[45\]/li_983_527# ANTENNA_user_to_mprj_oen_buffers\[63\]_A/li_63_n17#
+ PHY_299/li_0_527# user_to_mprj_in_buffers\[40\]/li_404_367# user_to_mprj_oen_buffers\[4\]/li_891_527#
+ mprj_dat_buf\[15\]/li_707_n17# FILLER_12_890/li_155_n17# la_buf\[26\]/li_63_527#
+ ANTENNA_user_to_mprj_in_gates\[107\]_B/li_63_527# user_to_mprj_in_gates\[54\]/li_615_527#
+ user_to_mprj_oen_buffers\[21\]/li_207_51# FILLER_23_489/li_155_n17# mprj_cyc_buf/li_707_527#
+ _358_/li_0_527# la_buf\[6\]/li_431_n17# mprj_sel_buf\[3\]/li_983_527# user_to_mprj_oen_buffers\[76\]/li_1075_527#
+ FILLER_9_1127/li_155_n17# user_to_mprj_in_gates\[93\]/li_18_51# user_to_mprj_oen_buffers\[60\]/li_0_n17#
+ _348_/li_155_n17# _397_/li_0_527# ANTENNA__332__A/li_63_n17# la_buf\[21\]/li_431_527#
+ _647_/li_155_n17# user_to_mprj_oen_buffers\[42\]/li_983_527# FILLER_5_857/li_155_527#
+ la_buf\[3\]/li_707_527# mprj_dat_buf\[20\]/li_1167_527# user_to_mprj_in_gates\[56\]/li_707_367#
+ _391_/li_247_527# user_to_mprj_in_gates\[61\]/li_339_527# user_to_mprj_oen_buffers\[85\]/li_1075_n17#
+ powergood_check/FILLER_1_8/li_641_n17# powergood_check/mprj_logic_high_lv/li_0_1611#
+ FILLER_10_463/li_0_527# FILLER_16_1421/li_155_n17# user_to_mprj_in_buffers\[72\]/li_615_n17#
+ la_buf\[21\]/li_0_527# mprj_adr_buf\[16\]/li_207_51# FILLER_11_1210/li_63_527# FILLER_19_56/li_0_n17#
+ user_to_mprj_in_gates\[117\]/li_707_367# mprj_adr_buf\[9\]/li_215_311# user_to_mprj_in_gates\[124\]/li_615_n17#
+ user_to_mprj_oen_buffers\[75\]/li_17_51# FILLER_15_2107/li_155_527# _350_/li_155_n17#
+ powergood_check/FILLER_1_236/li_161_n17# _437_/li_155_527# user_to_mprj_oen_buffers\[87\]/li_207_51#
+ FILLER_9_1179/li_0_527# PHY_840/li_0_527# powergood_check/FILLER_2_8/li_257_797#
+ FILLER_25_1827/li_0_527# user_to_mprj_in_gates\[46\]/li_247_527# la_buf\[87\]/li_17_51#
+ la_buf\[95\]/li_1535_527# la_buf\[114\]/li_431_n17# PHY_479/li_0_527# la_buf\[28\]/li_0_n17#
+ powergood_check/FILLER_1_32/li_641_n17# user_to_mprj_in_gates\[42\]/li_18_51# user_to_mprj_oen_buffers\[54\]/li_431_527#
+ user_to_mprj_oen_buffers\[40\]/li_1443_n17# la_buf\[94\]/li_63_527# powergood_check/FILLER_2_195/li_65_n17#
+ _527_/li_155_n17# user_to_mprj_in_gates\[44\]/li_707_367# mprj_dat_buf\[27\]/li_63_n17#
+ FILLER_10_471/li_0_n17# user_to_mprj_in_gates\[51\]/li_615_n17# powergood_check/FILLER_2_211/li_100_536#
+ FILLER_18_539/li_63_527# powergood_check/FILLER_1_212/li_115_72# user_to_mprj_oen_buffers\[22\]/li_707_527#
+ la_buf\[49\]/li_207_51# FILLER_17_1570/li_63_n17# _439_/li_247_527# user_to_mprj_oen_buffers\[53\]/li_795_379#
+ la_buf\[112\]/li_207_51# powergood_check/FILLER_1_131/li_0_797# FILLER_24_1758/li_0_n17#
+ ANTENNA_la_buf\[110\]_A/li_63_527# user_to_mprj_in_gates\[112\]/li_615_n17# user_to_mprj_oen_buffers\[63\]/li_431_n17#
+ user_to_mprj_in_gates\[110\]/li_339_527# powergood_check/FILLER_0_88/li_115_72#
+ user_to_mprj_oen_buffers\[24\]/li_17_51# FILLER_17_507/li_0_n17# powergood_check/FILLER_1_140/li_737_797#
+ powergood_check/FILLER_2_211/li_449_797# user_to_mprj_in_gates\[30\]/li_615_527#
+ la_buf\[36\]/li_17_51# _654_/li_247_527# la_buf\[51\]/li_207_51# user_to_mprj_oen_buffers\[30\]/li_983_n17#
+ user_to_mprj_oen_buffers\[39\]/li_0_n17# FILLER_10_785/li_63_n17# powergood_check/FILLER_0_232/li_100_536#
+ user_to_mprj_in_gates\[32\]/li_707_367# _560_/li_0_n17# FILLER_15_230/li_63_527#
+ la_buf\[40\]/li_1351_527# FILLER_19_1446/li_155_n17# ANTENNA_la_buf\[15\]_A/li_63_n17#
+ ANTENNA__349__A/li_0_527# powergood_check/FILLER_2_171/li_545_797# ANTENNA_la_buf\[127\]_A/li_63_n17#
+ powergood_check/FILLER_1_220/li_0_n17# _595_/li_155_n17# user_to_mprj_in_gates\[100\]/li_615_n17#
+ user_to_mprj_oen_buffers\[51\]/li_431_n17# powergood_check/FILLER_0_232/li_449_797#
+ PHY_268/li_0_527# FILLER_22_2092/li_155_527# _386_/li_0_n17# la_buf\[90\]/li_891_527#
+ user_to_mprj_oen_buffers\[124\]/li_779_17# FILLER_7_942/li_63_527# powergood_check/FILLER_2_203/li_257_n17#
+ la_buf\[26\]/li_1351_n17# mprj_cyc_buf/li_615_527# FILLER_11_1462/li_63_n17# mprj_adr_buf\[20\]/li_215_311#
+ user_to_mprj_oen_buffers\[68\]/li_1351_527# FILLER_15_335/li_0_n17# user_to_mprj_in_gates\[38\]/li_63_n17#
+ powergood_check/FILLER_0_272/li_737_797# mprj_dat_buf\[11\]/li_207_51# la_buf\[98\]/li_779_17#
+ FILLER_12_1623/li_0_n17# powergood_check/FILLER_2_259/li_115_72# _461_/li_247_527#
+ user_to_mprj_oen_buffers\[62\]/li_1167_n17# mprj_dat_buf\[13\]/li_1351_527# powergood_check/FILLER_2_243/li_545_n17#
+ ANTENNA_user_to_mprj_in_gates\[118\]_A/li_63_527# powergood_check/FILLER_1_62/li_257_n17#
+ powergood_check/FILLER_0_192/li_545_797# FILLER_6_1013/li_155_n17# user_to_mprj_in_gates\[59\]/li_155_n17#
+ mprj_sel_buf\[2\]/li_983_527# la_buf\[122\]/li_1167_n17# PHY_792/li_0_527# user_to_mprj_oen_buffers\[75\]/li_611_17#
+ powergood_check/FILLER_2_163/li_353_n17# user_to_mprj_in_gates\[40\]/li_63_n17#
+ user_to_mprj_oen_buffers\[16\]/li_707_n17# powergood_check/FILLER_2_227/li_0_797#
+ FILLER_15_1802/li_63_527# user_to_mprj_in_gates\[105\]/li_0_n17# user_to_mprj_oen_buffers\[26\]/li_207_51#
+ user_to_mprj_in_buffers\[69\]/li_615_n17# FILLER_12_1117/li_0_n17# FILLER_21_1448/li_63_527#
+ mprj_clk2_buf/li_63_527# user_to_mprj_in_gates\[61\]/li_615_527# user_to_mprj_in_buffers\[61\]/li_236_367#
+ la_buf\[14\]/li_0_n17# la_buf\[29\]/li_0_n17# user_to_mprj_in_buffers\[79\]/li_615_527#
+ FILLER_18_528/li_63_n17# user_to_mprj_in_gates\[60\]/li_431_527# user_to_mprj_oen_buffers\[93\]/li_1259_527#
+ _634_/li_0_527# mprj_adr_buf\[15\]/li_17_51# FILLER_17_1520/li_63_n17# la_buf\[123\]/li_0_n17#
+ mprj_stb_buf/li_983_527# user_to_mprj_in_buffers\[45\]/li_615_527# user_to_mprj_in_gates\[81\]/li_0_527#
+ user_to_mprj_in_buffers\[3\]/li_523_n17# user_to_mprj_oen_buffers\[44\]/li_523_n17#
+ user_to_mprj_in_gates\[47\]/li_155_n17# FILLER_7_1148/li_0_n17# ANTENNA_user_to_mprj_oen_buffers\[55\]_TE/li_63_n17#
+ powergood_check/FILLER_1_188/li_65_n17# FILLER_15_96/li_0_n17# _410_/li_0_527# user_to_mprj_in_gates\[43\]/li_247_527#
+ FILLER_9_1097/li_0_527# la_buf\[70\]/li_1075_n17# _355_/li_155_n17# FILLER_9_1273/li_63_527#
+ la_buf\[104\]/li_247_n17# FILLER_12_1931/li_155_527# user_to_mprj_in_gates\[78\]/li_0_n17#
+ _530_/li_0_527# FILLER_25_949/li_0_n17# user_to_mprj_in_gates\[28\]/li_431_n17#
+ powergood_check/FILLER_2_251/li_641_797# mprj_adr_buf\[23\]/li_207_51# user_to_mprj_oen_buffers\[56\]/li_247_527#
+ la_buf\[14\]/li_0_527# user_to_mprj_in_gates\[92\]/li_18_51# ANTENNA_user_to_mprj_in_gates\[36\]_A/li_63_n17#
+ user_to_mprj_oen_buffers\[94\]/li_207_51# la_buf\[109\]/li_891_527# mprj_adr_buf\[24\]/li_891_n17#
+ powergood_check/FILLER_0_8/li_65_797# la_buf\[90\]/li_215_311# user_to_mprj_oen_buffers\[103\]/li_1535_n17#
+ user_to_mprj_in_gates\[39\]/li_615_n17# powergood_check/FILLER_2_219/li_65_n17#
+ la_buf\[95\]/li_707_527# la_buf\[117\]/li_207_51# user_to_mprj_in_gates\[34\]/li_707_n17#
+ FILLER_11_1351/li_63_527# powergood_check/FILLER_2_107/li_65_n17# la_buf\[49\]/li_215_311#
+ user_to_mprj_oen_buffers\[74\]/li_17_51# _534_/li_155_n17# mprj_cyc_buf/li_1535_n17#
+ user_to_mprj_in_gates\[86\]/li_0_n17# la_buf\[86\]/li_17_51# user_to_mprj_in_gates\[88\]/li_523_n17#
+ la_buf\[56\]/li_207_51# FILLER_9_719/li_63_527# user_to_mprj_in_buffers\[109\]/li_236_17#
+ user_to_mprj_in_gates\[86\]/li_247_527# FILLER_21_1405/li_155_n17# powergood_check/FILLER_2_16/li_353_797#
+ powergood_check/FILLER_0_248/li_0_n17# _346_/li_0_527# user_to_mprj_in_gates\[41\]/li_18_51#
+ FILLER_20_1625/li_63_527# powergood_check/FILLER_1_164/li_161_n17# _623_/li_155_527#
+ FILLER_7_921/li_155_527# mprj_adr_buf\[7\]/li_1259_527# user_to_mprj_in_gates\[95\]/li_247_n17#
+ FILLER_10_578/li_63_n17# powergood_check/FILLER_0_272/li_65_797# la_buf\[52\]/li_615_527#
+ _337_/li_247_n17# la_buf\[37\]/li_523_n17# FILLER_23_1778/li_155_527# FILLER_25_1343/li_63_527#
+ powergood_check/FILLER_0_160/li_65_797# la_buf\[37\]/li_215_311# mprj_adr_buf\[11\]/li_795_379#
+ ANTENNA__563__A/li_63_527# FILLER_9_582/li_155_527# mprj_adr_buf\[11\]/li_779_17#
+ user_to_mprj_oen_buffers\[23\]/li_17_51# powergood_check/FILLER_0_24/li_161_797#
+ user_to_mprj_in_gates\[74\]/li_247_527# la_buf\[35\]/li_17_51# FILLER_9_600/li_155_n17#
+ mprj_dat_buf\[27\]/li_1167_n17# FILLER_13_699/li_155_527# FILLER_28_51/li_63_527#
+ mprj_dat_buf\[16\]/li_207_51# FILLER_25_819/li_155_n17# FILLER_25_1241/li_0_n17#
+ mprj_dat_buf\[9\]/li_215_311# powergood_check/FILLER_2_8/li_257_n17# FILLER_11_1749/li_63_n17#
+ _550_/li_0_n17# user_to_mprj_oen_buffers\[83\]/li_0_527# PHY_278/li_0_n17# FILLER_25_1648/li_155_n17#
+ user_to_mprj_in_gates\[83\]/li_247_n17# FILLER_22_1909/li_63_527# FILLER_13_1574/li_0_527#
+ _337_/li_0_n17# FILLER_24_1628/li_63_n17# user_to_mprj_in_gates\[45\]/li_63_n17#
+ mprj_adr_buf\[26\]/li_611_17# _392_/li_155_527# la_buf\[6\]/li_1075_n17# ANTENNA_la_buf\[109\]_TE/li_63_n17#
+ FILLER_21_1741/li_0_n17# mprj_dat_buf\[21\]/li_215_311# FILLER_11_1035/li_0_n17#
+ la_buf\[10\]/li_891_n17# FILLER_3_893/li_155_n17# FILLER_25_1096/li_63_527# la_buf\[25\]/li_215_311#
+ powergood_check/mprj_logic_high_lv/li_737_1611# la_buf\[127\]/li_1351_527# user_to_mprj_in_gates\[116\]/li_523_527#
+ la_buf\[50\]/li_1167_527# mprj_dat_buf\[29\]/li_63_n17# la_buf\[4\]/li_615_527#
+ powergood_check/FILLER_0_160/li_100_536# FILLER_25_849/li_0_n17# user_to_mprj_oen_buffers\[126\]/li_215_311#
+ la_buf\[109\]/li_215_311# PHY_467/li_0_527# mprj_logic_high_inst/m2_572_856# powergood_check/FILLER_1_131/li_0_n17#
+ FILLER_23_70/li_63_n17# FILLER_9_803/li_0_n17# PHY_240/li_0_n17# user_to_mprj_oen_buffers\[79\]/li_0_n17#
+ user_to_mprj_in_gates\[112\]/li_0_n17# ANTENNA_user_to_mprj_in_gates\[54\]_A/li_63_527#
+ powergood_check/FILLER_1_140/li_737_n17# powergood_check/FILLER_2_211/li_449_n17#
+ FILLER_13_1714/li_63_527# powergood_check/FILLER_0_160/li_449_797# user_to_mprj_in_gates\[123\]/li_247_527#
+ user_to_mprj_oen_buffers\[33\]/li_207_51# la_buf\[101\]/li_63_527# la_buf\[59\]/li_611_17#
+ la_buf\[26\]/li_1351_527# powergood_check/FILLER_2_107/li_100_536# FILLER_13_1199/li_155_n17#
+ FILLER_12_689/li_155_527# FILLER_13_925/li_0_n17# la_buf\[118\]/li_1259_527# mprj_adr_buf\[20\]/li_1167_n17#
+ la_buf\[7\]/li_1351_527# la_buf\[122\]/li_611_17# _660_/li_0_n17# powergood_check/FILLER_2_259/li_0_n17#
+ FILLER_22_1909/li_155_527# user_to_mprj_oen_buffers\[58\]/li_215_311# _571_/li_155_527#
+ la_buf\[13\]/li_215_311# powergood_check/FILLER_1_8/li_161_n17# la_buf\[40\]/li_63_527#
+ mprj_sel_buf\[2\]/li_207_51# FILLER_17_350/li_63_527# la_buf\[99\]/li_1443_527#
+ la_buf\[26\]/li_1259_527# user_to_mprj_oen_buffers\[7\]/li_707_n17# user_to_mprj_in_gates\[21\]/li_431_n17#
+ PHY_325/li_0_n17# powergood_check/FILLER_2_107/li_449_797# user_to_mprj_oen_buffers\[114\]/li_215_311#
+ powergood_check/FILLER_2_171/li_545_n17# user_to_mprj_in_gates\[50\]/li_247_527#
+ mprj_adr_buf\[28\]/li_207_51# FILLER_13_1428/li_63_527# FILLER_13_1816/li_0_527#
+ FILLER_13_2009/li_63_n17# powergood_check/FILLER_2_300/li_65_797# _449_/li_0_527#
+ _362_/li_155_n17# user_to_mprj_oen_buffers\[99\]/li_207_51# mprj_adr_buf\[28\]/li_523_n17#
+ ANTENNA__358__A/li_0_n17# mprj_adr_buf\[14\]/li_17_51# user_to_mprj_in_gates\[111\]/li_247_527#
+ user_to_mprj_oen_buffers\[48\]/li_1167_n17# mprj_adr_buf\[29\]/li_247_527# FILLER_14_1662/li_0_527#
+ powergood_check/FILLER_1_220/li_100_536# FILLER_16_1839/li_155_527# user_to_mprj_in_gates\[31\]/li_523_527#
+ powergood_check/mprj2_logic_high_hvl/li_43_635# powergood_check/FILLER_1_32/li_161_n17#
+ user_to_mprj_oen_buffers\[61\]/li_615_527# PHY_239/li_0_527# user_to_mprj_in_buffers\[48\]/li_404_367#
+ PHY_379/li_0_527# mprj_adr_buf\[30\]/li_207_51# powergood_check/FILLER_0_272/li_737_n17#
+ mprj_dat_buf\[19\]/li_611_17# user_to_mprj_oen_buffers\[46\]/li_215_311# PHY_461/li_0_n17#
+ mprj_dat_buf\[4\]/li_891_527# la_buf\[109\]/li_1075_n17# la_buf\[11\]/li_891_n17#
+ user_to_mprj_oen_buffers\[3\]/li_207_51# la_buf\[96\]/li_1443_527# user_to_mprj_in_gates\[40\]/li_523_n17#
+ user_to_mprj_oen_buffers\[102\]/li_215_311# mprj_dat_buf\[13\]/li_983_n17# mprj_dat_buf\[25\]/li_431_527#
+ la_buf\[124\]/li_207_51# la_buf\[29\]/li_431_527# user_to_mprj_oen_buffers\[82\]/li_779_17#
+ powergood_check/FILLER_1_140/li_257_797# powergood_check/FILLER_2_227/li_0_n17#
+ _441_/li_247_527# user_to_mprj_in_gates\[91\]/li_18_51# la_buf\[5\]/li_983_n17#
+ user_to_mprj_in_gates\[101\]/li_523_n17# user_to_mprj_in_gates\[69\]/li_339_527#
+ powergood_check/FILLER_1_48/li_641_797# _377_/li_0_527# FILLER_0_91/li_0_527# user_to_mprj_in_gates\[75\]/li_155_n17#
+ FILLER_25_945/li_63_n17# la_buf\[63\]/li_207_51# user_to_mprj_in_buffers\[36\]/li_404_367#
+ PHY_298/li_0_527# user_to_mprj_oen_buffers\[1\]/li_1351_527# la_buf\[38\]/li_431_n17#
+ ANTENNA_user_to_mprj_in_gates\[110\]_B/li_63_527# FILLER_13_1017/li_63_n17# user_to_mprj_oen_buffers\[34\]/li_215_311#
+ ANTENNA_user_to_mprj_in_gates\[57\]_B/li_63_n17# user_to_mprj_in_gates\[29\]/li_247_527#
+ _331_/li_155_527# user_to_mprj_in_gates\[78\]/li_339_n17# mprj_dat_buf\[7\]/li_1351_n17#
+ user_to_mprj_oen_buffers\[73\]/li_17_51# mprj_adr_buf\[2\]/li_63_n17# _585_/li_0_527#
+ mprj_dat_buf\[25\]/li_523_n17# la_buf\[85\]/li_17_51# powergood_check/FILLER_1_212/li_257_n17#
+ mprj_adr_buf\[15\]/li_983_527# user_to_mprj_oen_buffers\[25\]/li_1351_527# FILLER_11_1544/li_0_n17#
+ FILLER_20_129/li_0_527# user_to_mprj_oen_buffers\[90\]/li_1259_n17# ANTENNA_user_to_mprj_in_gates\[103\]_A/li_63_n17#
+ user_to_mprj_in_gates\[59\]/li_615_n17# ANTENNA__594__A/li_63_n17# user_to_mprj_in_gates\[40\]/li_18_51#
+ FILLER_15_1688/li_155_527# mprj_dat_buf\[7\]/li_707_527# FILLER_25_638/li_0_n17#
+ powergood_check/FILLER_2_24/li_545_797# user_to_mprj_oen_buffers\[63\]/li_523_n17#
+ powergood_check/FILLER_1_252/li_545_n17# mprj_dat_buf\[3\]/li_1167_527# user_to_mprj_in_buffers\[67\]/li_523_n17#
+ FILLER_14_1447/li_0_527# powergood_check/FILLER_0_272/li_257_797# FILLER_17_1424/li_0_n17#
+ la_buf\[22\]/li_707_527# _399_/li_247_527# user_to_mprj_in_gates\[77\]/li_0_527#
+ mprj_dat_buf\[22\]/li_431_n17# powergood_check/mprj2_logic_high_lv/li_1601_797#
+ _397_/li_155_527# mprj_dat_buf\[23\]/li_207_51# powergood_check/mprj_logic_high_lv/li_384_137#
+ user_to_mprj_in_gates\[103\]/li_63_n17# _650_/li_0_n17# user_to_mprj_in_gates\[118\]/li_339_527#
+ powergood_check/FILLER_0_176/li_0_n17# _394_/li_0_527# user_to_mprj_in_gates\[59\]/li_18_51#
+ user_to_mprj_oen_buffers\[22\]/li_215_311# FILLER_21_184/li_63_n17# user_to_mprj_in_gates\[38\]/li_615_527#
+ user_to_mprj_oen_buffers\[91\]/li_431_527# user_to_mprj_in_gates\[66\]/li_339_n17#
+ _510_/li_155_527# FILLER_3_763/li_63_527# mprj_adr_buf\[7\]/li_891_527# user_to_mprj_in_gates\[81\]/li_707_367#
+ user_to_mprj_oen_buffers\[22\]/li_17_51# PHY_354/li_0_527# user_to_mprj_oen_buffers\[38\]/li_983_n17#
+ FILLER_28_63/li_155_n17# user_to_mprj_oen_buffers\[83\]/li_63_527# la_buf\[34\]/li_17_51#
+ powergood_check/FILLER_2_219/li_257_797# mprj_stb_buf/li_1351_527# _360_/li_0_527#
+ _652_/li_0_n17# powergood_check/mprj2_logic_high_hvl/li_307_57# user_to_mprj_in_gates\[47\]/li_615_n17#
+ powergood_check/FILLER_0_32/li_353_797# FILLER_5_613/li_63_527# user_to_mprj_oen_buffers\[38\]/li_207_51#
+ _569_/li_247_n17# FILLER_9_338/li_0_527# la_buf\[106\]/li_0_527# mprj_dat_buf\[3\]/li_247_527#
+ user_to_mprj_oen_buffers\[6\]/li_611_17# powergood_check/FILLER_2_16/li_353_n17#
+ powergood_check/FILLER_2_259/li_545_797# user_to_mprj_in_gates\[99\]/li_155_527#
+ FILLER_23_1451/li_155_n17# user_to_mprj_oen_buffers\[59\]/li_431_n17# la_buf\[86\]/li_523_n17#
+ la_buf\[2\]/li_983_n17# user_to_mprj_oen_buffers\[105\]/li_795_379# user_to_mprj_in_gates\[106\]/li_339_527#
+ la_buf\[106\]/li_891_527# la_buf\[53\]/li_983_527# user_to_mprj_oen_buffers\[10\]/li_215_311#
+ la_buf\[108\]/li_1259_527# powergood_check/FILLER_1_131/li_34_73# powergood_check/FILLER_2_179/li_353_797#
+ FILLER_11_1666/li_63_n17# PHY_173/li_0_n17# user_to_mprj_oen_buffers\[40\]/li_207_51#
+ FILLER_18_1439/li_63_527# powergood_check/FILLER_1_24/li_65_n17# _366_/li_0_n17#
+ _584_/li_247_n17# FILLER_16_1421/li_63_527# mprj_adr_buf\[28\]/li_215_311# mprj_dat_buf\[28\]/li_0_n17#
+ FILLER_25_1315/li_155_n17# FILLER_13_1408/li_0_527# _367_/li_155_n17# FILLER_13_1816/li_63_527#
+ user_to_mprj_in_gates\[28\]/li_707_367# user_to_mprj_in_buffers\[75\]/li_51_367#
+ ANTENNA__570__A/li_63_n17# FILLER_16_1419/li_0_527# user_to_mprj_in_gates\[33\]/li_339_527#
+ FILLER_12_1338/li_0_527# powergood_check/FILLER_0_96/li_65_797# user_to_mprj_oen_buffers\[37\]/li_795_379#
+ user_to_mprj_in_gates\[87\]/li_155_527# FILLER_3_1383/li_63_527# la_buf\[74\]/li_523_n17#
+ mprj_adr_buf\[8\]/li_63_n17# _456_/li_155_527# user_to_mprj_in_gates\[42\]/li_339_n17#
+ user_to_mprj_oen_buffers\[8\]/li_207_51# FILLER_22_1663/li_0_527# user_to_mprj_oen_buffers\[71\]/li_1351_527#
+ mprj_adr_buf\[16\]/li_215_311# FILLER_10_1284/li_63_527# user_to_mprj_in_gates\[96\]/li_155_n17#
+ user_to_mprj_in_gates\[103\]/li_339_n17# user_to_mprj_in_gates\[16\]/li_707_367#
+ FILLER_11_897/li_155_n17# powergood_check/FILLER_1_0/li_115_72# _546_/li_155_n17#
+ user_to_mprj_in_gates\[95\]/li_707_n17# la_buf\[68\]/li_207_51# mprj_adr_buf\[13\]/li_17_51#
+ user_to_mprj_oen_buffers\[25\]/li_795_379# user_to_mprj_in_buffers\[34\]/li_236_17#
+ FILLER_12_967/li_63_527# FILLER_12_617/li_155_527# _336_/li_155_527# FILLER_9_440/li_63_n17#
+ FILLER_20_449/li_63_527# powergood_check/FILLER_1_115/li_0_n17# powergood_check/FILLER_1_268/li_0_797#
+ la_buf\[70\]/li_207_51# _331_/li_247_527# FILLER_21_1985/li_63_527# user_to_mprj_in_buffers\[123\]/li_236_17#
+ mprj_dat_buf\[29\]/li_891_527# FILLER_16_44/li_0_527# powergood_check/FILLER_1_156/li_0_797#
+ user_to_mprj_in_gates\[84\]/li_155_n17# user_to_mprj_in_buffers\[2\]/li_404_17#
+ user_to_mprj_oen_buffers\[22\]/li_63_527# powergood_check/FILLER_0_224/li_115_72#
+ la_buf\[83\]/li_891_n17# user_to_mprj_in_gates\[90\]/li_18_51# user_to_mprj_in_gates\[83\]/li_707_n17#
+ user_to_mprj_in_buffers\[13\]/li_404_17# la_buf\[98\]/li_215_311# la_buf\[51\]/li_779_17#
+ mprj_adr_buf\[2\]/li_1351_n17# powergood_check/FILLER_0_112/li_115_72# powergood_check/FILLER_2_107/li_449_n17#
+ _367_/li_0_527# _657_/li_0_n17# _658_/li_0_527# FILLER_21_1695/li_155_527# FILLER_24_90/li_0_n17#
+ user_to_mprj_in_gates\[65\]/li_431_n17# la_buf\[28\]/li_247_n17# user_to_mprj_in_gates\[63\]/li_155_527#
+ mprj_dat_buf\[28\]/li_207_51# powergood_check/FILLER_2_300/li_65_n17# user_to_mprj_oen_buffers\[95\]/li_523_n17#
+ FILLER_12_839/li_0_527# FILLER_13_837/li_0_n17# FILLER_13_1067/li_155_527# FILLER_25_823/li_63_n17#
+ FILLER_13_1704/li_155_527# la_buf\[72\]/li_707_n17# user_to_mprj_in_buffers\[118\]/li_404_367#
+ FILLER_25_1051/li_155_n17# FILLER_25_974/li_63_n17# user_to_mprj_oen_buffers\[72\]/li_17_51#
+ la_buf\[51\]/li_1075_n17# FILLER_26_1282/li_155_527# FILLER_11_1351/li_155_527#
+ la_buf\[84\]/li_17_51# user_to_mprj_in_gates\[57\]/li_63_n17# user_to_mprj_in_buffers\[3\]/li_51_367#
+ mprj_dat_buf\[30\]/li_207_51# FILLER_17_1520/li_0_n17# powergood_check/FILLER_1_131/li_353_797#
+ FILLER_12_1106/li_63_n17# powergood_check/mprj2_logic_high_lv/li_929_1611# _371_/li_247_527#
+ user_to_mprj_in_buffers\[29\]/li_615_527# FILLER_17_1580/li_0_527# powergood_check/FILLER_0_224/li_65_n17#
+ mprj_dat_buf\[7\]/li_523_n17# la_buf\[86\]/li_215_311# user_to_mprj_in_gates\[120\]/li_431_527#
+ PHY_705/li_0_n17# mprj_dat_buf\[11\]/li_779_17# mprj_adr_buf\[2\]/li_983_n17# powergood_check/FILLER_1_140/li_257_n17#
+ FILLER_26_721/li_155_527# user_to_mprj_oen_buffers\[83\]/li_523_n17# FILLER_13_1017/li_155_527#
+ powergood_check/FILLER_2_32/li_737_797# powergood_check/FILLER_1_268/li_0_n17# user_to_mprj_oen_buffers\[117\]/li_247_n17#
+ powergood_check/FILLER_1_48/li_641_n17# user_to_mprj_in_gates\[58\]/li_18_51# FILLER_5_763/li_63_n17#
+ user_to_mprj_in_buffers\[106\]/li_404_367# FILLER_20_263/li_0_527# user_to_mprj_in_buffers\[103\]/li_51_367#
+ user_to_mprj_oen_buffers\[45\]/li_207_51# FILLER_5_714/li_63_527# mprj_dat_buf\[27\]/li_431_n17#
+ FILLER_16_508/li_0_527# la_buf\[29\]/li_1167_527# FILLER_23_1413/li_0_n17# powergood_check/FILLER_2_227/li_100_536#
+ FILLER_26_1191/li_155_527# PHY_300/li_0_527# user_to_mprj_oen_buffers\[21\]/li_17_51#
+ powergood_check/FILLER_1_180/li_545_n17# powergood_check/FILLER_2_251/li_257_n17#
+ user_to_mprj_in_gates\[32\]/li_431_527# FILLER_21_1573/li_155_527# la_buf\[33\]/li_17_51#
+ ANTENNA_mprj_clk_buf_TE/li_63_n17# powergood_check/FILLER_1_260/li_115_72# mprj_cyc_buf/li_1075_n17#
+ _583_/li_155_527# FILLER_26_1082/li_0_527# FILLER_6_815/li_0_527# FILLER_25_1019/li_155_n17#
+ FILLER_19_52/li_0_527# FILLER_13_777/li_0_527# user_to_mprj_in_buffers\[71\]/li_51_17#
+ la_buf\[74\]/li_215_311# powergood_check/FILLER_2_227/li_449_797# user_to_mprj_oen_buffers\[74\]/li_1075_n17#
+ user_to_mprj_in_gates\[27\]/li_523_n17# FILLER_24_2090/li_0_527# mprj_adr_buf\[2\]/li_207_51#
+ la_buf\[48\]/li_615_527# la_buf\[73\]/li_611_17# la_buf\[58\]/li_1351_527# mprj_sel_buf\[3\]/li_1535_527#
+ la_buf\[109\]/li_1535_n17# mprj_dat_buf\[29\]/li_215_311# la_buf\[79\]/li_779_17#
+ FILLER_26_203/li_63_n17# la_buf\[12\]/li_1535_n17# FILLER_7_1035/li_0_n17# powergood_check/FILLER_2_24/li_545_n17#
+ _390_/li_247_527# FILLER_25_746/li_155_n17# FILLER_20_465/li_63_527# la_buf\[28\]/li_1443_n17#
+ user_to_mprj_in_gates\[1\]/li_431_527# powergood_check/FILLER_0_248/li_100_536#
+ FILLER_5_617/li_63_527# powergood_check/FILLER_2_267/li_737_797# FILLER_25_839/li_0_n17#
+ FILLER_26_1062/li_155_527# FILLER_27_798/li_0_n17# _356_/li_0_n17# ANTENNA__368__A/li_0_n17#
+ user_to_mprj_oen_buffers\[60\]/li_63_n17# la_buf\[7\]/li_891_527# powergood_check/FILLER_2_187/li_545_797#
+ mprj_dat_buf\[18\]/li_1075_527# FILLER_5_1176/li_0_527# FILLER_12_1557/li_63_n17#
+ mprj_cyc_buf/li_215_311# mprj_sel_buf\[2\]/li_215_311# powergood_check/FILLER_0_248/li_449_797#
+ user_to_mprj_in_gates\[98\]/li_615_527# la_buf\[62\]/li_215_311# la_buf\[70\]/li_523_n17#
+ user_to_mprj_in_gates\[79\]/li_247_n17# powergood_check/FILLER_2_219/li_257_n17#
+ user_to_mprj_oen_buffers\[101\]/li_207_51# powergood_check/FILLER_0_168/li_257_797#
+ FILLER_9_884/li_0_527# mprj_dat_buf\[17\]/li_215_311# powergood_check/FILLER_1_48/li_161_797#
+ PHY_325/li_0_527# la_buf\[2\]/li_611_17# la_buf\[22\]/li_63_n17# FILLER_25_1648/li_63_n17#
+ powergood_check/FILLER_0_200/li_353_797# user_to_mprj_in_gates\[58\]/li_247_527#
+ la_buf\[75\]/li_207_51# powergood_check/FILLER_2_259/li_545_n17# mprj_dat_buf\[1\]/li_63_527#
+ user_to_mprj_in_buffers\[97\]/li_615_n17# FILLER_23_625/li_0_527# mprj_vdd_pwrgood/li_155_527#
+ user_to_mprj_in_buffers\[7\]/li_404_17# la_buf\[89\]/li_795_379# FILLER_25_1481/li_0_527#
+ user_to_mprj_oen_buffers\[63\]/li_983_n17# user_to_mprj_in_buffers\[111\]/li_51_367#
+ powergood_check/FILLER_2_179/li_353_n17# powergood_check/FILLER_2_195/li_115_72#
+ la_buf\[99\]/li_431_n17# _343_/li_155_527# user_to_mprj_in_gates\[119\]/li_247_527#
+ FILLER_9_516/li_0_n17# user_to_mprj_in_buffers\[18\]/li_404_17# la_buf\[56\]/li_779_17#
+ user_to_mprj_oen_buffers\[95\]/li_215_311# user_to_mprj_in_gates\[39\]/li_523_527#
+ powergood_check/FILLER_0_240/li_641_797# FILLER_21_1448/li_0_n17# la_buf\[50\]/li_215_311#
+ powergood_check/FILLER_1_220/li_65_n17# PHY_350/li_0_527# la_buf\[24\]/li_615_527#
+ mprj_adr_buf\[12\]/li_17_51# FILLER_12_982/li_0_n17# ANTENNA_user_to_mprj_oen_buffers\[5\]_TE/li_63_n17#
+ FILLER_25_1200/li_63_n17# _643_/li_0_527# FILLER_23_1429/li_0_n17# FILLER_21_70/li_155_n17#
+ _531_/li_0_527# ANTENNA_mprj_rstn_buf_TE/li_63_n17# FILLER_12_1697/li_63_n17# FILLER_21_1331/li_63_n17#
+ la_buf\[4\]/li_207_51# user_to_mprj_in_gates\[109\]/li_523_n17# _505_/li_247_n17#
+ FILLER_9_1282/li_63_527# user_to_mprj_in_gates\[107\]/li_247_527# user_to_mprj_in_buffers\[44\]/li_0_527#
+ FILLER_11_629/li_63_527# user_to_mprj_oen_buffers\[83\]/li_215_311# user_to_mprj_in_gates\[99\]/li_615_527#
+ user_to_mprj_in_gates\[27\]/li_523_527# FILLER_11_1572/li_0_n17# FILLER_13_1812/li_155_n17#
+ user_to_mprj_oen_buffers\[57\]/li_707_527# user_to_mprj_in_gates\[55\]/li_247_n17#
+ mprj_dat_buf\[9\]/li_17_51# user_to_mprj_oen_buffers\[92\]/li_1075_527# FILLER_13_548/li_0_527#
+ user_to_mprj_oen_buffers\[50\]/li_707_527# la_buf\[86\]/li_891_527# FILLER_17_1632/li_0_527#
+ la_buf\[122\]/li_215_311# mprj_dat_buf\[0\]/li_1351_527# FILLER_12_886/li_63_n17#
+ FILLER_9_1142/li_155_527# _627_/li_247_527# la_buf\[2\]/li_215_311# powergood_check/mprj_logic_high_hvl/li_353_797#
+ FILLER_17_1925/li_63_527# FILLER_9_1347/li_0_527# la_buf\[118\]/li_0_527# FILLER_11_1584/li_63_527#
+ powergood_check/FILLER_0_208/li_641_797# user_to_mprj_in_buffers\[21\]/li_51_367#
+ FILLER_9_697/li_0_n17# user_to_mprj_in_gates\[36\]/li_523_n17# FILLER_25_693/li_0_n17#
+ FILLER_17_249/li_0_527# ANTENNA_user_to_mprj_oen_buffers\[108\]_A/li_63_n17# PHY_863/li_0_527#
+ user_to_mprj_in_gates\[34\]/li_247_527# user_to_mprj_oen_buffers\[71\]/li_17_51#
+ mprj_stb_buf/li_63_527# user_to_mprj_in_gates\[95\]/li_523_527# mprj_sel_buf\[2\]/li_779_17#
+ FILLER_16_1601/li_63_527# user_to_mprj_oen_buffers\[88\]/li_247_n17# la_buf\[83\]/li_17_51#
+ user_to_mprj_in_buffers\[73\]/li_404_367# user_to_mprj_oen_buffers\[22\]/li_1443_n17#
+ la_buf\[57\]/li_63_527# ANTENNA__368__A/li_0_527# FILLER_13_1071/li_0_n17# FILLER_19_1417/li_0_n17#
+ user_to_mprj_oen_buffers\[29\]/li_1259_527# la_buf\[118\]/li_707_527# powergood_check/FILLER_2_267/li_65_n17#
+ _402_/li_247_527# user_to_mprj_oen_buffers\[71\]/li_215_311# user_to_mprj_oen_buffers\[52\]/li_207_51#
+ FILLER_25_891/li_63_n17# FILLER_15_554/li_63_527# user_to_mprj_in_gates\[87\]/li_615_527#
+ FILLER_10_509/li_63_n17# user_to_mprj_oen_buffers\[57\]/li_983_527# user_to_mprj_oen_buffers\[38\]/li_1351_n17#
+ mprj_adr_buf\[7\]/li_207_51# la_buf\[72\]/li_707_527# powergood_check/FILLER_2_155/li_65_n17#
+ PHY_742/li_0_n17# FILLER_5_1775/li_63_527# la_buf\[110\]/li_215_311# mprj_dat_buf\[5\]/li_983_527#
+ powergood_check/FILLER_1_115/li_100_536# FILLER_17_156/li_0_527# ANTENNA_user_to_mprj_in_gates\[32\]_B/li_63_527#
+ user_to_mprj_in_gates\[64\]/li_615_n17# FILLER_12_1035/li_63_527# FILLER_12_689/li_0_n17#
+ powergood_check/FILLER_1_16/li_545_n17# ANTENNA__365__A/li_63_n17# FILLER_12_1186/li_63_527#
+ _590_/li_155_527# user_to_mprj_in_gates\[104\]/li_247_n17# la_buf\[109\]/li_0_n17#
+ user_to_mprj_in_gates\[96\]/li_615_n17# user_to_mprj_in_gates\[57\]/li_18_51# user_to_mprj_in_gates\[94\]/li_339_527#
+ FILLER_26_1176/li_155_527# la_buf\[6\]/li_983_n17# FILLER_25_1111/li_0_n17# la_buf\[14\]/li_207_51#
+ FILLER_9_596/li_155_n17# la_buf\[53\]/li_795_379# user_to_mprj_oen_buffers\[20\]/li_17_51#
+ _480_/li_0_n17# la_buf\[21\]/li_983_527# FILLER_17_1580/li_0_n17# user_to_mprj_in_buffers\[61\]/li_404_367#
+ _577_/li_0_527# _468_/li_155_527# la_buf\[32\]/li_17_51# la_buf\[63\]/li_431_n17#
+ PHY_841/li_0_n17# la_buf\[91\]/li_63_527# mprj_dat_buf\[29\]/li_0_527# FILLER_21_2101/li_0_n17#
+ FILLER_11_2012/li_0_527# FILLER_9_582/li_63_527# la_buf\[22\]/li_1351_527# user_to_mprj_oen_buffers\[39\]/li_17_51#
+ FILLER_9_1038/li_155_527# la_buf\[63\]/li_983_527# FILLER_11_1610/li_0_n17# user_to_mprj_oen_buffers\[106\]/li_207_51#
+ PHY_319/li_0_n17# powergood_check/FILLER_1_188/li_115_72# powergood_check/FILLER_2_155/li_100_536#
+ _572_/li_247_n17# powergood_check/FILLER_1_131/li_353_n17# mprj_adr_buf\[6\]/li_891_527#
+ FILLER_15_361/li_0_n17# user_to_mprj_oen_buffers\[18\]/li_215_311# user_to_mprj_oen_buffers\[87\]/li_431_527#
+ _558_/li_155_n17# la_buf\[21\]/li_0_n17# user_to_mprj_in_gates\[77\]/li_707_367#
+ mprj_dat_buf\[21\]/li_707_527# FILLER_14_2096/li_155_n17# user_to_mprj_in_gates\[82\]/li_339_527#
+ FILLER_13_1578/li_0_n17# user_to_mprj_in_buffers\[46\]/li_236_17# FILLER_11_1351/li_155_n17#
+ powergood_check/FILLER_2_155/li_449_797# user_to_mprj_in_buffers\[92\]/li_523_n17#
+ FILLER_9_1142/li_63_527# la_buf\[41\]/li_795_379# _346_/li_0_n17# powergood_check/FILLER_2_32/li_737_n17#
+ powergood_check/FILLER_1_107/li_257_n17# FILLER_18_1463/li_0_n17# user_to_mprj_oen_buffers\[119\]/li_63_n17#
+ _560_/li_155_n17# la_buf\[51\]/li_431_n17# la_buf\[28\]/li_707_n17# FILLER_21_66/li_0_527#
+ user_to_mprj_in_gates\[91\]/li_339_n17# FILLER_17_1428/li_0_527# la_buf\[82\]/li_207_51#
+ powergood_check/FILLER_0_176/li_100_536# powergood_check/FILLER_2_203/li_0_797#
+ powergood_check/FILLER_2_219/li_115_72# user_to_mprj_in_buffers\[7\]/li_155_n17#
+ FILLER_18_1529/li_63_527# PHY_339/li_0_527# FILLER_14_1500/li_63_n17# FILLER_13_659/li_0_527#
+ FILLER_5_747/li_0_527# PHY_330/li_0_n17# powergood_check/FILLER_2_107/li_115_72#
+ FILLER_9_596/li_0_n17# la_buf\[51\]/li_1535_n17# ANTENNA__341__A/li_63_n17# la_buf\[30\]/li_431_527#
+ _350_/li_155_527# user_to_mprj_in_buffers\[25\]/li_404_17# user_to_mprj_in_gates\[72\]/li_431_527#
+ mprj_cyc_buf/li_1351_n17# powergood_check/FILLER_1_164/li_0_n17# powergood_check/FILLER_2_227/li_449_n17#
+ FILLER_27_873/li_63_n17# FILLER_18_504/li_63_527# user_to_mprj_in_buffers\[38\]/li_51_17#
+ user_to_mprj_oen_buffers\[126\]/li_1167_527# powergood_check/FILLER_0_176/li_449_797#
+ mprj_dat_buf\[4\]/li_0_527# PHY_294/li_0_527# la_buf\[9\]/li_207_51# la_buf\[89\]/li_247_n17#
+ FILLER_12_1673/li_0_n17# FILLER_19_604/li_0_527# _527_/li_155_527# powergood_check/FILLER_2_267/li_737_n17#
+ ANTENNA__382__A/li_0_n17# powergood_check/FILLER_0_24/li_0_797# la_buf\[123\]/li_431_n17#
+ user_to_mprj_oen_buffers\[117\]/li_707_n17# mprj_adr_buf\[11\]/li_17_51# user_to_mprj_in_gates\[69\]/li_63_n17#
+ powergood_check/FILLER_2_187/li_545_n17# powergood_check/mprj_logic_high_hvl/li_43_635#
+ ANTENNA_user_to_mprj_in_gates\[53\]_B/li_63_n17# user_to_mprj_in_gates\[122\]/li_63_n17#
+ mprj_adr_buf\[27\]/li_615_527# FILLER_23_56/li_63_n17# powergood_check/FILLER_0_0/li_545_797#
+ user_to_mprj_oen_buffers\[5\]/li_247_527# FILLER_20_2087/li_0_527# FILLER_22_1982/li_63_527#
+ user_to_mprj_oen_buffers\[21\]/li_891_527# la_buf\[102\]/li_431_527# powergood_check/FILLER_1_236/li_100_536#
+ FILLER_13_1207/li_155_n17# powergood_check/FILLER_2_32/li_257_797# FILLER_9_586/li_0_527#
+ _657_/li_247_527# powergood_check/FILLER_1_48/li_161_n17# user_to_mprj_in_gates\[71\]/li_63_n17#
+ mprj_dat_buf\[30\]/li_983_527# user_to_mprj_in_gates\[109\]/li_18_51# FILLER_25_1922/li_155_n17#
+ user_to_mprj_oen_buffers\[4\]/li_63_527# user_to_mprj_in_gates\[114\]/li_707_367#
+ la_buf\[97\]/li_1535_n17# powergood_check/FILLER_0_232/li_0_797# user_to_mprj_oen_buffers\[74\]/li_1535_n17#
+ FILLER_12_693/li_63_n17# user_to_mprj_in_gates\[31\]/li_155_n17# mprj_adr_buf\[6\]/li_215_311#
+ user_to_mprj_oen_buffers\[72\]/li_431_n17# ANTENNA__554__A/li_63_n17# user_to_mprj_in_gates\[3\]/li_431_527#
+ FILLER_17_1405/li_0_n17# FILLER_11_436/li_0_527# _407_/li_155_527# user_to_mprj_oen_buffers\[57\]/li_207_51#
+ FILLER_14_491/li_0_527# FILLER_21_1451/li_155_527# FILLER_12_581/li_63_n17# FILLER_7_1035/li_0_527#
+ la_buf\[44\]/li_983_n17# FILLER_11_1472/li_0_n17# mprj_dat_buf\[8\]/li_17_51# _347_/li_0_527#
+ powergood_check/FILLER_2_115/li_641_797# FILLER_26_1555/li_0_527# la_buf\[56\]/li_247_527#
+ FILLER_12_1069/li_155_527# user_to_mprj_oen_buffers\[38\]/li_779_17# mprj_adr_buf\[15\]/li_615_527#
+ FILLER_20_1459/li_0_527# FILLER_18_1994/li_63_n17# user_to_mprj_in_gates\[5\]/li_339_527#
+ _386_/li_0_527# mprj_dat_buf\[18\]/li_1535_527# user_to_mprj_oen_buffers\[7\]/li_891_527#
+ la_buf\[19\]/li_207_51# powergood_check/mprj2_logic_high_hvl/li_161_797# user_to_mprj_oen_buffers\[70\]/li_17_51#
+ user_to_mprj_oen_buffers\[50\]/li_795_379# user_to_mprj_oen_buffers\[96\]/li_1351_527#
+ FILLER_12_1462/li_63_527# la_buf\[82\]/li_17_51# powergood_check/FILLER_2_267/li_257_797#
+ _386_/li_155_n17# PHY_458/li_0_527# user_to_mprj_in_gates\[79\]/li_707_n17# user_to_mprj_oen_buffers\[40\]/li_779_17#
+ FILLER_5_714/li_155_527# FILLER_7_1031/li_155_527# user_to_mprj_oen_buffers\[60\]/li_431_n17#
+ _660_/li_247_527# FILLER_25_730/li_63_n17# mprj_dat_buf\[16\]/li_1351_n17# powergood_check/FILLER_0_80/li_353_797#
+ mprj_dat_buf\[6\]/li_1351_527# user_to_mprj_oen_buffers\[89\]/li_17_51# user_to_mprj_in_buffers\[90\]/li_339_527#
+ powergood_check/mprj2_logic_high_lv/li_161_1611# FILLER_26_856/li_63_527# la_buf\[21\]/li_207_51#
+ powergood_check/FILLER_1_228/li_257_n17# user_to_mprj_oen_buffers\[72\]/li_63_n17#
+ user_to_mprj_in_gates\[81\]/li_431_527# la_buf\[44\]/li_247_527# ANTENNA__487__A/li_63_527#
+ FILLER_17_543/li_0_n17# powergood_check/FILLER_0_232/li_65_797# FILLER_19_1581/li_0_n17#
+ _430_/li_247_527# user_to_mprj_in_gates\[56\]/li_18_51# PHY_477/li_0_527# powergood_check/FILLER_1_268/li_545_n17#
+ FILLER_23_1774/li_155_527# user_to_mprj_oen_buffers\[113\]/li_207_51# powergood_check/mprj_logic_high_hvl/li_353_n17#
+ powergood_check/FILLER_2_195/li_0_797# FILLER_25_709/li_0_n17# la_buf\[67\]/li_891_n17#
+ _565_/li_155_n17# la_buf\[31\]/li_17_51# powergood_check/FILLER_0_192/li_0_n17#
+ la_buf\[123\]/li_0_527# powergood_check/FILLER_1_62/li_65_797# powergood_check/mprj_logic_high_hvl/li_307_57#
+ la_buf\[87\]/li_207_51# FILLER_25_815/li_155_n17# FILLER_1_929/li_63_527# user_to_mprj_in_buffers\[9\]/li_615_527#
+ user_to_mprj_in_buffers\[53\]/li_236_17# user_to_mprj_oen_buffers\[38\]/li_17_51#
+ user_to_mprj_oen_buffers\[110\]/li_983_n17# FILLER_22_1909/li_63_n17# FILLER_11_1709/li_63_n17#
+ FILLER_17_1512/li_155_527# _477_/li_247_527# FILLER_21_1985/li_0_n17# ANTENNA_user_to_mprj_in_gates\[71\]_B/li_63_527#
+ powergood_check/FILLER_0_240/li_161_797# ANTENNA_user_to_mprj_in_gates\[46\]_B/li_63_n17#
+ FILLER_14_1784/li_63_527# _654_/li_155_527# user_to_mprj_in_buffers\[29\]/li_236_367#
+ FILLER_24_512/li_0_527# FILLER_26_920/li_0_527# FILLER_21_1448/li_0_527# FILLER_26_995/li_0_527#
+ user_to_mprj_in_gates\[80\]/li_615_n17# user_to_mprj_oen_buffers\[14\]/li_1351_527#
+ FILLER_20_547/li_0_527# user_to_mprj_oen_buffers\[86\]/li_247_n17# user_to_mprj_oen_buffers\[42\]/li_0_527#
+ FILLER_5_1031/li_63_527# mprj_sel_buf\[3\]/li_431_527# _336_/li_0_n17# la_buf\[42\]/li_983_n17#
+ user_to_mprj_in_gates\[55\]/li_707_n17# FILLER_23_1520/li_63_n17# user_to_mprj_oen_buffers\[50\]/li_1167_527#
+ powergood_check/FILLER_0_88/li_641_797# la_buf\[70\]/li_779_17# FILLER_19_1451/li_155_n17#
+ FILLER_21_1947/li_63_527# FILLER_13_837/li_63_527# user_to_mprj_oen_buffers\[62\]/li_611_17#
+ FILLER_20_75/li_63_527# _375_/li_0_n17# FILLER_24_2040/li_155_527# powergood_check/FILLER_1_115/li_449_n17#
+ user_to_mprj_oen_buffers\[7\]/li_215_311# user_to_mprj_in_gates\[38\]/li_523_527#
+ user_to_mprj_in_gates\[116\]/li_707_n17# la_buf\[0\]/li_523_n17# FILLER_17_62/li_63_n17#
+ user_to_mprj_oen_buffers\[65\]/li_247_527# user_to_mprj_in_gates\[127\]/li_63_n17#
+ la_buf\[20\]/li_247_527# FILLER_9_563/li_63_527# mprj_stb_buf/li_247_n17# _534_/li_155_527#
+ FILLER_25_1241/li_155_n17# FILLER_26_986/li_0_527# user_to_mprj_in_gates\[88\]/li_523_527#
+ FILLER_22_294/li_0_527# user_to_mprj_in_gates\[16\]/li_431_527# la_buf\[50\]/li_1167_n17#
+ FILLER_27_802/li_63_n17# la_buf\[24\]/li_611_17# user_to_mprj_oen_buffers\[89\]/li_1351_527#
+ user_to_mprj_oen_buffers\[74\]/li_247_n17# FILLER_12_697/li_155_527# user_to_mprj_oen_buffers\[14\]/li_1259_n17#
+ powergood_check/FILLER_0_208/li_161_797# user_to_mprj_oen_buffers\[88\]/li_891_n17#
+ la_buf\[58\]/li_215_311# mprj_we_buf/li_207_51# FILLER_19_1577/li_0_n17# user_to_mprj_in_gates\[105\]/li_155_n17#
+ FILLER_13_1017/li_0_n17# user_to_mprj_in_gates\[25\]/li_431_n17# powergood_check/FILLER_2_155/li_449_n17#
+ FILLER_23_621/li_63_527# la_buf\[18\]/li_63_527# FILLER_27_877/li_0_n17# FILLER_13_850/li_155_527#
+ la_buf\[5\]/li_1443_n17# mprj_adr_buf\[10\]/li_17_51# user_to_mprj_in_gates\[125\]/li_615_527#
+ _337_/li_247_527# FILLER_13_2020/li_155_527# FILLER_28_1735/li_0_n17# powergood_check/FILLER_0_8/li_115_72#
+ user_to_mprj_oen_buffers\[64\]/li_207_51# powergood_check/FILLER_0_80/li_0_797#
+ powergood_check/FILLER_2_203/li_0_n17# FILLER_11_838/li_155_n17# FILLER_13_1203/li_63_527#
+ user_to_mprj_in_gates\[76\]/li_523_527# mprj_adr_buf\[29\]/li_17_51# PHY_334/li_0_n17#
+ user_to_mprj_oen_buffers\[62\]/li_247_n17# FILLER_26_819/li_155_527# user_to_mprj_oen_buffers\[45\]/li_779_17#
+ user_to_mprj_in_gates\[108\]/li_18_51# user_to_mprj_oen_buffers\[91\]/li_891_n17#
+ mprj_dat_buf\[7\]/li_63_n17# PHY_276/li_0_n17# FILLER_25_1269/li_63_n17# la_buf\[31\]/li_891_n17#
+ la_buf\[46\]/li_215_311# FILLER_12_1927/li_155_n17# FILLER_9_348/li_63_n17# mprj_dat_buf\[25\]/li_0_527#
+ FILLER_12_1927/li_0_n17# FILLER_26_1057/li_0_527# user_to_mprj_oen_buffers\[95\]/li_1351_527#
+ user_to_mprj_in_gates\[81\]/li_0_n17# FILLER_12_772/li_155_527# la_buf\[26\]/li_207_51#
+ la_buf\[92\]/li_611_17# FILLER_14_2092/li_155_n17# mprj_dat_buf\[7\]/li_17_51# powergood_check/FILLER_1_164/li_100_536#
+ user_to_mprj_in_buffers\[104\]/li_51_17# _393_/li_155_n17# la_buf\[6\]/li_1075_527#
+ ANTENNA_user_to_mprj_in_gates\[64\]_B/li_63_527# ANTENNA_la_buf\[7\]_TE/li_63_527#
+ mprj_dat_buf\[29\]/li_63_527# FILLER_8_1020/li_0_527# powergood_check/FILLER_1_24/li_115_72#
+ user_to_mprj_in_gates\[64\]/li_523_527# powergood_check/FILLER_0_272/li_115_72#
+ FILLER_23_1915/li_155_527# user_to_mprj_oen_buffers\[118\]/li_207_51# user_to_mprj_in_gates\[92\]/li_247_n17#
+ mprj_cyc_buf/li_0_527# la_buf\[82\]/li_1535_n17# FILLER_25_1337/li_0_527# FILLER_23_1425/li_0_n17#
+ powergood_check/FILLER_0_160/li_115_72# powergood_check/mprj2_logic_high_lv/li_179_1349#
+ ANTENNA__345__A/li_0_n17# mprj_dat_buf\[30\]/li_215_311# la_buf\[81\]/li_17_51#
+ user_to_mprj_oen_buffers\[79\]/li_215_311# la_buf\[87\]/li_0_n17# ANTENNA_user_to_mprj_in_gates\[110\]_A/li_63_527#
+ ANTENNA_user_to_mprj_in_gates\[82\]_A/li_63_527# user_to_mprj_in_buffers\[7\]/li_615_n17#
+ ANTENNA_user_to_mprj_in_gates\[57\]_A/li_63_n17# la_buf\[34\]/li_215_311# powergood_check/FILLER_0_104/li_545_797#
+ la_buf\[84\]/li_707_n17# powergood_check/FILLER_2_32/li_257_n17# user_to_mprj_in_gates\[73\]/li_523_n17#
+ la_buf\[118\]/li_215_311# user_to_mprj_oen_buffers\[88\]/li_17_51# la_buf\[0\]/li_63_527#
+ user_to_mprj_in_gates\[71\]/li_247_527# user_to_mprj_oen_buffers\[120\]/li_207_51#
+ FILLER_13_1704/li_63_527# FILLER_19_2000/li_155_527# user_to_mprj_oen_buffers\[43\]/li_891_527#
+ FILLER_14_359/li_63_527# la_buf\[70\]/li_983_527# FILLER_22_515/li_0_n17# _659_/li_155_527#
+ mprj_dat_buf\[6\]/li_215_311# la_buf\[86\]/li_1443_527# la_buf\[24\]/li_1443_n17#
+ powergood_check/FILLER_2_195/li_257_797# _658_/li_0_n17# la_buf\[89\]/li_707_n17#
+ FILLER_13_428/li_63_n17# powergood_check/FILLER_0_240/li_65_n17# la_buf\[94\]/li_207_51#
+ FILLER_7_1035/li_63_527# user_to_mprj_in_gates\[55\]/li_18_51# user_to_mprj_in_gates\[52\]/li_523_527#
+ powergood_check/FILLER_2_115/li_641_n17# la_buf\[29\]/li_983_527# user_to_mprj_in_gates\[80\]/li_247_n17#
+ FILLER_13_1672/li_0_n17# FILLER_11_2009/li_63_527# user_to_mprj_oen_buffers\[60\]/li_1259_n17#
+ powergood_check/FILLER_1_156/li_257_n17# user_to_mprj_oen_buffers\[67\]/li_215_311#
+ la_buf\[98\]/li_983_527# la_buf\[22\]/li_215_311# la_buf\[30\]/li_17_51# user_to_mprj_oen_buffers\[91\]/li_1167_n17#
+ powergood_check/mprj2_logic_high_hvl/li_161_n17# la_buf\[106\]/li_215_311# user_to_mprj_oen_buffers\[123\]/li_215_311#
+ FILLER_12_664/li_0_n17# user_to_mprj_oen_buffers\[37\]/li_17_51# powergood_check/FILLER_2_267/li_257_n17#
+ powergood_check/FILLER_1_196/li_545_n17# FILLER_14_359/li_0_n17# la_buf\[49\]/li_17_51#
+ FILLER_17_1909/li_63_527# FILLER_25_1291/li_155_n17# powergood_check/FILLER_0_16/li_257_797#
+ _651_/li_0_n17# user_to_mprj_in_gates\[122\]/li_523_n17# user_to_mprj_in_buffers\[2\]/li_339_n17#
+ FILLER_16_1421/li_63_n17# powergood_check/FILLER_2_8/li_0_797# mprj_dat_buf\[13\]/li_1351_n17#
+ la_buf\[29\]/li_611_17# la_buf\[121\]/li_1535_n17# powergood_check/FILLER_1_8/li_100_536#
+ FILLER_16_1644/li_63_527# _589_/li_0_n17# la_buf\[59\]/li_431_n17# user_to_mprj_oen_buffers\[40\]/li_891_n17#
+ user_to_mprj_oen_buffers\[55\]/li_215_311# FILLER_3_759/li_0_527# la_buf\[10\]/li_215_311#
+ la_buf\[6\]/li_63_527# user_to_mprj_oen_buffers\[29\]/li_615_527# ANTENNA__644__A/li_0_n17#
+ user_to_mprj_in_gates\[27\]/li_247_n17# FILLER_0_201/li_63_527# la_buf\[56\]/li_707_527#
+ FILLER_9_966/li_155_527# user_to_mprj_oen_buffers\[111\]/li_215_311# la_buf\[4\]/li_779_17#
+ powergood_check/FILLER_2_195/li_0_n17# FILLER_11_1553/li_63_n17# user_to_mprj_in_gates\[83\]/li_63_n17#
+ user_to_mprj_oen_buffers\[16\]/li_63_n17# ANTENNA__349__A/li_63_n17# ANTENNA_user_to_mprj_oen_buffers\[4\]_A/li_63_n17#
+ FILLER_11_451/li_155_n17# user_to_mprj_oen_buffers\[91\]/li_983_527# user_to_mprj_oen_buffers\[69\]/li_207_51#
+ FILLER_11_1441/li_63_n17# powergood_check/FILLER_1_32/li_100_536# powergood_check/FILLER_1_62/li_65_n17#
+ FILLER_20_547/li_63_527# FILLER_19_245/li_63_n17# powergood_check/FILLER_2_115/li_161_797#
+ FILLER_14_491/li_0_n17# FILLER_13_1931/li_155_n17# FILLER_17_1584/li_0_n17# user_to_mprj_oen_buffers\[53\]/li_1351_527#
+ user_to_mprj_oen_buffers\[28\]/li_1351_n17# mprj_dat_buf\[1\]/li_207_51# powergood_check/FILLER_2_235/li_641_797#
+ FILLER_11_1544/li_0_527# user_to_mprj_in_buffers\[45\]/li_404_367# PHY_218/li_0_527#
+ FILLER_10_621/li_0_527# user_to_mprj_oen_buffers\[43\]/li_215_311# FILLER_12_978/li_155_527#
+ user_to_mprj_oen_buffers\[71\]/li_207_51# FILLER_13_1627/li_0_n17# la_buf\[44\]/li_707_527#
+ FILLER_17_1921/li_63_n17# FILLER_17_1935/li_63_527# FILLER_11_1813/li_63_n17# user_to_mprj_oen_buffers\[59\]/li_983_n17#
+ powergood_check/FILLER_0_216/li_353_797# la_buf\[2\]/li_1535_n17# FILLER_14_2096/li_63_527#
+ PHY_3/li_0_527# mprj_clk2_buf/li_207_51# user_to_mprj_oen_buffers\[52\]/li_779_17#
+ la_buf\[26\]/li_431_527# FILLER_24_512/li_155_n17# mprj_adr_buf\[7\]/li_779_17#
+ la_buf\[67\]/li_707_527# mprj_adr_buf\[29\]/li_1075_527# FILLER_9_512/li_63_n17#
+ FILLER_4_895/li_63_527# mprj_dat_buf\[7\]/li_1443_527# powergood_check/FILLER_0_256/li_641_797#
+ user_to_mprj_in_gates\[0\]/li_247_527# la_buf\[33\]/li_207_51# user_to_mprj_in_buffers\[76\]/li_523_n17#
+ la_buf\[86\]/li_1351_n17# mprj_adr_buf\[28\]/li_17_51# powergood_check/FILLER_0_8/li_353_797#
+ user_to_mprj_in_buffers\[33\]/li_404_367# la_buf\[109\]/li_795_379# la_buf\[35\]/li_431_n17#
+ user_to_mprj_oen_buffers\[56\]/li_1167_n17# _352_/li_0_n17# _487_/li_155_527# user_to_mprj_oen_buffers\[31\]/li_215_311#
+ user_to_mprj_in_gates\[107\]/li_18_51# FILLER_12_673/li_63_n17# powergood_check/FILLER_1_24/li_257_n17#
+ powergood_check/FILLER_2_115/li_65_797# la_buf\[14\]/li_779_17# user_to_mprj_in_gates\[90\]/li_707_367#
+ la_buf\[5\]/li_63_527# _439_/li_0_527# user_to_mprj_oen_buffers\[125\]/li_207_51#
+ _335_/li_247_n17# powergood_check/FILLER_1_300/li_161_n17# mprj_dat_buf\[6\]/li_17_51#
+ FILLER_13_756/li_155_527# FILLER_25_1035/li_63_n17# mprj_dat_buf\[7\]/li_431_n17#
+ la_buf\[14\]/li_431_527# _577_/li_155_n17# user_to_mprj_in_gates\[49\]/li_707_367#
+ FILLER_10_467/li_0_n17# FILLER_21_2105/li_155_n17# _478_/li_0_527# user_to_mprj_in_gates\[56\]/li_615_n17#
+ la_buf\[76\]/li_1535_n17# powergood_check/FILLER_2_0/li_65_797# la_buf\[99\]/li_207_51#
+ user_to_mprj_in_gates\[54\]/li_339_527# user_to_mprj_oen_buffers\[86\]/li_707_n17#
+ user_to_mprj_oen_buffers\[106\]/li_779_17# la_buf\[41\]/li_707_n17# _584_/li_247_527#
+ FILLER_25_934/li_63_n17# user_to_mprj_in_buffers\[21\]/li_404_367# FILLER_22_1722/li_0_527#
+ _356_/li_0_527# user_to_mprj_oen_buffers\[114\]/li_795_379# FILLER_19_1335/li_0_527#
+ la_buf\[4\]/li_891_527# powergood_check/FILLER_0_80/li_0_n17# FILLER_11_1817/li_0_527#
+ la_buf\[80\]/li_17_51# mprj_dat_buf\[1\]/li_983_527# user_to_mprj_oen_buffers\[124\]/li_431_n17#
+ mprj_adr_buf\[22\]/li_891_n17# _551_/li_0_527# mprj_stb_buf/li_707_n17# user_to_mprj_oen_buffers\[87\]/li_17_51#
+ powergood_check/FILLER_0_88/li_161_797# user_to_mprj_in_gates\[36\]/li_0_n17# user_to_mprj_oen_buffers\[47\]/li_431_527#
+
XFILLER_27_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_501_ la_data_out_mprj[30] vssd vssd vccd vccd _501_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_432_ mprj_adr_o_core[25] vssd vssd vccd vccd _432_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_363_ la_oen_mprj[95] vssd vssd vccd vccd _363_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[36\] _507_/Y la_buf\[36\]/TE vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_9_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] mprj_logic_high_inst/HI[355] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[25\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_9_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[76\] _344_/Y mprj_logic_high_inst/HI[278] vssd vssd vccd
+ vccd la_oen_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_8_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[24\] _463_/Y mprj_dat_buf\[24\]/TE vssd vssd vccd vccd mprj_dat_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high_inst/HI[306] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_415_ mprj_adr_o_core[8] vssd vssd vccd vccd _415_/Y sky130_fd_sc_hd__inv_2
X_346_ la_oen_mprj[78] vssd vssd vccd vccd _346_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high_inst/HI[329] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[41\]_TE la_buf\[41\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[26\]_TE mprj_logic_high_inst/HI[228] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] mprj_logic_high_inst/HI[422] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[92\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[64\]_TE la_buf\[64\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high_inst/HI[251] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[109\] _377_/Y mprj_logic_high_inst/HI[311] vssd vssd vccd
+ vccd la_oen_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_28_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[39\] _638_/Y mprj_logic_high_inst/HI[241] vssd vssd vccd
+ vccd la_oen_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_18_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[13\]_TE mprj_dat_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__402__A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y vssd vssd vccd vccd la_data_in_mprj[62]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[87\]_TE la_buf\[87\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_594_ la_data_out_mprj[123] vssd vssd vccd vccd _594_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[66\] _537_/Y la_buf\[66\]/TE vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__einvp_8
XPHY_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[122\] _593_/Y la_buf\[122\]/TE vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[70\]_B mprj_logic_high_inst/HI[400] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] mprj_logic_high_inst/HI[385] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[55\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[61\]_B mprj_logic_high_inst/HI[391] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[52\]_B mprj_logic_high_inst/HI[382] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_646_ la_oen_mprj[47] vssd vssd vccd vccd _646_/Y sky130_fd_sc_hd__inv_2
X_577_ la_data_out_mprj[106] vssd vssd vccd vccd _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[6\]_A _445_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y vssd vssd vccd vccd la_data_in_mprj[25]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[43\]_B mprj_logic_high_inst/HI[373] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[112\]_TE la_buf\[112\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[27\]_TE mprj_adr_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_178 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[34\]_B mprj_logic_high_inst/HI[364] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[95\]_A user_to_mprj_in_gates\[95\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__500__A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_500_ la_data_out_mprj[29] vssd vssd vccd vccd _500_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[3\] _602_/Y mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd la_oen_core[3] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[21\] _620_/Y mprj_logic_high_inst/HI[223] vssd vssd vccd
+ vccd la_oen_core[21] sky130_fd_sc_hd__einvp_8
X_431_ mprj_adr_o_core[24] vssd vssd vccd vccd _431_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_362_ la_oen_mprj[94] vssd vssd vccd vccd _362_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[29\] _500_/Y la_buf\[29\]/TE vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_13_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[122\]_A _593_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[25\]_B mprj_logic_high_inst/HI[355] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[86\]_A user_to_mprj_in_gates\[86\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__410__A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_629_ la_oen_mprj[30] vssd vssd vccd vccd _629_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[10\]_A user_to_mprj_in_gates\[10\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[124\]_A user_to_mprj_in_gates\[124\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] mprj_logic_high_inst/HI[348] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[18\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[113\]_A _584_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[77\]_A user_to_mprj_in_gates\[77\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[16\]_B mprj_logic_high_inst/HI[346] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_B mprj_logic_high_inst/HI[430] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[50\]_A _521_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high_inst/HI[284] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[115\]_A user_to_mprj_in_gates\[115\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[104\]_A _575_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[68\]_A user_to_mprj_in_gates\[68\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[41\]_A _512_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[69\] _337_/Y mprj_logic_high_inst/HI[271] vssd vssd vccd
+ vccd la_oen_core[69] sky130_fd_sc_hd__einvp_8
XFILLER_4_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[17\] _456_/Y mprj_dat_buf\[17\]/TE vssd vssd vccd vccd mprj_dat_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_414_ mprj_adr_o_core[7] vssd vssd vccd vccd _414_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[106\]_A user_to_mprj_in_gates\[106\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_345_ la_oen_mprj[77] vssd vssd vccd vccd _345_/Y sky130_fd_sc_hd__inv_2
XANTENNA__405__A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[59\]_A user_to_mprj_in_gates\[59\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[32\]_A _503_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[12\] _419_/Y mprj_adr_buf\[12\]/TE vssd vssd vccd vccd mprj_adr_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[126] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y vssd vssd vccd vccd la_data_in_mprj[92]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[99\]_A _570_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[23\]_A _494_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[14\]_A _485_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[96\] _567_/Y la_buf\[96\]/TE vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__einvp_8
XFILLER_19_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_58 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] mprj_logic_high_inst/HI[415] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[85\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[92\]_A _360_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[83\]_A _351_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[7\] _478_/Y la_buf\[7\]/TE vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__einvp_8
XFILLER_4_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[11\] _482_/Y la_buf\[11\]/TE vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__einvp_8
XFILLER_26_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[4\] _411_/Y mprj_adr_buf\[4\]/TE vssd vssd vccd vccd mprj_adr_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y vssd vssd vccd vccd la_data_in_mprj[55]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high_inst/HI[319] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[74\]_A _342_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] mprj_logic_high_inst/HI[441] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[111\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[31\]_TE la_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high_inst/HI[218] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[65\]_A _333_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__503__A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[121\] _389_/Y mprj_logic_high_inst/HI[323] vssd vssd vccd
+ vccd la_oen_core[121] sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[2\] _405_/Y mprj_sel_buf\[2\]/TE vssd vssd vccd vccd mprj_sel_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[51\] _650_/Y mprj_logic_high_inst/HI[253] vssd vssd vccd
+ vccd la_oen_core[51] sky130_fd_sc_hd__einvp_8
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_593_ la_data_out_mprj[122] vssd vssd vccd vccd _593_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[59\] _530_/Y la_buf\[59\]/TE vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__einvp_8
XPHY_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[56\]_A _655_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__413__A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[115\] _586_/Y la_buf\[115\]/TE vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_3_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[54\]_TE la_buf\[54\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[39\]_TE mprj_logic_high_inst/HI[241] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] mprj_logic_high_inst/HI[378] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[48\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[47\]_A _646_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[38\]_A _637_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[99\] _367_/Y mprj_logic_high_inst/HI[301] vssd vssd vccd
+ vccd la_oen_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_11_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_vdd_pwrgood mprj2_vdd_pwrgood/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_1_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[77\]_TE la_buf\[77\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_645_ la_oen_mprj[46] vssd vssd vccd vccd _645_/Y sky130_fd_sc_hd__inv_2
X_576_ la_data_out_mprj[105] vssd vssd vccd vccd _576_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__408__A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[29\]_A _628_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y vssd vssd vccd vccd la_data_in_mprj[18]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_adr_buf\[25\]_A _432_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[26\]_TE mprj_dat_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[5\]_TE mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[2\]_A _601_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_A _423_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_430_ mprj_adr_o_core[23] vssd vssd vccd vccd _430_/Y sky130_fd_sc_hd__inv_2
X_361_ la_oen_mprj[93] vssd vssd vccd vccd _361_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[14\] _613_/Y mprj_logic_high_inst/HI[216] vssd vssd vccd
+ vccd la_oen_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_10_820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_628_ la_oen_mprj[29] vssd vssd vccd vccd _628_/Y sky130_fd_sc_hd__inv_2
X_559_ la_data_out_mprj[88] vssd vssd vccd vccd _559_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__601__A la_oen_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__511__A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_413_ mprj_adr_o_core[6] vssd vssd vccd vccd _413_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[102\]_TE la_buf\[102\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[41\] _512_/Y la_buf\[41\]/TE vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__einvp_8
X_344_ la_oen_mprj[76] vssd vssd vccd vccd _344_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_adr_buf\[17\]_TE mprj_adr_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__421__A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[119] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[29\]_A _468_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y vssd vssd vccd vccd la_data_in_mprj[85]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] mprj_logic_high_inst/HI[360] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[30\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_24_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[1\]_A _408_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__331__A la_oen_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[5\]_TE mprj_dat_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_TE la_buf\[125\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__506__A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[81\] _349_/Y mprj_logic_high_inst/HI[283] vssd vssd vccd
+ vccd la_oen_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_2_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[89\] _560_/Y la_buf\[89\]/TE vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[72\]_TE mprj_logic_high_inst/HI[274] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__416__A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] mprj_logic_high_inst/HI[408] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[78\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj2_pwrgood_A mprj2_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high_inst/HI[297] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[7\]_A _478_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y vssd vssd vccd vccd la_data_in_mprj[48]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] mprj_logic_high_inst/HI[434] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[104\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[1\]_B user_to_mprj_in_gates\[1\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[114\] _382_/Y mprj_logic_high_inst/HI[316] vssd vssd vccd
+ vccd la_oen_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_5_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[44\] _643_/Y mprj_logic_high_inst/HI[246] vssd vssd vccd
+ vccd la_oen_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_5_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_592_ la_data_out_mprj[121] vssd vssd vccd vccd _592_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[108\] _579_/Y la_buf\[108\]/TE vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[101] sky130_fd_sc_hd__inv_8
XFILLER_19_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[5\]_A user_to_mprj_in_gates\[5\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__604__A la_oen_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[0\] _439_/Y mprj_dat_buf\[0\]/TE vssd vssd vccd vccd mprj_dat_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_26_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__514__A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[107\]_TE mprj_logic_high_inst/HI[309] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_644_ la_oen_mprj[45] vssd vssd vccd vccd _644_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[71\] _542_/Y la_buf\[71\]/TE vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__einvp_8
X_575_ la_data_out_mprj[104] vssd vssd vccd vccd _575_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__424__A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_12_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[21\]_TE la_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] mprj_logic_high_inst/HI[390] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[60\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__334__A la_oen_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__509__A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_360_ la_oen_mprj[92] vssd vssd vccd vccd _360_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[44\]_TE la_buf\[44\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high_inst/HI[231] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__419__A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_627_ la_oen_mprj[28] vssd vssd vccd vccd _627_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_558_ la_data_out_mprj[87] vssd vssd vccd vccd _558_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_489_ la_data_out_mprj[18] vssd vssd vccd vccd _489_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y vssd vssd vccd vccd la_data_in_mprj[30]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[67\]_TE la_buf\[67\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_412_ mprj_adr_o_core[5] vssd vssd vccd vccd _412_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_343_ la_oen_mprj[75] vssd vssd vccd vccd _343_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[34\] _505_/Y la_buf\[34\]/TE vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__einvp_8
XFILLER_10_662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y vssd vssd vccd vccd la_data_in_mprj[78]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] mprj_logic_high_inst/HI[353] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[23\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__612__A la_oen_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__522__A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[74\] _342_/Y mprj_logic_high_inst/HI[276] vssd vssd vccd
+ vccd la_oen_core[74] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[22\] _461_/Y mprj_dat_buf\[22\]/TE vssd vssd vccd vccd mprj_dat_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__432__A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__607__A la_oen_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[91\]_B mprj_logic_high_inst/HI[421] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__342__A la_oen_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__517__A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_B mprj_logic_high_inst/HI[412] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__427__A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_B mprj_logic_high_inst/HI[403] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[115\]_TE la_buf\[115\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] mprj_logic_high_inst/HI[420] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[90\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__337__A la_oen_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_B mprj_logic_high_inst/HI[394] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[62\]_TE mprj_logic_high_inst/HI[264] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[107\] _375_/Y mprj_logic_high_inst/HI[309] vssd vssd vccd
+ vccd la_oen_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_5_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_660_ la_oen_mprj[61] vssd vssd vccd vccd _660_/Y sky130_fd_sc_hd__inv_2
X_591_ la_data_out_mprj[120] vssd vssd vccd vccd _591_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[37\] _636_/Y mprj_logic_high_inst/HI[239] vssd vssd vccd
+ vccd la_oen_core[37] sky130_fd_sc_hd__einvp_8
XFILLER_16_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[55\]_B mprj_logic_high_inst/HI[385] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[40\]_A user_to_mprj_in_gates\[40\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y vssd vssd vccd vccd la_data_in_mprj[60]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[9\]_A _448_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[46\]_B mprj_logic_high_inst/HI[376] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_A _551_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high_inst/HI[287] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__620__A la_oen_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[31\]_A user_to_mprj_in_gates\[31\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[98\]_A user_to_mprj_in_gates\[98\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_B mprj_logic_high_inst/HI[367] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_B mprj_logic_high_inst/HI[451] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_A _542_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__530__A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_643_ la_oen_mprj[44] vssd vssd vccd vccd _643_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[22\]_A user_to_mprj_in_gates\[22\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_574_ la_data_out_mprj[103] vssd vssd vccd vccd _574_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[64\] _535_/Y la_buf\[64\]/TE vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__einvp_8
XPHY_151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[125\]_A _596_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[89\]_A user_to_mprj_in_gates\[89\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[28\]_B mprj_logic_high_inst/HI[358] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B mprj_logic_high_inst/HI[442] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[62\]_A _533_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[28\] _435_/Y mprj_adr_buf\[28\]/TE vssd vssd vccd vccd mprj_adr_o_user[28]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[120\] _591_/Y la_buf\[120\]/TE vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__einvp_8
XFILLER_12_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__440__A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] mprj_logic_high_inst/HI[383] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[53\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[13\]_A user_to_mprj_in_gates\[13\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[127\]_A user_to_mprj_in_gates\[127\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__615__A la_oen_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[116\]_A _587_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[19\]_B mprj_logic_high_inst/HI[349] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B mprj_logic_high_inst/HI[433] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[53\]_A _524_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__350__A la_oen_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[118\]_A user_to_mprj_in_gates\[118\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__525__A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[107\]_A _578_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[44\]_A _515_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_626_ la_oen_mprj[27] vssd vssd vccd vccd _626_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_557_ la_data_out_mprj[86] vssd vssd vccd vccd _557_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[109\]_A user_to_mprj_in_gates\[109\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_488_ la_data_out_mprj[17] vssd vssd vccd vccd _488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__435__A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y vssd vssd vccd vccd la_data_in_mprj[23]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[35\]_A _506_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[120\]_A _388_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__345__A la_oen_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_A _497_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[111\]_A _379_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_411_ mprj_adr_o_core[4] vssd vssd vccd vccd _411_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[1\] _600_/Y mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd la_oen_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_26_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_342_ la_oen_mprj[74] vssd vssd vccd vccd _342_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[11\]_TE la_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[17\]_A _488_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[27\] _498_/Y la_buf\[27\]/TE vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__einvp_8
XFILLER_13_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[102\]_A _370_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_609_ la_oen_mprj[10] vssd vssd vccd vccd _609_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] mprj_logic_high_inst/HI[346] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[16\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] mprj_logic_high_inst/HI[457] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[127\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_2010 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[34\]_TE la_buf\[34\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high_inst/HI[221] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[95\]_A _363_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_35 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[67\] _335_/Y mprj_logic_high_inst/HI[269] vssd vssd vccd
+ vccd la_oen_core[67] sky130_fd_sc_hd__einvp_8
XFILLER_8_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[15\] _454_/Y mprj_dat_buf\[15\]/TE vssd vssd vccd vccd mprj_dat_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[86\]_A _354_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[2\]_TE la_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[10\] _417_/Y mprj_adr_buf\[10\]/TE vssd vssd vccd vccd mprj_adr_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[124] sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_oen_buffers\[10\]_A _609_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y vssd vssd vccd vccd la_data_in_mprj[90]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[57\]_TE la_buf\[57\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[77\]_A _345_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__623__A la_oen_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[68\]_A _336_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__533__A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[94\] _565_/Y la_buf\[94\]/TE vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_21_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[59\]_A _658_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__443__A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] mprj_logic_high_inst/HI[413] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[83\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__618__A la_oen_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__353__A la_oen_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_590_ la_data_out_mprj[119] vssd vssd vccd vccd _590_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__528__A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[5\] _476_/Y la_buf\[5\]/TE vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__einvp_8
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[2\] _409_/Y mprj_adr_buf\[2\]/TE vssd vssd vccd vccd mprj_adr_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__438__A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y vssd vssd vccd vccd la_data_in_mprj[53]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[10\]_A _449_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[28\]_A _435_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__348__A la_oen_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_A _604_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[19\]_A _426_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_sel_buf\[0\] _403_/Y mprj_sel_buf\[0\]/TE vssd vssd vccd vccd mprj_sel_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_27_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_642_ la_oen_mprj[43] vssd vssd vccd vccd _642_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_573_ la_data_out_mprj[102] vssd vssd vccd vccd _573_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[57\] _528_/Y la_buf\[57\]/TE vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[105\]_TE la_buf\[105\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[113\] _584_/Y la_buf\[113\]/TE vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] mprj_logic_high_inst/HI[376] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[46\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high_inst/HI[254] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__631__A la_oen_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[8\]_TE mprj_dat_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] user_to_mprj_in_gates\[8\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[8\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[97\] _365_/Y mprj_logic_high_inst/HI[299] vssd vssd vccd
+ vccd la_oen_core[97] sky130_fd_sc_hd__einvp_8
XANTENNA__541__A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[90\]_TE la_buf\[90\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_625_ la_oen_mprj[26] vssd vssd vccd vccd _625_/Y sky130_fd_sc_hd__inv_2
X_556_ la_data_out_mprj[85] vssd vssd vccd vccd _556_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high_inst/HI[277] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_487_ la_data_out_mprj[16] vssd vssd vccd vccd _487_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y vssd vssd vccd vccd la_data_in_mprj[16]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__451__A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__626__A la_oen_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[4\]_A _411_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__361__A la_oen_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high_inst/HI[300] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_410_ mprj_adr_o_core[3] vssd vssd vccd vccd _410_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__536__A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[12\] _611_/Y mprj_logic_high_inst/HI[214] vssd vssd vccd
+ vccd la_oen_core[12] sky130_fd_sc_hd__einvp_8
X_341_ la_oen_mprj[73] vssd vssd vccd vccd _341_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y vssd vssd vccd vccd la_data_in_mprj[8]
+ sky130_fd_sc_hd__inv_8
XFILLER_10_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_stb_buf _401_/Y mprj_stb_buf/TE vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__einvp_8
XFILLER_4_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_608_ la_oen_mprj[9] vssd vssd vccd vccd _608_/Y sky130_fd_sc_hd__inv_2
XANTENNA__446__A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_539_ la_data_out_mprj[68] vssd vssd vccd vccd _539_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__356__A la_oen_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_clk_buf_A _398_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[30\]_TE mprj_adr_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[117] sky130_fd_sc_hd__inv_8
XFILLER_2_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y vssd vssd vccd vccd la_data_in_mprj[83]
+ sky130_fd_sc_hd__inv_8
XFILLER_24_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_B user_to_mprj_in_gates\[4\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[87\] _558_/Y la_buf\[87\]/TE vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_21_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_90 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[24\]_TE la_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] mprj_logic_high_inst/HI[406] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[76\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[8\]_A user_to_mprj_in_gates\[8\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__634__A la_oen_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__544__A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[47\]_TE la_buf\[47\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y vssd vssd vccd vccd la_data_in_mprj[46]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XPHY_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__454__A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__629__A la_oen_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] mprj_logic_high_inst/HI[432] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[102\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__364__A la_oen_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[112\] _380_/Y mprj_logic_high_inst/HI[314] vssd vssd vccd
+ vccd la_oen_core[112] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[42\] _641_/Y mprj_logic_high_inst/HI[244] vssd vssd vccd
+ vccd la_oen_core[42] sky130_fd_sc_hd__einvp_8
XANTENNA__539__A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_641_ la_oen_mprj[42] vssd vssd vccd vccd _641_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_572_ la_data_out_mprj[101] vssd vssd vccd vccd _572_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[106\] _577_/Y la_buf\[106\]/TE vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__einvp_8
XFILLER_7_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__449__A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] mprj_logic_high_inst/HI[369] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[39\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__359__A la_oen_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high_inst/HI[322] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_624_ la_oen_mprj[25] vssd vssd vccd vccd _624_/Y sky130_fd_sc_hd__inv_2
X_555_ la_data_out_mprj[84] vssd vssd vccd vccd _555_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_486_ la_data_out_mprj[15] vssd vssd vccd vccd _486_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_we_buf _402_/Y mprj_we_buf/TE vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__einvp_8
XFILLER_9_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_pwrgood mprj_pwrgood/A vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_9_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__642__A la_oen_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_340_ la_oen_mprj[72] vssd vssd vccd vccd _340_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__552__A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[42\]_TE mprj_logic_high_inst/HI[244] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_607_ la_oen_mprj[8] vssd vssd vccd vccd _607_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_538_ la_data_out_mprj[67] vssd vssd vccd vccd _538_/Y sky130_fd_sc_hd__inv_2
X_469_ mprj_dat_o_core[30] vssd vssd vccd vccd _469_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__462__A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[118\]_TE la_buf\[118\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__637__A la_oen_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_B mprj_logic_high_inst/HI[424] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__372__A la_oen_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[80\]_TE la_buf\[80\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[65\]_TE mprj_logic_high_inst/HI[267] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__547__A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_we_buf_A _402_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[85\]_B mprj_logic_high_inst/HI[415] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[32\] _503_/Y la_buf\[32\]/TE vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__einvp_8
XFILLER_13_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[70\]_A user_to_mprj_in_gates\[70\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y vssd vssd vccd vccd la_data_in_mprj[76]
+ sky130_fd_sc_hd__inv_8
XANTENNA__457__A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] mprj_logic_high_inst/HI[351] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[21\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[76\]_B mprj_logic_high_inst/HI[406] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high_inst/HI[290] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[9\] _448_/Y mprj_dat_buf\[9\]/TE vssd vssd vccd vccd mprj_dat_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_25_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[61\]_A user_to_mprj_in_gates\[61\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__367__A la_oen_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[67\]_B mprj_logic_high_inst/HI[397] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[72\] _340_/Y mprj_logic_high_inst/HI[274] vssd vssd vccd
+ vccd la_oen_core[72] sky130_fd_sc_hd__einvp_8
XFILLER_8_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[20\] _459_/Y mprj_dat_buf\[20\]/TE vssd vssd vccd vccd mprj_dat_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[52\]_A user_to_mprj_in_gates\[52\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[58\]_B mprj_logic_high_inst/HI[388] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[92\]_A _563_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[43\]_A user_to_mprj_in_gates\[43\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] mprj_logic_high_inst/HI[399] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[69\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_B mprj_logic_high_inst/HI[379] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[83\]_A _554_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__650__A la_oen_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[34\]_A user_to_mprj_in_gates\[34\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[20\]_TE mprj_adr_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[124\]_B mprj_logic_high_inst/HI[454] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[74\]_A _545_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__560__A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[25\]_A user_to_mprj_in_gates\[25\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[115\]_B mprj_logic_high_inst/HI[445] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y vssd vssd vccd vccd la_data_in_mprj[39]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[65\]_A _536_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__470__A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[16\]_A user_to_mprj_in_gates\[16\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__645__A la_oen_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[119\]_A _590_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_B mprj_logic_high_inst/HI[436] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[56\]_A _527_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__380__A la_oen_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[105\] _373_/Y mprj_logic_high_inst/HI[307] vssd vssd vccd
+ vccd la_oen_core[105] sky130_fd_sc_hd__einvp_8
XFILLER_5_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_640_ la_oen_mprj[41] vssd vssd vccd vccd _640_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_571_ la_data_out_mprj[100] vssd vssd vccd vccd _571_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[35\] _634_/Y mprj_logic_high_inst/HI[237] vssd vssd vccd
+ vccd la_oen_core[35] sky130_fd_sc_hd__einvp_8
XFILLER_18_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__555__A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[14\]_TE la_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[47\]_A _518_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__465__A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[38\]_A _509_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[123\]_A _391_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[37\]_TE la_buf\[37\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__375__A la_oen_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[29\]_A _500_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[114\]_A _382_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_623_ la_oen_mprj[24] vssd vssd vccd vccd _623_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[62\] _533_/Y la_buf\[62\]/TE vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__einvp_8
X_554_ la_data_out_mprj[83] vssd vssd vccd vccd _554_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_485_ la_data_out_mprj[14] vssd vssd vccd vccd _485_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[5\]_TE la_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[26\] _433_/Y mprj_adr_buf\[26\]/TE vssd vssd vccd vccd mprj_adr_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[40\]_A _639_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[105\]_A _373_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] mprj_logic_high_inst/HI[381] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[51\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[31\]_A _630_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_A _366_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[22\]_A _621_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_A _357_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_606_ la_oen_mprj[7] vssd vssd vccd vccd _606_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_537_ la_data_out_mprj[66] vssd vssd vccd vccd _537_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_468_ mprj_dat_o_core[29] vssd vssd vccd vccd _468_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_399_ caravel_clk2 vssd vssd vccd vccd _399_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y vssd vssd vccd vccd la_data_in_mprj[21]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_oen_buffers\[13\]_A _612_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] mprj_logic_high_inst/HI[429] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[99\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__653__A la_oen_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[110\]_TE mprj_logic_high_inst/HI[312] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__563__A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[25\] _496_/Y la_buf\[25\]/TE vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__einvp_8
XFILLER_6_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y vssd vssd vccd vccd la_data_in_mprj[69]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__473__A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] mprj_logic_high_inst/HI[344] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[14\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] mprj_logic_high_inst/HI[455] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[125\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__648__A la_oen_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[31\]_A _470_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__383__A la_oen_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[32\]_TE mprj_logic_high_inst/HI[234] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[65\] _333_/Y mprj_logic_high_inst/HI[267] vssd vssd vccd
+ vccd la_oen_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_8_1020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[13\] _452_/Y mprj_dat_buf\[13\]/TE vssd vssd vccd vccd mprj_dat_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__558__A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[108\]_TE la_buf\[108\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[22\]_A _461_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[7\]_TE mprj_adr_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[122] sky130_fd_sc_hd__inv_8
XFILLER_3_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__468__A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[70\]_TE la_buf\[70\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[13\]_A _452_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[55\]_TE mprj_logic_high_inst/HI[257] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__378__A la_oen_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[8\]_A _607_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[92\] _563_/Y la_buf\[92\]/TE vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[93\]_TE la_buf\[93\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high_inst/HI[280] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] mprj_logic_high_inst/HI[411] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[81\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_570_ la_data_out_mprj[99] vssd vssd vccd vccd _570_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[28\] _627_/Y mprj_logic_high_inst/HI[230] vssd vssd vccd
+ vccd la_oen_core[28] sky130_fd_sc_hd__einvp_8
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[0\]_A _471_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__571__A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[3\] _474_/Y la_buf\[3\]/TE vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__einvp_8
XFILLER_10_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[0\] _407_/Y mprj_adr_buf\[0\]/TE vssd vssd vccd vccd mprj_adr_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y vssd vssd vccd vccd la_data_in_mprj[51]
+ sky130_fd_sc_hd__inv_8
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__481__A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__656__A la_oen_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[7\]_A _414_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__391__A la_oen_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_622_ la_oen_mprj[23] vssd vssd vccd vccd _622_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__566__A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_553_ la_data_out_mprj[82] vssd vssd vccd vccd _553_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_484_ la_data_out_mprj[13] vssd vssd vccd vccd _484_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[55\] _526_/Y la_buf\[55\]/TE vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__einvp_8
XFILLER_18_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[19\] _426_/Y mprj_adr_buf\[19\]/TE vssd vssd vccd vccd mprj_adr_o_user[19]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[111\] _582_/Y la_buf\[111\]/TE vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__einvp_8
XFILLER_25_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y vssd vssd vccd vccd la_data_in_mprj[99]
+ sky130_fd_sc_hd__inv_8
XFILLER_23_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__476__A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] mprj_logic_high_inst/HI[374] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[44\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] user_to_mprj_in_gates\[6\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[6\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__386__A la_oen_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[95\] _363_/Y mprj_logic_high_inst/HI[297] vssd vssd vccd
+ vccd la_oen_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_5_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_81 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_605_ la_oen_mprj[6] vssd vssd vccd vccd _605_/Y sky130_fd_sc_hd__inv_2
X_536_ la_data_out_mprj[65] vssd vssd vccd vccd _536_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_467_ mprj_dat_o_core[28] vssd vssd vccd vccd _467_/Y sky130_fd_sc_hd__inv_2
X_398_ caravel_clk vssd vssd vccd vccd _398_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y vssd vssd vccd vccd la_data_in_mprj[14]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[27\]_TE la_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[7\]_B user_to_mprj_in_gates\[7\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[10\] _609_/Y mprj_logic_high_inst/HI[212] vssd vssd vccd
+ vccd la_oen_core[10] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y vssd vssd vccd vccd la_data_in_mprj[6]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[18\] _489_/Y la_buf\[18\]/TE vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_13_1498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_519_ la_data_out_mprj[48] vssd vssd vccd vccd _519_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] mprj_logic_high_inst/HI[448] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[118\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[58\] _657_/Y mprj_logic_high_inst/HI[260] vssd vssd vccd
+ vccd la_oen_core[58] sky130_fd_sc_hd__einvp_8
XFILLER_5_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__574__A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[115] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y vssd vssd vccd vccd la_data_in_mprj[81]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high_inst/HI[302] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__484__A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_1_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__659__A la_oen_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__394__A la_oen_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_51 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__569__A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high_inst/HI[325] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[85\] _556_/Y la_buf\[85\]/TE vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_19_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__479__A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] mprj_logic_high_inst/HI[404] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[74\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[22\]_TE mprj_logic_high_inst/HI[224] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__389__A la_oen_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[60\]_TE la_buf\[60\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[45\]_TE mprj_logic_high_inst/HI[247] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y vssd vssd vccd vccd la_data_in_mprj[44]
+ sky130_fd_sc_hd__inv_8
XPHY_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_sel_buf\[1\]_A _404_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] mprj_logic_high_inst/HI[430] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[100\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[83\]_TE la_buf\[83\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[68\]_TE mprj_logic_high_inst/HI[270] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[110\] _378_/Y mprj_logic_high_inst/HI[312] vssd vssd vccd
+ vccd la_oen_core[110] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[40\] _639_/Y mprj_logic_high_inst/HI[242] vssd vssd vccd
+ vccd la_oen_core[40] sky130_fd_sc_hd__einvp_8
X_621_ la_oen_mprj[22] vssd vssd vccd vccd _621_/Y sky130_fd_sc_hd__inv_2
X_552_ la_data_out_mprj[81] vssd vssd vccd vccd _552_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_483_ la_data_out_mprj[12] vssd vssd vccd vccd _483_/Y sky130_fd_sc_hd__inv_2
XANTENNA__582__A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[48\] _519_/Y la_buf\[48\]/TE vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_9_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[2\]_A _441_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[104\] _575_/Y la_buf\[104\]/TE vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_23_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] mprj_logic_high_inst/HI[367] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[37\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__492__A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[91\]_A user_to_mprj_in_gates\[91\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[30\]_B mprj_logic_high_inst/HI[360] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_B mprj_logic_high_inst/HI[427] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[88\] _356_/Y mprj_logic_high_inst/HI[290] vssd vssd vccd
+ vccd la_oen_core[88] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[21\]_B mprj_logic_high_inst/HI[351] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[82\]_A user_to_mprj_in_gates\[82\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__577__A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_604_ la_oen_mprj[5] vssd vssd vccd vccd _604_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_535_ la_data_out_mprj[64] vssd vssd vccd vccd _535_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[88\]_B mprj_logic_high_inst/HI[418] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_466_ mprj_dat_o_core[27] vssd vssd vccd vccd _466_/Y sky130_fd_sc_hd__inv_2
X_397_ user_resetn vssd vssd vccd vccd user_reset sky130_fd_sc_hd__inv_2
XFILLER_9_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[31\] _438_/Y mprj_adr_buf\[31\]/TE vssd vssd vccd vccd mprj_adr_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[120\]_A user_to_mprj_in_gates\[120\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[73\]_A user_to_mprj_in_gates\[73\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_B mprj_logic_high_inst/HI[342] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__487__A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[79\]_B mprj_logic_high_inst/HI[409] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[111\]_A user_to_mprj_in_gates\[111\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[100\]_A _571_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[64\]_A user_to_mprj_in_gates\[64\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__397__A user_resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[23\]_TE mprj_adr_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[102\]_A user_to_mprj_in_gates\[102\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[55\]_A user_to_mprj_in_gates\[55\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_518_ la_data_out_mprj[47] vssd vssd vccd vccd _518_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[95\]_A _566_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_449_ mprj_dat_o_core[10] vssd vssd vccd vccd _449_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[46\]_A user_to_mprj_in_gates\[46\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[86\]_A _557_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[37\]_A user_to_mprj_in_gates\[37\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[10\]_A _481_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[17\]_TE la_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_B mprj_logic_high_inst/HI[457] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[77\]_A _548_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__590__A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[30\] _501_/Y la_buf\[30\]/TE vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[28\]_A user_to_mprj_in_gates\[28\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[108] sky130_fd_sc_hd__inv_8
XFILLER_26_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y vssd vssd vccd vccd la_data_in_mprj[74]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[118\]_B mprj_logic_high_inst/HI[448] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[68\]_A _539_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_2010 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[19\]_A user_to_mprj_in_gates\[19\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[7\] _446_/Y mprj_dat_buf\[7\]/TE vssd vssd vccd vccd mprj_dat_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[109\]_B mprj_logic_high_inst/HI[439] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[59\]_A _530_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[70\] _338_/Y mprj_logic_high_inst/HI[272] vssd vssd vccd
+ vccd la_oen_core[70] sky130_fd_sc_hd__einvp_8
XFILLER_10_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[78\] _549_/Y la_buf\[78\]/TE vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__einvp_8
XANTENNA__585__A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[8\]_TE la_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[70\]_A _338_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] mprj_logic_high_inst/HI[397] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[67\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__495__A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[126\]_A _394_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[61\]_A _660_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[52\]_A _651_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_A _385_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y vssd vssd vccd vccd la_data_in_mprj[37]
+ sky130_fd_sc_hd__inv_8
XPHY_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[108\]_A _376_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[43\]_A _642_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high_inst/HI[315] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[34\]_A _633_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[103\] _371_/Y mprj_logic_high_inst/HI[305] vssd vssd vccd
+ vccd la_oen_core[103] sky130_fd_sc_hd__einvp_8
X_620_ la_oen_mprj[21] vssd vssd vccd vccd _620_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_551_ la_data_out_mprj[80] vssd vssd vccd vccd _551_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[33\] _632_/Y mprj_logic_high_inst/HI[235] vssd vssd vccd
+ vccd la_oen_core[33] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[30\]_A _437_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_482_ la_data_out_mprj[11] vssd vssd vccd vccd _482_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high_inst/HI[214] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[25\]_A _624_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[21\]_A _428_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj2_vdd_pwrgood_A mprj2_vdd_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_A _615_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[12\]_A _419_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[50\]_TE la_buf\[50\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high_inst/HI[237] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[29\] _468_/Y mprj_dat_buf\[29\]/TE vssd vssd vccd vccd mprj_dat_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_603_ la_oen_mprj[4] vssd vssd vccd vccd _603_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_534_ la_data_out_mprj[63] vssd vssd vccd vccd _534_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[60\] _531_/Y la_buf\[60\]/TE vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__einvp_8
X_465_ mprj_dat_o_core[26] vssd vssd vccd vccd _465_/Y sky130_fd_sc_hd__inv_2
XANTENNA__593__A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_396_ caravel_rstn vssd vssd vccd vccd _396_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[24\] _431_/Y mprj_adr_buf\[24\]/TE vssd vssd vccd vccd mprj_adr_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[73\]_TE la_buf\[73\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[58\]_TE mprj_logic_high_inst/HI[260] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[1\]_TE mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__588__A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[96\]_TE la_buf\[96\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[25\]_A _464_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_517_ la_data_out_mprj[46] vssd vssd vccd vccd _517_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_448_ mprj_dat_o_core[9] vssd vssd vccd vccd _448_/Y sky130_fd_sc_hd__inv_2
X_379_ la_oen_mprj[111] vssd vssd vccd vccd _379_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] mprj_logic_high_inst/HI[427] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[97\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__498__A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[16\]_A _455_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[23\] _494_/Y la_buf\[23\]/TE vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__einvp_8
XFILLER_3_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y vssd vssd vccd vccd la_data_in_mprj[67]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] mprj_logic_high_inst/HI[342] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[12\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_TE mprj_adr_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] mprj_logic_high_inst/HI[453] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[123\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[63\] _331_/Y mprj_logic_high_inst/HI[265] vssd vssd vccd
+ vccd la_oen_core[63] sky130_fd_sc_hd__einvp_8
XFILLER_27_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[11\] _450_/Y mprj_dat_buf\[11\]/TE vssd vssd vccd vccd mprj_dat_o_user[11]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[1\]_TE mprj_dat_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_A _474_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[121\]_TE la_buf\[121\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[127\] _598_/Y la_buf\[127\]/TE vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[120] sky130_fd_sc_hd__inv_8
XFILLER_18_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__596__A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[90\] _561_/Y la_buf\[90\]/TE vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_21_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high_inst/HI[293] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[1\]_A user_to_mprj_in_gates\[1\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_550_ la_data_out_mprj[79] vssd vssd vccd vccd _550_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[8\] _607_/Y mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd la_oen_core[8] sky130_fd_sc_hd__einvp_8
X_481_ la_data_out_mprj[10] vssd vssd vccd vccd _481_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[26\] _625_/Y mprj_logic_high_inst/HI[228] vssd vssd vccd
+ vccd la_oen_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_25_450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[1\] _472_/Y la_buf\[1\]/TE vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_10_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_602_ la_oen_mprj[3] vssd vssd vccd vccd _602_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_533_ la_data_out_mprj[62] vssd vssd vccd vccd _533_/Y sky130_fd_sc_hd__inv_2
X_464_ mprj_dat_o_core[25] vssd vssd vccd vccd _464_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[53\] _524_/Y la_buf\[53\]/TE vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__einvp_8
X_395_ la_oen_mprj[127] vssd vssd vccd vccd _395_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[17\] _424_/Y mprj_adr_buf\[17\]/TE vssd vssd vccd vccd mprj_adr_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y vssd vssd vccd vccd la_data_in_mprj[97]
+ sky130_fd_sc_hd__inv_8
XFILLER_27_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high_inst/HI[305] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] mprj_logic_high_inst/HI[372] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[42\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] user_to_mprj_in_gates\[4\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[4\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[93\] _361_/Y mprj_logic_high_inst/HI[295] vssd vssd vccd
+ vccd la_oen_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_2_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high_inst/HI[328] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_516_ la_data_out_mprj[45] vssd vssd vccd vccd _516_/Y sky130_fd_sc_hd__inv_2
X_447_ mprj_dat_o_core[8] vssd vssd vccd vccd _447_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_378_ la_oen_mprj[110] vssd vssd vccd vccd _378_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y vssd vssd vccd vccd la_data_in_mprj[12]
+ sky130_fd_sc_hd__inv_8
XFILLER_6_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[40\]_TE la_buf\[40\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[25\]_TE mprj_logic_high_inst/HI[227] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y vssd vssd vccd vccd la_data_in_mprj[4]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[63\]_TE la_buf\[63\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[16\] _487_/Y la_buf\[16\]/TE vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[48\]_TE mprj_logic_high_inst/HI[250] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__599__A la_oen_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[9\] _416_/Y mprj_adr_buf\[9\]/TE vssd vssd vccd vccd mprj_adr_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] mprj_logic_high_inst/HI[446] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[116\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[86\]_TE la_buf\[86\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[126\] _394_/Y mprj_logic_high_inst/HI[328] vssd vssd vccd
+ vccd la_oen_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_0_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[56\] _655_/Y mprj_logic_high_inst/HI[258] vssd vssd vccd
+ vccd la_oen_core[56] sky130_fd_sc_hd__einvp_8
XFILLER_19_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[113] sky130_fd_sc_hd__inv_8
XFILLER_26_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[60\]_B mprj_logic_high_inst/HI[390] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[51\]_B mprj_logic_high_inst/HI[381] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[83\] _554_/Y la_buf\[83\]/TE vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__einvp_8
XFILLER_21_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[5\]_A _444_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[42\]_B mprj_logic_high_inst/HI[372] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] mprj_logic_high_inst/HI[402] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[72\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[94\]_A user_to_mprj_in_gates\[94\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[33\]_B mprj_logic_high_inst/HI[363] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[111\]_TE la_buf\[111\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[26\]_TE mprj_adr_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_480_ la_data_out_mprj[9] vssd vssd vccd vccd _480_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[19\] _618_/Y mprj_logic_high_inst/HI[221] vssd vssd vccd
+ vccd la_oen_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_25_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[121\]_A _592_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[85\]_A user_to_mprj_in_gates\[85\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[24\]_B mprj_logic_high_inst/HI[354] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__400__A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y vssd vssd vccd vccd la_data_in_mprj[42]
+ sky130_fd_sc_hd__inv_8
XPHY_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[123\]_A user_to_mprj_in_gates\[123\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[112\]_A _583_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_B mprj_logic_high_inst/HI[345] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[76\]_A user_to_mprj_in_gates\[76\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[114\]_A user_to_mprj_in_gates\[114\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[103\]_A _574_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[67\]_A user_to_mprj_in_gates\[67\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[40\]_A _511_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high_inst/HI[283] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_601_ la_oen_mprj[2] vssd vssd vccd vccd _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_532_ la_data_out_mprj[61] vssd vssd vccd vccd _532_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_463_ mprj_dat_o_core[24] vssd vssd vccd vccd _463_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_394_ la_oen_mprj[126] vssd vssd vccd vccd _394_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[46\] _517_/Y la_buf\[46\]/TE vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[105\]_A user_to_mprj_in_gates\[105\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[58\]_A user_to_mprj_in_gates\[58\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[31\]_A _502_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[102\] _573_/Y la_buf\[102\]/TE vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_1_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[98\]_A _569_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] mprj_logic_high_inst/HI[365] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[35\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[49\]_A user_to_mprj_in_gates\[49\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[22\]_A _493_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[89\]_A _560_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[86\] _354_/Y mprj_logic_high_inst/HI[288] vssd vssd vccd
+ vccd la_oen_core[86] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[13\]_A _484_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_515_ la_data_out_mprj[44] vssd vssd vccd vccd _515_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_446_ mprj_dat_o_core[7] vssd vssd vccd vccd _446_/Y sky130_fd_sc_hd__inv_2
X_377_ la_oen_mprj[109] vssd vssd vccd vccd _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[91\]_A _359_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_A _350_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_429_ mprj_adr_o_core[22] vssd vssd vccd vccd _429_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[73\]_A _341_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] mprj_logic_high_inst/HI[439] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[109\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high_inst/HI[318] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[64\]_A _332_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[119\] _387_/Y mprj_logic_high_inst/HI[321] vssd vssd vccd
+ vccd la_oen_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_0_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[49\] _648_/Y mprj_logic_high_inst/HI[251] vssd vssd vccd
+ vccd la_oen_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_15_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[30\]_TE la_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high_inst/HI[217] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[55\]_A _654_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__403__A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[106] sky130_fd_sc_hd__inv_8
XFILLER_4_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y vssd vssd vccd vccd la_data_in_mprj[72]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[46\]_A _645_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[5\] _444_/Y mprj_dat_buf\[5\]/TE vssd vssd vccd vccd mprj_dat_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[53\]_TE la_buf\[53\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[38\]_TE mprj_logic_high_inst/HI[240] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[37\]_A _636_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[76\] _547_/Y la_buf\[76\]/TE vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__einvp_8
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[28\]_A _627_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[76\]_TE la_buf\[76\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[24\]_A _431_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] mprj_logic_high_inst/HI[395] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[65\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[19\]_A _618_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[1\]_A _600_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[15\]_A _422_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[99\]_TE la_buf\[99\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y vssd vssd vccd vccd la_data_in_mprj[35]
+ sky130_fd_sc_hd__inv_8
XPHY_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__501__A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _369_/Y mprj_logic_high_inst/HI[303] vssd vssd vccd
+ vccd la_oen_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_24_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_600_ la_oen_mprj[1] vssd vssd vccd vccd _600_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[31\] _630_/Y mprj_logic_high_inst/HI[233] vssd vssd vccd
+ vccd la_oen_core[31] sky130_fd_sc_hd__einvp_8
X_531_ la_data_out_mprj[60] vssd vssd vccd vccd _531_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_462_ mprj_dat_o_core[23] vssd vssd vccd vccd _462_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_393_ la_oen_mprj[125] vssd vssd vccd vccd _393_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[39\] _510_/Y la_buf\[39\]/TE vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_12_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__411__A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[28\]_A _467_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] mprj_logic_high_inst/HI[358] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[28\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[101\]_TE la_buf\[101\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[0\]_A _407_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_A _458_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_66 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[79\] _347_/Y mprj_logic_high_inst/HI[281] vssd vssd vccd
+ vccd la_oen_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_1_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[27\] _466_/Y mprj_dat_buf\[27\]/TE vssd vssd vccd vccd mprj_dat_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[4\]_TE mprj_dat_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_514_ la_data_out_mprj[43] vssd vssd vccd vccd _514_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[124\]_TE la_buf\[124\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_445_ mprj_dat_o_core[6] vssd vssd vccd vccd _445_/Y sky130_fd_sc_hd__inv_2
X_376_ la_oen_mprj[108] vssd vssd vccd vccd _376_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__406__A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[22\] _429_/Y mprj_adr_buf\[22\]/TE vssd vssd vccd vccd mprj_adr_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high_inst/HI[273] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[6\]_A _477_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high_inst/HI[296] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_428_ mprj_adr_o_core[21] vssd vssd vccd vccd _428_/Y sky130_fd_sc_hd__inv_2
X_359_ la_oen_mprj[91] vssd vssd vccd vccd _359_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] mprj_logic_high_inst/HI[425] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[95\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[0\]_B user_to_mprj_in_gates\[0\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[21\] _492_/Y la_buf\[21\]/TE vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__einvp_8
XFILLER_10_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[4\]_A user_to_mprj_in_gates\[4\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y vssd vssd vccd vccd la_data_in_mprj[65]
+ sky130_fd_sc_hd__inv_8
XFILLER_21_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] mprj_logic_high_inst/HI[340] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[10\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] mprj_logic_high_inst/HI[451] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[121\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__504__A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_66 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[61\] _660_/Y mprj_logic_high_inst/HI[263] vssd vssd vccd
+ vccd la_oen_core[61] sky130_fd_sc_hd__einvp_8
XFILLER_21_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[69\] _540_/Y la_buf\[69\]/TE vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__einvp_8
XPHY_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__414__A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[125\] _596_/Y la_buf\[125\]/TE vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_10_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high_inst/HI[308] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] mprj_logic_high_inst/HI[388] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[58\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[20\]_TE la_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_88 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__409__A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y vssd vssd vccd vccd la_data_in_mprj[28]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[43\]_TE la_buf\[43\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[28\]_TE mprj_logic_high_inst/HI[230] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_530_ la_data_out_mprj[59] vssd vssd vccd vccd _530_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[24\] _623_/Y mprj_logic_high_inst/HI[226] vssd vssd vccd
+ vccd la_oen_core[24] sky130_fd_sc_hd__einvp_8
X_461_ mprj_dat_o_core[22] vssd vssd vccd vccd _461_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[6\] _605_/Y mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd la_oen_core[6] sky130_fd_sc_hd__einvp_8
X_392_ la_oen_mprj[124] vssd vssd vccd vccd _392_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[66\]_TE la_buf\[66\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_659_ la_oen_mprj[60] vssd vssd vccd vccd _659_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[15\]_TE mprj_dat_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__602__A la_oen_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[89\]_TE la_buf\[89\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__512__A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_513_ la_data_out_mprj[42] vssd vssd vccd vccd _513_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_444_ mprj_dat_o_core[5] vssd vssd vccd vccd _444_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[51\] _522_/Y la_buf\[51\]/TE vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__einvp_8
X_375_ la_oen_mprj[107] vssd vssd vccd vccd _375_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__422__A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[15\] _422_/Y mprj_adr_buf\[15\]/TE vssd vssd vccd vccd mprj_adr_o_user[15]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y vssd vssd vccd vccd la_data_in_mprj[95]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] mprj_logic_high_inst/HI[370] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[40\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[90\]_B mprj_logic_high_inst/HI[420] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__332__A la_oen_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] user_to_mprj_in_gates\[2\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[2\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__507__A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[81\]_B mprj_logic_high_inst/HI[411] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[91\] _359_/Y mprj_logic_high_inst/HI[293] vssd vssd vccd
+ vccd la_oen_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_26_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[99\] _570_/Y la_buf\[99\]/TE vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_24_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__417__A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_427_ mprj_adr_o_core[20] vssd vssd vccd vccd _427_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_358_ la_oen_mprj[90] vssd vssd vccd vccd _358_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[72\]_B mprj_logic_high_inst/HI[402] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y vssd vssd vccd vccd la_data_in_mprj[10]
+ sky130_fd_sc_hd__inv_8
XFILLER_5_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] mprj_logic_high_inst/HI[418] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[88\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_B mprj_logic_high_inst/HI[393] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[114\]_TE la_buf\[114\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_TE mprj_adr_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y vssd vssd vccd vccd la_data_in_mprj[2]
+ sky130_fd_sc_hd__inv_8
XPHY_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[54\]_B mprj_logic_high_inst/HI[384] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[14\] _485_/Y la_buf\[14\]/TE vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_10_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[61\]_TE mprj_logic_high_inst/HI[263] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[7\] _414_/Y mprj_adr_buf\[7\]/TE vssd vssd vccd vccd mprj_adr_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y vssd vssd vccd vccd la_data_in_mprj[58]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[8\]_A _447_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[45\]_B mprj_logic_high_inst/HI[375] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__610__A la_oen_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] mprj_logic_high_inst/HI[444] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[114\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[30\]_A user_to_mprj_in_gates\[30\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[120\]_B mprj_logic_high_inst/HI[450] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_B mprj_logic_high_inst/HI[366] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[97\]_A user_to_mprj_in_gates\[97\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[70\]_A _541_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high_inst/HI[286] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[124\] _392_/Y mprj_logic_high_inst/HI[326] vssd vssd vccd
+ vccd la_oen_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_7_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__520__A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[54\] _653_/Y mprj_logic_high_inst/HI[256] vssd vssd vccd
+ vccd la_oen_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_21_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[21\]_A user_to_mprj_in_gates\[21\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[124\]_A _595_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B mprj_logic_high_inst/HI[441] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[88\]_A user_to_mprj_in_gates\[88\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_B mprj_logic_high_inst/HI[357] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[61\]_A _532_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[118\] _589_/Y la_buf\[118\]/TE vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_10_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[111] sky130_fd_sc_hd__inv_8
XANTENNA__430__A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[12\]_A user_to_mprj_in_gates\[12\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[126\]_A user_to_mprj_in_gates\[126\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__605__A la_oen_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[115\]_A _586_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[79\]_A user_to_mprj_in_gates\[79\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_B mprj_logic_high_inst/HI[348] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_B mprj_logic_high_inst/HI[432] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[52\]_A _523_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__340__A la_oen_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[117\]_A user_to_mprj_in_gates\[117\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__515__A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[106\]_A _577_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_A _514_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[81\] _552_/Y la_buf\[81\]/TE vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_5_2084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[108\]_A user_to_mprj_in_gates\[108\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__425__A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[34\]_A _505_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] mprj_logic_high_inst/HI[400] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[70\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_clk_buf _398_/Y mprj_clk_buf/TE vssd vssd vccd vccd user_clock sky130_fd_sc_hd__einvp_8
XFILLER_22_446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__335__A la_oen_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[25\]_A _496_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[110\]_A _378_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_460_ mprj_dat_o_core[21] vssd vssd vccd vccd _460_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_391_ la_oen_mprj[123] vssd vssd vccd vccd _391_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[17\] _616_/Y mprj_logic_high_inst/HI[219] vssd vssd vccd
+ vccd la_oen_core[17] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[16\]_A _487_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[101\]_A _369_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_658_ la_oen_mprj[59] vssd vssd vccd vccd _658_/Y sky130_fd_sc_hd__inv_2
X_589_ la_data_out_mprj[118] vssd vssd vccd vccd _589_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[10\]_TE la_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y vssd vssd vccd vccd la_data_in_mprj[40]
+ sky130_fd_sc_hd__inv_8
XPHY_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high_inst/HI[321] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_A _362_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_512_ la_data_out_mprj[41] vssd vssd vccd vccd _512_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[33\]_TE la_buf\[33\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_443_ mprj_dat_o_core[4] vssd vssd vccd vccd _443_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high_inst/HI[220] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_A _353_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_374_ la_oen_mprj[106] vssd vssd vccd vccd _374_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[44\] _515_/Y la_buf\[44\]/TE vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_9_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[100\] _571_/Y la_buf\[100\]/TE vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_0_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y vssd vssd vccd vccd la_data_in_mprj[88]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] mprj_logic_high_inst/HI[363] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[33\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[76\]_A _344_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[1\]_TE la_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__613__A la_oen_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[56\]_TE la_buf\[56\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[67\]_A _335_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__523__A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[84\] _352_/Y mprj_logic_high_inst/HI[286] vssd vssd vccd
+ vccd la_oen_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_3_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[58\]_A _657_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_426_ mprj_adr_o_core[19] vssd vssd vccd vccd _426_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_357_ la_oen_mprj[89] vssd vssd vccd vccd _357_/Y sky130_fd_sc_hd__inv_2
XANTENNA__433__A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[79\]_TE la_buf\[79\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__608__A la_oen_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[49\]_A _648_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__343__A la_oen_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[7\]_TE mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__428__A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_409_ mprj_adr_o_core[2] vssd vssd vccd vccd _409_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_adr_buf\[27\]_A _434_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_sel_buf\[2\]_TE mprj_sel_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] mprj_logic_high_inst/HI[437] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[107\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__338__A la_oen_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[4\]_A _603_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[18\]_A _425_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[117\] _385_/Y mprj_logic_high_inst/HI[319] vssd vssd vccd
+ vccd la_oen_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_21_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[47\] _646_/Y mprj_logic_high_inst/HI[249] vssd vssd vccd
+ vccd la_oen_core[47] sky130_fd_sc_hd__einvp_8
XPHY_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[104] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y vssd vssd vccd vccd la_data_in_mprj[70]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[104\]_TE la_buf\[104\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[19\]_TE mprj_adr_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__621__A la_oen_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[3\] _442_/Y mprj_dat_buf\[3\]/TE vssd vssd vccd vccd mprj_dat_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_22_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[51\]_TE mprj_logic_high_inst/HI[253] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__531__A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[7\]_TE mprj_dat_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[127\]_TE la_buf\[127\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[74\] _545_/Y la_buf\[74\]/TE vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__einvp_8
XFILLER_16_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__441__A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] mprj_logic_high_inst/HI[393] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[63\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high_inst/HI[276] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__616__A la_oen_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[3\]_A _410_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__351__A la_oen_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_390_ la_oen_mprj[122] vssd vssd vccd vccd _390_/Y sky130_fd_sc_hd__inv_2
XANTENNA__526__A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high_inst/HI[299] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_657_ la_oen_mprj[58] vssd vssd vccd vccd _657_/Y sky130_fd_sc_hd__inv_2
X_588_ la_data_out_mprj[117] vssd vssd vccd vccd _588_/Y sky130_fd_sc_hd__inv_2
XANTENNA__436__A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y vssd vssd vccd vccd la_data_in_mprj[33]
+ sky130_fd_sc_hd__inv_8
XPHY_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__346__A la_oen_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_511_ la_data_out_mprj[40] vssd vssd vccd vccd _511_/Y sky130_fd_sc_hd__inv_2
X_442_ mprj_dat_o_core[3] vssd vssd vccd vccd _442_/Y sky130_fd_sc_hd__inv_2
X_373_ la_oen_mprj[105] vssd vssd vccd vccd _373_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[37\] _508_/Y la_buf\[37\]/TE vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_A _480_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] mprj_logic_high_inst/HI[356] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[26\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_B user_to_mprj_in_gates\[3\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[77\] _345_/Y mprj_logic_high_inst/HI[279] vssd vssd vccd
+ vccd la_oen_core[77] sky130_fd_sc_hd__einvp_8
XFILLER_3_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[25\] _464_/Y mprj_dat_buf\[25\]/TE vssd vssd vccd vccd mprj_dat_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_425_ mprj_adr_o_core[18] vssd vssd vccd vccd _425_/Y sky130_fd_sc_hd__inv_2
X_356_ la_oen_mprj[88] vssd vssd vccd vccd _356_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[20\] _427_/Y mprj_adr_buf\[20\]/TE vssd vssd vccd vccd mprj_adr_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high_inst/HI[311] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[7\]_A user_to_mprj_in_gates\[7\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__624__A la_oen_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_TE la_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__534__A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_408_ mprj_adr_o_core[1] vssd vssd vccd vccd _408_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__444__A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_339_ la_oen_mprj[71] vssd vssd vccd vccd _339_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[46\]_TE la_buf\[46\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] mprj_logic_high_inst/HI[423] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[93\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__619__A la_oen_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__354__A la_oen_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_14_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__529__A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[69\]_TE la_buf\[69\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__439__A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y vssd vssd vccd vccd la_data_in_mprj[63]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_TE mprj_dat_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__349__A la_oen_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[67\] _538_/Y la_buf\[67\]/TE vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__einvp_8
XPHY_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[123\] _594_/Y la_buf\[123\]/TE vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__einvp_8
XFILLER_26_1066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] mprj_logic_high_inst/HI[386] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[56\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__632__A la_oen_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__542__A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_656_ la_oen_mprj[57] vssd vssd vccd vccd _656_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_587_ la_data_out_mprj[116] vssd vssd vccd vccd _587_/Y sky130_fd_sc_hd__inv_2
XPHY_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y vssd vssd vccd vccd la_data_in_mprj[26]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__452__A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[41\]_TE mprj_logic_high_inst/HI[243] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__627__A la_oen_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[93\]_B mprj_logic_high_inst/HI[423] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__362__A la_oen_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[117\]_TE la_buf\[117\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_510_ la_data_out_mprj[39] vssd vssd vccd vccd _510_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[4\] _603_/Y mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd la_oen_core[4] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[22\] _621_/Y mprj_logic_high_inst/HI[224] vssd vssd vccd
+ vccd la_oen_core[22] sky130_fd_sc_hd__einvp_8
XANTENNA__537__A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_441_ mprj_dat_o_core[2] vssd vssd vccd vccd _441_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_372_ la_oen_mprj[104] vssd vssd vccd vccd _372_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B mprj_logic_high_inst/HI[414] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[64\]_TE mprj_logic_high_inst/HI[266] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__447__A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_639_ la_oen_mprj[40] vssd vssd vccd vccd _639_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] mprj_logic_high_inst/HI[349] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[19\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[75\]_B mprj_logic_high_inst/HI[405] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[60\]_A user_to_mprj_in_gates\[60\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__357__A la_oen_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_B mprj_logic_high_inst/HI[396] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high_inst/HI[289] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[18\] _457_/Y mprj_dat_buf\[18\]/TE vssd vssd vccd vccd mprj_dat_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[51\]_A user_to_mprj_in_gates\[51\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_424_ mprj_adr_o_core[17] vssd vssd vccd vccd _424_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_355_ la_oen_mprj[87] vssd vssd vccd vccd _355_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_B mprj_logic_high_inst/HI[387] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[91\]_A _562_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[13\] _420_/Y mprj_adr_buf\[13\]/TE vssd vssd vccd vccd mprj_adr_o_user[13]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[127] sky130_fd_sc_hd__inv_8
XFILLER_9_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y vssd vssd vccd vccd la_data_in_mprj[93]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_buffers\[42\]_A user_to_mprj_in_gates\[42\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[48\]_B mprj_logic_high_inst/HI[378] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[82\]_A _553_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__640__A la_oen_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] user_to_mprj_in_gates\[0\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[0\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[33\]_A user_to_mprj_in_gates\[33\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[123\]_B mprj_logic_high_inst/HI[453] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[39\]_B mprj_logic_high_inst/HI[369] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[73\]_A _544_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__550__A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[24\]_A user_to_mprj_in_gates\[24\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[97\] _568_/Y la_buf\[97\]/TE vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__einvp_8
XFILLER_4_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_407_ mprj_adr_o_core[0] vssd vssd vccd vccd _407_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[127\]_A _598_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_B mprj_logic_high_inst/HI[444] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_14_395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_338_ la_oen_mprj[70] vssd vssd vccd vccd _338_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[64\]_A _535_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__460__A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] mprj_logic_high_inst/HI[416] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[86\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[15\]_A user_to_mprj_in_gates\[15\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__635__A la_oen_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[118\]_A _589_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_B mprj_logic_high_inst/HI[435] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[55\]_A _526_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__370__A la_oen_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__545__A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y vssd vssd vccd vccd la_data_in_mprj[0]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[109\]_A _580_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[46\]_A _517_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[8\] _479_/Y la_buf\[8\]/TE vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__einvp_8
Xla_buf\[12\] _483_/Y la_buf\[12\]/TE vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__einvp_8
XFILLER_10_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[5\] _412_/Y mprj_adr_buf\[5\]/TE vssd vssd vccd vccd mprj_adr_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y vssd vssd vccd vccd la_data_in_mprj[56]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[13\]_TE la_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__455__A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[37\]_A _508_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[122\]_A _390_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] mprj_logic_high_inst/HI[442] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[112\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__365__A la_oen_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[28\]_A _499_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[122\] _390_/Y mprj_logic_high_inst/HI[324] vssd vssd vccd
+ vccd la_oen_core[122] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[113\]_A _381_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_sel_buf\[3\] _406_/Y mprj_sel_buf\[3\]/TE vssd vssd vccd vccd mprj_sel_o_user[3]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[52\] _651_/Y mprj_logic_high_inst/HI[254] vssd vssd vccd
+ vccd la_oen_core[52] sky130_fd_sc_hd__einvp_8
XFILLER_5_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[36\]_TE la_buf\[36\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[19\]_A _490_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[116\] _587_/Y la_buf\[116\]/TE vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[104\]_A _372_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk2_buf_A _399_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] mprj_logic_high_inst/HI[379] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[49\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[4\]_TE la_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_A _629_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[59\]_TE la_buf\[59\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_A _365_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[21\]_A _620_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_655_ la_oen_mprj[56] vssd vssd vccd vccd _655_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[88\]_A _356_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_586_ la_data_out_mprj[115] vssd vssd vccd vccd _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y vssd vssd vccd vccd la_data_in_mprj[19]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[12\]_A _611_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[79\]_A _347_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__643__A la_oen_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_440_ mprj_dat_o_core[1] vssd vssd vccd vccd _440_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[15\] _614_/Y mprj_logic_high_inst/HI[217] vssd vssd vccd
+ vccd la_oen_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_13_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_371_ la_oen_mprj[103] vssd vssd vccd vccd _371_/Y sky130_fd_sc_hd__inv_2
XANTENNA__553__A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_638_ la_oen_mprj[39] vssd vssd vccd vccd _638_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_569_ la_data_out_mprj[98] vssd vssd vccd vccd _569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__463__A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__638__A la_oen_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[30\]_A _469_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__373__A la_oen_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__548__A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_423_ mprj_adr_o_core[16] vssd vssd vccd vccd _423_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[21\]_A _460_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[42\] _513_/Y la_buf\[42\]/TE vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__einvp_8
X_354_ la_oen_mprj[86] vssd vssd vccd vccd _354_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[31\]_TE mprj_logic_high_inst/HI[233] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y vssd vssd vccd vccd la_data_in_mprj[86]
+ sky130_fd_sc_hd__inv_8
XFILLER_24_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__458__A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[107\]_TE la_buf\[107\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] mprj_logic_high_inst/HI[361] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[31\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[12\]_A _451_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[6\]_TE mprj_adr_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__368__A la_oen_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[7\]_A _606_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[54\]_TE mprj_logic_high_inst/HI[256] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[82\] _350_/Y mprj_logic_high_inst/HI[284] vssd vssd vccd
+ vccd la_oen_core[82] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[30\] _469_/Y mprj_dat_buf\[30\]/TE vssd vssd vccd vccd mprj_dat_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_406_ mprj_sel_o_core[3] vssd vssd vccd vccd _406_/Y sky130_fd_sc_hd__inv_2
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_337_ la_oen_mprj[69] vssd vssd vccd vccd _337_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] mprj_logic_high_inst/HI[409] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[79\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[92\]_TE la_buf\[92\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high_inst/HI[279] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__651__A la_oen_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_cyc_buf_TE mprj_cyc_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__561__A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y vssd vssd vccd vccd la_data_in_mprj[49]
+ sky130_fd_sc_hd__inv_8
XANTENNA__471__A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] mprj_logic_high_inst/HI[435] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[105\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__646__A la_oen_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[6\]_A _413_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj2_logic_high_inst mprj2_pwrgood/A vccd2 vssd2 mprj2_logic_high
XFILLER_25_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__381__A la_oen_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[115\] _383_/Y mprj_logic_high_inst/HI[317] vssd vssd vccd
+ vccd la_oen_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_28_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[45\] _644_/Y mprj_logic_high_inst/HI[247] vssd vssd vccd
+ vccd la_oen_core[45] sky130_fd_sc_hd__einvp_8
XFILLER_5_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__556__A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[109\] _580_/Y la_buf\[109\]/TE vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_26_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[102] sky130_fd_sc_hd__inv_8
XFILLER_23_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__466__A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[1\] _440_/Y mprj_dat_buf\[1\]/TE vssd vssd vccd vccd mprj_dat_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_22_1400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_logic_high_inst mprj_rstn_buf/TE la_buf\[26\]/TE la_buf\[27\]/TE la_buf\[28\]/TE
+ la_buf\[29\]/TE la_buf\[30\]/TE la_buf\[31\]/TE la_buf\[32\]/TE la_buf\[33\]/TE
+ la_buf\[34\]/TE la_buf\[35\]/TE mprj_adr_buf\[0\]/TE la_buf\[36\]/TE la_buf\[37\]/TE
+ la_buf\[38\]/TE la_buf\[39\]/TE la_buf\[40\]/TE la_buf\[41\]/TE la_buf\[42\]/TE
+ la_buf\[43\]/TE la_buf\[44\]/TE la_buf\[45\]/TE mprj_adr_buf\[1\]/TE la_buf\[46\]/TE
+ la_buf\[47\]/TE la_buf\[48\]/TE la_buf\[49\]/TE la_buf\[50\]/TE la_buf\[51\]/TE
+ la_buf\[52\]/TE la_buf\[53\]/TE la_buf\[54\]/TE la_buf\[55\]/TE mprj_adr_buf\[2\]/TE
+ la_buf\[56\]/TE la_buf\[57\]/TE la_buf\[58\]/TE la_buf\[59\]/TE la_buf\[60\]/TE
+ la_buf\[61\]/TE la_buf\[62\]/TE la_buf\[63\]/TE la_buf\[64\]/TE la_buf\[65\]/TE
+ mprj_adr_buf\[3\]/TE la_buf\[66\]/TE la_buf\[67\]/TE la_buf\[68\]/TE la_buf\[69\]/TE
+ la_buf\[70\]/TE la_buf\[71\]/TE la_buf\[72\]/TE la_buf\[73\]/TE la_buf\[74\]/TE
+ la_buf\[75\]/TE mprj_adr_buf\[4\]/TE la_buf\[76\]/TE la_buf\[77\]/TE la_buf\[78\]/TE
+ la_buf\[79\]/TE la_buf\[80\]/TE la_buf\[81\]/TE la_buf\[82\]/TE la_buf\[83\]/TE
+ la_buf\[84\]/TE la_buf\[85\]/TE mprj_adr_buf\[5\]/TE la_buf\[86\]/TE la_buf\[87\]/TE
+ la_buf\[88\]/TE la_buf\[89\]/TE la_buf\[90\]/TE la_buf\[91\]/TE la_buf\[92\]/TE
+ la_buf\[93\]/TE la_buf\[94\]/TE la_buf\[95\]/TE mprj_adr_buf\[6\]/TE la_buf\[96\]/TE
+ la_buf\[97\]/TE la_buf\[98\]/TE la_buf\[99\]/TE la_buf\[100\]/TE la_buf\[101\]/TE
+ la_buf\[102\]/TE la_buf\[103\]/TE la_buf\[104\]/TE la_buf\[105\]/TE mprj_adr_buf\[7\]/TE
+ la_buf\[106\]/TE la_buf\[107\]/TE la_buf\[108\]/TE la_buf\[109\]/TE la_buf\[110\]/TE
+ la_buf\[111\]/TE la_buf\[112\]/TE la_buf\[113\]/TE la_buf\[114\]/TE la_buf\[115\]/TE
+ mprj_adr_buf\[8\]/TE la_buf\[116\]/TE la_buf\[117\]/TE la_buf\[118\]/TE la_buf\[119\]/TE
+ la_buf\[120\]/TE la_buf\[121\]/TE la_buf\[122\]/TE la_buf\[123\]/TE la_buf\[124\]/TE
+ la_buf\[125\]/TE mprj_adr_buf\[9\]/TE mprj_clk_buf/TE la_buf\[126\]/TE la_buf\[127\]/TE
+ mprj_logic_high_inst/HI[202] mprj_logic_high_inst/HI[203] mprj_logic_high_inst/HI[204]
+ mprj_logic_high_inst/HI[205] mprj_logic_high_inst/HI[206] mprj_logic_high_inst/HI[207]
+ mprj_logic_high_inst/HI[208] mprj_logic_high_inst/HI[209] mprj_adr_buf\[10\]/TE
+ mprj_logic_high_inst/HI[210] mprj_logic_high_inst/HI[211] mprj_logic_high_inst/HI[212]
+ mprj_logic_high_inst/HI[213] mprj_logic_high_inst/HI[214] mprj_logic_high_inst/HI[215]
+ mprj_logic_high_inst/HI[216] mprj_logic_high_inst/HI[217] mprj_logic_high_inst/HI[218]
+ mprj_logic_high_inst/HI[219] mprj_adr_buf\[11\]/TE mprj_logic_high_inst/HI[220]
+ mprj_logic_high_inst/HI[221] mprj_logic_high_inst/HI[222] mprj_logic_high_inst/HI[223]
+ mprj_logic_high_inst/HI[224] mprj_logic_high_inst/HI[225] mprj_logic_high_inst/HI[226]
+ mprj_logic_high_inst/HI[227] mprj_logic_high_inst/HI[228] mprj_logic_high_inst/HI[229]
+ mprj_adr_buf\[12\]/TE mprj_logic_high_inst/HI[230] mprj_logic_high_inst/HI[231]
+ mprj_logic_high_inst/HI[232] mprj_logic_high_inst/HI[233] mprj_logic_high_inst/HI[234]
+ mprj_logic_high_inst/HI[235] mprj_logic_high_inst/HI[236] mprj_logic_high_inst/HI[237]
+ mprj_logic_high_inst/HI[238] mprj_logic_high_inst/HI[239] mprj_adr_buf\[13\]/TE
+ mprj_logic_high_inst/HI[240] mprj_logic_high_inst/HI[241] mprj_logic_high_inst/HI[242]
+ mprj_logic_high_inst/HI[243] mprj_logic_high_inst/HI[244] mprj_logic_high_inst/HI[245]
+ mprj_logic_high_inst/HI[246] mprj_logic_high_inst/HI[247] mprj_logic_high_inst/HI[248]
+ mprj_logic_high_inst/HI[249] mprj_adr_buf\[14\]/TE mprj_logic_high_inst/HI[250]
+ mprj_logic_high_inst/HI[251] mprj_logic_high_inst/HI[252] mprj_logic_high_inst/HI[253]
+ mprj_logic_high_inst/HI[254] mprj_logic_high_inst/HI[255] mprj_logic_high_inst/HI[256]
+ mprj_logic_high_inst/HI[257] mprj_logic_high_inst/HI[258] mprj_logic_high_inst/HI[259]
+ mprj_adr_buf\[15\]/TE mprj_logic_high_inst/HI[260] mprj_logic_high_inst/HI[261]
+ mprj_logic_high_inst/HI[262] mprj_logic_high_inst/HI[263] mprj_logic_high_inst/HI[264]
+ mprj_logic_high_inst/HI[265] mprj_logic_high_inst/HI[266] mprj_logic_high_inst/HI[267]
+ mprj_logic_high_inst/HI[268] mprj_logic_high_inst/HI[269] mprj_adr_buf\[16\]/TE
+ mprj_logic_high_inst/HI[270] mprj_logic_high_inst/HI[271] mprj_logic_high_inst/HI[272]
+ mprj_logic_high_inst/HI[273] mprj_logic_high_inst/HI[274] mprj_logic_high_inst/HI[275]
+ mprj_logic_high_inst/HI[276] mprj_logic_high_inst/HI[277] mprj_logic_high_inst/HI[278]
+ mprj_logic_high_inst/HI[279] mprj_adr_buf\[17\]/TE mprj_logic_high_inst/HI[280]
+ mprj_logic_high_inst/HI[281] mprj_logic_high_inst/HI[282] mprj_logic_high_inst/HI[283]
+ mprj_logic_high_inst/HI[284] mprj_logic_high_inst/HI[285] mprj_logic_high_inst/HI[286]
+ mprj_logic_high_inst/HI[287] mprj_logic_high_inst/HI[288] mprj_logic_high_inst/HI[289]
+ mprj_adr_buf\[18\]/TE mprj_logic_high_inst/HI[290] mprj_logic_high_inst/HI[291]
+ mprj_logic_high_inst/HI[292] mprj_logic_high_inst/HI[293] mprj_logic_high_inst/HI[294]
+ mprj_logic_high_inst/HI[295] mprj_logic_high_inst/HI[296] mprj_logic_high_inst/HI[297]
+ mprj_logic_high_inst/HI[298] mprj_logic_high_inst/HI[299] mprj_adr_buf\[19\]/TE
+ mprj_clk2_buf/TE mprj_logic_high_inst/HI[300] mprj_logic_high_inst/HI[301] mprj_logic_high_inst/HI[302]
+ mprj_logic_high_inst/HI[303] mprj_logic_high_inst/HI[304] mprj_logic_high_inst/HI[305]
+ mprj_logic_high_inst/HI[306] mprj_logic_high_inst/HI[307] mprj_logic_high_inst/HI[308]
+ mprj_logic_high_inst/HI[309] mprj_adr_buf\[20\]/TE mprj_logic_high_inst/HI[310]
+ mprj_logic_high_inst/HI[311] mprj_logic_high_inst/HI[312] mprj_logic_high_inst/HI[313]
+ mprj_logic_high_inst/HI[314] mprj_logic_high_inst/HI[315] mprj_logic_high_inst/HI[316]
+ mprj_logic_high_inst/HI[317] mprj_logic_high_inst/HI[318] mprj_logic_high_inst/HI[319]
+ mprj_adr_buf\[21\]/TE mprj_logic_high_inst/HI[320] mprj_logic_high_inst/HI[321]
+ mprj_logic_high_inst/HI[322] mprj_logic_high_inst/HI[323] mprj_logic_high_inst/HI[324]
+ mprj_logic_high_inst/HI[325] mprj_logic_high_inst/HI[326] mprj_logic_high_inst/HI[327]
+ mprj_logic_high_inst/HI[328] mprj_logic_high_inst/HI[329] mprj_adr_buf\[22\]/TE
+ user_to_mprj_in_gates\[0\]/B user_to_mprj_in_gates\[1\]/B user_to_mprj_in_gates\[2\]/B
+ user_to_mprj_in_gates\[3\]/B user_to_mprj_in_gates\[4\]/B user_to_mprj_in_gates\[5\]/B
+ user_to_mprj_in_gates\[6\]/B user_to_mprj_in_gates\[7\]/B user_to_mprj_in_gates\[8\]/B
+ user_to_mprj_in_gates\[9\]/B mprj_adr_buf\[23\]/TE mprj_logic_high_inst/HI[340]
+ mprj_logic_high_inst/HI[341] mprj_logic_high_inst/HI[342] mprj_logic_high_inst/HI[343]
+ mprj_logic_high_inst/HI[344] mprj_logic_high_inst/HI[345] mprj_logic_high_inst/HI[346]
+ mprj_logic_high_inst/HI[347] mprj_logic_high_inst/HI[348] mprj_logic_high_inst/HI[349]
+ mprj_adr_buf\[24\]/TE mprj_logic_high_inst/HI[350] mprj_logic_high_inst/HI[351]
+ mprj_logic_high_inst/HI[352] mprj_logic_high_inst/HI[353] mprj_logic_high_inst/HI[354]
+ mprj_logic_high_inst/HI[355] mprj_logic_high_inst/HI[356] mprj_logic_high_inst/HI[357]
+ mprj_logic_high_inst/HI[358] mprj_logic_high_inst/HI[359] mprj_adr_buf\[25\]/TE
+ mprj_logic_high_inst/HI[360] mprj_logic_high_inst/HI[361] mprj_logic_high_inst/HI[362]
+ mprj_logic_high_inst/HI[363] mprj_logic_high_inst/HI[364] mprj_logic_high_inst/HI[365]
+ mprj_logic_high_inst/HI[366] mprj_logic_high_inst/HI[367] mprj_logic_high_inst/HI[368]
+ mprj_logic_high_inst/HI[369] mprj_adr_buf\[26\]/TE mprj_logic_high_inst/HI[370]
+ mprj_logic_high_inst/HI[371] mprj_logic_high_inst/HI[372] mprj_logic_high_inst/HI[373]
+ mprj_logic_high_inst/HI[374] mprj_logic_high_inst/HI[375] mprj_logic_high_inst/HI[376]
+ mprj_logic_high_inst/HI[377] mprj_logic_high_inst/HI[378] mprj_logic_high_inst/HI[379]
+ mprj_adr_buf\[27\]/TE mprj_logic_high_inst/HI[380] mprj_logic_high_inst/HI[381]
+ mprj_logic_high_inst/HI[382] mprj_logic_high_inst/HI[383] mprj_logic_high_inst/HI[384]
+ mprj_logic_high_inst/HI[385] mprj_logic_high_inst/HI[386] mprj_logic_high_inst/HI[387]
+ mprj_logic_high_inst/HI[388] mprj_logic_high_inst/HI[389] mprj_adr_buf\[28\]/TE
+ mprj_logic_high_inst/HI[390] mprj_logic_high_inst/HI[391] mprj_logic_high_inst/HI[392]
+ mprj_logic_high_inst/HI[393] mprj_logic_high_inst/HI[394] mprj_logic_high_inst/HI[395]
+ mprj_logic_high_inst/HI[396] mprj_logic_high_inst/HI[397] mprj_logic_high_inst/HI[398]
+ mprj_logic_high_inst/HI[399] mprj_adr_buf\[29\]/TE mprj_cyc_buf/TE mprj_logic_high_inst/HI[400]
+ mprj_logic_high_inst/HI[401] mprj_logic_high_inst/HI[402] mprj_logic_high_inst/HI[403]
+ mprj_logic_high_inst/HI[404] mprj_logic_high_inst/HI[405] mprj_logic_high_inst/HI[406]
+ mprj_logic_high_inst/HI[407] mprj_logic_high_inst/HI[408] mprj_logic_high_inst/HI[409]
+ mprj_adr_buf\[30\]/TE mprj_logic_high_inst/HI[410] mprj_logic_high_inst/HI[411]
+ mprj_logic_high_inst/HI[412] mprj_logic_high_inst/HI[413] mprj_logic_high_inst/HI[414]
+ mprj_logic_high_inst/HI[415] mprj_logic_high_inst/HI[416] mprj_logic_high_inst/HI[417]
+ mprj_logic_high_inst/HI[418] mprj_logic_high_inst/HI[419] mprj_adr_buf\[31\]/TE
+ mprj_logic_high_inst/HI[420] mprj_logic_high_inst/HI[421] mprj_logic_high_inst/HI[422]
+ mprj_logic_high_inst/HI[423] mprj_logic_high_inst/HI[424] mprj_logic_high_inst/HI[425]
+ mprj_logic_high_inst/HI[426] mprj_logic_high_inst/HI[427] mprj_logic_high_inst/HI[428]
+ mprj_logic_high_inst/HI[429] mprj_dat_buf\[0\]/TE mprj_logic_high_inst/HI[430] mprj_logic_high_inst/HI[431]
+ mprj_logic_high_inst/HI[432] mprj_logic_high_inst/HI[433] mprj_logic_high_inst/HI[434]
+ mprj_logic_high_inst/HI[435] mprj_logic_high_inst/HI[436] mprj_logic_high_inst/HI[437]
+ mprj_logic_high_inst/HI[438] mprj_logic_high_inst/HI[439] mprj_dat_buf\[1\]/TE mprj_logic_high_inst/HI[440]
+ mprj_logic_high_inst/HI[441] mprj_logic_high_inst/HI[442] mprj_logic_high_inst/HI[443]
+ mprj_logic_high_inst/HI[444] mprj_logic_high_inst/HI[445] mprj_logic_high_inst/HI[446]
+ mprj_logic_high_inst/HI[447] mprj_logic_high_inst/HI[448] mprj_logic_high_inst/HI[449]
+ mprj_dat_buf\[2\]/TE mprj_logic_high_inst/HI[450] mprj_logic_high_inst/HI[451] mprj_logic_high_inst/HI[452]
+ mprj_logic_high_inst/HI[453] mprj_logic_high_inst/HI[454] mprj_logic_high_inst/HI[455]
+ mprj_logic_high_inst/HI[456] mprj_logic_high_inst/HI[457] mprj_pwrgood/A mprj_dat_buf\[3\]/TE
+ mprj_dat_buf\[4\]/TE mprj_dat_buf\[5\]/TE mprj_dat_buf\[6\]/TE mprj_dat_buf\[7\]/TE
+ mprj_stb_buf/TE mprj_dat_buf\[8\]/TE mprj_dat_buf\[9\]/TE mprj_dat_buf\[10\]/TE
+ mprj_dat_buf\[11\]/TE mprj_dat_buf\[12\]/TE mprj_dat_buf\[13\]/TE mprj_dat_buf\[14\]/TE
+ mprj_dat_buf\[15\]/TE mprj_dat_buf\[16\]/TE mprj_dat_buf\[17\]/TE mprj_we_buf/TE
+ mprj_dat_buf\[18\]/TE mprj_dat_buf\[19\]/TE mprj_dat_buf\[20\]/TE mprj_dat_buf\[21\]/TE
+ mprj_dat_buf\[22\]/TE mprj_dat_buf\[23\]/TE mprj_dat_buf\[24\]/TE mprj_dat_buf\[25\]/TE
+ mprj_dat_buf\[26\]/TE mprj_dat_buf\[27\]/TE mprj_sel_buf\[0\]/TE mprj_dat_buf\[28\]/TE
+ mprj_dat_buf\[29\]/TE mprj_dat_buf\[30\]/TE mprj_dat_buf\[31\]/TE la_buf\[0\]/TE
+ la_buf\[1\]/TE la_buf\[2\]/TE la_buf\[3\]/TE la_buf\[4\]/TE la_buf\[5\]/TE mprj_sel_buf\[1\]/TE
+ la_buf\[6\]/TE la_buf\[7\]/TE la_buf\[8\]/TE la_buf\[9\]/TE la_buf\[10\]/TE la_buf\[11\]/TE
+ la_buf\[12\]/TE la_buf\[13\]/TE la_buf\[14\]/TE la_buf\[15\]/TE mprj_sel_buf\[2\]/TE
+ la_buf\[16\]/TE la_buf\[17\]/TE la_buf\[18\]/TE la_buf\[19\]/TE la_buf\[20\]/TE
+ la_buf\[21\]/TE la_buf\[22\]/TE la_buf\[23\]/TE la_buf\[24\]/TE la_buf\[25\]/TE
+ mprj_sel_buf\[3\]/TE vccd1 vssd1 mprj_logic_high
XFILLER_27_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__376__A la_oen_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_654_ la_oen_mprj[55] vssd vssd vccd vccd _654_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[72\] _543_/Y la_buf\[72\]/TE vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__einvp_8
X_585_ la_data_out_mprj[114] vssd vssd vccd vccd _585_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] mprj_logic_high_inst/HI[391] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[61\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[26\]_TE la_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[6\]_B user_to_mprj_in_gates\[6\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_370_ la_oen_mprj[102] vssd vssd vccd vccd _370_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_637_ la_oen_mprj[38] vssd vssd vccd vccd _637_/Y sky130_fd_sc_hd__inv_2
X_568_ la_data_out_mprj[97] vssd vssd vccd vccd _568_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y vssd vssd vccd vccd la_data_in_mprj[31]
+ sky130_fd_sc_hd__inv_8
X_499_ la_data_out_mprj[28] vssd vssd vccd vccd _499_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[49\]_TE la_buf\[49\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__654__A la_oen_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_422_ mprj_adr_o_core[15] vssd vssd vccd vccd _422_/Y sky130_fd_sc_hd__inv_2
XANTENNA__564__A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
X_353_ la_oen_mprj[85] vssd vssd vccd vccd _353_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[35\] _506_/Y la_buf\[35\]/TE vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__einvp_8
XFILLER_6_711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y vssd vssd vccd vccd la_data_in_mprj[79]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__474__A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] mprj_logic_high_inst/HI[354] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[24\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__649__A la_oen_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XPHY_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__384__A la_oen_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[75\] _343_/Y mprj_logic_high_inst/HI[277] vssd vssd vccd
+ vccd la_oen_core[75] sky130_fd_sc_hd__einvp_8
XFILLER_8_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[23\] _462_/Y mprj_dat_buf\[23\]/TE vssd vssd vccd vccd mprj_dat_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__559__A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_405_ mprj_sel_o_core[2] vssd vssd vccd vccd _405_/Y sky130_fd_sc_hd__inv_2
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_336_ la_oen_mprj[68] vssd vssd vccd vccd _336_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__469__A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high_inst/HI[324] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__379__A la_oen_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[21\]_TE mprj_logic_high_inst/HI[223] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xpowergood_check mprj2_vdd_pwrgood/A mprj_vdd_pwrgood/A vccd vssd vdda1 vssd vdda2
+ vssd powergood_check/FILLER_2_300/li_65_797# powergood_check/FILLER_1_260/li_65_797#
+ powergood_check/FILLER_2_115/li_737_n17# powergood_check/FILLER_1_131/li_0_n17#
+ powergood_check/FILLER_1_32/li_161_n17# powergood_check/FILLER_1_8/li_161_n17# powergood_check/FILLER_1_48/li_641_797#
+ powergood_check/FILLER_2_243/li_0_797# powergood_check/FILLER_2_115/li_257_797#
+ powergood_check/FILLER_0_216/li_100_536# powergood_check/FILLER_2_155/li_545_797#
+ powergood_check/FILLER_2_24/li_545_797# powergood_check/FILLER_0_216/li_449_797#
+ powergood_check/mprj2_logic_high_lv/li_514_79# powergood_check/FILLER_1_107/li_353_n17#
+ powergood_check/FILLER_0_264/li_0_797# powergood_check/FILLER_2_227/li_545_n17#
+ powergood_check/mprj2_logic_high_hvl/li_161_797# powergood_check/FILLER_0_32/li_353_797#
+ powergood_check/FILLER_0_176/li_545_797# powergood_check/FILLER_2_187/li_641_n17#
+ powergood_check/mprj2_logic_high_lv/li_161_1611# powergood_check/FILLER_2_16/li_353_n17#
+ powergood_check/FILLER_1_131/li_353_n17# powergood_check/FILLER_1_180/li_161_n17#
+ powergood_check/FILLER_1_24/li_65_n17# powergood_check/FILLER_1_131/li_34_73# powergood_check/FILLER_2_267/li_353_797#
+ powergood_check/FILLER_1_268/li_0_797# powergood_check/FILLER_1_188/li_65_797# powergood_check/FILLER_0_232/li_0_n17#
+ powergood_check/FILLER_0_96/li_65_797# powergood_check/FILLER_2_259/li_161_n17#
+ powergood_check/FILLER_1_156/li_0_797# powergood_check/FILLER_1_268/li_641_n17#
+ powergood_check/FILLER_0_224/li_115_72# powergood_check/FILLER_0_112/li_115_72#
+ powergood_check/FILLER_2_300/li_65_n17# powergood_check/mprj2_logic_high_lv/li_34_216#
+ powergood_check/FILLER_2_171/li_0_797# powergood_check/FILLER_2_32/li_737_797# powergood_check/FILLER_1_48/li_641_n17#
+ powergood_check/FILLER_1_115/li_545_n17# powergood_check/FILLER_2_115/li_257_n17#
+ powergood_check/FILLER_1_260/li_115_72# powergood_check/FILLER_2_243/li_0_n17# powergood_check/FILLER_2_155/li_545_n17#
+ powergood_check/mprj2_logic_high_lv/li_179_1349# powergood_check/FILLER_2_24/li_545_n17#
+ powergood_check/FILLER_1_204/li_100_536# powergood_check/mprj_logic_high_lv/li_545_1611#
+ powergood_check/FILLER_0_264/li_0_n17# powergood_check/FILLER_1_48/li_161_797# powergood_check/mprj2_logic_high_hvl/li_161_n17#
+ powergood_check/FILLER_2_235/li_257_797# powergood_check/FILLER_2_195/li_115_72#
+ powergood_check/FILLER_2_8/li_65_797# powergood_check/FILLER_1_220/li_65_n17# powergood_check/FILLER_0_104/li_641_797#
+ powergood_check/FILLER_2_195/li_353_797# powergood_check/FILLER_0_256/li_257_797#
+ powergood_check/FILLER_1_236/li_545_n17# powergood_check/FILLER_0_160/li_0_n17#
+ powergood_check/FILLER_2_267/li_353_n17# powergood_check/FILLER_1_196/li_641_n17#
+ powergood_check/FILLER_2_187/li_161_n17# powergood_check/FILLER_2_267/li_65_n17#
+ powergood_check/FILLER_2_155/li_65_n17# powergood_check/FILLER_1_16/li_545_n17#
+ powergood_check/FILLER_2_171/li_0_n17# powergood_check/mprj2_logic_high_lv/li_26_452#
+ powergood_check/FILLER_1_188/li_115_72# powergood_check/FILLER_2_32/li_737_n17#
+ powergood_check/mprj_logic_high_lv/m1_0_n23# powergood_check/FILLER_2_219/li_115_72#
+ powergood_check/FILLER_2_107/li_115_72# powergood_check/FILLER_1_268/li_161_n17#
+ powergood_check/FILLER_2_243/li_100_536# powergood_check/FILLER_2_243/li_449_797#
+ powergood_check/FILLER_0_24/li_0_797# powergood_check/FILLER_2_163/li_257_797# powergood_check/FILLER_2_32/li_257_797#
+ powergood_check/FILLER_0_264/li_100_536# powergood_check/FILLER_0_208/li_65_n17#
+ powergood_check/FILLER_1_48/li_161_n17# powergood_check/FILLER_0_264/li_449_797#
+ powergood_check/FILLER_2_235/li_257_n17# powergood_check/FILLER_2_8/li_65_n17# powergood_check/FILLER_0_0/li_545_797#
+ powergood_check/FILLER_1_164/li_545_n17# powergood_check/FILLER_0_184/li_257_797#
+ powergood_check/FILLER_2_195/li_353_n17# powergood_check/FILLER_0_232/li_0_797#
+ powergood_check/FILLER_0_80/li_353_797# powergood_check/mprj2_logic_high_lv/li_1313_1611#
+ powergood_check/FILLER_0_232/li_65_797# powergood_check/FILLER_2_203/li_641_797#
+ powergood_check/FILLER_1_32/li_0_n17# powergood_check/FILLER_0_224/li_641_797# powergood_check/FILLER_0_104/li_161_797#
+ powergood_check/mprj_logic_high_lv/li_1505_797# powergood_check/FILLER_2_195/li_0_797#
+ powergood_check/FILLER_1_62/li_65_797# powergood_check/FILLER_0_88/li_641_797# powergood_check/FILLER_1_196/li_161_n17#
+ powergood_check/FILLER_2_171/li_100_536# powergood_check/FILLER_2_171/li_449_797#
+ powergood_check/FILLER_2_0/li_0_797# powergood_check/FILLER_0_192/li_100_536# powergood_check/FILLER_2_243/li_449_n17#
+ powergood_check/FILLER_2_163/li_257_n17# powergood_check/mprj2_logic_high_lv/li_34_1244#
+ powergood_check/FILLER_0_272/li_115_72# powergood_check/FILLER_0_192/li_449_797#
+ powergood_check/FILLER_0_160/li_115_72# powergood_check/FILLER_1_180/li_0_n17# powergood_check/FILLER_2_32/li_257_n17#
+ powergood_check/FILLER_2_187/li_0_797# powergood_check/FILLER_1_252/li_100_536#
+ powergood_check/FILLER_1_24/li_115_72# powergood_check/FILLER_2_251/li_545_797#
+ powergood_check/FILLER_0_16/li_257_797# powergood_check/FILLER_2_203/li_641_n17#
+ powergood_check/FILLER_0_112/li_353_797# powergood_check/FILLER_1_244/li_257_n17#
+ powergood_check/FILLER_1_32/li_100_536# powergood_check/FILLER_2_8/li_0_797# powergood_check/FILLER_1_8/li_100_536#
+ powergood_check/FILLER_0_104/li_161_n17# powergood_check/FILLER_2_195/li_0_n17#
+ powergood_check/FILLER_1_62/li_65_n17# powergood_check/FILLER_1_204/li_65_797# powergood_check/FILLER_2_115/li_65_797#
+ powergood_check/FILLER_1_24/li_257_n17# powergood_check/FILLER_2_171/li_449_n17#
+ powergood_check/FILLER_0_224/li_161_797# powergood_check/FILLER_0_8/li_353_797#
+ powergood_check/FILLER_0_88/li_161_797# powergood_check/FILLER_2_32/li_0_797# powergood_check/FILLER_2_0/li_0_n17#
+ powergood_check/FILLER_1_140/li_0_797# powergood_check/FILLER_1_220/li_115_72# powergood_check/FILLER_0_24/li_100_536#
+ powergood_check/FILLER_1_180/li_100_536# powergood_check/FILLER_0_208/li_0_797#
+ powergood_check/mprj_logic_high_lv/m1_0_51# powergood_check/FILLER_0_24/li_449_797#
+ powergood_check/FILLER_2_187/li_0_n17# powergood_check/FILLER_2_267/li_115_72# powergood_check/FILLER_0_256/li_65_n17#
+ powergood_check/FILLER_0_96/li_115_72# powergood_check/FILLER_2_259/li_100_536#
+ powergood_check/FILLER_2_155/li_115_72# powergood_check/FILLER_1_62/li_545_797#
+ powergood_check/FILLER_1_172/li_257_n17# powergood_check/FILLER_2_259/li_449_797#
+ powergood_check/FILLER_2_179/li_257_797# powergood_check/FILLER_0_0/li_0_797# powergood_check/FILLER_2_211/li_353_797#
+ powergood_check/FILLER_1_140/li_641_797# powergood_check/FILLER_2_8/li_0_n17# powergood_check/FILLER_1_32/li_449_n17#
+ powergood_check/FILLER_1_196/li_65_n17# powergood_check/FILLER_1_8/li_449_n17# powergood_check/FILLER_2_227/li_65_n17#
+ powergood_check/FILLER_2_203/li_161_n17# powergood_check/FILLER_2_115/li_65_n17#
+ powergood_check/FILLER_0_232/li_353_797# powergood_check/FILLER_1_212/li_641_n17#
+ powergood_check/FILLER_1_0/li_0_n17# powergood_check/FILLER_0_96/li_353_797# powergood_check/FILLER_0_272/li_641_797#
+ powergood_check/FILLER_1_0/li_641_n17# powergood_check/FILLER_2_219/li_641_797#
+ powergood_check/FILLER_2_0/li_257_797# powergood_check/FILLER_1_62/li_0_797# powergood_check/FILLER_2_32/li_0_n17#
+ powergood_check/FILLER_1_140/li_0_n17# powergood_check/mprj_logic_high_lv/li_449_1611#
+ powergood_check/FILLER_2_8/li_115_72# powergood_check/FILLER_2_8/li_545_797# powergood_check/FILLER_0_208/li_0_n17#
+ powergood_check/FILLER_1_16/li_0_n17# powergood_check/FILLER_0_184/li_65_n17# powergood_check/FILLER_2_187/li_100_536#
+ powergood_check/FILLER_2_187/li_449_797# powergood_check/FILLER_1_62/li_545_n17#
+ powergood_check/FILLER_2_259/li_449_n17# powergood_check/FILLER_0_200/li_257_797#
+ powergood_check/mprj_logic_high_lv/li_833_1611# powergood_check/FILLER_2_211/li_353_n17#
+ powergood_check/FILLER_2_179/li_257_n17# powergood_check/FILLER_0_240/li_545_797#
+ powergood_check/FILLER_1_140/li_641_n17# powergood_check/FILLER_2_251/li_641_n17#
+ powergood_check/FILLER_0_160/li_353_797# powergood_check/FILLER_2_107/li_353_797#
+ powergood_check/FILLER_1_268/li_100_536# powergood_check/FILLER_2_16/li_641_797#
+ powergood_check/FILLER_0_272/li_641_n17# powergood_check/FILLER_0_208/li_545_797#
+ powergood_check/FILLER_0_96/li_353_n17# powergood_check/FILLER_2_0/li_257_n17# powergood_check/FILLER_2_219/li_641_n17#
+ powergood_check/FILLER_1_140/li_161_797# powergood_check/mprj2_logic_high_lv/m1_0_51#
+ powergood_check/FILLER_1_48/li_100_536# powergood_check/FILLER_0_168/li_641_797#
+ powergood_check/FILLER_1_48/li_449_797# powergood_check/FILLER_1_212/li_161_n17#
+ powergood_check/mprj2_logic_high_lv/li_1455_797# powergood_check/FILLER_1_32/li_65_n17#
+ powergood_check/FILLER_1_62/li_0_n17# powergood_check/FILLER_0_272/li_161_797# powergood_check/FILLER_1_0/li_161_n17#
+ powergood_check/FILLER_1_220/li_65_797# powergood_check/FILLER_1_164/li_0_797# powergood_check/FILLER_2_8/li_545_n17#
+ powergood_check/FILLER_0_232/li_115_72# powergood_check/FILLER_2_187/li_449_n17#
+ powergood_check/mprj2_logic_high_lv/li_1217_1611# powergood_check/FILLER_1_62/li_115_72#
+ powergood_check/mprj_logic_high_lv/li_34_1244# powergood_check/FILLER_2_115/li_545_797#
+ powergood_check/FILLER_1_196/li_100_536# powergood_check/FILLER_0_224/li_0_797#
+ powergood_check/FILLER_1_107/li_641_n17# powergood_check/mprj_logic_high_lv/li_1121_1611#
+ powergood_check/FILLER_2_107/li_353_n17# powergood_check/FILLER_0_272/li_65_n17#
+ powergood_check/FILLER_0_32/li_641_797# powergood_check/mprj2_logic_high_lv/li_1601_1611#
+ powergood_check/FILLER_2_16/li_641_n17# powergood_check/FILLER_0_16/li_65_797# powergood_check/FILLER_1_188/li_257_n17#
+ powergood_check/mprj_logic_high_lv/li_179_79# powergood_check/FILLER_0_224/li_0_n17#
+ powergood_check/FILLER_1_140/li_161_n17# powergood_check/FILLER_2_251/li_161_n17#
+ powergood_check/FILLER_1_260/li_641_n17# powergood_check/FILLER_2_227/li_353_797#
+ powergood_check/FILLER_1_48/li_449_n17# powergood_check/FILLER_2_267/li_641_797#
+ powergood_check/FILLER_2_16/li_161_797# powergood_check/FILLER_0_248/li_353_797#
+ powergood_check/FILLER_1_228/li_641_n17# powergood_check/FILLER_2_219/li_161_n17#
+ powergood_check/FILLER_2_163/li_65_n17# powergood_check/mprj2_logic_high_lv/li_26_893#
+ powergood_check/FILLER_0_168/li_161_797# powergood_check/FILLER_0_104/li_100_536#
+ powergood_check/FILLER_1_196/li_115_72# powergood_check/FILLER_0_104/li_449_797#
+ powergood_check/FILLER_2_227/li_115_72# powergood_check/FILLER_2_115/li_545_n17#
+ powergood_check/FILLER_2_115/li_115_72# powergood_check/FILLER_0_200/li_65_n17#
+ powergood_check/FILLER_1_268/li_65_n17# powergood_check/mprj2_logic_high_lv/li_384_137#
+ powergood_check/FILLER_1_156/li_65_n17# powergood_check/FILLER_2_235/li_545_797#
+ powergood_check/FILLER_2_155/li_353_797# powergood_check/FILLER_2_24/li_353_797#
+ powergood_check/FILLER_0_216/li_257_797# powergood_check/FILLER_1_107/li_161_n17#
+ powergood_check/FILLER_2_195/li_641_797# powergood_check/FILLER_0_256/li_545_797#
+ powergood_check/FILLER_2_227/li_353_n17# powergood_check/FILLER_0_240/li_65_797#
+ powergood_check/FILLER_0_32/li_161_797# powergood_check/FILLER_1_156/li_641_n17#
+ powergood_check/FILLER_0_176/li_353_797# powergood_check/FILLER_2_267/li_641_n17#
+ powergood_check/FILLER_2_16/li_161_n17# powergood_check/FILLER_1_196/li_0_n17# powergood_check/FILLER_1_268/li_65_797#
+ powergood_check/FILLER_1_228/li_161_n17# powergood_check/FILLER_1_107/li_65_n17#
+ powergood_check/FILLER_2_203/li_100_536# powergood_check/FILLER_2_203/li_449_797#
+ powergood_check/FILLER_2_251/li_0_797# powergood_check/mprj2_logic_high_lv/li_353_1611#
+ powergood_check/FILLER_0_224/li_100_536# powergood_check/FILLER_2_163/li_545_797#
+ powergood_check/FILLER_2_32/li_545_797# powergood_check/FILLER_0_224/li_449_797#
+ powergood_check/FILLER_0_88/li_100_536# powergood_check/FILLER_1_115/li_353_n17#
+ powergood_check/FILLER_0_88/li_449_797# powergood_check/FILLER_2_235/li_545_n17#
+ powergood_check/FILLER_2_155/li_353_n17# powergood_check/FILLER_1_32/li_115_72#
+ powergood_check/FILLER_0_168/li_65_797# powergood_check/FILLER_0_184/li_545_797#
+ powergood_check/FILLER_2_195/li_641_n17# powergood_check/FILLER_2_24/li_353_n17#
+ powergood_check/FILLER_0_80/li_641_797# powergood_check/FILLER_1_260/li_161_n17#
+ powergood_check/FILLER_1_196/li_65_797# powergood_check/FILLER_0_240/li_0_n17# powergood_check/FILLER_1_236/li_0_797#
+ powergood_check/FILLER_1_156/li_161_n17# powergood_check/FILLER_2_267/li_161_n17#
+ powergood_check/mprj_logic_high_lv/li_737_1611# powergood_check/FILLER_2_179/li_0_797#
+ powergood_check/FILLER_1_16/li_353_n17# powergood_check/FILLER_2_203/li_449_n17#
+ powergood_check/FILLER_2_251/li_0_n17# powergood_check/FILLER_0_200/li_0_797# powergood_check/FILLER_2_163/li_545_n17#
+ powergood_check/mprj2_logic_high_hvl/li_43_635# powergood_check/FILLER_2_32/li_545_n17#
+ powergood_check/FILLER_0_216/li_0_797# powergood_check/FILLER_1_212/li_100_536#
+ powergood_check/FILLER_1_0/li_100_536# powergood_check/FILLER_1_260/li_0_797# powergood_check/FILLER_2_243/li_257_797#
+ powergood_check/FILLER_0_16/li_545_797# powergood_check/FILLER_2_163/li_115_72#
+ powergood_check/FILLER_1_300/li_65_n17# powergood_check/FILLER_0_112/li_641_797#
+ powergood_check/FILLER_0_264/li_257_797# powergood_check/FILLER_1_244/li_545_n17#
+ powergood_check/FILLER_0_0/li_353_797# powergood_check/FILLER_0_168/li_0_n17# powergood_check/FILLER_2_195/li_161_n17#
+ powergood_check/mprj2_logic_high_hvl/li_307_57# powergood_check/FILLER_0_80/li_161_797#
+ powergood_check/FILLER_2_235/li_65_n17# powergood_check/FILLER_1_24/li_545_n17#
+ powergood_check/FILLER_1_268/li_115_72# powergood_check/FILLER_0_8/li_641_797# powergood_check/FILLER_1_156/li_115_72#
+ powergood_check/FILLER_2_179/li_0_n17# powergood_check/mprj_logic_high_lv/li_1025_1611#
+ powergood_check/FILLER_0_16/li_115_72# powergood_check/FILLER_1_140/li_100_536#
+ powergood_check/FILLER_0_160/li_0_797# powergood_check/FILLER_2_251/li_100_536#
+ powergood_check/FILLER_1_140/li_449_797# powergood_check/FILLER_1_131/li_257_797#
+ powergood_check/FILLER_1_188/li_0_797# powergood_check/mprj2_logic_high_lv/li_1505_1611#
+ powergood_check/FILLER_0_32/li_0_797# powergood_check/FILLER_2_171/li_257_797# powergood_check/FILLER_0_272/li_100_536#
+ powergood_check/FILLER_1_228/li_65_n17# powergood_check/FILLER_0_216/li_65_n17#
+ powergood_check/FILLER_0_272/li_449_797# powergood_check/FILLER_1_260/li_0_n17#
+ powergood_check/FILLER_2_243/li_257_n17# powergood_check/FILLER_2_219/li_100_536#
+ powergood_check/FILLER_0_192/li_257_797# powergood_check/FILLER_1_0/li_449_n17#
+ powergood_check/FILLER_1_172/li_545_n17# powergood_check/FILLER_2_219/li_449_797#
+ powergood_check/FILLER_2_267/li_0_797# powergood_check/FILLER_2_179/li_545_797#
+ powergood_check/FILLER_2_251/li_353_797# powergood_check/FILLER_2_211/li_641_797#
+ powergood_check/mprj_logic_high_lv/li_384_137# powergood_check/FILLER_0_200/li_65_797#
+ powergood_check/FILLER_1_32/li_737_n17# powergood_check/FILLER_1_107/li_115_72#
+ powergood_check/FILLER_0_232/li_641_797# powergood_check/FILLER_0_112/li_161_797#
+ powergood_check/FILLER_2_16/li_0_797# powergood_check/FILLER_0_96/li_641_797# powergood_check/FILLER_2_0/li_545_797#
+ powergood_check/mprj_logic_high_hvl/li_353_797# powergood_check/FILLER_1_107/li_100_536#
+ powergood_check/FILLER_1_131/li_257_n17# powergood_check/FILLER_1_140/li_449_n17#
+ powergood_check/FILLER_2_251/li_449_n17# powergood_check/FILLER_2_171/li_257_n17#
+ powergood_check/FILLER_0_240/li_115_72# powergood_check/FILLER_0_8/li_161_797# powergood_check/FILLER_1_188/li_0_n17#
+ powergood_check/FILLER_2_16/li_100_536# powergood_check/FILLER_2_16/li_449_797#
+ powergood_check/FILLER_0_272/li_449_n17# powergood_check/FILLER_1_260/li_100_536#
+ powergood_check/FILLER_0_168/li_100_536# powergood_check/FILLER_2_219/li_449_n17#
+ powergood_check/FILLER_0_168/li_449_797# powergood_check/FILLER_2_267/li_0_n17#
+ powergood_check/FILLER_0_200/li_545_797# powergood_check/FILLER_0_24/li_257_797#
+ powergood_check/FILLER_2_179/li_545_n17# powergood_check/FILLER_2_211/li_641_n17#
+ powergood_check/FILLER_1_252/li_257_n17# powergood_check/FILLER_1_228/li_100_536#
+ powergood_check/FILLER_0_160/li_641_797# powergood_check/FILLER_2_107/li_641_797#
+ powergood_check/FILLER_1_62/li_353_797# powergood_check/FILLER_1_268/li_737_797#
+ powergood_check/FILLER_2_259/li_257_797# powergood_check/FILLER_2_16/li_0_n17# powergood_check/FILLER_0_96/li_641_n17#
+ powergood_check/FILLER_0_24/li_65_797# powergood_check/FILLER_1_212/li_65_797# powergood_check/FILLER_2_0/li_545_n17#
+ powergood_check/FILLER_1_32/li_257_n17# powergood_check/mprj_logic_high_hvl/li_353_n17#
+ powergood_check/FILLER_1_8/li_257_n17# powergood_check/FILLER_0_0/li_65_797# powergood_check/mprj_logic_high_lv/li_65_797#
+ powergood_check/mprj2_logic_high_lv/li_257_1611# powergood_check/FILLER_1_48/li_737_797#
+ powergood_check/FILLER_0_232/li_161_797# powergood_check/FILLER_0_168/li_115_72#
+ powergood_check/FILLER_1_48/li_0_797# powergood_check/FILLER_0_96/li_161_797# powergood_check/FILLER_0_112/li_0_n17#
+ powergood_check/FILLER_2_171/li_65_n17# powergood_check/FILLER_0_32/li_100_536#
+ powergood_check/mprj2_logic_high_hvl/li_257_797# powergood_check/FILLER_2_16/li_449_n17#
+ powergood_check/FILLER_0_32/li_449_797# powergood_check/mprj2_logic_high_lv/li_641_1611#
+ powergood_check/FILLER_2_8/li_353_797# powergood_check/FILLER_0_264/li_65_n17# powergood_check/FILLER_2_235/li_115_72#
+ powergood_check/FILLER_1_156/li_100_536# powergood_check/FILLER_1_180/li_257_n17#
+ powergood_check/FILLER_1_204/li_161_n17# powergood_check/FILLER_2_267/li_100_536#
+ powergood_check/FILLER_2_267/li_449_797# powergood_check/FILLER_1_204/li_0_797#
+ powergood_check/FILLER_2_187/li_257_797# powergood_check/mprj_logic_high_hvl/li_43_635#
+ powergood_check/FILLER_0_232/li_65_n17# powergood_check/FILLER_2_107/li_641_n17#
+ powergood_check/FILLER_1_268/li_737_n17# powergood_check/FILLER_1_62/li_353_n17#
+ powergood_check/FILLER_1_164/li_65_n17# powergood_check/FILLER_2_259/li_257_n17#
+ powergood_check/FILLER_1_188/li_545_n17# powergood_check/FILLER_2_211/li_161_n17#
+ powergood_check/FILLER_0_240/li_353_797# powergood_check/FILLER_1_220/li_641_n17#
+ powergood_check/FILLER_0_160/li_161_797# powergood_check/FILLER_2_227/li_641_797#
+ powergood_check/FILLER_2_107/li_161_797# powergood_check/FILLER_1_48/li_737_n17#
+ powergood_check/FILLER_1_228/li_115_72# powergood_check/FILLER_0_208/li_353_797#
+ powergood_check/mprj_logic_high_hvl/li_307_57# powergood_check/FILLER_0_248/li_641_797#
+ powergood_check/FILLER_1_48/li_0_n17# powergood_check/FILLER_1_48/li_257_797# powergood_check/mprj2_logic_high_hvl/li_257_n17#
+ powergood_check/FILLER_2_195/li_100_536# powergood_check/mprj2_logic_high_lv/li_384_1039#
+ powergood_check/FILLER_0_112/li_0_797# powergood_check/FILLER_2_195/li_449_797#
+ powergood_check/FILLER_2_8/li_353_n17# powergood_check/FILLER_1_115/li_65_n17# powergood_check/FILLER_0_160/li_65_n17#
+ powergood_check/FILLER_2_267/li_449_n17# powergood_check/FILLER_1_204/li_0_n17#
+ powergood_check/FILLER_2_187/li_257_n17# powergood_check/FILLER_2_107/li_0_797#
+ powergood_check/FILLER_2_115/li_353_797# powergood_check/mprj_logic_high_lv/li_826_79#
+ powergood_check/FILLER_2_155/li_641_797# powergood_check/FILLER_0_216/li_545_797#
+ powergood_check/FILLER_0_176/li_65_797# powergood_check/FILLER_2_24/li_641_797#
+ powergood_check/FILLER_2_227/li_641_n17# powergood_check/FILLER_2_107/li_161_n17#
+ powergood_check/FILLER_1_268/li_257_n17# powergood_check/FILLER_0_176/li_641_797#
+ powergood_check/mprj2_logic_high_lv/li_1409_1611# powergood_check/FILLER_1_220/li_161_n17#
+ powergood_check/FILLER_1_228/li_65_797# powergood_check/FILLER_1_48/li_257_n17#
+ powergood_check/FILLER_0_200/li_115_72# powergood_check/mprj_logic_high_lv/li_1313_1611#
+ powergood_check/FILLER_0_248/li_161_797# powergood_check/FILLER_0_80/li_100_536#
+ powergood_check/FILLER_2_195/li_449_n17# powergood_check/FILLER_0_80/li_449_797#
+ powergood_check/FILLER_2_107/li_0_n17# powergood_check/FILLER_0_104/li_257_797#
+ powergood_check/FILLER_1_115/li_641_n17# powergood_check/mprj2_logic_high_lv/li_506_1123#
+ powergood_check/FILLER_0_96/li_0_797# powergood_check/FILLER_2_155/li_0_797# powergood_check/FILLER_2_115/li_353_n17#
+ powergood_check/mprj_logic_high_lv/li_514_79# powergood_check/FILLER_2_155/li_641_n17#
+ powergood_check/FILLER_2_24/li_641_n17# powergood_check/FILLER_1_196/li_257_n17#
+ powergood_check/FILLER_2_171/li_115_72# powergood_check/FILLER_2_235/li_353_797#
+ powergood_check/FILLER_1_156/li_65_797# powergood_check/FILLER_2_24/li_161_797#
+ powergood_check/FILLER_0_256/li_353_797# powergood_check/FILLER_1_236/li_641_n17#
+ powergood_check/FILLER_2_243/li_65_n17# powergood_check/FILLER_2_227/li_161_n17#
+ powergood_check/FILLER_0_176/li_161_797# powergood_check/FILLER_2_16/li_65_797#
+ powergood_check/FILLER_0_112/li_100_536# powergood_check/mprj_logic_high_lv/li_34_216#
+ powergood_check/FILLER_1_16/li_641_n17# powergood_check/FILLER_0_112/li_449_797#
+ powergood_check/FILLER_1_164/li_115_72# powergood_check/FILLER_0_24/li_115_72# powergood_check/FILLER_0_0/li_115_72#
+ powergood_check/FILLER_2_155/li_0_n17# powergood_check/FILLER_2_203/li_257_797#
+ powergood_check/mprj2_logic_high_lv/li_0_1611# powergood_check/FILLER_1_236/li_65_n17#
+ powergood_check/FILLER_2_243/li_545_797# powergood_check/FILLER_0_8/li_100_536#
+ powergood_check/FILLER_2_163/li_353_797# powergood_check/FILLER_2_32/li_353_797#
+ powergood_check/FILLER_0_224/li_257_797# powergood_check/FILLER_1_204/li_545_n17#
+ powergood_check/FILLER_0_8/li_449_797# powergood_check/FILLER_1_115/li_161_n17#
+ powergood_check/FILLER_0_264/li_545_797# powergood_check/FILLER_0_88/li_257_797#
+ powergood_check/FILLER_2_235/li_353_n17# powergood_check/FILLER_2_155/li_161_n17#
+ powergood_check/FILLER_1_164/li_641_n17# powergood_check/FILLER_0_184/li_353_797#
+ powergood_check/FILLER_2_24/li_161_n17# powergood_check/FILLER_0_0/li_641_797# powergood_check/FILLER_1_115/li_115_72#
+ powergood_check/mprj2_logic_high_lv/li_545_1611# powergood_check/FILLER_2_16/li_65_n17#
+ powergood_check/FILLER_2_300/li_0_797# powergood_check/FILLER_1_236/li_161_n17#
+ powergood_check/mprj_logic_high_lv/li_26_452# powergood_check/FILLER_2_211/li_100_536#
+ powergood_check/FILLER_2_211/li_449_797# powergood_check/FILLER_1_140/li_737_797#
+ powergood_check/FILLER_0_232/li_100_536# powergood_check/FILLER_2_171/li_545_797#
+ powergood_check/FILLER_1_220/li_0_n17# powergood_check/FILLER_1_16/li_161_n17# powergood_check/FILLER_0_96/li_100_536#
+ powergood_check/FILLER_2_203/li_257_n17# powergood_check/FILLER_0_272/li_737_797#
+ powergood_check/FILLER_0_232/li_449_797# powergood_check/FILLER_0_96/li_449_797#
+ powergood_check/FILLER_2_243/li_545_n17# powergood_check/FILLER_0_248/li_65_797#
+ powergood_check/FILLER_0_192/li_545_797# powergood_check/FILLER_1_8/li_0_n17# powergood_check/FILLER_2_227/li_0_797#
+ powergood_check/FILLER_2_163/li_353_n17# powergood_check/FILLER_2_32/li_353_n17#
+ powergood_check/FILLER_2_251/li_641_797# powergood_check/FILLER_0_16/li_353_797#
+ powergood_check/mprj_logic_high_lv/li_929_1611# powergood_check/mprj2_logic_high_lv/li_756_683#
+ powergood_check/FILLER_0_248/li_0_n17# powergood_check/FILLER_0_32/li_65_797# powergood_check/FILLER_1_164/li_161_n17#
+ powergood_check/FILLER_1_252/li_0_797# powergood_check/FILLER_0_0/li_161_797# powergood_check/FILLER_1_24/li_353_n17#
+ powergood_check/FILLER_0_160/li_100_536# powergood_check/FILLER_0_176/li_115_72#
+ powergood_check/FILLER_2_211/li_449_n17# powergood_check/FILLER_1_140/li_737_n17#
+ powergood_check/FILLER_0_160/li_449_797# powergood_check/FILLER_2_259/li_0_n17#
+ powergood_check/FILLER_2_107/li_100_536# powergood_check/FILLER_2_171/li_545_n17#
+ powergood_check/FILLER_2_107/li_449_797# powergood_check/FILLER_2_24/li_0_797# powergood_check/FILLER_0_272/li_737_n17#
+ powergood_check/FILLER_1_220/li_100_536# powergood_check/FILLER_0_96/li_449_n17#
+ powergood_check/FILLER_2_227/li_0_n17# powergood_check/FILLER_1_140/li_257_797#
+ powergood_check/mprj2_logic_high_lv/li_1505_797# powergood_check/FILLER_0_24/li_545_797#
+ powergood_check/FILLER_2_243/li_115_72# powergood_check/FILLER_1_212/li_257_n17#
+ powergood_check/FILLER_0_272/li_257_797# powergood_check/FILLER_1_252/li_545_n17#
+ powergood_check/FILLER_1_62/li_641_797# powergood_check/FILLER_1_0/li_257_n17# powergood_check/FILLER_0_176/li_0_n17#
+ powergood_check/FILLER_2_219/li_257_797# powergood_check/mprj2_logic_high_hvl/li_0_797#
+ powergood_check/FILLER_1_172/li_65_n17# powergood_check/mprj_logic_high_lv/li_1217_1611#
+ powergood_check/FILLER_2_259/li_545_797# powergood_check/FILLER_2_179/li_353_797#
+ powergood_check/FILLER_2_203/li_65_n17# powergood_check/FILLER_1_252/li_0_n17# powergood_check/FILLER_1_32/li_545_n17#
+ powergood_check/FILLER_0_192/li_0_797# powergood_check/FILLER_1_8/li_545_n17# powergood_check/FILLER_1_236/li_115_72#
+ powergood_check/FILLER_2_0/li_353_797# powergood_check/FILLER_1_115/li_0_n17# powergood_check/FILLER_2_300/li_0_n17#
+ powergood_check/mprj_logic_high_hvl/li_161_797# powergood_check/FILLER_2_107/li_449_n17#
+ powergood_check/mprj_logic_high_lv/li_161_1611# powergood_check/FILLER_0_32/li_737_797#
+ powergood_check/FILLER_2_24/li_0_n17# powergood_check/FILLER_0_224/li_65_n17# powergood_check/FILLER_2_8/li_641_797#
+ powergood_check/FILLER_1_268/li_0_n17# powergood_check/FILLER_1_140/li_257_n17#
+ powergood_check/FILLER_2_251/li_257_n17# powergood_check/FILLER_2_227/li_100_536#
+ powergood_check/FILLER_1_180/li_545_n17# powergood_check/FILLER_2_227/li_449_797#
+ powergood_check/FILLER_2_16/li_115_72# powergood_check/FILLER_2_267/li_737_797#
+ powergood_check/FILLER_2_187/li_545_797# powergood_check/FILLER_2_16/li_257_797#
+ powergood_check/FILLER_0_248/li_100_536# powergood_check/FILLER_2_219/li_257_n17#
+ powergood_check/FILLER_0_248/li_449_797# powergood_check/FILLER_1_236/li_0_n17#
+ powergood_check/FILLER_1_62/li_641_n17# powergood_check/FILLER_0_168/li_257_797#
+ powergood_check/FILLER_2_259/li_545_n17# powergood_check/FILLER_0_200/li_353_797#
+ powergood_check/mprj2_logic_high_hvl/li_0_n17# powergood_check/FILLER_2_179/li_353_n17#
+ powergood_check/FILLER_0_240/li_641_797# powergood_check/FILLER_0_184/li_65_797#
+ powergood_check/FILLER_1_62/li_161_797# powergood_check/mprj_logic_high_lv/li_179_1349#
+ powergood_check/FILLER_1_48/li_65_797# powergood_check/FILLER_0_208/li_641_797#
+ powergood_check/FILLER_2_0/li_353_n17# powergood_check/FILLER_1_115/li_100_536#
+ powergood_check/FILLER_0_80/li_65_797# powergood_check/mprj_logic_high_hvl/li_161_n17#
+ powergood_check/FILLER_2_155/li_100_536# powergood_check/FILLER_1_48/li_545_797#
+ powergood_check/FILLER_2_24/li_100_536# powergood_check/FILLER_2_155/li_449_797#
+ powergood_check/FILLER_2_24/li_449_797# powergood_check/FILLER_2_8/li_641_n17# powergood_check/FILLER_1_107/li_257_n17#
+ powergood_check/FILLER_2_227/li_449_n17# powergood_check/FILLER_2_203/li_0_797#
+ powergood_check/FILLER_0_208/li_65_797# powergood_check/FILLER_1_0/li_65_n17# powergood_check/FILLER_1_164/li_0_n17#
+ powergood_check/FILLER_0_176/li_100_536# powergood_check/FILLER_2_267/li_737_n17#
+ powergood_check/FILLER_2_16/li_257_n17# powergood_check/FILLER_0_32/li_257_797#
+ powergood_check/FILLER_0_176/li_449_797# powergood_check/FILLER_2_187/li_545_n17#
+ powergood_check/FILLER_1_156/li_0_n17# powergood_check/FILLER_2_8/li_161_797# powergood_check/FILLER_1_236/li_100_536#
+ powergood_check/FILLER_2_115/li_641_797# powergood_check/mprj2_logic_high_lv/li_449_1611#
+ powergood_check/FILLER_2_235/li_0_797# powergood_check/FILLER_2_267/li_257_797#
+ powergood_check/FILLER_1_228/li_257_n17# powergood_check/FILLER_1_268/li_545_n17#
+ powergood_check/FILLER_1_16/li_100_536# powergood_check/FILLER_1_48/li_65_n17# powergood_check/FILLER_1_62/li_161_n17#
+ powergood_check/FILLER_0_192/li_0_n17# powergood_check/FILLER_1_180/li_0_797# powergood_check/FILLER_0_240/li_161_797#
+ powergood_check/mprj_logic_high_lv/m1_0_689# powergood_check/mprj_logic_high_lv/li_756_683#
+ powergood_check/mprj2_logic_high_lv/li_833_1611# powergood_check/mprj2_logic_high_hvl/li_65_797#
+ powergood_check/FILLER_0_248/li_115_72# powergood_check/FILLER_1_48/li_545_n17#
+ powergood_check/FILLER_0_80/li_65_n17# powergood_check/FILLER_1_115/li_449_n17#
+ powergood_check/FILLER_2_251/li_65_n17# powergood_check/FILLER_0_208/li_161_797#
+ powergood_check/FILLER_2_155/li_449_n17# powergood_check/FILLER_2_24/li_65_797#
+ powergood_check/FILLER_2_203/li_0_n17# powergood_check/FILLER_2_24/li_449_n17# powergood_check/FILLER_0_88/li_0_797#
+ powergood_check/FILLER_1_172/li_115_72# powergood_check/FILLER_0_32/li_115_72# powergood_check/FILLER_1_164/li_100_536#
+ powergood_check/FILLER_2_203/li_115_72# powergood_check/FILLER_0_104/li_545_797#
+ powergood_check/FILLER_2_195/li_257_797# powergood_check/FILLER_2_8/li_161_n17#
+ powergood_check/FILLER_2_235/li_0_n17# powergood_check/FILLER_2_115/li_641_n17#
+ powergood_check/FILLER_1_244/li_65_n17# powergood_check/FILLER_0_240/li_65_n17#
+ powergood_check/FILLER_1_156/li_257_n17# powergood_check/FILLER_2_267/li_257_n17#
+ powergood_check/FILLER_0_8/li_65_797# powergood_check/FILLER_1_196/li_545_n17# powergood_check/mprj2_logic_high_lv/li_161_797#
+ powergood_check/FILLER_1_16/li_449_n17# powergood_check/FILLER_2_235/li_641_797#
+ powergood_check/FILLER_2_115/li_161_797# powergood_check/FILLER_2_179/li_65_n17#
+ powergood_check/mprj2_logic_high_hvl/li_65_n17# powergood_check/FILLER_0_216/li_353_797#
+ powergood_check/FILLER_0_256/li_641_797# powergood_check/FILLER_2_24/li_65_n17#
+ powergood_check/FILLER_1_300/li_161_n17# powergood_check/mprj_logic_high_lv/li_26_893#
+ powergood_check/FILLER_0_112/li_737_797# powergood_check/FILLER_0_0/li_100_536#
+ powergood_check/FILLER_0_168/li_65_n17# powergood_check/FILLER_0_0/li_449_797# powergood_check/FILLER_2_195/li_257_n17#
+ powergood_check/FILLER_0_80/li_257_797# powergood_check/FILLER_2_203/li_545_797#
+ powergood_check/FILLER_2_163/li_641_797# powergood_check/FILLER_0_256/li_65_797#
+ powergood_check/mprj2_logic_high_lv/li_65_1611# powergood_check/FILLER_2_32/li_641_797#
+ powergood_check/FILLER_0_224/li_545_797# powergood_check/FILLER_0_88/li_545_797#
+ powergood_check/FILLER_2_235/li_641_n17# powergood_check/FILLER_2_115/li_161_n17#
+ powergood_check/FILLER_0_184/li_641_797# powergood_check/mprj_logic_high_lv/li_1505_1611#
+ powergood_check/FILLER_1_260/li_257_n17# powergood_check/FILLER_1_0/li_115_72# powergood_check/FILLER_1_236/li_65_797#
+ powergood_check/FILLER_1_212/li_0_797# powergood_check/FILLER_0_256/li_161_797#
+ powergood_check/FILLER_0_184/li_115_72# powergood_check/FILLER_2_219/li_0_797# powergood_check/FILLER_1_48/li_115_72#
+ powergood_check/FILLER_0_112/li_257_797# powergood_check/FILLER_2_203/li_545_n17#
+ powergood_check/FILLER_0_240/li_0_797# powergood_check/FILLER_0_104/li_0_797# powergood_check/FILLER_2_163/li_641_n17#
+ powergood_check/FILLER_2_32/li_641_n17# powergood_check/FILLER_2_251/li_115_72#
+ powergood_check/FILLER_1_131/li_65_797# powergood_check/FILLER_0_80/li_115_72# powergood_check/mprj2_logic_high_lv/m1_0_689#
+ powergood_check/FILLER_2_243/li_353_797# powergood_check/FILLER_0_16/li_641_797#
+ powergood_check/FILLER_1_164/li_65_797# powergood_check/FILLER_0_8/li_257_797# powergood_check/FILLER_1_180/li_65_n17#
+ powergood_check/FILLER_2_32/li_161_797# powergood_check/FILLER_0_264/li_353_797#
+ powergood_check/FILLER_1_244/li_641_n17# powergood_check/FILLER_0_208/li_115_72#
+ powergood_check/FILLER_2_235/li_161_n17# powergood_check/FILLER_0_184/li_161_797#
+ powergood_check/FILLER_2_211/li_65_n17# powergood_check/FILLER_0_272/li_0_797# powergood_check/mprj_logic_high_lv/li_0_797#
+ powergood_check/mprj_logic_high_hvl/li_65_797# powergood_check/FILLER_1_244/li_115_72#
+ powergood_check/FILLER_1_24/li_641_n17# powergood_check/FILLER_2_219/li_0_n17# powergood_check/FILLER_0_168/li_0_797#
+ powergood_check/FILLER_1_62/li_100_536# powergood_check/FILLER_2_115/li_0_797# powergood_check/FILLER_1_62/li_449_797#
+ powergood_check/FILLER_0_104/li_0_n17# powergood_check/FILLER_1_228/li_0_797# powergood_check/FILLER_2_179/li_115_72#
+ powergood_check/FILLER_2_211/li_257_797# powergood_check/FILLER_1_140/li_545_797#
+ powergood_check/FILLER_1_131/li_65_n17# powergood_check/mprj_logic_high_lv/li_1455_797#
+ powergood_check/FILLER_2_171/li_353_797# powergood_check/FILLER_1_212/li_545_n17#
+ powergood_check/mprj2_logic_high_lv/li_737_1611# powergood_check/FILLER_2_24/li_115_72#
+ powergood_check/FILLER_0_232/li_257_797# powergood_check/FILLER_0_96/li_257_797#
+ powergood_check/FILLER_2_243/li_353_n17# powergood_check/FILLER_0_272/li_545_797#
+ powergood_check/FILLER_0_192/li_353_797# powergood_check/FILLER_1_0/li_545_n17#
+ powergood_check/FILLER_1_172/li_641_n17# powergood_check/FILLER_2_219/li_545_797#
+ powergood_check/FILLER_2_163/li_161_n17# powergood_check/FILLER_2_32/li_161_n17#
+ powergood_check/mprj_logic_high_lv/li_161_797# powergood_check/FILLER_2_179/li_641_797#
+ powergood_check/FILLER_0_192/li_65_797# powergood_check/FILLER_2_251/li_449_797#
+ powergood_check/FILLER_2_8/li_100_536# powergood_check/FILLER_1_300/li_0_n17# powergood_check/FILLER_0_16/li_161_797#
+ powergood_check/FILLER_2_8/li_449_797# powergood_check/FILLER_1_244/li_161_n17#
+ powergood_check/mprj_logic_high_hvl/li_65_n17# powergood_check/FILLER_2_0/li_641_797#
+ powergood_check/FILLER_0_8/li_115_72# powergood_check/FILLER_0_80/li_0_797# powergood_check/FILLER_2_115/li_0_n17#
+ powergood_check/FILLER_1_62/li_449_n17# powergood_check/FILLER_0_240/li_100_536#
+ powergood_check/FILLER_1_228/li_0_n17# powergood_check/FILLER_1_24/li_161_n17# powergood_check/FILLER_2_211/li_257_n17#
+ powergood_check/FILLER_0_240/li_449_797# powergood_check/FILLER_1_140/li_545_n17#
+ powergood_check/FILLER_0_160/li_257_797# powergood_check/FILLER_2_251/li_545_n17#
+ powergood_check/FILLER_2_171/li_353_n17# powergood_check/FILLER_2_107/li_257_797#
+ powergood_check/FILLER_0_216/li_65_797# powergood_check/FILLER_0_208/li_100_536#
+ powergood_check/FILLER_0_104/li_65_797# powergood_check/FILLER_2_211/li_0_797# powergood_check/FILLER_2_16/li_545_797#
+ powergood_check/FILLER_0_272/li_545_n17# powergood_check/FILLER_0_208/li_449_797#
+ powergood_check/FILLER_2_219/li_545_n17# powergood_check/FILLER_0_176/li_0_797#
+ powergood_check/FILLER_0_200/li_641_797# powergood_check/FILLER_0_24/li_353_797#
+ powergood_check/mprj2_logic_high_lv/li_179_79# powergood_check/FILLER_0_168/li_545_797#
+ powergood_check/FILLER_1_252/li_65_797# powergood_check/FILLER_2_179/li_641_n17#
+ powergood_check/mprj_logic_high_lv/li_65_1611# powergood_check/FILLER_1_140/li_65_797#
+ powergood_check/FILLER_0_256/li_0_n17# powergood_check/FILLER_2_8/li_449_n17# powergood_check/FILLER_1_172/li_161_n17#
+ powergood_check/FILLER_2_0/li_65_797# powergood_check/FILLER_2_259/li_353_797# powergood_check/FILLER_1_180/li_65_797#
+ powergood_check/FILLER_0_80/li_0_n17# powergood_check/FILLER_2_0/li_641_n17# powergood_check/FILLER_0_256/li_115_72#
+ powergood_check/FILLER_1_32/li_353_n17# powergood_check/FILLER_1_8/li_353_n17# powergood_check/FILLER_2_115/li_100_536#
+ powergood_check/FILLER_2_115/li_449_797# powergood_check/FILLER_2_32/li_65_797#
+ powergood_check/FILLER_2_163/li_0_797# powergood_check/FILLER_2_0/li_161_797# powergood_check/FILLER_0_112/li_65_n17#
+ powergood_check/FILLER_2_107/li_257_n17# powergood_check/FILLER_1_180/li_115_72#
+ powergood_check/mprj2_logic_high_hvl/li_353_797# powergood_check/FILLER_0_32/li_545_797#
+ powergood_check/FILLER_0_104/li_65_n17# powergood_check/FILLER_0_184/li_0_797# powergood_check/mprj_logic_high_lv/li_1409_1611#
+ powergood_check/FILLER_2_211/li_115_72# powergood_check/FILLER_2_211/li_0_n17# powergood_check/FILLER_2_16/li_545_n17#
+ powergood_check/FILLER_1_220/li_257_n17# powergood_check/FILLER_1_260/li_545_n17#
+ powergood_check/FILLER_1_244/li_0_797# powergood_check/FILLER_0_184/li_0_n17# powergood_check/FILLER_1_204/li_257_n17#
+ powergood_check/FILLER_2_227/li_257_797# powergood_check/FILLER_1_252/li_65_n17#
+ powergood_check/FILLER_1_140/li_65_n17# powergood_check/FILLER_2_267/li_545_797#
+ powergood_check/FILLER_2_187/li_353_797# powergood_check/mprj2_logic_high_lv/li_0_797#
+ powergood_check/FILLER_0_248/li_257_797# powergood_check/FILLER_1_228/li_545_n17#
+ powergood_check/mprj_logic_high_lv/li_353_1611# powergood_check/FILLER_2_259/li_353_n17#
+ powergood_check/FILLER_2_0/li_65_n17# powergood_check/FILLER_0_200/li_161_797# powergood_check/FILLER_1_188/li_641_n17#
+ powergood_check/FILLER_2_179/li_161_n17# powergood_check/FILLER_2_187/li_65_n17#
+ powergood_check/FILLER_1_204/li_115_72# powergood_check/FILLER_1_115/li_737_n17#
+ powergood_check/FILLER_2_115/li_449_n17# powergood_check/FILLER_2_163/li_0_n17#
+ powergood_check/FILLER_2_32/li_65_n17# powergood_check/FILLER_2_300/li_161_797#
+ powergood_check/FILLER_2_0/li_161_n17# powergood_check/FILLER_1_107/li_0_n17# powergood_check/FILLER_2_235/li_100_536#
+ powergood_check/FILLER_1_48/li_353_797# powergood_check/mprj2_logic_high_hvl/li_353_n17#
+ powergood_check/FILLER_2_235/li_449_797# powergood_check/FILLER_1_172/li_0_797#
+ powergood_check/FILLER_2_155/li_257_797# powergood_check/FILLER_2_24/li_257_797#
+ powergood_check/FILLER_0_256/li_100_536# powergood_check/FILLER_2_227/li_257_n17#
+ powergood_check/FILLER_2_195/li_545_797# powergood_check/FILLER_0_256/li_449_797#
+ powergood_check/FILLER_1_244/li_0_n17# powergood_check/FILLER_1_156/li_545_n17#
+ powergood_check/FILLER_2_267/li_545_n17# powergood_check/FILLER_0_176/li_257_797#
+ powergood_check/FILLER_2_187/li_353_n17# powergood_check/FILLER_0_96/li_0_n17# powergood_check/FILLER_0_264/li_65_797#
+ powergood_check/FILLER_1_24/li_0_n17# powergood_check/FILLER_0_216/li_641_797# powergood_check/mprj2_logic_high_lv/li_1121_1611#
+ powergood_check/FILLER_0_272/li_0_n17# powergood_check/FILLER_1_188/li_161_n17#
+ powergood_check/FILLER_2_300/li_161_n17# powergood_check/FILLER_2_163/li_100_536#
+ powergood_check/FILLER_2_32/li_100_536# powergood_check/FILLER_2_163/li_449_797#
+ powergood_check/FILLER_2_32/li_449_797# powergood_check/FILLER_1_48/li_353_n17#
+ powergood_check/FILLER_1_115/li_257_n17# powergood_check/FILLER_0_184/li_100_536#
+ powergood_check/FILLER_0_192/li_115_72# powergood_check/FILLER_2_235/li_449_n17#
+ powergood_check/FILLER_2_155/li_257_n17# powergood_check/FILLER_0_8/li_0_797# powergood_check/FILLER_1_172/li_0_n17#
+ powergood_check/FILLER_0_184/li_449_797# powergood_check/FILLER_2_195/li_545_n17#
+ powergood_check/FILLER_2_24/li_257_n17# powergood_check/FILLER_0_80/li_545_797#
+ powergood_check/FILLER_1_260/li_65_n17# powergood_check/FILLER_1_244/li_100_536#
+ powergood_check/FILLER_0_104/li_353_797# powergood_check/FILLER_1_236/li_257_n17#
+ powergood_check/FILLER_1_24/li_100_536# powergood_check/FILLER_1_16/li_65_n17# powergood_check/FILLER_0_200/li_0_n17#
+ powergood_check/FILLER_0_88/li_65_797# powergood_check/FILLER_1_131/li_50_537# powergood_check/FILLER_0_216/li_115_72#
+ powergood_check/FILLER_1_16/li_257_n17# powergood_check/FILLER_0_104/li_115_72#
+ powergood_check/FILLER_1_8/li_65_n17# powergood_check/FILLER_2_163/li_449_n17# powergood_check/FILLER_0_216/li_161_797#
+ powergood_check/FILLER_2_32/li_449_n17# powergood_check/FILLER_1_252/li_115_72#
+ powergood_check/FILLER_1_140/li_115_72# powergood_check/FILLER_0_16/li_100_536#
+ powergood_check/FILLER_1_172/li_100_536# powergood_check/FILLER_0_16/li_449_797#
+ powergood_check/FILLER_2_0/li_115_72# powergood_check/FILLER_0_112/li_545_797# powergood_check/FILLER_2_187/li_115_72#
+ powergood_check/FILLER_0_248/li_65_n17# powergood_check/FILLER_1_164/li_257_n17#
+ powergood_check/FILLER_1_212/li_65_n17# powergood_check/FILLER_0_0/li_257_797# powergood_check/FILLER_1_24/li_449_n17#
+ powergood_check/FILLER_2_203/li_353_797# powergood_check/FILLER_2_32/li_115_72#
+ powergood_check/FILLER_2_259/li_65_n17# powergood_check/FILLER_2_243/li_641_797#
+ powergood_check/FILLER_1_204/li_641_n17# powergood_check/FILLER_0_224/li_353_797#
+ powergood_check/FILLER_0_8/li_545_797# powergood_check/FILLER_0_88/li_353_797# powergood_check/FILLER_0_264/li_641_797#
+ powergood_check/FILLER_0_176/li_65_n17# powergood_check/FILLER_1_62/li_737_797#
+ powergood_check/FILLER_2_179/li_100_536# powergood_check/FILLER_2_179/li_449_797#
+ powergood_check/mprj_logic_high_lv/li_257_1611# powergood_check/FILLER_2_211/li_545_797#
+ powergood_check/mprj_logic_high_lv/li_0_1611# powergood_check/FILLER_2_171/li_641_797#
+ powergood_check/FILLER_1_212/li_0_n17# powergood_check/FILLER_2_203/li_353_n17#
+ powergood_check/FILLER_0_232/li_545_797# powergood_check/FILLER_0_224/li_65_797#
+ powergood_check/FILLER_0_96/li_545_797# powergood_check/FILLER_0_112/li_65_797#
+ powergood_check/FILLER_2_243/li_641_n17# powergood_check/FILLER_2_0/li_100_536#
+ powergood_check/FILLER_0_256/li_0_797# powergood_check/FILLER_0_192/li_641_797#
+ powergood_check/FILLER_2_0/li_449_797# powergood_check/mprj_logic_high_hvl/li_257_797#
+ powergood_check/FILLER_0_16/li_0_797# powergood_check/mprj_logic_high_lv/li_641_1611#
+ powergood_check/FILLER_2_259/li_0_797# powergood_check/FILLER_1_244/li_65_797# powergood_check/mprj2_logic_high_lv/li_65_797#
+ powergood_check/FILLER_0_264/li_161_797# powergood_check/FILLER_1_196/li_0_797#
+ powergood_check/FILLER_0_264/li_115_72# powergood_check/FILLER_1_62/li_737_n17#
+ powergood_check/FILLER_0_200/li_100_536# powergood_check/FILLER_0_200/li_449_797#
+ powergood_check/FILLER_1_16/li_115_72# powergood_check/FILLER_2_211/li_545_n17#
+ powergood_check/FILLER_2_179/li_449_n17# powergood_check/FILLER_0_248/li_0_797#
+ powergood_check/FILLER_0_160/li_545_797# powergood_check/FILLER_2_171/li_641_n17#
+ powergood_check/FILLER_2_107/li_545_797# powergood_check/FILLER_1_62/li_257_797#
+ powergood_check/FILLER_1_188/li_100_536# powergood_check/FILLER_0_96/li_545_n17#
+ powergood_check/FILLER_1_131/li_161_797# powergood_check/mprj2_logic_high_lv/li_1601_797#
+ powergood_check/FILLER_2_0/li_449_n17# powergood_check/FILLER_1_8/li_115_72# powergood_check/FILLER_1_140/li_353_797#
+ powergood_check/mprj2_logic_high_lv/li_1025_1611# powergood_check/FILLER_0_24/li_641_797#
+ powergood_check/mprj_logic_high_hvl/li_257_n17# powergood_check/mprj_logic_high_lv/li_384_1039#
+ powergood_check/FILLER_1_220/li_0_797# powergood_check/FILLER_1_172/li_65_797# powergood_check/FILLER_0_216/li_0_n17#
+ powergood_check/FILLER_2_107/li_65_797# powergood_check/FILLER_1_252/li_641_n17#
+ powergood_check/FILLER_2_243/li_161_n17# powergood_check/FILLER_0_272/li_353_797#
+ powergood_check/FILLER_1_0/li_353_n17# powergood_check/FILLER_0_192/li_161_797#
+ powergood_check/FILLER_2_219/li_353_797# powergood_check/FILLER_2_259/li_641_797#
+ powergood_check/FILLER_2_195/li_65_n17# powergood_check/FILLER_1_32/li_641_n17#
+ powergood_check/FILLER_2_251/li_257_797# powergood_check/FILLER_1_212/li_115_72#
+ powergood_check/FILLER_1_8/li_641_n17# powergood_check/FILLER_2_8/li_257_797# powergood_check/FILLER_1_204/li_65_n17#
+ powergood_check/FILLER_2_115/li_737_797# powergood_check/mprj2_logic_high_lv/li_929_1611#
+ powergood_check/FILLER_1_131/li_0_797# powergood_check/FILLER_0_88/li_115_72# powergood_check/FILLER_2_259/li_115_72#
+ powergood_check/FILLER_2_107/li_545_n17# powergood_check/FILLER_1_62/li_257_n17#
+ powergood_check/FILLER_0_192/li_65_n17# powergood_check/FILLER_0_240/li_257_797#
+ powergood_check/FILLER_1_220/li_545_n17# powergood_check/mprj2_logic_high_lv/li_826_79#
+ powergood_check/FILLER_1_131/li_161_n17# powergood_check/FILLER_1_140/li_353_n17#
+ powergood_check/FILLER_1_188/li_65_n17# powergood_check/FILLER_2_251/li_353_n17#
+ powergood_check/FILLER_1_180/li_641_n17# powergood_check/FILLER_2_227/li_545_797#
+ powergood_check/FILLER_2_219/li_65_n17# powergood_check/FILLER_2_171/li_161_n17#
+ powergood_check/FILLER_2_107/li_65_n17# powergood_check/FILLER_2_16/li_353_797#
+ powergood_check/FILLER_0_208/li_257_797# powergood_check/FILLER_2_187/li_641_797#
+ powergood_check/FILLER_1_131/li_353_797# powergood_check/FILLER_0_272/li_65_797#
+ powergood_check/FILLER_0_248/li_545_797# powergood_check/FILLER_2_219/li_353_n17#
+ powergood_check/FILLER_0_24/li_161_797# powergood_check/FILLER_0_160/li_65_797#
+ powergood_check/FILLER_0_168/li_353_797# powergood_check/FILLER_2_259/li_641_n17#
+ powergood_check/FILLER_1_252/li_161_n17# powergood_check/mprj_logic_high_lv/li_506_1123#
+ powergood_check/FILLER_2_8/li_257_n17# mgmt_protect_hv
XFILLER_19_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] mprj_logic_high_inst/HI[421] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[91\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[44\]_TE mprj_logic_high_inst/HI[246] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_sel_buf\[0\]_A _403_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[108\] _376_/Y mprj_logic_high_inst/HI[310] vssd vssd vccd
+ vccd la_oen_core[108] sky130_fd_sc_hd__einvp_8
XFILLER_28_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[38\] _637_/Y mprj_logic_high_inst/HI[240] vssd vssd vccd
+ vccd la_oen_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_16_459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__572__A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[82\]_TE la_buf\[82\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[1\]_A _440_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[67\]_TE mprj_logic_high_inst/HI[269] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y vssd vssd vccd vccd la_data_in_mprj[61]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__482__A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[90\]_A user_to_mprj_in_gates\[90\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__657__A la_oen_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B mprj_logic_high_inst/HI[426] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__392__A la_oen_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[81\]_A user_to_mprj_in_gates\[81\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[20\]_B mprj_logic_high_inst/HI[350] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__567__A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_653_ la_oen_mprj[54] vssd vssd vccd vccd _653_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_584_ la_data_out_mprj[113] vssd vssd vccd vccd _584_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[65\] _536_/Y la_buf\[65\]/TE vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_16_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[87\]_B mprj_logic_high_inst/HI[417] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[29\] _436_/Y mprj_adr_buf\[29\]/TE vssd vssd vccd vccd mprj_adr_o_user[29]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[121\] _592_/Y la_buf\[121\]/TE vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__einvp_8
XFILLER_12_1669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[72\]_A user_to_mprj_in_gates\[72\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_B mprj_logic_high_inst/HI[341] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__477__A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] mprj_logic_high_inst/HI[384] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[54\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[78\]_B mprj_logic_high_inst/HI[408] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[110\]_A user_to_mprj_in_gates\[110\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[63\]_A user_to_mprj_in_gates\[63\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__387__A la_oen_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_B mprj_logic_high_inst/HI[399] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[101\]_A user_to_mprj_in_gates\[101\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[54\]_A user_to_mprj_in_gates\[54\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_636_ la_oen_mprj[37] vssd vssd vccd vccd _636_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_567_ la_data_out_mprj[96] vssd vssd vccd vccd _567_/Y sky130_fd_sc_hd__inv_2
X_498_ la_data_out_mprj[27] vssd vssd vccd vccd _498_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[94\]_A _565_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y vssd vssd vccd vccd la_data_in_mprj[24]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[45\]_A user_to_mprj_in_gates\[45\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[85\]_A _556_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[36\]_A user_to_mprj_in_gates\[36\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_421_ mprj_adr_o_core[14] vssd vssd vccd vccd _421_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[2\] _601_/Y mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd la_oen_core[2] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[20\] _619_/Y mprj_logic_high_inst/HI[222] vssd vssd vccd
+ vccd la_oen_core[20] sky130_fd_sc_hd__einvp_8
X_352_ la_oen_mprj[84] vssd vssd vccd vccd _352_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[126\]_B mprj_logic_high_inst/HI[456] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[76\]_A _547_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__580__A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[28\] _499_/Y la_buf\[28\]/TE vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__einvp_8
XFILLER_10_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[27\]_A user_to_mprj_in_gates\[27\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[16\]_TE la_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_619_ la_oen_mprj[20] vssd vssd vccd vccd _619_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[117\]_B mprj_logic_high_inst/HI[447] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[67\]_A _538_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] mprj_logic_high_inst/HI[347] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[17\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__490__A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[18\]_A user_to_mprj_in_gates\[18\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[108\]_B mprj_logic_high_inst/HI[438] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[58\]_A _529_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[68\] _336_/Y mprj_logic_high_inst/HI[270] vssd vssd vccd
+ vccd la_oen_core[68] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[16\] _455_/Y mprj_dat_buf\[16\]/TE vssd vssd vccd vccd mprj_dat_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[39\]_TE la_buf\[39\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__575__A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_404_ mprj_sel_o_core[1] vssd vssd vccd vccd _404_/Y sky130_fd_sc_hd__inv_2
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[49\]_A _520_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_335_ la_oen_mprj[67] vssd vssd vccd vccd _335_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[11\] _418_/Y mprj_adr_buf\[11\]/TE vssd vssd vccd vccd mprj_adr_o_user[11]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[125] sky130_fd_sc_hd__inv_8
XFILLER_2_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y vssd vssd vccd vccd la_data_in_mprj[91]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__485__A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[7\]_TE la_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[125\]_A _393_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[60\]_A _659_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__395__A la_oen_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[51\]_A _650_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[116\]_A _384_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[95\] _566_/Y la_buf\[95\]/TE vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_19_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[42\]_A _641_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[107\]_A _375_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] mprj_logic_high_inst/HI[414] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[84\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[33\]_A _632_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[24\]_A _623_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[112\]_TE mprj_logic_high_inst/HI[314] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[6\] _477_/Y la_buf\[6\]/TE vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__einvp_8
Xla_buf\[10\] _481_/Y la_buf\[10\]/TE vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_26_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[3\] _410_/Y mprj_adr_buf\[3\]/TE vssd vssd vccd vccd mprj_adr_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_we_buf_TE mprj_we_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[20\]_A _427_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y vssd vssd vccd vccd la_data_in_mprj[54]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high_inst/HI[213] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[15\]_A _614_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] mprj_logic_high_inst/HI[440] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[110\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[11\]_A _418_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[120\] _388_/Y mprj_logic_high_inst/HI[322] vssd vssd vccd
+ vccd la_oen_core[120] sky130_fd_sc_hd__einvp_8
XFILLER_1_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[1\] _404_/Y mprj_sel_buf\[1\]/TE vssd vssd vccd vccd mprj_sel_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_27_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[50\] _649_/Y mprj_logic_high_inst/HI[252] vssd vssd vccd
+ vccd la_oen_core[50] sky130_fd_sc_hd__einvp_8
XFILLER_5_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_652_ la_oen_mprj[53] vssd vssd vccd vccd _652_/Y sky130_fd_sc_hd__inv_2
X_583_ la_data_out_mprj[112] vssd vssd vccd vccd _583_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__583__A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[58\] _529_/Y la_buf\[58\]/TE vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__einvp_8
XPHY_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[34\]_TE mprj_logic_high_inst/HI[236] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[114\] _585_/Y la_buf\[114\]/TE vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_3_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] mprj_logic_high_inst/HI[377] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[47\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__493__A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[9\]_TE mprj_adr_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] user_to_mprj_in_gates\[9\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[9\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[72\]_TE la_buf\[72\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[57\]_TE mprj_logic_high_inst/HI[259] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[98\] _366_/Y mprj_logic_high_inst/HI[300] vssd vssd vccd
+ vccd la_oen_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_1_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__578__A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_635_ la_oen_mprj[36] vssd vssd vccd vccd _635_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[24\]_A _463_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_566_ la_data_out_mprj[95] vssd vssd vccd vccd _566_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_497_ la_data_out_mprj[26] vssd vssd vccd vccd _497_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[0\]_TE mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y vssd vssd vccd vccd la_data_in_mprj[17]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_TE la_buf\[95\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__488__A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[15\]_A _454_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__398__A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_420_ mprj_adr_o_core[13] vssd vssd vccd vccd _420_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[13\] _612_/Y mprj_logic_high_inst/HI[215] vssd vssd vccd
+ vccd la_oen_core[13] sky130_fd_sc_hd__einvp_8
X_351_ la_oen_mprj[83] vssd vssd vccd vccd _351_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y vssd vssd vccd vccd la_data_in_mprj[9]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_618_ la_oen_mprj[19] vssd vssd vccd vccd _618_/Y sky130_fd_sc_hd__inv_2
X_549_ la_data_out_mprj[78] vssd vssd vccd vccd _549_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_403_ mprj_sel_o_core[0] vssd vssd vccd vccd _403_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[2\]_A _473_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[40\] _511_/Y la_buf\[40\]/TE vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__einvp_8
X_334_ la_oen_mprj[66] vssd vssd vccd vccd _334_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__591__A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[118] sky130_fd_sc_hd__inv_8
XFILLER_2_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y vssd vssd vccd vccd la_data_in_mprj[84]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[0\]_TE mprj_dat_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[120\]_TE la_buf\[120\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_A _416_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[80\] _348_/Y mprj_logic_high_inst/HI[282] vssd vssd vccd
+ vccd la_oen_core[80] sky130_fd_sc_hd__einvp_8
XFILLER_11_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__586__A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[88\] _559_/Y la_buf\[88\]/TE vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__einvp_8
XFILLER_21_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[0\]_A user_to_mprj_in_gates\[0\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] mprj_logic_high_inst/HI[407] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[77\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__496__A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high_inst/HI[292] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[29\]_TE la_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y vssd vssd vccd vccd la_data_in_mprj[47]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_2111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] mprj_logic_high_inst/HI[433] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[103\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[113\] _381_/Y mprj_logic_high_inst/HI[315] vssd vssd vccd
+ vccd la_oen_core[113] sky130_fd_sc_hd__einvp_8
Xmprj_clk2_buf _399_/Y mprj_clk2_buf/TE vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[9\]_B user_to_mprj_in_gates\[9\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_651_ la_oen_mprj[52] vssd vssd vccd vccd _651_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[43\] _642_/Y mprj_logic_high_inst/HI[245] vssd vssd vccd
+ vccd la_oen_core[43] sky130_fd_sc_hd__einvp_8
XFILLER_25_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_582_ la_data_out_mprj[111] vssd vssd vccd vccd _582_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[107\] _578_/Y la_buf\[107\]/TE vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_27_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[100] sky130_fd_sc_hd__inv_8
XFILLER_3_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high_inst/HI[304] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_634_ la_oen_mprj[35] vssd vssd vccd vccd _634_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__594__A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[70\] _541_/Y la_buf\[70\]/TE vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__einvp_8
XFILLER_2_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_565_ la_data_out_mprj[94] vssd vssd vccd vccd _565_/Y sky130_fd_sc_hd__inv_2
X_496_ la_data_out_mprj[25] vssd vssd vccd vccd _496_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high_inst/HI[327] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[24\]_TE mprj_logic_high_inst/HI[226] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_350_ la_oen_mprj[82] vssd vssd vccd vccd _350_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__589__A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_617_ la_oen_mprj[18] vssd vssd vccd vccd _617_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_548_ la_data_out_mprj[77] vssd vssd vccd vccd _548_/Y sky130_fd_sc_hd__inv_2
X_479_ la_data_out_mprj[8] vssd vssd vccd vccd _479_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[62\]_TE la_buf\[62\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high_inst/HI[249] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__499__A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_402_ mprj_we_o_core vssd vssd vccd vccd _402_/Y sky130_fd_sc_hd__inv_2
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_333_ la_oen_mprj[65] vssd vssd vccd vccd _333_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[85\]_TE la_buf\[85\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[33\] _504_/Y la_buf\[33\]/TE vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__einvp_8
XFILLER_13_1574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y vssd vssd vccd vccd la_data_in_mprj[77]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] mprj_logic_high_inst/HI[352] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[22\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_A _406_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[50\]_B mprj_logic_high_inst/HI[380] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[73\] _341_/Y mprj_logic_high_inst/HI[275] vssd vssd vccd
+ vccd la_oen_core[73] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[21\] _460_/Y mprj_dat_buf\[21\]/TE vssd vssd vccd vccd mprj_dat_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[4\]_A _443_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[41\]_B mprj_logic_high_inst/HI[371] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[93\]_A user_to_mprj_in_gates\[93\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[32\]_B mprj_logic_high_inst/HI[362] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[99\]_B mprj_logic_high_inst/HI[429] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[120\]_A _591_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[84\]_A user_to_mprj_in_gates\[84\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[23\]_B mprj_logic_high_inst/HI[353] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__597__A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[110\]_TE la_buf\[110\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[122\]_A user_to_mprj_in_gates\[122\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[111\]_A _582_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[75\]_A user_to_mprj_in_gates\[75\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B mprj_logic_high_inst/HI[344] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[113\]_A user_to_mprj_in_gates\[113\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[102\]_A _573_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[66\]_A user_to_mprj_in_gates\[66\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _374_/Y mprj_logic_high_inst/HI[308] vssd vssd vccd
+ vccd la_oen_core[106] sky130_fd_sc_hd__einvp_8
X_650_ la_oen_mprj[51] vssd vssd vccd vccd _650_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[36\] _635_/Y mprj_logic_high_inst/HI[238] vssd vssd vccd
+ vccd la_oen_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_5_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_581_ la_data_out_mprj[110] vssd vssd vccd vccd _581_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[104\]_A user_to_mprj_in_gates\[104\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[57\]_A user_to_mprj_in_gates\[57\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[30\]_A _501_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high_inst/HI[282] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[19\]_TE la_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[97\]_A _568_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[48\]_A user_to_mprj_in_gates\[48\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[21\]_A _492_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_A _559_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[39\]_A user_to_mprj_in_gates\[39\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[12\]_A _483_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_51 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_633_ la_oen_mprj[34] vssd vssd vccd vccd _633_/Y sky130_fd_sc_hd__inv_2
X_564_ la_data_out_mprj[93] vssd vssd vccd vccd _564_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[79\]_A _550_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[63\] _534_/Y la_buf\[63\]/TE vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__einvp_8
X_495_ la_data_out_mprj[24] vssd vssd vccd vccd _495_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[27\] _434_/Y mprj_adr_buf\[27\]/TE vssd vssd vccd vccd mprj_adr_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] mprj_logic_high_inst/HI[382] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[52\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[90\]_A _358_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[81\]_A _349_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_616_ la_oen_mprj[17] vssd vssd vccd vccd _616_/Y sky130_fd_sc_hd__inv_2
X_547_ la_data_out_mprj[76] vssd vssd vccd vccd _547_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_478_ la_data_out_mprj[7] vssd vssd vccd vccd _478_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[72\]_A _340_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y vssd vssd vccd vccd la_data_in_mprj[22]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[63\]_A _331_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[0\] _599_/Y mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd la_oen_core[0] sky130_fd_sc_hd__einvp_8
X_401_ mprj_stb_o_core vssd vssd vccd vccd _401_/Y sky130_fd_sc_hd__inv_2
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_332_ la_oen_mprj[64] vssd vssd vccd vccd _332_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_A _653_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[119\]_A _387_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high_inst/HI[317] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[26\] _497_/Y la_buf\[26\]/TE vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_26_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] mprj_logic_high_inst/HI[345] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[15\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[45\]_A _644_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high_inst/HI[216] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] mprj_logic_high_inst/HI[456] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[126\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[36\]_A _635_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[66\] _334_/Y mprj_logic_high_inst/HI[268] vssd vssd vccd
+ vccd la_oen_core[66] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[14\] _453_/Y mprj_dat_buf\[14\]/TE vssd vssd vccd vccd mprj_dat_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[52\]_TE la_buf\[52\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[37\]_TE mprj_logic_high_inst/HI[239] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[27\]_A _626_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[123] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_adr_buf\[23\]_A _430_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[0\]_A _599_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[18\]_A _617_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_A _421_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[75\]_TE la_buf\[75\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[93\] _564_/Y la_buf\[93\]/TE vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_5_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[98\]_TE la_buf\[98\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] mprj_logic_high_inst/HI[412] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[82\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_580_ la_data_out_mprj[109] vssd vssd vccd vccd _580_/Y sky130_fd_sc_hd__inv_2
XPHY_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[29\] _628_/Y mprj_logic_high_inst/HI[231] vssd vssd vccd
+ vccd la_oen_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_25_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[4\] _475_/Y la_buf\[4\]/TE vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__einvp_8
XFILLER_4_632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__401__A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[1\] _408_/Y mprj_adr_buf\[1\]/TE vssd vssd vccd vccd mprj_adr_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[27\]_A _466_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y vssd vssd vccd vccd la_data_in_mprj[52]
+ sky130_fd_sc_hd__inv_8
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_A _457_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[100\]_TE la_buf\[100\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_632_ la_oen_mprj[33] vssd vssd vccd vccd _632_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_563_ la_data_out_mprj[92] vssd vssd vccd vccd _563_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_494_ la_data_out_mprj[23] vssd vssd vccd vccd _494_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[56\] _527_/Y la_buf\[56\]/TE vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__einvp_8
XFILLER_9_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[112\] _583_/Y la_buf\[112\]/TE vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__einvp_8
XFILLER_5_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[3\]_TE mprj_dat_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] mprj_logic_high_inst/HI[375] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[45\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[123\]_TE la_buf\[123\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] user_to_mprj_in_gates\[7\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[7\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[70\]_TE mprj_logic_high_inst/HI[272] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[96\] _364_/Y mprj_logic_high_inst/HI[298] vssd vssd vccd
+ vccd la_oen_core[96] sky130_fd_sc_hd__einvp_8
XFILLER_6_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[5\]_A _476_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_615_ la_oen_mprj[16] vssd vssd vccd vccd _615_/Y sky130_fd_sc_hd__inv_2
X_546_ la_data_out_mprj[75] vssd vssd vccd vccd _546_/Y sky130_fd_sc_hd__inv_2
X_477_ la_data_out_mprj[6] vssd vssd vccd vccd _477_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y vssd vssd vccd vccd la_data_in_mprj[15]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high_inst/HI[295] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj2_pwrgood mprj2_pwrgood/A vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_28_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_400_ mprj_cyc_o_core vssd vssd vccd vccd _400_/Y sky130_fd_sc_hd__inv_2
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[11\] _610_/Y mprj_logic_high_inst/HI[213] vssd vssd vccd
+ vccd la_oen_core[11] sky130_fd_sc_hd__einvp_8
X_331_ la_oen_mprj[63] vssd vssd vccd vccd _331_/Y sky130_fd_sc_hd__inv_2
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y vssd vssd vccd vccd la_data_in_mprj[7]
+ sky130_fd_sc_hd__inv_8
XFILLER_10_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[19\] _490_/Y la_buf\[19\]/TE vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_13_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[3\]_A user_to_mprj_in_gates\[3\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_529_ la_data_out_mprj[58] vssd vssd vccd vccd _529_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_vdd_pwrgood_A mprj_vdd_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] mprj_logic_high_inst/HI[449] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[119\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[59\] _658_/Y mprj_logic_high_inst/HI[261] vssd vssd vccd
+ vccd la_oen_core[59] sky130_fd_sc_hd__einvp_8
XFILLER_21_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__404__A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[116] sky130_fd_sc_hd__inv_8
XFILLER_6_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y vssd vssd vccd vccd la_data_in_mprj[82]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_A _396_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_25_1200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[105\]_TE mprj_logic_high_inst/HI[307] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[86\] _557_/Y la_buf\[86\]/TE vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_5_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] mprj_logic_high_inst/HI[405] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[75\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[42\]_TE la_buf\[42\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high_inst/HI[229] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y vssd vssd vccd vccd la_data_in_mprj[45]
+ sky130_fd_sc_hd__inv_8
XPHY_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[65\]_TE la_buf\[65\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] mprj_logic_high_inst/HI[431] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[101\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_10_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[14\]_TE mprj_dat_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__502__A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[111\] _379_/Y mprj_logic_high_inst/HI[313] vssd vssd vccd
+ vccd la_oen_core[111] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[41\] _640_/Y mprj_logic_high_inst/HI[243] vssd vssd vccd
+ vccd la_oen_core[41] sky130_fd_sc_hd__einvp_8
X_631_ la_oen_mprj[32] vssd vssd vccd vccd _631_/Y sky130_fd_sc_hd__inv_2
X_562_ la_data_out_mprj[91] vssd vssd vccd vccd _562_/Y sky130_fd_sc_hd__inv_2
X_493_ la_data_out_mprj[22] vssd vssd vccd vccd _493_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[88\]_TE la_buf\[88\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[49\] _520_/Y la_buf\[49\]/TE vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_16_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__412__A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[105\] _576_/Y la_buf\[105\]/TE vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__einvp_8
XFILLER_23_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] mprj_logic_high_inst/HI[368] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[38\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[80\]_B mprj_logic_high_inst/HI[410] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[89\] _357_/Y mprj_logic_high_inst/HI[291] vssd vssd vccd
+ vccd la_oen_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_2_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_614_ la_oen_mprj[15] vssd vssd vccd vccd _614_/Y sky130_fd_sc_hd__inv_2
X_545_ la_data_out_mprj[74] vssd vssd vccd vccd _545_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__407__A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_476_ la_data_out_mprj[5] vssd vssd vccd vccd _476_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B mprj_logic_high_inst/HI[401] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_B mprj_logic_high_inst/HI[392] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_330_ la_oen_mprj[62] vssd vssd vccd vccd _330_/Y sky130_fd_sc_hd__inv_2
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[53\]_B mprj_logic_high_inst/HI[383] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[113\]_TE la_buf\[113\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[28\]_TE mprj_adr_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[7\]_A _446_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_528_ la_data_out_mprj[57] vssd vssd vccd vccd _528_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_459_ mprj_dat_o_core[20] vssd vssd vccd vccd _459_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[44\]_B mprj_logic_high_inst/HI[374] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__600__A la_oen_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_TE mprj_logic_high_inst/HI[262] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[96\]_A user_to_mprj_in_gates\[96\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[35\]_B mprj_logic_high_inst/HI[365] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__510__A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[20\]_A user_to_mprj_in_gates\[20\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[31\] _502_/Y la_buf\[31\]/TE vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[123\]_A _594_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[87\]_A user_to_mprj_in_gates\[87\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[26\]_B mprj_logic_high_inst/HI[356] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_B mprj_logic_high_inst/HI[440] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[60\]_A _531_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high_inst/HI[285] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__420__A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[109] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y vssd vssd vccd vccd la_data_in_mprj[75]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[11\]_A user_to_mprj_in_gates\[11\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] mprj_logic_high_inst/HI[350] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[20\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[125\]_A user_to_mprj_in_gates\[125\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[114\]_A _585_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[17\]_B mprj_logic_high_inst/HI[347] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_B mprj_logic_high_inst/HI[431] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[78\]_A user_to_mprj_in_gates\[78\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[51\]_A _522_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[8\] _447_/Y mprj_dat_buf\[8\]/TE vssd vssd vccd vccd mprj_dat_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__330__A la_oen_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[116\]_A user_to_mprj_in_gates\[116\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[105\]_A _576_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__505__A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[69\]_A user_to_mprj_in_gates\[69\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[42\]_A _513_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[71\] _339_/Y mprj_logic_high_inst/HI[273] vssd vssd vccd
+ vccd la_oen_core[71] sky130_fd_sc_hd__einvp_8
XFILLER_23_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[79\] _550_/Y la_buf\[79\]/TE vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_27_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[107\]_A user_to_mprj_in_gates\[107\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__415__A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[33\]_A _504_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] mprj_logic_high_inst/HI[398] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[68\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[24\]_A _495_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[15\]_A _486_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[100\]_A _368_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y vssd vssd vccd vccd la_data_in_mprj[38]
+ sky130_fd_sc_hd__inv_8
XPHY_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[93\]_A _361_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[104\] _372_/Y mprj_logic_high_inst/HI[306] vssd vssd vccd
+ vccd la_oen_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_28_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_630_ la_oen_mprj[31] vssd vssd vccd vccd _630_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[34\] _633_/Y mprj_logic_high_inst/HI[236] vssd vssd vccd
+ vccd la_oen_core[34] sky130_fd_sc_hd__einvp_8
XFILLER_22_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_561_ la_data_out_mprj[90] vssd vssd vccd vccd _561_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_492_ la_data_out_mprj[21] vssd vssd vccd vccd _492_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[84\]_A _352_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high_inst/HI[320] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[32\]_TE la_buf\[32\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[17\]_TE mprj_logic_high_inst/HI[219] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[75\]_A _343_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__603__A la_oen_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[66\]_A _334_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_45 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[0\]_TE la_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__513__A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_613_ la_oen_mprj[14] vssd vssd vccd vccd _613_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[55\]_TE la_buf\[55\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_544_ la_data_out_mprj[73] vssd vssd vccd vccd _544_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[61\] _532_/Y la_buf\[61\]/TE vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__einvp_8
XFILLER_18_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_475_ la_data_out_mprj[4] vssd vssd vccd vccd _475_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[57\]_A _656_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[25\] _432_/Y mprj_adr_buf\[25\]/TE vssd vssd vccd vccd mprj_adr_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__423__A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] mprj_logic_high_inst/HI[380] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[50\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[48\]_A _647_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__333__A la_oen_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[78\]_TE la_buf\[78\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__508__A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[39\]_A _638_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_TE mprj_dat_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__418__A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_527_ la_data_out_mprj[56] vssd vssd vccd vccd _527_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[6\]_TE mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_458_ mprj_dat_o_core[19] vssd vssd vccd vccd _458_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_389_ la_oen_mprj[121] vssd vssd vccd vccd _389_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y vssd vssd vccd vccd la_data_in_mprj[20]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] mprj_logic_high_inst/HI[428] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[98\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[26\]_A _433_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[3\]_A _602_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[17\]_A _424_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[24\] _495_/Y la_buf\[24\]/TE vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__einvp_8
XFILLER_11_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y vssd vssd vccd vccd la_data_in_mprj[68]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] mprj_logic_high_inst/HI[343] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[13\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__611__A la_oen_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] mprj_logic_high_inst/HI[454] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[124\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[103\]_TE la_buf\[103\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__521__A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[64\] _332_/Y mprj_logic_high_inst/HI[266] vssd vssd vccd
+ vccd la_oen_core[64] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[12\] _451_/Y mprj_dat_buf\[12\]/TE vssd vssd vccd vccd mprj_dat_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_cyc_buf_A _400_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[50\]_TE mprj_logic_high_inst/HI[252] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__431__A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[121] sky130_fd_sc_hd__inv_8
XFILLER_3_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[6\]_TE mprj_dat_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[126\]_TE la_buf\[126\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__606__A la_oen_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[2\]_A _409_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__341__A la_oen_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[73\]_TE mprj_logic_high_inst/HI[275] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__516__A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[91\] _562_/Y la_buf\[91\]/TE vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_15_230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__426__A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] mprj_logic_high_inst/HI[410] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[80\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high_inst/HI[298] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__336__A la_oen_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_560_ la_data_out_mprj[89] vssd vssd vccd vccd _560_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[27\] _626_/Y mprj_logic_high_inst/HI[229] vssd vssd vccd
+ vccd la_oen_core[27] sky130_fd_sc_hd__einvp_8
X_491_ la_data_out_mprj[20] vssd vssd vccd vccd _491_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[9\] _608_/Y mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd la_oen_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_25_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[2\] _473_/Y la_buf\[2\]/TE vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__einvp_8
XFILLER_5_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[8\]_A _479_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y vssd vssd vccd vccd la_data_in_mprj[50]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[2\]_B user_to_mprj_in_gates\[2\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_612_ la_oen_mprj[13] vssd vssd vccd vccd _612_/Y sky130_fd_sc_hd__inv_2
X_543_ la_data_out_mprj[72] vssd vssd vccd vccd _543_/Y sky130_fd_sc_hd__inv_2
X_474_ la_data_out_mprj[3] vssd vssd vccd vccd _474_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[54\] _525_/Y la_buf\[54\]/TE vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_9_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[18\] _425_/Y mprj_adr_buf\[18\]/TE vssd vssd vccd vccd mprj_adr_o_user[18]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[110\] _581_/Y la_buf\[110\]/TE vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__einvp_8
XFILLER_9_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y vssd vssd vccd vccd la_data_in_mprj[98]
+ sky130_fd_sc_hd__inv_8
XFILLER_23_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[6\]_A user_to_mprj_in_gates\[6\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] mprj_logic_high_inst/HI[373] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[43\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__A la_oen_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] user_to_mprj_in_gates\[5\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[5\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[108\]_TE mprj_logic_high_inst/HI[310] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__524__A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[94\] _362_/Y mprj_logic_high_inst/HI[296] vssd vssd vccd
+ vccd la_oen_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_2_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[22\]_TE la_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_526_ la_data_out_mprj[55] vssd vssd vccd vccd _526_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_457_ mprj_dat_o_core[18] vssd vssd vccd vccd _457_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_388_ la_oen_mprj[120] vssd vssd vccd vccd _388_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_9_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__434__A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y vssd vssd vccd vccd la_data_in_mprj[13]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__609__A la_oen_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__344__A la_oen_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[45\]_TE la_buf\[45\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__519__A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y vssd vssd vccd vccd la_data_in_mprj[5]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[17\] _488_/Y la_buf\[17\]/TE vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__einvp_8
XFILLER_26_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__429__A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_509_ la_data_out_mprj[38] vssd vssd vccd vccd _509_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[68\]_TE la_buf\[68\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] mprj_logic_high_inst/HI[447] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[117\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__339__A la_oen_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[127\] _395_/Y mprj_logic_high_inst/HI[329] vssd vssd vccd
+ vccd la_oen_core[127] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[57\] _656_/Y mprj_logic_high_inst/HI[259] vssd vssd vccd
+ vccd la_oen_core[57] sky130_fd_sc_hd__einvp_8
XFILLER_25_1770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[114] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y vssd vssd vccd vccd la_data_in_mprj[80]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__622__A la_oen_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__532__A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[84\] _555_/Y la_buf\[84\]/TE vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_15_242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__442__A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] mprj_logic_high_inst/HI[403] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[73\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__617__A la_oen_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[92\]_B mprj_logic_high_inst/HI[422] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__352__A la_oen_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high_inst/HI[242] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_490_ la_data_out_mprj[19] vssd vssd vccd vccd _490_/Y sky130_fd_sc_hd__inv_2
XANTENNA__527__A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[83\]_B mprj_logic_high_inst/HI[413] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[116\]_TE la_buf\[116\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__437__A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y vssd vssd vccd vccd la_data_in_mprj[43]
+ sky130_fd_sc_hd__inv_8
XPHY_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[74\]_B mprj_logic_high_inst/HI[404] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[63\]_TE mprj_logic_high_inst/HI[265] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__347__A la_oen_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[65\]_B mprj_logic_high_inst/HI[395] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[50\]_A user_to_mprj_in_gates\[50\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_611_ la_oen_mprj[12] vssd vssd vccd vccd _611_/Y sky130_fd_sc_hd__inv_2
X_542_ la_data_out_mprj[71] vssd vssd vccd vccd _542_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_473_ la_data_out_mprj[2] vssd vssd vccd vccd _473_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[47\] _518_/Y la_buf\[47\]/TE vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[56\]_B mprj_logic_high_inst/HI[386] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[90\]_A _561_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high_inst/HI[288] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[103\] _574_/Y la_buf\[103\]/TE vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__einvp_8
XFILLER_9_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[41\]_A user_to_mprj_in_gates\[41\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] mprj_logic_high_inst/HI[366] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[36\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[47\]_B mprj_logic_high_inst/HI[377] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[81\]_A _552_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__630__A la_oen_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[32\]_A user_to_mprj_in_gates\[32\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[99\]_A user_to_mprj_in_gates\[99\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[38\]_B mprj_logic_high_inst/HI[368] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_B mprj_logic_high_inst/HI[452] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[72\]_A _543_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[87\] _355_/Y mprj_logic_high_inst/HI[289] vssd vssd vccd
+ vccd la_oen_core[87] sky130_fd_sc_hd__einvp_8
XANTENNA__540__A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[23\]_A user_to_mprj_in_gates\[23\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_525_ la_data_out_mprj[54] vssd vssd vccd vccd _525_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_456_ mprj_dat_o_core[17] vssd vssd vccd vccd _456_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[126\]_A _597_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_387_ la_oen_mprj[119] vssd vssd vccd vccd _387_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[113\]_B mprj_logic_high_inst/HI[443] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_B mprj_logic_high_inst/HI[359] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[30\] _437_/Y mprj_adr_buf\[30\]/TE vssd vssd vccd vccd mprj_adr_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[63\]_A _534_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__450__A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[14\]_A user_to_mprj_in_gates\[14\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[117\]_A _588_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__625__A la_oen_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_B mprj_logic_high_inst/HI[434] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[54\]_A _525_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__360__A la_oen_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_stb_buf_A _401_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[119\]_A user_to_mprj_in_gates\[119\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[108\]_A _579_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__535__A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[45\]_A _516_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_508_ la_data_out_mprj[37] vssd vssd vccd vccd _508_/Y sky130_fd_sc_hd__inv_2
XANTENNA__445__A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_439_ mprj_dat_o_core[0] vssd vssd vccd vccd _439_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[36\]_A _507_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_A _389_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_71 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[12\]_TE la_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__355__A la_oen_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[27\]_A _498_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[112\]_A _380_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_49 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[18\]_A _489_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[103\]_A _371_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[107] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y vssd vssd vccd vccd la_data_in_mprj[73]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[35\]_TE la_buf\[35\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _445_/Y mprj_dat_buf\[6\]/TE vssd vssd vccd vccd mprj_dat_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_25_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[96\]_A _364_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_TE la_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[20\]_A _619_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[58\]_TE la_buf\[58\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[77\] _548_/Y la_buf\[77\]/TE vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__einvp_8
XFILLER_28_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[87\]_A _355_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[11\]_A _610_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] mprj_logic_high_inst/HI[396] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[66\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[78\]_A _346_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__633__A la_oen_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[69\]_A _337_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__543__A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y vssd vssd vccd vccd la_data_in_mprj[36]
+ sky130_fd_sc_hd__inv_8
XPHY_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__453__A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__628__A la_oen_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__363__A la_oen_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[102\] _370_/Y mprj_logic_high_inst/HI[304] vssd vssd vccd
+ vccd la_oen_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_4_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_610_ la_oen_mprj[11] vssd vssd vccd vccd _610_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_541_ la_data_out_mprj[70] vssd vssd vccd vccd _541_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[32\] _631_/Y mprj_logic_high_inst/HI[234] vssd vssd vccd
+ vccd la_oen_core[32] sky130_fd_sc_hd__einvp_8
X_472_ la_data_out_mprj[1] vssd vssd vccd vccd _472_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[20\]_A _459_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__448__A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[11\]_A _450_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] mprj_logic_high_inst/HI[359] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[29\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high_inst/HI[232] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_A _436_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__358__A la_oen_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[6\]_A _605_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[106\]_TE la_buf\[106\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[28\] _467_/Y mprj_dat_buf\[28\]/TE vssd vssd vccd vccd mprj_dat_o_user[28]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_524_ la_data_out_mprj[53] vssd vssd vccd vccd _524_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_455_ mprj_dat_o_core[16] vssd vssd vccd vccd _455_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[53\]_TE mprj_logic_high_inst/HI[255] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_386_ la_oen_mprj[118] vssd vssd vccd vccd _386_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[23\] _430_/Y mprj_adr_buf\[23\]/TE vssd vssd vccd vccd mprj_adr_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[9\]_TE mprj_dat_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__641__A la_oen_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[91\]_TE la_buf\[91\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[76\]_TE mprj_logic_high_inst/HI[278] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__551__A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_507_ la_data_out_mprj[36] vssd vssd vccd vccd _507_/Y sky130_fd_sc_hd__inv_2
X_438_ mprj_adr_o_core[31] vssd vssd vccd vccd _438_/Y sky130_fd_sc_hd__inv_2
X_369_ la_oen_mprj[101] vssd vssd vccd vccd _369_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__461__A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] mprj_logic_high_inst/HI[426] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[96\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high_inst/HI[301] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__636__A la_oen_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[5\]_A _412_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__371__A la_oen_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[22\] _493_/Y la_buf\[22\]/TE vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__einvp_8
XFILLER_13_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_stb_buf_TE mprj_stb_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y vssd vssd vccd vccd la_data_in_mprj[66]
+ sky130_fd_sc_hd__inv_8
XANTENNA__456__A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] mprj_logic_high_inst/HI[341] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[11\]/Y sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] mprj_logic_high_inst/HI[452] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[122\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__366__A la_oen_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_TE mprj_adr_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[62\] _330_/Y mprj_logic_high_inst/HI[264] vssd vssd vccd
+ vccd la_oen_core[62] sky130_fd_sc_hd__einvp_8
XFILLER_27_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[10\] _449_/Y mprj_dat_buf\[10\]/TE vssd vssd vccd vccd mprj_dat_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[126\] _597_/Y la_buf\[126\]/TE vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_10_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] mprj_logic_high_inst/HI[389] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[59\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[5\]_B user_to_mprj_in_gates\[5\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[25\]_TE la_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y vssd vssd vccd vccd la_data_in_mprj[29]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__644__A la_oen_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[48\]_TE la_buf\[48\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_540_ la_data_out_mprj[69] vssd vssd vccd vccd _540_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[25\] _624_/Y mprj_logic_high_inst/HI[227] vssd vssd vccd
+ vccd la_oen_core[25] sky130_fd_sc_hd__einvp_8
X_471_ la_data_out_mprj[0] vssd vssd vccd vccd _471_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[7\] _606_/Y mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd la_oen_core[7] sky130_fd_sc_hd__einvp_8
XFILLER_26_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__554__A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xla_buf\[0\] _471_/Y la_buf\[0\]/TE vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__einvp_8
XFILLER_5_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__464__A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_6_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__639__A la_oen_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__374__A la_oen_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_17_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__549__A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_523_ la_data_out_mprj[52] vssd vssd vccd vccd _523_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_454_ mprj_dat_o_core[15] vssd vssd vccd vccd _454_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[52\] _523_/Y la_buf\[52\]/TE vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__einvp_8
X_385_ la_oen_mprj[117] vssd vssd vccd vccd _385_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[16\] _423_/Y mprj_adr_buf\[16\]/TE vssd vssd vccd vccd mprj_adr_o_user[16]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y vssd vssd vccd vccd la_data_in_mprj[96]
+ sky130_fd_sc_hd__inv_8
XFILLER_27_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__459__A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_rstn_buf _396_/Y mprj_rstn_buf/TE vssd vssd vccd vccd user_resetn sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] mprj_logic_high_inst/HI[371] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[41\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] user_to_mprj_in_gates\[3\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[3\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__369__A la_oen_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_TE mprj_logic_high_inst/HI[323] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[92\] _360_/Y mprj_logic_high_inst/HI[294] vssd vssd vccd
+ vccd la_oen_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_24_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[20\]_TE mprj_logic_high_inst/HI[222] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_506_ la_data_out_mprj[35] vssd vssd vccd vccd _506_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_437_ mprj_adr_o_core[30] vssd vssd vccd vccd _437_/Y sky130_fd_sc_hd__inv_2
X_368_ la_oen_mprj[100] vssd vssd vccd vccd _368_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y vssd vssd vccd vccd la_data_in_mprj[11]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] mprj_logic_high_inst/HI[419] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[89\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__652__A la_oen_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[43\]_TE mprj_logic_high_inst/HI[245] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_cyc_buf _400_/Y mprj_cyc_buf/TE vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__einvp_8
XFILLER_15_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y vssd vssd vccd vccd la_data_in_mprj[3]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__562__A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[15\] _486_/Y la_buf\[15\]/TE vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[119\]_TE la_buf\[119\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_A _439_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[8\] _415_/Y mprj_adr_buf\[8\]/TE vssd vssd vccd vccd mprj_adr_o_user[8]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y vssd vssd vccd vccd la_data_in_mprj[59]
+ sky130_fd_sc_hd__inv_8
XANTENNA__472__A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[81\]_TE la_buf\[81\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[66\]_TE mprj_logic_high_inst/HI[268] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] mprj_logic_high_inst/HI[445] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[115\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__647__A la_oen_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_746 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[95\]_B mprj_logic_high_inst/HI[425] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__382__A la_oen_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_clk2_buf_TE mprj_clk2_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[30\]_TE mprj_dat_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[125\] _393_/Y mprj_logic_high_inst/HI[327] vssd vssd vccd
+ vccd la_oen_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_0_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[55\] _654_/Y mprj_logic_high_inst/HI[257] vssd vssd vccd
+ vccd la_oen_core[55] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[80\]_A user_to_mprj_in_gates\[80\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__557__A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[86\]_B mprj_logic_high_inst/HI[416] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high_inst/HI[291] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[119\] _590_/Y la_buf\[119\]/TE vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_3_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[112] sky130_fd_sc_hd__inv_8
XFILLER_6_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[71\]_A user_to_mprj_in_gates\[71\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[10\]_B mprj_logic_high_inst/HI[340] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__467__A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_B mprj_logic_high_inst/HI[407] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[62\]_A user_to_mprj_in_gates\[62\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__377__A la_oen_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[68\]_B mprj_logic_high_inst/HI[398] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[100\]_A user_to_mprj_in_gates\[100\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[53\]_A user_to_mprj_in_gates\[53\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[82\] _553_/Y la_buf\[82\]/TE vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__einvp_8
XFILLER_1_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_B mprj_logic_high_inst/HI[389] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[93\]_A _564_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[44\]_A user_to_mprj_in_gates\[44\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] mprj_logic_high_inst/HI[401] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[71\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[84\]_A _555_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__660__A la_oen_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[35\]_A user_to_mprj_in_gates\[35\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_470_ mprj_dat_o_core[31] vssd vssd vccd vccd _470_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[18\] _617_/Y mprj_logic_high_inst/HI[220] vssd vssd vccd
+ vccd la_oen_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_25_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_B mprj_logic_high_inst/HI[455] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[75\]_A _546_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[26\]_A user_to_mprj_in_gates\[26\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_599_ la_oen_mprj[0] vssd vssd vccd vccd _599_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y vssd vssd vccd vccd la_data_in_mprj[41]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[116\]_B mprj_logic_high_inst/HI[446] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[66\]_A _537_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__480__A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[17\]_A user_to_mprj_in_gates\[17\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[15\]_TE la_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__655__A la_oen_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[107\]_B mprj_logic_high_inst/HI[437] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[57\]_A _528_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__390__A la_oen_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_522_ la_data_out_mprj[51] vssd vssd vccd vccd _522_/Y sky130_fd_sc_hd__inv_2
X_453_ mprj_dat_o_core[14] vssd vssd vccd vccd _453_/Y sky130_fd_sc_hd__inv_2
XANTENNA__565__A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_384_ la_oen_mprj[116] vssd vssd vccd vccd _384_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[45\] _516_/Y la_buf\[45\]/TE vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[48\]_A _519_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[101\] _572_/Y la_buf\[101\]/TE vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_0_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y vssd vssd vccd vccd la_data_in_mprj[89]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[38\]_TE la_buf\[38\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__475__A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] mprj_logic_high_inst/HI[364] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[34\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[39\]_A _510_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[124\]_A _392_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__385__A la_oen_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[6\]_TE la_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[85\] _353_/Y mprj_logic_high_inst/HI[287] vssd vssd vccd
+ vccd la_oen_core[85] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[50\]_A _649_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_A _383_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_505_ la_data_out_mprj[34] vssd vssd vccd vccd _505_/Y sky130_fd_sc_hd__inv_2
X_436_ mprj_adr_o_core[29] vssd vssd vccd vccd _436_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_367_ la_oen_mprj[99] vssd vssd vccd vccd _367_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[41\]_A _640_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[106\]_A _374_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_A _631_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[99\]_A _367_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_A _622_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_419_ mprj_adr_o_core[12] vssd vssd vccd vccd _419_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high_inst/HI[313] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[14\]_A _613_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] mprj_logic_high_inst/HI[438] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[108\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[10\]_A _417_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high_inst/HI[212] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[118\] _386_/Y mprj_logic_high_inst/HI[320] vssd vssd vccd
+ vccd la_oen_core[118] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[48\] _647_/Y mprj_logic_high_inst/HI[250] vssd vssd vccd
+ vccd la_oen_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_28_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__573__A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[105] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y vssd vssd vccd vccd la_data_in_mprj[71]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[33\]_TE mprj_logic_high_inst/HI[235] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_84 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[4\] _443_/Y mprj_dat_buf\[4\]/TE vssd vssd vccd vccd mprj_dat_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__658__A la_oen_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[109\]_TE la_buf\[109\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__393__A la_oen_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__568__A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_TE la_buf\[71\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_A _462_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[75\] _546_/Y la_buf\[75\]/TE vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[56\]_TE mprj_logic_high_inst/HI[258] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__478__A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] mprj_logic_high_inst/HI[394] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[64\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[14\]_A _453_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[94\]_TE la_buf\[94\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__388__A la_oen_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[79\]_TE mprj_logic_high_inst/HI[281] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[9\]_A _608_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_598_ la_data_out_mprj[127] vssd vssd vccd vccd _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y vssd vssd vccd vccd la_data_in_mprj[34]
+ sky130_fd_sc_hd__inv_8
XPHY_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[100\] _368_/Y mprj_logic_high_inst/HI[302] vssd vssd vccd
+ vccd la_oen_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_8_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[30\] _629_/Y mprj_logic_high_inst/HI[232] vssd vssd vccd
+ vccd la_oen_core[30] sky130_fd_sc_hd__einvp_8
X_521_ la_data_out_mprj[50] vssd vssd vccd vccd _521_/Y sky130_fd_sc_hd__inv_2
X_452_ mprj_dat_o_core[13] vssd vssd vccd vccd _452_/Y sky130_fd_sc_hd__inv_2
X_383_ la_oen_mprj[115] vssd vssd vccd vccd _383_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[1\]_A _472_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__581__A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[38\] _509_/Y la_buf\[38\]/TE vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_12_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] mprj_logic_high_inst/HI[357] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[27\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__491__A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_A _415_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[78\] _346_/Y mprj_logic_high_inst/HI[280] vssd vssd vccd
+ vccd la_oen_core[78] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[26\] _465_/Y mprj_dat_buf\[26\]/TE vssd vssd vccd vccd mprj_dat_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__576__A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_504_ la_data_out_mprj[33] vssd vssd vccd vccd _504_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_435_ mprj_adr_o_core[28] vssd vssd vccd vccd _435_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_366_ la_oen_mprj[98] vssd vssd vccd vccd _366_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[21\] _428_/Y mprj_adr_buf\[21\]/TE vssd vssd vccd vccd mprj_adr_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__486__A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__396__A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[28\]_TE la_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_418_ mprj_adr_o_core[11] vssd vssd vccd vccd _418_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_349_ la_oen_mprj[81] vssd vssd vccd vccd _349_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] mprj_logic_high_inst/HI[424] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[94\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[8\]_B user_to_mprj_in_gates\[8\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[20\] _491_/Y la_buf\[20\]/TE vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__einvp_8
XFILLER_3_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_87 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y vssd vssd vccd vccd la_data_in_mprj[64]
+ sky130_fd_sc_hd__inv_8
XFILLER_21_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_41 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] mprj_logic_high_inst/HI[450] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[120\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[60\] _659_/Y mprj_logic_high_inst/HI[262] vssd vssd vccd
+ vccd la_oen_core[60] sky130_fd_sc_hd__einvp_8
XFILLER_0_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high_inst/HI[303] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__584__A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[68\] _539_/Y la_buf\[68\]/TE vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__einvp_8
XPHY_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[124\] _595_/Y la_buf\[124\]/TE vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_4_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] mprj_logic_high_inst/HI[387] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[57\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__494__A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_22_515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high_inst/HI[326] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__579__A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_TE mprj_logic_high_inst/HI[225] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_597_ la_data_out_mprj[126] vssd vssd vccd vccd _597_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y vssd vssd vccd vccd la_data_in_mprj[27]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__489__A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[61\]_TE la_buf\[61\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high_inst/HI[248] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__399__A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_520_ la_data_out_mprj[49] vssd vssd vccd vccd _520_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[5\] _604_/Y mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd la_oen_core[5] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[23\] _622_/Y mprj_logic_high_inst/HI[225] vssd vssd vccd
+ vccd la_oen_core[23] sky130_fd_sc_hd__einvp_8
X_451_ mprj_dat_o_core[12] vssd vssd vccd vccd _451_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_382_ la_oen_mprj[114] vssd vssd vccd vccd _382_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[10\]_TE mprj_dat_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_649_ la_oen_mprj[50] vssd vssd vccd vccd _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[84\]_TE la_buf\[84\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[69\]_TE mprj_logic_high_inst/HI[271] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[2\]_A _405_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[19\] _458_/Y mprj_dat_buf\[19\]/TE vssd vssd vccd vccd mprj_dat_o_user[19]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_503_ la_data_out_mprj[32] vssd vssd vccd vccd _503_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_434_ mprj_adr_o_core[27] vssd vssd vccd vccd _434_/Y sky130_fd_sc_hd__inv_2
XANTENNA__592__A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[50\] _521_/Y la_buf\[50\]/TE vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__einvp_8
X_365_ la_oen_mprj[97] vssd vssd vccd vccd _365_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_A _442_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[14\] _421_/Y mprj_adr_buf\[14\]/TE vssd vssd vccd vccd mprj_adr_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[40\]_B mprj_logic_high_inst/HI[370] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y vssd vssd vccd vccd la_data_in_mprj[94]
+ sky130_fd_sc_hd__inv_8
XFILLER_3_76 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] user_to_mprj_in_gates\[1\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[1\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[92\]_A user_to_mprj_in_gates\[92\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[31\]_B mprj_logic_high_inst/HI[361] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_B mprj_logic_high_inst/HI[428] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[90\] _358_/Y mprj_logic_high_inst/HI[292] vssd vssd vccd
+ vccd la_oen_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_3_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[83\]_A user_to_mprj_in_gates\[83\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[22\]_B mprj_logic_high_inst/HI[352] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[98\] _569_/Y la_buf\[98\]/TE vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_4_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__587__A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[89\]_B mprj_logic_high_inst/HI[419] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_417_ mprj_adr_o_core[10] vssd vssd vccd vccd _417_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_348_ la_oen_mprj[80] vssd vssd vccd vccd _348_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[121\]_A user_to_mprj_in_gates\[121\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[110\]_A _581_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[74\]_A user_to_mprj_in_gates\[74\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[13\]_B mprj_logic_high_inst/HI[343] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] mprj_logic_high_inst/HI[417] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[87\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__497__A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[112\]_A user_to_mprj_in_gates\[112\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[101\]_A _572_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[65\]_A user_to_mprj_in_gates\[65\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y vssd vssd vccd vccd la_data_in_mprj[1]
+ sky130_fd_sc_hd__inv_8
XPHY_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[103\]_A user_to_mprj_in_gates\[103\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[13\] _484_/Y la_buf\[13\]/TE vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__einvp_8
Xla_buf\[9\] _480_/Y la_buf\[9\]/TE vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_10_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[56\]_A user_to_mprj_in_gates\[56\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[6\] _413_/Y mprj_adr_buf\[6\]/TE vssd vssd vccd vccd mprj_adr_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y vssd vssd vccd vccd la_data_in_mprj[57]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[96\]_A _567_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[47\]_A user_to_mprj_in_gates\[47\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[20\]_A _491_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] mprj_logic_high_inst/HI[443] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[113\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[18\]_TE la_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[87\]_A _558_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[38\]_A user_to_mprj_in_gates\[38\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[123\] _391_/Y mprj_logic_high_inst/HI[325] vssd vssd vccd
+ vccd la_oen_core[123] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[11\]_A _482_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[53\] _652_/Y mprj_logic_high_inst/HI[255] vssd vssd vccd
+ vccd la_oen_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_1_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[78\]_A _549_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[29\]_A user_to_mprj_in_gates\[29\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[117\] _588_/Y la_buf\[117\]/TE vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_4_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[110] sky130_fd_sc_hd__inv_8
XFILLER_19_362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_B mprj_logic_high_inst/HI[449] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[69\]_A _540_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_TE la_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[80\]_A _348_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[80\] _551_/Y la_buf\[80\]/TE vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__einvp_8
XANTENNA__595__A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_596_ la_data_out_mprj[125] vssd vssd vccd vccd _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[71\]_A _339_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[62\]_A _330_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[127\]_A _395_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_450_ mprj_dat_o_core[11] vssd vssd vccd vccd _450_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[16\] _615_/Y mprj_logic_high_inst/HI[218] vssd vssd vccd
+ vccd la_oen_core[16] sky130_fd_sc_hd__einvp_8
X_381_ la_oen_mprj[113] vssd vssd vccd vccd _381_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[53\]_A _652_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[118\]_A _386_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_648_ la_oen_mprj[49] vssd vssd vccd vccd _648_/Y sky130_fd_sc_hd__inv_2
X_579_ la_data_out_mprj[108] vssd vssd vccd vccd _579_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[114\]_TE mprj_logic_high_inst/HI[316] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[44\]_A _643_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[109\]_A _377_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high_inst/HI[215] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[35\]_A _634_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_A _438_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_502_ la_data_out_mprj[31] vssd vssd vccd vccd _502_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_433_ mprj_adr_o_core[26] vssd vssd vccd vccd _433_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_364_ la_oen_mprj[96] vssd vssd vccd vccd _364_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[43\] _514_/Y la_buf\[43\]/TE vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__einvp_8
XFILLER_9_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[26\]_A _625_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[22\]_A _429_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y vssd vssd vccd vccd la_data_in_mprj[87]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[51\]_TE la_buf\[51\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] mprj_logic_high_inst/HI[362] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[32\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high_inst/HI[238] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[17\]_A _616_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_A _420_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[83\] _351_/Y mprj_logic_high_inst/HI[285] vssd vssd vccd
+ vccd la_oen_core[83] sky130_fd_sc_hd__einvp_8
XFILLER_3_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[31\] _470_/Y mprj_dat_buf\[31\]/TE vssd vssd vccd vccd mprj_dat_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[74\]_TE la_buf\[74\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[59\]_TE mprj_logic_high_inst/HI[261] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_416_ mprj_adr_o_core[9] vssd vssd vccd vccd _416_/Y sky130_fd_sc_hd__inv_2
X_347_ la_oen_mprj[79] vssd vssd vccd vccd _347_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[97\]_TE la_buf\[97\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__598__A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[26\]_A _465_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[17\]_A _456_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] mprj_logic_high_inst/HI[436] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[106\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[116\] _384_/Y mprj_logic_high_inst/HI[318] vssd vssd vccd
+ vccd la_oen_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_5_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[46\] _645_/Y mprj_logic_high_inst/HI[248] vssd vssd vccd
+ vccd la_oen_core[46] sky130_fd_sc_hd__einvp_8
XFILLER_1_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[14\]_TE mprj_adr_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[103] sky130_fd_sc_hd__inv_8
XFILLER_19_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[2\] _441_/Y mprj_dat_buf\[2\]/TE vssd vssd vccd vccd mprj_dat_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[2\]_TE mprj_dat_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[122\]_TE la_buf\[122\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[4\]_A _475_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[73\] _544_/Y la_buf\[73\]/TE vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__einvp_8
X_595_ la_data_out_mprj[124] vssd vssd vccd vccd _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] mprj_logic_high_inst/HI[392] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[62\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_380_ la_oen_mprj[112] vssd vssd vccd vccd _380_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high_inst/HI[294] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_647_ la_oen_mprj[48] vssd vssd vccd vccd _647_/Y sky130_fd_sc_hd__inv_2
X_578_ la_data_out_mprj[107] vssd vssd vccd vccd _578_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[2\]_A user_to_mprj_in_gates\[2\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y vssd vssd vccd vccd la_data_in_mprj[32]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_1808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__diode_2 abstract view
.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped A X VPWR VGND LVPWR LVGND FILLER_0_28/li_65_797#
+ lvlshiftdown/li_1313_1611# lvlshiftdown/li_353_1611# FILLER_1_8/li_161_n17# FILLER_1_8/li_50_537#
+ FILLER_0_28/li_0_n17# lvlshiftdown/li_65_797# FILLER_0_24/li_0_797# FILLER_0_0/li_545_797#
+ FILLER_2_8/li_65_n17# lvlshiftdown/li_826_79# FILLER_0_16/li_257_797# FILLER_1_0/li_545_n17#
+ lvlshiftdown/li_514_79# lvlshiftdown/li_257_1611# FILLER_0_8/li_353_797# FILLER_2_0/li_0_797#
+ FILLER_2_0/li_641_797# lvlshiftdown/li_1217_1611# FILLER_2_0/li_0_n17# lvlshiftdown/li_34_216#
+ lvlshiftdown/li_1601_1611# lvlshiftdown/li_641_1611# FILLER_0_0/li_0_797# FILLER_2_0/li_161_797#
+ lvlshiftdown/li_384_1039# lvlshiftdown/li_26_452# FILLER_1_0/li_0_n17# FILLER_2_8/li_0_797#
+ lvlshiftdown/li_756_683# FILLER_2_0/li_257_n17# FILLER_2_8/li_0_n17# lvlshiftdown/li_506_1123#
+ FILLER_1_8/li_0_n17# FILLER_0_16/li_65_797# FILLER_1_8/li_34_73# lvlshiftdown/li_545_1611#
+ lvlshiftdown/li_1505_1611# lvlshiftdown/m1_0_n23# lvlshiftdown/li_1505_797# FILLER_0_16/li_545_797#
+ FILLER_2_0/li_449_797# lvlshiftdown/li_161_797# FILLER_1_0/li_100_536# FILLER_0_0/li_353_797#
+ FILLER_0_8/li_641_797# lvlshiftdown/li_26_893# ANTENNA_lvlshiftdown_A/li_65_n17#
+ FILLER_0_16/li_115_72# lvlshiftdown/li_65_1611# FILLER_1_0/li_353_n17# FILLER_1_8/li_257_797#
+ FILLER_0_8/li_161_797# lvlshiftdown/li_0_797# FILLER_0_24/li_257_797# lvlshiftdown/li_1409_1611#
+ lvlshiftdown/li_449_1611# FILLER_0_24/li_65_797# lvlshiftdown/li_833_1611# FILLER_2_0/li_545_n17#
+ FILLER_0_0/li_65_797# lvlshiftdown/li_0_1611# FILLER_0_24/li_34_73# FILLER_1_8/li_257_n17#
+ FILLER_1_0/li_65_n17# FILLER_0_0/li_115_72# FILLER_0_8/li_449_797# lvlshiftdown/li_737_1611#
+ FILLER_0_8/li_100_536# FILLER_0_0/li_641_797# lvlshiftdown/m1_0_51# FILLER_0_16/li_353_797#
+ FILLER_2_0/li_257_797# FILLER_1_0/li_641_n17# FILLER_0_0/li_161_797# FILLER_0_24/li_50_537#
+ FILLER_1_0/li_161_n17# FILLER_2_0/li_65_797# FILLER_2_0/li_353_n17# FILLER_0_8/li_65_797#
+ FILLER_2_8/li_161_n17# FILLER_0_0/li_449_797# FILLER_0_0/li_100_536# FILLER_0_16/li_0_797#
+ FILLER_1_0/li_115_72# FILLER_1_0/li_449_n17# lvlshiftdown/li_1601_797# FILLER_0_8/li_257_797#
+ FILLER_0_16/li_641_797# FILLER_2_0/li_545_797# lvlshiftdown/li_929_1611# FILLER_0_16/li_161_797#
+ FILLER_0_8/li_115_72# FILLER_1_8/li_353_797# lvlshiftdown/li_34_1244# lvlshiftdown/li_161_1611#
+ FILLER_0_28/li_0_797# lvlshiftdown/li_1121_1611# FILLER_2_0/li_641_n17# FILLER_1_8/li_353_n17#
+ lvlshiftdown/li_179_1349# FILLER_2_0/li_65_n17# lvlshiftdown/m1_0_689# FILLER_2_0/li_161_n17#
+ FILLER_0_8/li_0_797# FILLER_2_8/li_65_797# ANTENNA_lvlshiftdown_A/li_0_n17# lvlshiftdown/li_179_79#
+ FILLER_1_8/li_65_n17# FILLER_0_16/li_449_797# lvlshiftdown/li_1025_1611# FILLER_0_16/li_100_536#
+ FILLER_0_0/li_257_797# lvlshiftdown/li_384_137# FILLER_2_0/li_115_72# FILLER_0_8/li_545_797#
+ FILLER_0_28/li_161_797# FILLER_1_0/li_257_n17# FILLER_2_0/li_100_536# lvlshiftdown/li_1455_797#
+ FILLER_2_0/li_353_797# FILLER_2_0/li_449_n17#
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_2
XFILLER_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
XFILLER_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
XANTENNA_lvlshiftdown_A A VGND VGND VPWR VPWR sky130_fd_sc_hvl__diode_2
XFILLER_2_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
XFILLER_0_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_8 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_2
Xlvlshiftdown A LVPWR VGND VGND VPWR VPWR X sky130_fd_sc_hvl__lsbufhv2lv_1
XFILLER_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
.ends

* Black-box entry subcircuit for user_project_wrapper abstract view
.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[29]
+ analog_io[2] analog_io[30] analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7]
+ analog_io[8] analog_io[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] user_clock2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2
.ends

* Black-box entry subcircuit for storage abstract view
.subckt storage mgmt_addr[0] mgmt_addr[1] mgmt_addr[2] mgmt_addr[3] mgmt_addr[4] mgmt_addr[5]
+ mgmt_addr[6] mgmt_addr[7] mgmt_addr_ro[0] mgmt_addr_ro[1] mgmt_addr_ro[2] mgmt_addr_ro[3]
+ mgmt_addr_ro[4] mgmt_addr_ro[5] mgmt_addr_ro[6] mgmt_addr_ro[7] mgmt_clk mgmt_ena[0]
+ mgmt_ena[1] mgmt_ena_ro mgmt_rdata[0] mgmt_rdata[10] mgmt_rdata[11] mgmt_rdata[12]
+ mgmt_rdata[13] mgmt_rdata[14] mgmt_rdata[15] mgmt_rdata[16] mgmt_rdata[17] mgmt_rdata[18]
+ mgmt_rdata[19] mgmt_rdata[1] mgmt_rdata[20] mgmt_rdata[21] mgmt_rdata[22] mgmt_rdata[23]
+ mgmt_rdata[24] mgmt_rdata[25] mgmt_rdata[26] mgmt_rdata[27] mgmt_rdata[28] mgmt_rdata[29]
+ mgmt_rdata[2] mgmt_rdata[30] mgmt_rdata[31] mgmt_rdata[32] mgmt_rdata[33] mgmt_rdata[34]
+ mgmt_rdata[35] mgmt_rdata[36] mgmt_rdata[37] mgmt_rdata[38] mgmt_rdata[39] mgmt_rdata[3]
+ mgmt_rdata[40] mgmt_rdata[41] mgmt_rdata[42] mgmt_rdata[43] mgmt_rdata[44] mgmt_rdata[45]
+ mgmt_rdata[46] mgmt_rdata[47] mgmt_rdata[48] mgmt_rdata[49] mgmt_rdata[4] mgmt_rdata[50]
+ mgmt_rdata[51] mgmt_rdata[52] mgmt_rdata[53] mgmt_rdata[54] mgmt_rdata[55] mgmt_rdata[56]
+ mgmt_rdata[57] mgmt_rdata[58] mgmt_rdata[59] mgmt_rdata[5] mgmt_rdata[60] mgmt_rdata[61]
+ mgmt_rdata[62] mgmt_rdata[63] mgmt_rdata[6] mgmt_rdata[7] mgmt_rdata[8] mgmt_rdata[9]
+ mgmt_rdata_ro[0] mgmt_rdata_ro[10] mgmt_rdata_ro[11] mgmt_rdata_ro[12] mgmt_rdata_ro[13]
+ mgmt_rdata_ro[14] mgmt_rdata_ro[15] mgmt_rdata_ro[16] mgmt_rdata_ro[17] mgmt_rdata_ro[18]
+ mgmt_rdata_ro[19] mgmt_rdata_ro[1] mgmt_rdata_ro[20] mgmt_rdata_ro[21] mgmt_rdata_ro[22]
+ mgmt_rdata_ro[23] mgmt_rdata_ro[24] mgmt_rdata_ro[25] mgmt_rdata_ro[26] mgmt_rdata_ro[27]
+ mgmt_rdata_ro[28] mgmt_rdata_ro[29] mgmt_rdata_ro[2] mgmt_rdata_ro[30] mgmt_rdata_ro[31]
+ mgmt_rdata_ro[3] mgmt_rdata_ro[4] mgmt_rdata_ro[5] mgmt_rdata_ro[6] mgmt_rdata_ro[7]
+ mgmt_rdata_ro[8] mgmt_rdata_ro[9] mgmt_wdata[0] mgmt_wdata[10] mgmt_wdata[11] mgmt_wdata[12]
+ mgmt_wdata[13] mgmt_wdata[14] mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17] mgmt_wdata[18]
+ mgmt_wdata[19] mgmt_wdata[1] mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23]
+ mgmt_wdata[24] mgmt_wdata[25] mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29]
+ mgmt_wdata[2] mgmt_wdata[30] mgmt_wdata[31] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5]
+ mgmt_wdata[6] mgmt_wdata[7] mgmt_wdata[8] mgmt_wdata[9] mgmt_wen[0] mgmt_wen[1]
+ mgmt_wen_mask[0] mgmt_wen_mask[1] mgmt_wen_mask[2] mgmt_wen_mask[3] mgmt_wen_mask[4]
+ mgmt_wen_mask[5] mgmt_wen_mask[6] mgmt_wen_mask[7] VPWR VGND
.ends

.subckt caravel clock flash_clk flash_csb flash_io0 flash_io1 gpio mprj_io[0] mprj_io[10]
+ mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16] mprj_io[17]
+ mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22] mprj_io[23]
+ mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29] mprj_io[2]
+ mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35] mprj_io[36]
+ mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9]
+ resetb vddio pwr_ctrl_out[0] pwr_ctrl_out[1] pwr_ctrl_out[2] pwr_ctrl_out[3] vccd1_pad
+ vccd2_pad vccd_pad vdda1_pad vdda2_pad vdda_pad vssa1_pad vssa2_pad vssa_pad vssd1_pad
+ vssd2_pad vssd_pad vssio_pad2
Xgpio_control_in\[28\] soc/mgmt_in_data[28] gpio_control_in\[28\]/one soc/mgmt_in_data[28]
+ gpio_control_in\[28\]/one padframe/mprj_io_analog_en[28] padframe/mprj_io_analog_pol[28]
+ padframe/mprj_io_analog_sel[28] padframe/mprj_io_dm[84] padframe/mprj_io_dm[85]
+ padframe/mprj_io_dm[86] padframe/mprj_io_holdover[28] padframe/mprj_io_ib_mode_sel[28]
+ padframe/mprj_io_in[28] padframe/mprj_io_inp_dis[28] padframe/mprj_io_out[28] padframe/mprj_io_oeb[28]
+ padframe/mprj_io_slow_sel[28] padframe/mprj_io_vtrip_sel[28] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[28\]/serial_data_in gpio_control_in\[29\]/serial_data_in
+ gpio_control_in\[28\]/user_gpio_in gpio_control_in\[28\]/user_gpio_oeb gpio_control_in\[28\]/user_gpio_out
+ gpio_control_in\[28\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[10\] soc/mgmt_in_data[10] gpio_control_in\[10\]/one soc/mgmt_in_data[10]
+ gpio_control_in\[10\]/one padframe/mprj_io_analog_en[10] padframe/mprj_io_analog_pol[10]
+ padframe/mprj_io_analog_sel[10] padframe/mprj_io_dm[30] padframe/mprj_io_dm[31]
+ padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10] padframe/mprj_io_ib_mode_sel[10]
+ padframe/mprj_io_in[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_out[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[9\]/serial_data_out gpio_control_in\[11\]/serial_data_in
+ gpio_control_in\[10\]/user_gpio_in gpio_control_in\[10\]/user_gpio_oeb gpio_control_in\[10\]/user_gpio_out
+ gpio_control_in\[10\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xpadframe clock soc/clock por/por_l flash_clk soc/flash_clk soc/flash_clk_ieb soc/flash_clk_oeb
+ flash_csb soc/flash_csb soc/flash_csb_ieb soc/flash_csb_oeb flash_io0 soc/flash_io0_di
+ soc/flash_io0_do padframe/flash_io0_ieb_core padframe/flash_io0_oeb_core flash_io1
+ soc/flash_io1_di soc/flash_io1_do padframe/flash_io1_ieb_core padframe/flash_io1_oeb_core
+ gpio soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad padframe/gpio_mode1_core
+ soc/gpio_out_pad soc/gpio_outenb_pad mprj_io[0] padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0]
+ padframe/mprj_io_analog_sel[0] padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2]
+ por/porb_h vddio padframe/mprj_io_holdover[0] padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_inp_dis[0]
+ padframe/mprj_io_oeb[0] padframe/mprj_io_out[0] padframe/mprj_io_slow_sel[0] padframe/mprj_io_vtrip_sel[0]
+ padframe/mprj_io_in[0] padframe/mprj_analog_io[3] mprj_io[10] padframe/mprj_io_analog_en[10]
+ padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10] padframe/mprj_io_dm[30]
+ padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] por/porb_h vddio padframe/mprj_io_holdover[10]
+ padframe/mprj_io_ib_mode_sel[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_out[10] padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10]
+ padframe/mprj_io_in[10] padframe/mprj_analog_io[4] mprj_io[11] padframe/mprj_io_analog_en[11]
+ padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11] padframe/mprj_io_dm[33]
+ padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] por/porb_h vddio padframe/mprj_io_holdover[11]
+ padframe/mprj_io_ib_mode_sel[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_out[11] padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11]
+ padframe/mprj_io_in[11] padframe/mprj_analog_io[5] mprj_io[12] padframe/mprj_io_analog_en[12]
+ padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12] padframe/mprj_io_dm[36]
+ padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] por/porb_h vddio padframe/mprj_io_holdover[12]
+ padframe/mprj_io_ib_mode_sel[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_out[12] padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12]
+ padframe/mprj_io_in[12] padframe/mprj_analog_io[6] mprj_io[13] padframe/mprj_io_analog_en[13]
+ padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13] padframe/mprj_io_dm[39]
+ padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] por/porb_h vddio padframe/mprj_io_holdover[13]
+ padframe/mprj_io_ib_mode_sel[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_out[13] padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13]
+ padframe/mprj_io_in[13] padframe/mprj_analog_io[7] mprj_io[14] padframe/mprj_io_analog_en[14]
+ padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14] padframe/mprj_io_dm[42]
+ padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] por/porb_h vddio padframe/mprj_io_holdover[14]
+ padframe/mprj_io_ib_mode_sel[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_out[14] padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14]
+ padframe/mprj_io_in[14] padframe/mprj_analog_io[8] mprj_io[15] padframe/mprj_io_analog_en[15]
+ padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15] padframe/mprj_io_dm[45]
+ padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] por/porb_h vddio padframe/mprj_io_holdover[15]
+ padframe/mprj_io_ib_mode_sel[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_out[15] padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15]
+ padframe/mprj_io_in[15] padframe/mprj_analog_io[9] mprj_io[16] padframe/mprj_io_analog_en[16]
+ padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16] padframe/mprj_io_dm[48]
+ padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] por/porb_h vddio padframe/mprj_io_holdover[16]
+ padframe/mprj_io_ib_mode_sel[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_out[16] padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16]
+ padframe/mprj_io_in[16] padframe/mprj_analog_io[10] mprj_io[17] padframe/mprj_io_analog_en[17]
+ padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17] padframe/mprj_io_dm[51]
+ padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] por/porb_h vddio padframe/mprj_io_holdover[17]
+ padframe/mprj_io_ib_mode_sel[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_out[17] padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17]
+ padframe/mprj_io_in[17] mprj_io[1] padframe/mprj_io_analog_en[1] padframe/mprj_io_analog_pol[1]
+ padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3] padframe/mprj_io_dm[4] padframe/mprj_io_dm[5]
+ por/porb_h vddio padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1] padframe/mprj_io_inp_dis[1]
+ padframe/mprj_io_oeb[1] padframe/mprj_io_out[1] padframe/mprj_io_slow_sel[1] padframe/mprj_io_vtrip_sel[1]
+ padframe/mprj_io_in[1] mprj_io[2] padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2]
+ padframe/mprj_io_analog_sel[2] padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8]
+ por/porb_h vddio padframe/mprj_io_holdover[2] padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_inp_dis[2]
+ padframe/mprj_io_oeb[2] padframe/mprj_io_out[2] padframe/mprj_io_slow_sel[2] padframe/mprj_io_vtrip_sel[2]
+ padframe/mprj_io_in[2] mprj_io[3] padframe/mprj_io_analog_en[3] padframe/mprj_io_analog_pol[3]
+ padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[10] padframe/mprj_io_dm[11] padframe/mprj_io_dm[9]
+ por/porb_h vddio padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3] padframe/mprj_io_inp_dis[3]
+ padframe/mprj_io_oeb[3] padframe/mprj_io_out[3] padframe/mprj_io_slow_sel[3] padframe/mprj_io_vtrip_sel[3]
+ padframe/mprj_io_in[3] mprj_io[4] padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4]
+ padframe/mprj_io_analog_sel[4] padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14]
+ por/porb_h vddio padframe/mprj_io_holdover[4] padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_inp_dis[4]
+ padframe/mprj_io_oeb[4] padframe/mprj_io_out[4] padframe/mprj_io_slow_sel[4] padframe/mprj_io_vtrip_sel[4]
+ padframe/mprj_io_in[4] mprj_io[5] padframe/mprj_io_analog_en[5] padframe/mprj_io_analog_pol[5]
+ padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15] padframe/mprj_io_dm[16] padframe/mprj_io_dm[17]
+ por/porb_h vddio padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5] padframe/mprj_io_inp_dis[5]
+ padframe/mprj_io_oeb[5] padframe/mprj_io_out[5] padframe/mprj_io_slow_sel[5] padframe/mprj_io_vtrip_sel[5]
+ padframe/mprj_io_in[5] mprj_io[6] padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6]
+ padframe/mprj_io_analog_sel[6] padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20]
+ por/porb_h vddio padframe/mprj_io_holdover[6] padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_inp_dis[6]
+ padframe/mprj_io_oeb[6] padframe/mprj_io_out[6] padframe/mprj_io_slow_sel[6] padframe/mprj_io_vtrip_sel[6]
+ padframe/mprj_io_in[6] padframe/mprj_analog_io[0] mprj_io[7] padframe/mprj_io_analog_en[7]
+ padframe/mprj_io_analog_pol[7] padframe/mprj_io_analog_sel[7] padframe/mprj_io_dm[21]
+ padframe/mprj_io_dm[22] padframe/mprj_io_dm[23] por/porb_h vddio padframe/mprj_io_holdover[7]
+ padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_inp_dis[7] padframe/mprj_io_oeb[7]
+ padframe/mprj_io_out[7] padframe/mprj_io_slow_sel[7] padframe/mprj_io_vtrip_sel[7]
+ padframe/mprj_io_in[7] padframe/mprj_analog_io[1] mprj_io[8] padframe/mprj_io_analog_en[8]
+ padframe/mprj_io_analog_pol[8] padframe/mprj_io_analog_sel[8] padframe/mprj_io_dm[24]
+ padframe/mprj_io_dm[25] padframe/mprj_io_dm[26] por/porb_h vddio padframe/mprj_io_holdover[8]
+ padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_inp_dis[8] padframe/mprj_io_oeb[8]
+ padframe/mprj_io_out[8] padframe/mprj_io_slow_sel[8] padframe/mprj_io_vtrip_sel[8]
+ padframe/mprj_io_in[8] padframe/mprj_analog_io[2] mprj_io[9] padframe/mprj_io_analog_en[9]
+ padframe/mprj_io_analog_pol[9] padframe/mprj_io_analog_sel[9] padframe/mprj_io_dm[27]
+ padframe/mprj_io_dm[28] padframe/mprj_io_dm[29] por/porb_h vddio padframe/mprj_io_holdover[9]
+ padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_inp_dis[9] padframe/mprj_io_oeb[9]
+ padframe/mprj_io_out[9] padframe/mprj_io_slow_sel[9] padframe/mprj_io_vtrip_sel[9]
+ padframe/mprj_io_in[9] padframe/mprj_analog_io[11] mprj_io[18] padframe/mprj_io_analog_en[18]
+ padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18] padframe/mprj_io_dm[54]
+ padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] por/porb_h vddio padframe/mprj_io_holdover[18]
+ padframe/mprj_io_ib_mode_sel[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_out[18] padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18]
+ padframe/mprj_io_in[18] padframe/mprj_analog_io[21] mprj_io[28] padframe/mprj_io_analog_en[28]
+ padframe/mprj_io_analog_pol[28] padframe/mprj_io_analog_sel[28] padframe/mprj_io_dm[84]
+ padframe/mprj_io_dm[85] padframe/mprj_io_dm[86] por/porb_h vddio padframe/mprj_io_holdover[28]
+ padframe/mprj_io_ib_mode_sel[28] padframe/mprj_io_inp_dis[28] padframe/mprj_io_oeb[28]
+ padframe/mprj_io_out[28] padframe/mprj_io_slow_sel[28] padframe/mprj_io_vtrip_sel[28]
+ padframe/mprj_io_in[28] padframe/mprj_analog_io[22] mprj_io[29] padframe/mprj_io_analog_en[29]
+ padframe/mprj_io_analog_pol[29] padframe/mprj_io_analog_sel[29] padframe/mprj_io_dm[87]
+ padframe/mprj_io_dm[88] padframe/mprj_io_dm[89] por/porb_h vddio padframe/mprj_io_holdover[29]
+ padframe/mprj_io_ib_mode_sel[29] padframe/mprj_io_inp_dis[29] padframe/mprj_io_oeb[29]
+ padframe/mprj_io_out[29] padframe/mprj_io_slow_sel[29] padframe/mprj_io_vtrip_sel[29]
+ padframe/mprj_io_in[29] padframe/mprj_analog_io[23] mprj_io[30] padframe/mprj_io_analog_en[30]
+ padframe/mprj_io_analog_pol[30] padframe/mprj_io_analog_sel[30] padframe/mprj_io_dm[90]
+ padframe/mprj_io_dm[91] padframe/mprj_io_dm[92] por/porb_h vddio padframe/mprj_io_holdover[30]
+ padframe/mprj_io_ib_mode_sel[30] padframe/mprj_io_inp_dis[30] padframe/mprj_io_oeb[30]
+ padframe/mprj_io_out[30] padframe/mprj_io_slow_sel[30] padframe/mprj_io_vtrip_sel[30]
+ padframe/mprj_io_in[30] padframe/mprj_analog_io[24] mprj_io[31] padframe/mprj_io_analog_en[31]
+ padframe/mprj_io_analog_pol[31] padframe/mprj_io_analog_sel[31] padframe/mprj_io_dm[93]
+ padframe/mprj_io_dm[94] padframe/mprj_io_dm[95] por/porb_h vddio padframe/mprj_io_holdover[31]
+ padframe/mprj_io_ib_mode_sel[31] padframe/mprj_io_inp_dis[31] padframe/mprj_io_oeb[31]
+ padframe/mprj_io_out[31] padframe/mprj_io_slow_sel[31] padframe/mprj_io_vtrip_sel[31]
+ padframe/mprj_io_in[31] padframe/mprj_analog_io[25] mprj_io[32] padframe/mprj_io_analog_en[32]
+ padframe/mprj_io_analog_pol[32] padframe/mprj_io_analog_sel[32] padframe/mprj_io_dm[96]
+ padframe/mprj_io_dm[97] padframe/mprj_io_dm[98] por/porb_h vddio padframe/mprj_io_holdover[32]
+ padframe/mprj_io_ib_mode_sel[32] padframe/mprj_io_inp_dis[32] padframe/mprj_io_oeb[32]
+ padframe/mprj_io_out[32] padframe/mprj_io_slow_sel[32] padframe/mprj_io_vtrip_sel[32]
+ padframe/mprj_io_in[32] padframe/mprj_analog_io[26] mprj_io[33] padframe/mprj_io_analog_en[33]
+ padframe/mprj_io_analog_pol[33] padframe/mprj_io_analog_sel[33] padframe/mprj_io_dm[100]
+ padframe/mprj_io_dm[101] padframe/mprj_io_dm[99] por/porb_h vddio padframe/mprj_io_holdover[33]
+ padframe/mprj_io_ib_mode_sel[33] padframe/mprj_io_inp_dis[33] padframe/mprj_io_oeb[33]
+ padframe/mprj_io_out[33] padframe/mprj_io_slow_sel[33] padframe/mprj_io_vtrip_sel[33]
+ padframe/mprj_io_in[33] padframe/mprj_analog_io[27] mprj_io[34] padframe/mprj_io_analog_en[34]
+ padframe/mprj_io_analog_pol[34] padframe/mprj_io_analog_sel[34] padframe/mprj_io_dm[102]
+ padframe/mprj_io_dm[103] padframe/mprj_io_dm[104] por/porb_h vddio padframe/mprj_io_holdover[34]
+ padframe/mprj_io_ib_mode_sel[34] padframe/mprj_io_inp_dis[34] padframe/mprj_io_oeb[34]
+ padframe/mprj_io_out[34] padframe/mprj_io_slow_sel[34] padframe/mprj_io_vtrip_sel[34]
+ padframe/mprj_io_in[34] padframe/mprj_analog_io[28] mprj_io[35] padframe/mprj_io_analog_en[35]
+ padframe/mprj_io_analog_pol[35] padframe/mprj_io_analog_sel[35] padframe/mprj_io_dm[105]
+ padframe/mprj_io_dm[106] padframe/mprj_io_dm[107] por/porb_h vddio padframe/mprj_io_holdover[35]
+ padframe/mprj_io_ib_mode_sel[35] padframe/mprj_io_inp_dis[35] padframe/mprj_io_oeb[35]
+ padframe/mprj_io_out[35] padframe/mprj_io_slow_sel[35] padframe/mprj_io_vtrip_sel[35]
+ padframe/mprj_io_in[35] padframe/mprj_analog_io[29] mprj_io[36] padframe/mprj_io_analog_en[36]
+ padframe/mprj_io_analog_pol[36] padframe/mprj_io_analog_sel[36] padframe/mprj_io_dm[108]
+ padframe/mprj_io_dm[109] padframe/mprj_io_dm[110] por/porb_h vddio padframe/mprj_io_holdover[36]
+ padframe/mprj_io_ib_mode_sel[36] padframe/mprj_io_inp_dis[36] padframe/mprj_io_oeb[36]
+ padframe/mprj_io_out[36] padframe/mprj_io_slow_sel[36] padframe/mprj_io_vtrip_sel[36]
+ padframe/mprj_io_in[36] padframe/mprj_analog_io[30] mprj_io[37] padframe/mprj_io_analog_en[37]
+ padframe/mprj_io_analog_pol[37] padframe/mprj_io_analog_sel[37] padframe/mprj_io_dm[111]
+ padframe/mprj_io_dm[112] padframe/mprj_io_dm[113] por/porb_h vddio padframe/mprj_io_holdover[37]
+ padframe/mprj_io_ib_mode_sel[37] padframe/mprj_io_inp_dis[37] padframe/mprj_io_oeb[37]
+ padframe/mprj_io_out[37] padframe/mprj_io_slow_sel[37] padframe/mprj_io_vtrip_sel[37]
+ padframe/mprj_io_in[37] padframe/mprj_analog_io[12] mprj_io[19] padframe/mprj_io_analog_en[19]
+ padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19] padframe/mprj_io_dm[57]
+ padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] por/porb_h vddio padframe/mprj_io_holdover[19]
+ padframe/mprj_io_ib_mode_sel[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_out[19] padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19]
+ padframe/mprj_io_in[19] padframe/mprj_analog_io[13] mprj_io[20] padframe/mprj_io_analog_en[20]
+ padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20] padframe/mprj_io_dm[60]
+ padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] por/porb_h vddio padframe/mprj_io_holdover[20]
+ padframe/mprj_io_ib_mode_sel[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_out[20] padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20]
+ padframe/mprj_io_in[20] padframe/mprj_analog_io[14] mprj_io[21] padframe/mprj_io_analog_en[21]
+ padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21] padframe/mprj_io_dm[63]
+ padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] por/porb_h vddio padframe/mprj_io_holdover[21]
+ padframe/mprj_io_ib_mode_sel[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_out[21] padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21]
+ padframe/mprj_io_in[21] padframe/mprj_analog_io[15] mprj_io[22] padframe/mprj_io_analog_en[22]
+ padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22] padframe/mprj_io_dm[66]
+ padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] por/porb_h vddio padframe/mprj_io_holdover[22]
+ padframe/mprj_io_ib_mode_sel[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_out[22] padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22]
+ padframe/mprj_io_in[22] padframe/mprj_analog_io[16] mprj_io[23] padframe/mprj_io_analog_en[23]
+ padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23] padframe/mprj_io_dm[69]
+ padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] por/porb_h vddio padframe/mprj_io_holdover[23]
+ padframe/mprj_io_ib_mode_sel[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_out[23] padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23]
+ padframe/mprj_io_in[23] padframe/mprj_analog_io[17] mprj_io[24] padframe/mprj_io_analog_en[24]
+ padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24] padframe/mprj_io_dm[72]
+ padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] por/porb_h vddio padframe/mprj_io_holdover[24]
+ padframe/mprj_io_ib_mode_sel[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_out[24] padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24]
+ padframe/mprj_io_in[24] padframe/mprj_analog_io[18] mprj_io[25] padframe/mprj_io_analog_en[25]
+ padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] por/porb_h vddio padframe/mprj_io_holdover[25]
+ padframe/mprj_io_ib_mode_sel[25] padframe/mprj_io_inp_dis[25] padframe/mprj_io_oeb[25]
+ padframe/mprj_io_out[25] padframe/mprj_io_slow_sel[25] padframe/mprj_io_vtrip_sel[25]
+ padframe/mprj_io_in[25] padframe/mprj_analog_io[19] mprj_io[26] padframe/mprj_io_analog_en[26]
+ padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26] padframe/mprj_io_dm[78]
+ padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] por/porb_h vddio padframe/mprj_io_holdover[26]
+ padframe/mprj_io_ib_mode_sel[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_out[26] padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26]
+ padframe/mprj_io_in[26] padframe/mprj_analog_io[20] mprj_io[27] padframe/mprj_io_analog_en[27]
+ padframe/mprj_io_analog_pol[27] padframe/mprj_io_analog_sel[27] padframe/mprj_io_dm[81]
+ padframe/mprj_io_dm[82] padframe/mprj_io_dm[83] por/porb_h vddio padframe/mprj_io_holdover[27]
+ padframe/mprj_io_ib_mode_sel[27] padframe/mprj_io_inp_dis[27] padframe/mprj_io_oeb[27]
+ padframe/mprj_io_out[27] padframe/mprj_io_slow_sel[27] padframe/mprj_io_vtrip_sel[27]
+ padframe/mprj_io_in[27] resetb padframe/porb_h rstb_level/A soc/VPWR mprj/vccd1
+ vccd1_pad mprj/vccd2 vccd2_pad vccd_pad padframe/vdda mprj/vdda1 vdda1_pad mprj/vdda2
+ vdda2_pad vdda_pad vddio padframe/vddio_pad padframe/vssa por/vss vssa1_pad por/vss
+ vssa2_pad vssa_pad por/vss mprj/vssd1 vssd1_pad mprj/vssd2 vssd2_pad vssd_pad por/vss
+ padframe/vssio_pad vssio_pad2 padframe/vddio_pad2 padframe/vssa1_pad2 padframe/vdda1_pad2
+ chip_io
Xgpio_control_in\[26\] soc/mgmt_in_data[26] gpio_control_in\[26\]/one soc/mgmt_in_data[26]
+ gpio_control_in\[26\]/one padframe/mprj_io_analog_en[26] padframe/mprj_io_analog_pol[26]
+ padframe/mprj_io_analog_sel[26] padframe/mprj_io_dm[78] padframe/mprj_io_dm[79]
+ padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26] padframe/mprj_io_ib_mode_sel[26]
+ padframe/mprj_io_in[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_out[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[26\]/serial_data_in gpio_control_in\[27\]/serial_data_in
+ gpio_control_in\[26\]/user_gpio_in gpio_control_in\[26\]/user_gpio_oeb gpio_control_in\[26\]/user_gpio_out
+ gpio_control_in\[26\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[33\] soc/mgmt_in_data[33] gpio_control_in\[33\]/one soc/mgmt_in_data[33]
+ gpio_control_in\[33\]/one padframe/mprj_io_analog_en[33] padframe/mprj_io_analog_pol[33]
+ padframe/mprj_io_analog_sel[33] padframe/mprj_io_dm[99] padframe/mprj_io_dm[100]
+ padframe/mprj_io_dm[101] padframe/mprj_io_holdover[33] padframe/mprj_io_ib_mode_sel[33]
+ padframe/mprj_io_in[33] padframe/mprj_io_inp_dis[33] padframe/mprj_io_out[33] padframe/mprj_io_oeb[33]
+ padframe/mprj_io_slow_sel[33] padframe/mprj_io_vtrip_sel[33] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[33\]/serial_data_in gpio_control_in\[34\]/serial_data_in
+ gpio_control_in\[33\]/user_gpio_in gpio_control_in\[33\]/user_gpio_oeb gpio_control_in\[33\]/user_gpio_out
+ gpio_control_in\[33\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xsoc soc/clock soc/user_clk soc/resetb soc/flash_clk soc/flash_clk_ieb soc/flash_clk_oeb
+ soc/flash_csb soc/flash_csb_ieb soc/flash_csb_oeb soc/flash_io0_di soc/flash_io0_do
+ soc/flash_io0_ieb soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_ieb
+ soc/flash_io1_oeb soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad soc/gpio_mode1_pad
+ soc/gpio_out_pad soc/gpio_outenb_pad soc/jtag_out soc/jtag_outenb soc/la_input[0]
+ soc/la_input[100] soc/la_input[101] soc/la_input[102] soc/la_input[103] soc/la_input[104]
+ soc/la_input[105] soc/la_input[106] soc/la_input[107] soc/la_input[108] soc/la_input[109]
+ soc/la_input[10] soc/la_input[110] soc/la_input[111] soc/la_input[112] soc/la_input[113]
+ soc/la_input[114] soc/la_input[115] soc/la_input[116] soc/la_input[117] soc/la_input[118]
+ soc/la_input[119] soc/la_input[11] soc/la_input[120] soc/la_input[121] soc/la_input[122]
+ soc/la_input[123] soc/la_input[124] soc/la_input[125] soc/la_input[126] soc/la_input[127]
+ soc/la_input[12] soc/la_input[13] soc/la_input[14] soc/la_input[15] soc/la_input[16]
+ soc/la_input[17] soc/la_input[18] soc/la_input[19] soc/la_input[1] soc/la_input[20]
+ soc/la_input[21] soc/la_input[22] soc/la_input[23] soc/la_input[24] soc/la_input[25]
+ soc/la_input[26] soc/la_input[27] soc/la_input[28] soc/la_input[29] soc/la_input[2]
+ soc/la_input[30] soc/la_input[31] soc/la_input[32] soc/la_input[33] soc/la_input[34]
+ soc/la_input[35] soc/la_input[36] soc/la_input[37] soc/la_input[38] soc/la_input[39]
+ soc/la_input[3] soc/la_input[40] soc/la_input[41] soc/la_input[42] soc/la_input[43]
+ soc/la_input[44] soc/la_input[45] soc/la_input[46] soc/la_input[47] soc/la_input[48]
+ soc/la_input[49] soc/la_input[4] soc/la_input[50] soc/la_input[51] soc/la_input[52]
+ soc/la_input[53] soc/la_input[54] soc/la_input[55] soc/la_input[56] soc/la_input[57]
+ soc/la_input[58] soc/la_input[59] soc/la_input[5] soc/la_input[60] soc/la_input[61]
+ soc/la_input[62] soc/la_input[63] soc/la_input[64] soc/la_input[65] soc/la_input[66]
+ soc/la_input[67] soc/la_input[68] soc/la_input[69] soc/la_input[6] soc/la_input[70]
+ soc/la_input[71] soc/la_input[72] soc/la_input[73] soc/la_input[74] soc/la_input[75]
+ soc/la_input[76] soc/la_input[77] soc/la_input[78] soc/la_input[79] soc/la_input[7]
+ soc/la_input[80] soc/la_input[81] soc/la_input[82] soc/la_input[83] soc/la_input[84]
+ soc/la_input[85] soc/la_input[86] soc/la_input[87] soc/la_input[88] soc/la_input[89]
+ soc/la_input[8] soc/la_input[90] soc/la_input[91] soc/la_input[92] soc/la_input[93]
+ soc/la_input[94] soc/la_input[95] soc/la_input[96] soc/la_input[97] soc/la_input[98]
+ soc/la_input[99] soc/la_input[9] soc/la_oen[0] soc/la_oen[100] soc/la_oen[101] soc/la_oen[102]
+ soc/la_oen[103] soc/la_oen[104] soc/la_oen[105] soc/la_oen[106] soc/la_oen[107]
+ soc/la_oen[108] soc/la_oen[109] soc/la_oen[10] soc/la_oen[110] soc/la_oen[111] soc/la_oen[112]
+ soc/la_oen[113] soc/la_oen[114] soc/la_oen[115] soc/la_oen[116] soc/la_oen[117]
+ soc/la_oen[118] soc/la_oen[119] soc/la_oen[11] soc/la_oen[120] soc/la_oen[121] soc/la_oen[122]
+ soc/la_oen[123] soc/la_oen[124] soc/la_oen[125] soc/la_oen[126] soc/la_oen[127]
+ soc/la_oen[12] soc/la_oen[13] soc/la_oen[14] soc/la_oen[15] soc/la_oen[16] soc/la_oen[17]
+ soc/la_oen[18] soc/la_oen[19] soc/la_oen[1] soc/la_oen[20] soc/la_oen[21] soc/la_oen[22]
+ soc/la_oen[23] soc/la_oen[24] soc/la_oen[25] soc/la_oen[26] soc/la_oen[27] soc/la_oen[28]
+ soc/la_oen[29] soc/la_oen[2] soc/la_oen[30] soc/la_oen[31] soc/la_oen[32] soc/la_oen[33]
+ soc/la_oen[34] soc/la_oen[35] soc/la_oen[36] soc/la_oen[37] soc/la_oen[38] soc/la_oen[39]
+ soc/la_oen[3] soc/la_oen[40] soc/la_oen[41] soc/la_oen[42] soc/la_oen[43] soc/la_oen[44]
+ soc/la_oen[45] soc/la_oen[46] soc/la_oen[47] soc/la_oen[48] soc/la_oen[49] soc/la_oen[4]
+ soc/la_oen[50] soc/la_oen[51] soc/la_oen[52] soc/la_oen[53] soc/la_oen[54] soc/la_oen[55]
+ soc/la_oen[56] soc/la_oen[57] soc/la_oen[58] soc/la_oen[59] soc/la_oen[5] soc/la_oen[60]
+ soc/la_oen[61] soc/la_oen[62] soc/la_oen[63] soc/la_oen[64] soc/la_oen[65] soc/la_oen[66]
+ soc/la_oen[67] soc/la_oen[68] soc/la_oen[69] soc/la_oen[6] soc/la_oen[70] soc/la_oen[71]
+ soc/la_oen[72] soc/la_oen[73] soc/la_oen[74] soc/la_oen[75] soc/la_oen[76] soc/la_oen[77]
+ soc/la_oen[78] soc/la_oen[79] soc/la_oen[7] soc/la_oen[80] soc/la_oen[81] soc/la_oen[82]
+ soc/la_oen[83] soc/la_oen[84] soc/la_oen[85] soc/la_oen[86] soc/la_oen[87] soc/la_oen[88]
+ soc/la_oen[89] soc/la_oen[8] soc/la_oen[90] soc/la_oen[91] soc/la_oen[92] soc/la_oen[93]
+ soc/la_oen[94] soc/la_oen[95] soc/la_oen[96] soc/la_oen[97] soc/la_oen[98] soc/la_oen[99]
+ soc/la_oen[9] soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102]
+ soc/la_output[103] soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107]
+ soc/la_output[108] soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111]
+ soc/la_output[112] soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116]
+ soc/la_output[117] soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120]
+ soc/la_output[121] soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125]
+ soc/la_output[126] soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14]
+ soc/la_output[15] soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19]
+ soc/la_output[1] soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23]
+ soc/la_output[24] soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28]
+ soc/la_output[29] soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32]
+ soc/la_output[33] soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37]
+ soc/la_output[38] soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41]
+ soc/la_output[42] soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46]
+ soc/la_output[47] soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50]
+ soc/la_output[51] soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55]
+ soc/la_output[56] soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5]
+ soc/la_output[60] soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64]
+ soc/la_output[65] soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69]
+ soc/la_output[6] soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73]
+ soc/la_output[74] soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78]
+ soc/la_output[79] soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82]
+ soc/la_output[83] soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87]
+ soc/la_output[88] soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91]
+ soc/la_output[92] soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96]
+ soc/la_output[97] soc/la_output[98] soc/la_output[99] soc/la_output[9] soc/mask_rev[0]
+ soc/mask_rev[10] soc/mask_rev[11] soc/mask_rev[12] soc/mask_rev[13] soc/mask_rev[14]
+ soc/mask_rev[15] soc/mask_rev[16] soc/mask_rev[17] soc/mask_rev[18] soc/mask_rev[19]
+ soc/mask_rev[1] soc/mask_rev[20] soc/mask_rev[21] soc/mask_rev[22] soc/mask_rev[23]
+ soc/mask_rev[24] soc/mask_rev[25] soc/mask_rev[26] soc/mask_rev[27] soc/mask_rev[28]
+ soc/mask_rev[29] soc/mask_rev[2] soc/mask_rev[30] soc/mask_rev[31] soc/mask_rev[3]
+ soc/mask_rev[4] soc/mask_rev[5] soc/mask_rev[6] soc/mask_rev[7] soc/mask_rev[8]
+ soc/mask_rev[9] soc/mgmt_addr[0] soc/mgmt_addr[1] soc/mgmt_addr[2] soc/mgmt_addr[3]
+ soc/mgmt_addr[4] soc/mgmt_addr[5] soc/mgmt_addr[6] soc/mgmt_addr[7] soc/mgmt_addr_ro[0]
+ soc/mgmt_addr_ro[1] soc/mgmt_addr_ro[2] soc/mgmt_addr_ro[3] soc/mgmt_addr_ro[4]
+ soc/mgmt_addr_ro[5] soc/mgmt_addr_ro[6] soc/mgmt_addr_ro[7] soc/mgmt_ena[0] soc/mgmt_ena[1]
+ soc/mgmt_ena_ro soc/mgmt_in_data[0] soc/mgmt_in_data[10] soc/mgmt_in_data[11] soc/mgmt_in_data[12]
+ soc/mgmt_in_data[13] soc/mgmt_in_data[14] soc/mgmt_in_data[15] soc/mgmt_in_data[16]
+ soc/mgmt_in_data[17] soc/mgmt_in_data[18] soc/mgmt_in_data[19] soc/mgmt_in_data[1]
+ soc/mgmt_in_data[20] soc/mgmt_in_data[21] soc/mgmt_in_data[22] soc/mgmt_in_data[23]
+ soc/mgmt_in_data[24] soc/mgmt_in_data[25] soc/mgmt_in_data[26] soc/mgmt_in_data[27]
+ soc/mgmt_in_data[28] soc/mgmt_in_data[29] soc/mgmt_in_data[2] soc/mgmt_in_data[30]
+ soc/mgmt_in_data[31] soc/mgmt_in_data[32] soc/mgmt_in_data[33] soc/mgmt_in_data[34]
+ soc/mgmt_in_data[35] soc/mgmt_in_data[36] soc/mgmt_in_data[37] soc/mgmt_in_data[3]
+ soc/mgmt_in_data[4] soc/mgmt_in_data[5] soc/mgmt_in_data[6] soc/mgmt_in_data[7]
+ soc/mgmt_in_data[8] soc/mgmt_in_data[9] soc/mgmt_out_data[0] soc/mgmt_in_data[10]
+ soc/mgmt_in_data[11] soc/mgmt_in_data[12] soc/mgmt_in_data[13] soc/mgmt_in_data[14]
+ soc/mgmt_in_data[15] soc/mgmt_in_data[16] soc/mgmt_in_data[17] soc/mgmt_in_data[18]
+ soc/mgmt_in_data[19] soc/mgmt_out_data[1] soc/mgmt_in_data[20] soc/mgmt_in_data[21]
+ soc/mgmt_in_data[22] soc/mgmt_in_data[23] soc/mgmt_in_data[24] soc/mgmt_in_data[25]
+ soc/mgmt_in_data[26] soc/mgmt_in_data[27] soc/mgmt_in_data[28] soc/mgmt_in_data[29]
+ soc/mgmt_in_data[2] soc/mgmt_in_data[30] soc/mgmt_in_data[31] soc/mgmt_in_data[32]
+ soc/mgmt_in_data[33] soc/mgmt_in_data[34] soc/mgmt_in_data[35] soc/mgmt_in_data[36]
+ soc/mgmt_in_data[37] soc/mgmt_in_data[3] soc/mgmt_in_data[4] soc/mgmt_in_data[5]
+ soc/mgmt_in_data[6] soc/mgmt_in_data[7] soc/mgmt_in_data[8] soc/mgmt_in_data[9]
+ soc/mgmt_rdata[0] soc/mgmt_rdata[10] soc/mgmt_rdata[11] soc/mgmt_rdata[12] soc/mgmt_rdata[13]
+ soc/mgmt_rdata[14] soc/mgmt_rdata[15] soc/mgmt_rdata[16] soc/mgmt_rdata[17] soc/mgmt_rdata[18]
+ soc/mgmt_rdata[19] soc/mgmt_rdata[1] soc/mgmt_rdata[20] soc/mgmt_rdata[21] soc/mgmt_rdata[22]
+ soc/mgmt_rdata[23] soc/mgmt_rdata[24] soc/mgmt_rdata[25] soc/mgmt_rdata[26] soc/mgmt_rdata[27]
+ soc/mgmt_rdata[28] soc/mgmt_rdata[29] soc/mgmt_rdata[2] soc/mgmt_rdata[30] soc/mgmt_rdata[31]
+ soc/mgmt_rdata[32] soc/mgmt_rdata[33] soc/mgmt_rdata[34] soc/mgmt_rdata[35] soc/mgmt_rdata[36]
+ soc/mgmt_rdata[37] soc/mgmt_rdata[38] soc/mgmt_rdata[39] soc/mgmt_rdata[3] soc/mgmt_rdata[40]
+ soc/mgmt_rdata[41] soc/mgmt_rdata[42] soc/mgmt_rdata[43] soc/mgmt_rdata[44] soc/mgmt_rdata[45]
+ soc/mgmt_rdata[46] soc/mgmt_rdata[47] soc/mgmt_rdata[48] soc/mgmt_rdata[49] soc/mgmt_rdata[4]
+ soc/mgmt_rdata[50] soc/mgmt_rdata[51] soc/mgmt_rdata[52] soc/mgmt_rdata[53] soc/mgmt_rdata[54]
+ soc/mgmt_rdata[55] soc/mgmt_rdata[56] soc/mgmt_rdata[57] soc/mgmt_rdata[58] soc/mgmt_rdata[59]
+ soc/mgmt_rdata[5] soc/mgmt_rdata[60] soc/mgmt_rdata[61] soc/mgmt_rdata[62] soc/mgmt_rdata[63]
+ soc/mgmt_rdata[6] soc/mgmt_rdata[7] soc/mgmt_rdata[8] soc/mgmt_rdata[9] soc/mgmt_rdata_ro[0]
+ soc/mgmt_rdata_ro[10] soc/mgmt_rdata_ro[11] soc/mgmt_rdata_ro[12] soc/mgmt_rdata_ro[13]
+ soc/mgmt_rdata_ro[14] soc/mgmt_rdata_ro[15] soc/mgmt_rdata_ro[16] soc/mgmt_rdata_ro[17]
+ soc/mgmt_rdata_ro[18] soc/mgmt_rdata_ro[19] soc/mgmt_rdata_ro[1] soc/mgmt_rdata_ro[20]
+ soc/mgmt_rdata_ro[21] soc/mgmt_rdata_ro[22] soc/mgmt_rdata_ro[23] soc/mgmt_rdata_ro[24]
+ soc/mgmt_rdata_ro[25] soc/mgmt_rdata_ro[26] soc/mgmt_rdata_ro[27] soc/mgmt_rdata_ro[28]
+ soc/mgmt_rdata_ro[29] soc/mgmt_rdata_ro[2] soc/mgmt_rdata_ro[30] soc/mgmt_rdata_ro[31]
+ soc/mgmt_rdata_ro[3] soc/mgmt_rdata_ro[4] soc/mgmt_rdata_ro[5] soc/mgmt_rdata_ro[6]
+ soc/mgmt_rdata_ro[7] soc/mgmt_rdata_ro[8] soc/mgmt_rdata_ro[9] soc/mgmt_wdata[0]
+ soc/mgmt_wdata[10] soc/mgmt_wdata[11] soc/mgmt_wdata[12] soc/mgmt_wdata[13] soc/mgmt_wdata[14]
+ soc/mgmt_wdata[15] soc/mgmt_wdata[16] soc/mgmt_wdata[17] soc/mgmt_wdata[18] soc/mgmt_wdata[19]
+ soc/mgmt_wdata[1] soc/mgmt_wdata[20] soc/mgmt_wdata[21] soc/mgmt_wdata[22] soc/mgmt_wdata[23]
+ soc/mgmt_wdata[24] soc/mgmt_wdata[25] soc/mgmt_wdata[26] soc/mgmt_wdata[27] soc/mgmt_wdata[28]
+ soc/mgmt_wdata[29] soc/mgmt_wdata[2] soc/mgmt_wdata[30] soc/mgmt_wdata[31] soc/mgmt_wdata[3]
+ soc/mgmt_wdata[4] soc/mgmt_wdata[5] soc/mgmt_wdata[6] soc/mgmt_wdata[7] soc/mgmt_wdata[8]
+ soc/mgmt_wdata[9] soc/mgmt_wen[0] soc/mgmt_wen[1] soc/mgmt_wen_mask[0] soc/mgmt_wen_mask[1]
+ soc/mgmt_wen_mask[2] soc/mgmt_wen_mask[3] soc/mgmt_wen_mask[4] soc/mgmt_wen_mask[5]
+ soc/mgmt_wen_mask[6] soc/mgmt_wen_mask[7] soc/mprj2_vcc_pwrgood soc/mprj2_vdd_pwrgood
+ soc/mprj_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12]
+ soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17]
+ soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21]
+ soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26]
+ soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30]
+ soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6]
+ soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9] soc/mprj_cyc_o soc/mprj_dat_i[0]
+ soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14]
+ soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19]
+ soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23]
+ soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28]
+ soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3]
+ soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8]
+ soc/mprj_dat_i[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12]
+ soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17]
+ soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21]
+ soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26]
+ soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30]
+ soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6]
+ soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/mprj_io_loader_clock soc/mprj_io_loader_data
+ soc/mprj_io_loader_resetn soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2]
+ soc/mprj_sel_o[3] soc/mprj_stb_o soc/mprj_vcc_pwrgood soc/mprj_vdd_pwrgood soc/mprj_we_o
+ soc/porb pwr_ctrl_out[0] pwr_ctrl_out[1] pwr_ctrl_out[2] pwr_ctrl_out[3] soc/resetb
+ soc/sdo_out soc/sdo_outenb soc/user_clk soc/VPWR por/vss mgmt_core
Xgpio_control_in\[19\] soc/mgmt_in_data[19] gpio_control_in\[19\]/one soc/mgmt_in_data[19]
+ gpio_control_in\[19\]/one padframe/mprj_io_analog_en[19] padframe/mprj_io_analog_pol[19]
+ padframe/mprj_io_analog_sel[19] padframe/mprj_io_dm[57] padframe/mprj_io_dm[58]
+ padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19] padframe/mprj_io_ib_mode_sel[19]
+ padframe/mprj_io_in[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_out[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[19\]/serial_data_in gpio_control_in\[20\]/serial_data_in
+ gpio_control_in\[19\]/user_gpio_in gpio_control_in\[19\]/user_gpio_oeb gpio_control_in\[19\]/user_gpio_out
+ gpio_control_in\[19\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[31\] soc/mgmt_in_data[31] gpio_control_in\[31\]/one soc/mgmt_in_data[31]
+ gpio_control_in\[31\]/one padframe/mprj_io_analog_en[31] padframe/mprj_io_analog_pol[31]
+ padframe/mprj_io_analog_sel[31] padframe/mprj_io_dm[93] padframe/mprj_io_dm[94]
+ padframe/mprj_io_dm[95] padframe/mprj_io_holdover[31] padframe/mprj_io_ib_mode_sel[31]
+ padframe/mprj_io_in[31] padframe/mprj_io_inp_dis[31] padframe/mprj_io_out[31] padframe/mprj_io_oeb[31]
+ padframe/mprj_io_slow_sel[31] padframe/mprj_io_vtrip_sel[31] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[31\]/serial_data_in gpio_control_in\[32\]/serial_data_in
+ gpio_control_in\[31\]/user_gpio_in gpio_control_in\[31\]/user_gpio_oeb gpio_control_in\[31\]/user_gpio_out
+ gpio_control_in\[31\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xpor vddio soc/VPWR por/vss por/porb_h por/por_l soc/porb simple_por
Xgpio_control_in\[24\] soc/mgmt_in_data[24] gpio_control_in\[24\]/one soc/mgmt_in_data[24]
+ gpio_control_in\[24\]/one padframe/mprj_io_analog_en[24] padframe/mprj_io_analog_pol[24]
+ padframe/mprj_io_analog_sel[24] padframe/mprj_io_dm[72] padframe/mprj_io_dm[73]
+ padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24] padframe/mprj_io_ib_mode_sel[24]
+ padframe/mprj_io_in[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_out[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[24\]/serial_data_in gpio_control_in\[25\]/serial_data_in
+ gpio_control_in\[24\]/user_gpio_in gpio_control_in\[24\]/user_gpio_oeb gpio_control_in\[24\]/user_gpio_out
+ gpio_control_in\[24\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_bidir\[1\] soc/mgmt_in_data[1] soc/sdo_outenb soc/sdo_out gpio_control_bidir\[1\]/one
+ padframe/mprj_io_analog_en[1] padframe/mprj_io_analog_pol[1] padframe/mprj_io_analog_sel[1]
+ padframe/mprj_io_dm[3] padframe/mprj_io_dm[4] padframe/mprj_io_dm[5] padframe/mprj_io_holdover[1]
+ padframe/mprj_io_ib_mode_sel[1] padframe/mprj_io_in[1] padframe/mprj_io_inp_dis[1]
+ padframe/mprj_io_out[1] padframe/mprj_io_oeb[1] padframe/mprj_io_slow_sel[1] padframe/mprj_io_vtrip_sel[1]
+ soc/mprj_io_loader_resetn soc/mprj_io_loader_clock gpio_control_bidir\[1\]/serial_data_in
+ gpio_control_in\[2\]/serial_data_in gpio_control_bidir\[1\]/user_gpio_in gpio_control_bidir\[1\]/user_gpio_oeb
+ gpio_control_bidir\[1\]/user_gpio_out gpio_control_bidir\[1\]/zero soc/VPWR por/vss
+ mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[17\] soc/mgmt_in_data[17] gpio_control_in\[17\]/one soc/mgmt_in_data[17]
+ gpio_control_in\[17\]/one padframe/mprj_io_analog_en[17] padframe/mprj_io_analog_pol[17]
+ padframe/mprj_io_analog_sel[17] padframe/mprj_io_dm[51] padframe/mprj_io_dm[52]
+ padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17] padframe/mprj_io_ib_mode_sel[17]
+ padframe/mprj_io_in[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_out[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[17\]/serial_data_in gpio_control_in\[18\]/serial_data_in
+ gpio_control_in\[17\]/user_gpio_in gpio_control_in\[17\]/user_gpio_oeb gpio_control_in\[17\]/user_gpio_out
+ gpio_control_in\[17\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[22\] soc/mgmt_in_data[22] gpio_control_in\[22\]/one soc/mgmt_in_data[22]
+ gpio_control_in\[22\]/one padframe/mprj_io_analog_en[22] padframe/mprj_io_analog_pol[22]
+ padframe/mprj_io_analog_sel[22] padframe/mprj_io_dm[66] padframe/mprj_io_dm[67]
+ padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22] padframe/mprj_io_ib_mode_sel[22]
+ padframe/mprj_io_in[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_out[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[22\]/serial_data_in gpio_control_in\[23\]/serial_data_in
+ gpio_control_in\[22\]/user_gpio_in gpio_control_in\[22\]/user_gpio_oeb gpio_control_in\[22\]/user_gpio_out
+ gpio_control_in\[22\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[8\] soc/mgmt_in_data[8] gpio_control_in\[8\]/one soc/mgmt_in_data[8]
+ gpio_control_in\[8\]/one padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8]
+ padframe/mprj_io_analog_sel[8] padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26]
+ padframe/mprj_io_holdover[8] padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_in[8]
+ padframe/mprj_io_inp_dis[8] padframe/mprj_io_out[8] padframe/mprj_io_oeb[8] padframe/mprj_io_slow_sel[8]
+ padframe/mprj_io_vtrip_sel[8] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[8\]/serial_data_in gpio_control_in\[9\]/serial_data_in gpio_control_in\[8\]/user_gpio_in
+ gpio_control_in\[8\]/user_gpio_oeb gpio_control_in\[8\]/user_gpio_out gpio_control_in\[8\]/zero
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[15\] soc/mgmt_in_data[15] gpio_control_in\[15\]/one soc/mgmt_in_data[15]
+ gpio_control_in\[15\]/one padframe/mprj_io_analog_en[15] padframe/mprj_io_analog_pol[15]
+ padframe/mprj_io_analog_sel[15] padframe/mprj_io_dm[45] padframe/mprj_io_dm[46]
+ padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15] padframe/mprj_io_ib_mode_sel[15]
+ padframe/mprj_io_in[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_out[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[15\]/serial_data_in gpio_control_in\[16\]/serial_data_in
+ gpio_control_in\[15\]/user_gpio_in gpio_control_in\[15\]/user_gpio_oeb gpio_control_in\[15\]/user_gpio_out
+ gpio_control_in\[15\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xuser_id_value soc/mask_rev[0] soc/mask_rev[10] soc/mask_rev[11] soc/mask_rev[12]
+ soc/mask_rev[13] soc/mask_rev[14] soc/mask_rev[15] soc/mask_rev[16] soc/mask_rev[17]
+ soc/mask_rev[18] soc/mask_rev[19] soc/mask_rev[1] soc/mask_rev[20] soc/mask_rev[21]
+ soc/mask_rev[22] soc/mask_rev[23] soc/mask_rev[24] soc/mask_rev[25] soc/mask_rev[26]
+ soc/mask_rev[27] soc/mask_rev[28] soc/mask_rev[29] soc/mask_rev[2] soc/mask_rev[30]
+ soc/mask_rev[31] soc/mask_rev[3] soc/mask_rev[4] soc/mask_rev[5] soc/mask_rev[6]
+ soc/mask_rev[7] soc/mask_rev[8] soc/mask_rev[9] soc/VPWR por/vss user_id_programming
Xgpio_control_in\[20\] soc/mgmt_in_data[20] gpio_control_in\[20\]/one soc/mgmt_in_data[20]
+ gpio_control_in\[20\]/one padframe/mprj_io_analog_en[20] padframe/mprj_io_analog_pol[20]
+ padframe/mprj_io_analog_sel[20] padframe/mprj_io_dm[60] padframe/mprj_io_dm[61]
+ padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20] padframe/mprj_io_ib_mode_sel[20]
+ padframe/mprj_io_in[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_out[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[20\]/serial_data_in gpio_control_in\[21\]/serial_data_in
+ gpio_control_in\[20\]/user_gpio_in gpio_control_in\[20\]/user_gpio_oeb gpio_control_in\[20\]/user_gpio_out
+ gpio_control_in\[20\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[6\] soc/mgmt_in_data[6] gpio_control_in\[6\]/one soc/mgmt_in_data[6]
+ gpio_control_in\[6\]/one padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6]
+ padframe/mprj_io_analog_sel[6] padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20]
+ padframe/mprj_io_holdover[6] padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_in[6]
+ padframe/mprj_io_inp_dis[6] padframe/mprj_io_out[6] padframe/mprj_io_oeb[6] padframe/mprj_io_slow_sel[6]
+ padframe/mprj_io_vtrip_sel[6] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[6\]/serial_data_in gpio_control_in\[7\]/serial_data_in gpio_control_in\[6\]/user_gpio_in
+ gpio_control_in\[6\]/user_gpio_oeb gpio_control_in\[6\]/user_gpio_out gpio_control_in\[6\]/zero
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[13\] soc/mgmt_in_data[13] gpio_control_in\[13\]/one soc/mgmt_in_data[13]
+ gpio_control_in\[13\]/one padframe/mprj_io_analog_en[13] padframe/mprj_io_analog_pol[13]
+ padframe/mprj_io_analog_sel[13] padframe/mprj_io_dm[39] padframe/mprj_io_dm[40]
+ padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13] padframe/mprj_io_ib_mode_sel[13]
+ padframe/mprj_io_in[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_out[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[13\]/serial_data_in gpio_control_in\[14\]/serial_data_in
+ gpio_control_in\[13\]/user_gpio_in gpio_control_in\[13\]/user_gpio_oeb gpio_control_in\[13\]/user_gpio_out
+ gpio_control_in\[13\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[36\] soc/mgmt_in_data[36] gpio_control_in\[36\]/one soc/mgmt_in_data[36]
+ gpio_control_in\[36\]/one padframe/mprj_io_analog_en[36] padframe/mprj_io_analog_pol[36]
+ padframe/mprj_io_analog_sel[36] padframe/mprj_io_dm[108] padframe/mprj_io_dm[109]
+ padframe/mprj_io_dm[110] padframe/mprj_io_holdover[36] padframe/mprj_io_ib_mode_sel[36]
+ padframe/mprj_io_in[36] padframe/mprj_io_inp_dis[36] padframe/mprj_io_out[36] padframe/mprj_io_oeb[36]
+ padframe/mprj_io_slow_sel[36] padframe/mprj_io_vtrip_sel[36] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[36\]/serial_data_in gpio_control_in\[37\]/serial_data_in
+ gpio_control_in\[36\]/user_gpio_in gpio_control_in\[36\]/user_gpio_oeb gpio_control_in\[36\]/user_gpio_out
+ gpio_control_in\[36\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[29\] soc/mgmt_in_data[29] gpio_control_in\[29\]/one soc/mgmt_in_data[29]
+ gpio_control_in\[29\]/one padframe/mprj_io_analog_en[29] padframe/mprj_io_analog_pol[29]
+ padframe/mprj_io_analog_sel[29] padframe/mprj_io_dm[87] padframe/mprj_io_dm[88]
+ padframe/mprj_io_dm[89] padframe/mprj_io_holdover[29] padframe/mprj_io_ib_mode_sel[29]
+ padframe/mprj_io_in[29] padframe/mprj_io_inp_dis[29] padframe/mprj_io_out[29] padframe/mprj_io_oeb[29]
+ padframe/mprj_io_slow_sel[29] padframe/mprj_io_vtrip_sel[29] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[29\]/serial_data_in gpio_control_in\[30\]/serial_data_in
+ gpio_control_in\[29\]/user_gpio_in gpio_control_in\[29\]/user_gpio_oeb gpio_control_in\[29\]/user_gpio_out
+ gpio_control_in\[29\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[4\] soc/mgmt_in_data[4] gpio_control_in\[4\]/one soc/mgmt_in_data[4]
+ gpio_control_in\[4\]/one padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4]
+ padframe/mprj_io_analog_sel[4] padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14]
+ padframe/mprj_io_holdover[4] padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_in[4]
+ padframe/mprj_io_inp_dis[4] padframe/mprj_io_out[4] padframe/mprj_io_oeb[4] padframe/mprj_io_slow_sel[4]
+ padframe/mprj_io_vtrip_sel[4] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[4\]/serial_data_in gpio_control_in\[5\]/serial_data_in gpio_control_in\[4\]/user_gpio_in
+ gpio_control_in\[4\]/user_gpio_oeb gpio_control_in\[4\]/user_gpio_out gpio_control_in\[4\]/zero
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[11\] soc/mgmt_in_data[11] gpio_control_in\[11\]/one soc/mgmt_in_data[11]
+ gpio_control_in\[11\]/one padframe/mprj_io_analog_en[11] padframe/mprj_io_analog_pol[11]
+ padframe/mprj_io_analog_sel[11] padframe/mprj_io_dm[33] padframe/mprj_io_dm[34]
+ padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11] padframe/mprj_io_ib_mode_sel[11]
+ padframe/mprj_io_in[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_out[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[11\]/serial_data_in gpio_control_in\[12\]/serial_data_in
+ gpio_control_in\[11\]/user_gpio_in gpio_control_in\[11\]/user_gpio_oeb gpio_control_in\[11\]/user_gpio_out
+ gpio_control_in\[11\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[34\] soc/mgmt_in_data[34] gpio_control_in\[34\]/one soc/mgmt_in_data[34]
+ gpio_control_in\[34\]/one padframe/mprj_io_analog_en[34] padframe/mprj_io_analog_pol[34]
+ padframe/mprj_io_analog_sel[34] padframe/mprj_io_dm[102] padframe/mprj_io_dm[103]
+ padframe/mprj_io_dm[104] padframe/mprj_io_holdover[34] padframe/mprj_io_ib_mode_sel[34]
+ padframe/mprj_io_in[34] padframe/mprj_io_inp_dis[34] padframe/mprj_io_out[34] padframe/mprj_io_oeb[34]
+ padframe/mprj_io_slow_sel[34] padframe/mprj_io_vtrip_sel[34] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[34\]/serial_data_in gpio_control_in\[35\]/serial_data_in
+ gpio_control_in\[34\]/user_gpio_in gpio_control_in\[34\]/user_gpio_oeb gpio_control_in\[34\]/user_gpio_out
+ gpio_control_in\[34\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xmgmt_buffers soc/user_clk soc/user_clk soc/resetb mgmt_buffers/la_data_in_core[0]
+ mgmt_buffers/la_data_in_core[100] mgmt_buffers/la_data_in_core[101] mgmt_buffers/la_data_in_core[102]
+ mgmt_buffers/la_data_in_core[103] mgmt_buffers/la_data_in_core[104] mgmt_buffers/la_data_in_core[105]
+ mgmt_buffers/la_data_in_core[106] mgmt_buffers/la_data_in_core[107] mgmt_buffers/la_data_in_core[108]
+ mgmt_buffers/la_data_in_core[109] mgmt_buffers/la_data_in_core[10] mgmt_buffers/la_data_in_core[110]
+ mgmt_buffers/la_data_in_core[111] mgmt_buffers/la_data_in_core[112] mgmt_buffers/la_data_in_core[113]
+ mgmt_buffers/la_data_in_core[114] mgmt_buffers/la_data_in_core[115] mgmt_buffers/la_data_in_core[116]
+ mgmt_buffers/la_data_in_core[117] mgmt_buffers/la_data_in_core[118] mgmt_buffers/la_data_in_core[119]
+ mgmt_buffers/la_data_in_core[11] mgmt_buffers/la_data_in_core[120] mgmt_buffers/la_data_in_core[121]
+ mgmt_buffers/la_data_in_core[122] mgmt_buffers/la_data_in_core[123] mgmt_buffers/la_data_in_core[124]
+ mgmt_buffers/la_data_in_core[125] mgmt_buffers/la_data_in_core[126] mgmt_buffers/la_data_in_core[127]
+ mgmt_buffers/la_data_in_core[12] mgmt_buffers/la_data_in_core[13] mgmt_buffers/la_data_in_core[14]
+ mgmt_buffers/la_data_in_core[15] mgmt_buffers/la_data_in_core[16] mgmt_buffers/la_data_in_core[17]
+ mgmt_buffers/la_data_in_core[18] mgmt_buffers/la_data_in_core[19] mgmt_buffers/la_data_in_core[1]
+ mgmt_buffers/la_data_in_core[20] mgmt_buffers/la_data_in_core[21] mgmt_buffers/la_data_in_core[22]
+ mgmt_buffers/la_data_in_core[23] mgmt_buffers/la_data_in_core[24] mgmt_buffers/la_data_in_core[25]
+ mgmt_buffers/la_data_in_core[26] mgmt_buffers/la_data_in_core[27] mgmt_buffers/la_data_in_core[28]
+ mgmt_buffers/la_data_in_core[29] mgmt_buffers/la_data_in_core[2] mgmt_buffers/la_data_in_core[30]
+ mgmt_buffers/la_data_in_core[31] mgmt_buffers/la_data_in_core[32] mgmt_buffers/la_data_in_core[33]
+ mgmt_buffers/la_data_in_core[34] mgmt_buffers/la_data_in_core[35] mgmt_buffers/la_data_in_core[36]
+ mgmt_buffers/la_data_in_core[37] mgmt_buffers/la_data_in_core[38] mgmt_buffers/la_data_in_core[39]
+ mgmt_buffers/la_data_in_core[3] mgmt_buffers/la_data_in_core[40] mgmt_buffers/la_data_in_core[41]
+ mgmt_buffers/la_data_in_core[42] mgmt_buffers/la_data_in_core[43] mgmt_buffers/la_data_in_core[44]
+ mgmt_buffers/la_data_in_core[45] mgmt_buffers/la_data_in_core[46] mgmt_buffers/la_data_in_core[47]
+ mgmt_buffers/la_data_in_core[48] mgmt_buffers/la_data_in_core[49] mgmt_buffers/la_data_in_core[4]
+ mgmt_buffers/la_data_in_core[50] mgmt_buffers/la_data_in_core[51] mgmt_buffers/la_data_in_core[52]
+ mgmt_buffers/la_data_in_core[53] mgmt_buffers/la_data_in_core[54] mgmt_buffers/la_data_in_core[55]
+ mgmt_buffers/la_data_in_core[56] mgmt_buffers/la_data_in_core[57] mgmt_buffers/la_data_in_core[58]
+ mgmt_buffers/la_data_in_core[59] mgmt_buffers/la_data_in_core[5] mgmt_buffers/la_data_in_core[60]
+ mgmt_buffers/la_data_in_core[61] mgmt_buffers/la_data_in_core[62] mgmt_buffers/la_data_in_core[63]
+ mgmt_buffers/la_data_in_core[64] mgmt_buffers/la_data_in_core[65] mgmt_buffers/la_data_in_core[66]
+ mgmt_buffers/la_data_in_core[67] mgmt_buffers/la_data_in_core[68] mgmt_buffers/la_data_in_core[69]
+ mgmt_buffers/la_data_in_core[6] mgmt_buffers/la_data_in_core[70] mgmt_buffers/la_data_in_core[71]
+ mgmt_buffers/la_data_in_core[72] mgmt_buffers/la_data_in_core[73] mgmt_buffers/la_data_in_core[74]
+ mgmt_buffers/la_data_in_core[75] mgmt_buffers/la_data_in_core[76] mgmt_buffers/la_data_in_core[77]
+ mgmt_buffers/la_data_in_core[78] mgmt_buffers/la_data_in_core[79] mgmt_buffers/la_data_in_core[7]
+ mgmt_buffers/la_data_in_core[80] mgmt_buffers/la_data_in_core[81] mgmt_buffers/la_data_in_core[82]
+ mgmt_buffers/la_data_in_core[83] mgmt_buffers/la_data_in_core[84] mgmt_buffers/la_data_in_core[85]
+ mgmt_buffers/la_data_in_core[86] mgmt_buffers/la_data_in_core[87] mgmt_buffers/la_data_in_core[88]
+ mgmt_buffers/la_data_in_core[89] mgmt_buffers/la_data_in_core[8] mgmt_buffers/la_data_in_core[90]
+ mgmt_buffers/la_data_in_core[91] mgmt_buffers/la_data_in_core[92] mgmt_buffers/la_data_in_core[93]
+ mgmt_buffers/la_data_in_core[94] mgmt_buffers/la_data_in_core[95] mgmt_buffers/la_data_in_core[96]
+ mgmt_buffers/la_data_in_core[97] mgmt_buffers/la_data_in_core[98] mgmt_buffers/la_data_in_core[99]
+ mgmt_buffers/la_data_in_core[9] soc/la_input[0] soc/la_input[100] soc/la_input[101]
+ soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105] soc/la_input[106]
+ soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10] soc/la_input[110]
+ soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114] soc/la_input[115]
+ soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119] soc/la_input[11]
+ soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123] soc/la_input[124]
+ soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67] soc/la_input[68]
+ soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71] soc/la_input[72]
+ soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76] soc/la_input[77]
+ soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80] soc/la_input[81]
+ soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85] soc/la_input[86]
+ soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8] soc/la_input[90]
+ soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94] soc/la_input[95]
+ soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99] soc/la_input[9]
+ mgmt_buffers/la_data_out_core[0] mgmt_buffers/la_data_out_core[100] mgmt_buffers/la_data_out_core[101]
+ mgmt_buffers/la_data_out_core[102] mgmt_buffers/la_data_out_core[103] mgmt_buffers/la_data_out_core[104]
+ mgmt_buffers/la_data_out_core[105] mgmt_buffers/la_data_out_core[106] mgmt_buffers/la_data_out_core[107]
+ mgmt_buffers/la_data_out_core[108] mgmt_buffers/la_data_out_core[109] mgmt_buffers/la_data_out_core[10]
+ mgmt_buffers/la_data_out_core[110] mgmt_buffers/la_data_out_core[111] mgmt_buffers/la_data_out_core[112]
+ mgmt_buffers/la_data_out_core[113] mgmt_buffers/la_data_out_core[114] mgmt_buffers/la_data_out_core[115]
+ mgmt_buffers/la_data_out_core[116] mgmt_buffers/la_data_out_core[117] mgmt_buffers/la_data_out_core[118]
+ mgmt_buffers/la_data_out_core[119] mgmt_buffers/la_data_out_core[11] mgmt_buffers/la_data_out_core[120]
+ mgmt_buffers/la_data_out_core[121] mgmt_buffers/la_data_out_core[122] mgmt_buffers/la_data_out_core[123]
+ mgmt_buffers/la_data_out_core[124] mgmt_buffers/la_data_out_core[125] mgmt_buffers/la_data_out_core[126]
+ mgmt_buffers/la_data_out_core[127] mgmt_buffers/la_data_out_core[12] mgmt_buffers/la_data_out_core[13]
+ mgmt_buffers/la_data_out_core[14] mgmt_buffers/la_data_out_core[15] mgmt_buffers/la_data_out_core[16]
+ mgmt_buffers/la_data_out_core[17] mgmt_buffers/la_data_out_core[18] mgmt_buffers/la_data_out_core[19]
+ mgmt_buffers/la_data_out_core[1] mgmt_buffers/la_data_out_core[20] mgmt_buffers/la_data_out_core[21]
+ mgmt_buffers/la_data_out_core[22] mgmt_buffers/la_data_out_core[23] mgmt_buffers/la_data_out_core[24]
+ mgmt_buffers/la_data_out_core[25] mgmt_buffers/la_data_out_core[26] mgmt_buffers/la_data_out_core[27]
+ mgmt_buffers/la_data_out_core[28] mgmt_buffers/la_data_out_core[29] mgmt_buffers/la_data_out_core[2]
+ mgmt_buffers/la_data_out_core[30] mgmt_buffers/la_data_out_core[31] mgmt_buffers/la_data_out_core[32]
+ mgmt_buffers/la_data_out_core[33] mgmt_buffers/la_data_out_core[34] mgmt_buffers/la_data_out_core[35]
+ mgmt_buffers/la_data_out_core[36] mgmt_buffers/la_data_out_core[37] mgmt_buffers/la_data_out_core[38]
+ mgmt_buffers/la_data_out_core[39] mgmt_buffers/la_data_out_core[3] mgmt_buffers/la_data_out_core[40]
+ mgmt_buffers/la_data_out_core[41] mgmt_buffers/la_data_out_core[42] mgmt_buffers/la_data_out_core[43]
+ mgmt_buffers/la_data_out_core[44] mgmt_buffers/la_data_out_core[45] mgmt_buffers/la_data_out_core[46]
+ mgmt_buffers/la_data_out_core[47] mgmt_buffers/la_data_out_core[48] mgmt_buffers/la_data_out_core[49]
+ mgmt_buffers/la_data_out_core[4] mgmt_buffers/la_data_out_core[50] mgmt_buffers/la_data_out_core[51]
+ mgmt_buffers/la_data_out_core[52] mgmt_buffers/la_data_out_core[53] mgmt_buffers/la_data_out_core[54]
+ mgmt_buffers/la_data_out_core[55] mgmt_buffers/la_data_out_core[56] mgmt_buffers/la_data_out_core[57]
+ mgmt_buffers/la_data_out_core[58] mgmt_buffers/la_data_out_core[59] mgmt_buffers/la_data_out_core[5]
+ mgmt_buffers/la_data_out_core[60] mgmt_buffers/la_data_out_core[61] mgmt_buffers/la_data_out_core[62]
+ mgmt_buffers/la_data_out_core[63] mgmt_buffers/la_data_out_core[64] mgmt_buffers/la_data_out_core[65]
+ mgmt_buffers/la_data_out_core[66] mgmt_buffers/la_data_out_core[67] mgmt_buffers/la_data_out_core[68]
+ mgmt_buffers/la_data_out_core[69] mgmt_buffers/la_data_out_core[6] mgmt_buffers/la_data_out_core[70]
+ mgmt_buffers/la_data_out_core[71] mgmt_buffers/la_data_out_core[72] mgmt_buffers/la_data_out_core[73]
+ mgmt_buffers/la_data_out_core[74] mgmt_buffers/la_data_out_core[75] mgmt_buffers/la_data_out_core[76]
+ mgmt_buffers/la_data_out_core[77] mgmt_buffers/la_data_out_core[78] mgmt_buffers/la_data_out_core[79]
+ mgmt_buffers/la_data_out_core[7] mgmt_buffers/la_data_out_core[80] mgmt_buffers/la_data_out_core[81]
+ mgmt_buffers/la_data_out_core[82] mgmt_buffers/la_data_out_core[83] mgmt_buffers/la_data_out_core[84]
+ mgmt_buffers/la_data_out_core[85] mgmt_buffers/la_data_out_core[86] mgmt_buffers/la_data_out_core[87]
+ mgmt_buffers/la_data_out_core[88] mgmt_buffers/la_data_out_core[89] mgmt_buffers/la_data_out_core[8]
+ mgmt_buffers/la_data_out_core[90] mgmt_buffers/la_data_out_core[91] mgmt_buffers/la_data_out_core[92]
+ mgmt_buffers/la_data_out_core[93] mgmt_buffers/la_data_out_core[94] mgmt_buffers/la_data_out_core[95]
+ mgmt_buffers/la_data_out_core[96] mgmt_buffers/la_data_out_core[97] mgmt_buffers/la_data_out_core[98]
+ mgmt_buffers/la_data_out_core[99] mgmt_buffers/la_data_out_core[9] soc/la_output[0]
+ soc/la_output[100] soc/la_output[101] soc/la_output[102] soc/la_output[103] soc/la_output[104]
+ soc/la_output[105] soc/la_output[106] soc/la_output[107] soc/la_output[108] soc/la_output[109]
+ soc/la_output[10] soc/la_output[110] soc/la_output[111] soc/la_output[112] soc/la_output[113]
+ soc/la_output[114] soc/la_output[115] soc/la_output[116] soc/la_output[117] soc/la_output[118]
+ soc/la_output[119] soc/la_output[11] soc/la_output[120] soc/la_output[121] soc/la_output[122]
+ soc/la_output[123] soc/la_output[124] soc/la_output[125] soc/la_output[126] soc/la_output[127]
+ soc/la_output[12] soc/la_output[13] soc/la_output[14] soc/la_output[15] soc/la_output[16]
+ soc/la_output[17] soc/la_output[18] soc/la_output[19] soc/la_output[1] soc/la_output[20]
+ soc/la_output[21] soc/la_output[22] soc/la_output[23] soc/la_output[24] soc/la_output[25]
+ soc/la_output[26] soc/la_output[27] soc/la_output[28] soc/la_output[29] soc/la_output[2]
+ soc/la_output[30] soc/la_output[31] soc/la_output[32] soc/la_output[33] soc/la_output[34]
+ soc/la_output[35] soc/la_output[36] soc/la_output[37] soc/la_output[38] soc/la_output[39]
+ soc/la_output[3] soc/la_output[40] soc/la_output[41] soc/la_output[42] soc/la_output[43]
+ soc/la_output[44] soc/la_output[45] soc/la_output[46] soc/la_output[47] soc/la_output[48]
+ soc/la_output[49] soc/la_output[4] soc/la_output[50] soc/la_output[51] soc/la_output[52]
+ soc/la_output[53] soc/la_output[54] soc/la_output[55] soc/la_output[56] soc/la_output[57]
+ soc/la_output[58] soc/la_output[59] soc/la_output[5] soc/la_output[60] soc/la_output[61]
+ soc/la_output[62] soc/la_output[63] soc/la_output[64] soc/la_output[65] soc/la_output[66]
+ soc/la_output[67] soc/la_output[68] soc/la_output[69] soc/la_output[6] soc/la_output[70]
+ soc/la_output[71] soc/la_output[72] soc/la_output[73] soc/la_output[74] soc/la_output[75]
+ soc/la_output[76] soc/la_output[77] soc/la_output[78] soc/la_output[79] soc/la_output[7]
+ soc/la_output[80] soc/la_output[81] soc/la_output[82] soc/la_output[83] soc/la_output[84]
+ soc/la_output[85] soc/la_output[86] soc/la_output[87] soc/la_output[88] soc/la_output[89]
+ soc/la_output[8] soc/la_output[90] soc/la_output[91] soc/la_output[92] soc/la_output[93]
+ soc/la_output[94] soc/la_output[95] soc/la_output[96] soc/la_output[97] soc/la_output[98]
+ soc/la_output[99] soc/la_output[9] mgmt_buffers/la_oen_core[0] mgmt_buffers/la_oen_core[100]
+ mgmt_buffers/la_oen_core[101] mgmt_buffers/la_oen_core[102] mgmt_buffers/la_oen_core[103]
+ mgmt_buffers/la_oen_core[104] mgmt_buffers/la_oen_core[105] mgmt_buffers/la_oen_core[106]
+ mgmt_buffers/la_oen_core[107] mgmt_buffers/la_oen_core[108] mgmt_buffers/la_oen_core[109]
+ mgmt_buffers/la_oen_core[10] mgmt_buffers/la_oen_core[110] mgmt_buffers/la_oen_core[111]
+ mgmt_buffers/la_oen_core[112] mgmt_buffers/la_oen_core[113] mgmt_buffers/la_oen_core[114]
+ mgmt_buffers/la_oen_core[115] mgmt_buffers/la_oen_core[116] mgmt_buffers/la_oen_core[117]
+ mgmt_buffers/la_oen_core[118] mgmt_buffers/la_oen_core[119] mgmt_buffers/la_oen_core[11]
+ mgmt_buffers/la_oen_core[120] mgmt_buffers/la_oen_core[121] mgmt_buffers/la_oen_core[122]
+ mgmt_buffers/la_oen_core[123] mgmt_buffers/la_oen_core[124] mgmt_buffers/la_oen_core[125]
+ mgmt_buffers/la_oen_core[126] mgmt_buffers/la_oen_core[127] mgmt_buffers/la_oen_core[12]
+ mgmt_buffers/la_oen_core[13] mgmt_buffers/la_oen_core[14] mgmt_buffers/la_oen_core[15]
+ mgmt_buffers/la_oen_core[16] mgmt_buffers/la_oen_core[17] mgmt_buffers/la_oen_core[18]
+ mgmt_buffers/la_oen_core[19] mgmt_buffers/la_oen_core[1] mgmt_buffers/la_oen_core[20]
+ mgmt_buffers/la_oen_core[21] mgmt_buffers/la_oen_core[22] mgmt_buffers/la_oen_core[23]
+ mgmt_buffers/la_oen_core[24] mgmt_buffers/la_oen_core[25] mgmt_buffers/la_oen_core[26]
+ mgmt_buffers/la_oen_core[27] mgmt_buffers/la_oen_core[28] mgmt_buffers/la_oen_core[29]
+ mgmt_buffers/la_oen_core[2] mgmt_buffers/la_oen_core[30] mgmt_buffers/la_oen_core[31]
+ mgmt_buffers/la_oen_core[32] mgmt_buffers/la_oen_core[33] mgmt_buffers/la_oen_core[34]
+ mgmt_buffers/la_oen_core[35] mgmt_buffers/la_oen_core[36] mgmt_buffers/la_oen_core[37]
+ mgmt_buffers/la_oen_core[38] mgmt_buffers/la_oen_core[39] mgmt_buffers/la_oen_core[3]
+ mgmt_buffers/la_oen_core[40] mgmt_buffers/la_oen_core[41] mgmt_buffers/la_oen_core[42]
+ mgmt_buffers/la_oen_core[43] mgmt_buffers/la_oen_core[44] mgmt_buffers/la_oen_core[45]
+ mgmt_buffers/la_oen_core[46] mgmt_buffers/la_oen_core[47] mgmt_buffers/la_oen_core[48]
+ mgmt_buffers/la_oen_core[49] mgmt_buffers/la_oen_core[4] mgmt_buffers/la_oen_core[50]
+ mgmt_buffers/la_oen_core[51] mgmt_buffers/la_oen_core[52] mgmt_buffers/la_oen_core[53]
+ mgmt_buffers/la_oen_core[54] mgmt_buffers/la_oen_core[55] mgmt_buffers/la_oen_core[56]
+ mgmt_buffers/la_oen_core[57] mgmt_buffers/la_oen_core[58] mgmt_buffers/la_oen_core[59]
+ mgmt_buffers/la_oen_core[5] mgmt_buffers/la_oen_core[60] mgmt_buffers/la_oen_core[61]
+ mgmt_buffers/la_oen_core[62] mgmt_buffers/la_oen_core[63] mgmt_buffers/la_oen_core[64]
+ mgmt_buffers/la_oen_core[65] mgmt_buffers/la_oen_core[66] mgmt_buffers/la_oen_core[67]
+ mgmt_buffers/la_oen_core[68] mgmt_buffers/la_oen_core[69] mgmt_buffers/la_oen_core[6]
+ mgmt_buffers/la_oen_core[70] mgmt_buffers/la_oen_core[71] mgmt_buffers/la_oen_core[72]
+ mgmt_buffers/la_oen_core[73] mgmt_buffers/la_oen_core[74] mgmt_buffers/la_oen_core[75]
+ mgmt_buffers/la_oen_core[76] mgmt_buffers/la_oen_core[77] mgmt_buffers/la_oen_core[78]
+ mgmt_buffers/la_oen_core[79] mgmt_buffers/la_oen_core[7] mgmt_buffers/la_oen_core[80]
+ mgmt_buffers/la_oen_core[81] mgmt_buffers/la_oen_core[82] mgmt_buffers/la_oen_core[83]
+ mgmt_buffers/la_oen_core[84] mgmt_buffers/la_oen_core[85] mgmt_buffers/la_oen_core[86]
+ mgmt_buffers/la_oen_core[87] mgmt_buffers/la_oen_core[88] mgmt_buffers/la_oen_core[89]
+ mgmt_buffers/la_oen_core[8] mgmt_buffers/la_oen_core[90] mgmt_buffers/la_oen_core[91]
+ mgmt_buffers/la_oen_core[92] mgmt_buffers/la_oen_core[93] mgmt_buffers/la_oen_core[94]
+ mgmt_buffers/la_oen_core[95] mgmt_buffers/la_oen_core[96] mgmt_buffers/la_oen_core[97]
+ mgmt_buffers/la_oen_core[98] mgmt_buffers/la_oen_core[99] mgmt_buffers/la_oen_core[9]
+ soc/la_oen[0] soc/la_oen[100] soc/la_oen[101] soc/la_oen[102] soc/la_oen[103] soc/la_oen[104]
+ soc/la_oen[105] soc/la_oen[106] soc/la_oen[107] soc/la_oen[108] soc/la_oen[109]
+ soc/la_oen[10] soc/la_oen[110] soc/la_oen[111] soc/la_oen[112] soc/la_oen[113] soc/la_oen[114]
+ soc/la_oen[115] soc/la_oen[116] soc/la_oen[117] soc/la_oen[118] soc/la_oen[119]
+ soc/la_oen[11] soc/la_oen[120] soc/la_oen[121] soc/la_oen[122] soc/la_oen[123] soc/la_oen[124]
+ soc/la_oen[125] soc/la_oen[126] soc/la_oen[127] soc/la_oen[12] soc/la_oen[13] soc/la_oen[14]
+ soc/la_oen[15] soc/la_oen[16] soc/la_oen[17] soc/la_oen[18] soc/la_oen[19] soc/la_oen[1]
+ soc/la_oen[20] soc/la_oen[21] soc/la_oen[22] soc/la_oen[23] soc/la_oen[24] soc/la_oen[25]
+ soc/la_oen[26] soc/la_oen[27] soc/la_oen[28] soc/la_oen[29] soc/la_oen[2] soc/la_oen[30]
+ soc/la_oen[31] soc/la_oen[32] soc/la_oen[33] soc/la_oen[34] soc/la_oen[35] soc/la_oen[36]
+ soc/la_oen[37] soc/la_oen[38] soc/la_oen[39] soc/la_oen[3] soc/la_oen[40] soc/la_oen[41]
+ soc/la_oen[42] soc/la_oen[43] soc/la_oen[44] soc/la_oen[45] soc/la_oen[46] soc/la_oen[47]
+ soc/la_oen[48] soc/la_oen[49] soc/la_oen[4] soc/la_oen[50] soc/la_oen[51] soc/la_oen[52]
+ soc/la_oen[53] soc/la_oen[54] soc/la_oen[55] soc/la_oen[56] soc/la_oen[57] soc/la_oen[58]
+ soc/la_oen[59] soc/la_oen[5] soc/la_oen[60] soc/la_oen[61] soc/la_oen[62] soc/la_oen[63]
+ soc/la_oen[64] soc/la_oen[65] soc/la_oen[66] soc/la_oen[67] soc/la_oen[68] soc/la_oen[69]
+ soc/la_oen[6] soc/la_oen[70] soc/la_oen[71] soc/la_oen[72] soc/la_oen[73] soc/la_oen[74]
+ soc/la_oen[75] soc/la_oen[76] soc/la_oen[77] soc/la_oen[78] soc/la_oen[79] soc/la_oen[7]
+ soc/la_oen[80] soc/la_oen[81] soc/la_oen[82] soc/la_oen[83] soc/la_oen[84] soc/la_oen[85]
+ soc/la_oen[86] soc/la_oen[87] soc/la_oen[88] soc/la_oen[89] soc/la_oen[8] soc/la_oen[90]
+ soc/la_oen[91] soc/la_oen[92] soc/la_oen[93] soc/la_oen[94] soc/la_oen[95] soc/la_oen[96]
+ soc/la_oen[97] soc/la_oen[98] soc/la_oen[99] soc/la_oen[9] soc/mprj_adr_o[0] soc/mprj_adr_o[10]
+ soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15]
+ soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1]
+ soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24]
+ soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29]
+ soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4]
+ soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9]
+ mgmt_buffers/mprj_adr_o_user[0] mgmt_buffers/mprj_adr_o_user[10] mgmt_buffers/mprj_adr_o_user[11]
+ mgmt_buffers/mprj_adr_o_user[12] mgmt_buffers/mprj_adr_o_user[13] mgmt_buffers/mprj_adr_o_user[14]
+ mgmt_buffers/mprj_adr_o_user[15] mgmt_buffers/mprj_adr_o_user[16] mgmt_buffers/mprj_adr_o_user[17]
+ mgmt_buffers/mprj_adr_o_user[18] mgmt_buffers/mprj_adr_o_user[19] mgmt_buffers/mprj_adr_o_user[1]
+ mgmt_buffers/mprj_adr_o_user[20] mgmt_buffers/mprj_adr_o_user[21] mgmt_buffers/mprj_adr_o_user[22]
+ mgmt_buffers/mprj_adr_o_user[23] mgmt_buffers/mprj_adr_o_user[24] mgmt_buffers/mprj_adr_o_user[25]
+ mgmt_buffers/mprj_adr_o_user[26] mgmt_buffers/mprj_adr_o_user[27] mgmt_buffers/mprj_adr_o_user[28]
+ mgmt_buffers/mprj_adr_o_user[29] mgmt_buffers/mprj_adr_o_user[2] mgmt_buffers/mprj_adr_o_user[30]
+ mgmt_buffers/mprj_adr_o_user[31] mgmt_buffers/mprj_adr_o_user[3] mgmt_buffers/mprj_adr_o_user[4]
+ mgmt_buffers/mprj_adr_o_user[5] mgmt_buffers/mprj_adr_o_user[6] mgmt_buffers/mprj_adr_o_user[7]
+ mgmt_buffers/mprj_adr_o_user[8] mgmt_buffers/mprj_adr_o_user[9] soc/mprj_cyc_o mgmt_buffers/mprj_cyc_o_user
+ soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13]
+ soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18]
+ soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22]
+ soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27]
+ soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31]
+ soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7]
+ soc/mprj_dat_o[8] soc/mprj_dat_o[9] mgmt_buffers/mprj_dat_o_user[0] mgmt_buffers/mprj_dat_o_user[10]
+ mgmt_buffers/mprj_dat_o_user[11] mgmt_buffers/mprj_dat_o_user[12] mgmt_buffers/mprj_dat_o_user[13]
+ mgmt_buffers/mprj_dat_o_user[14] mgmt_buffers/mprj_dat_o_user[15] mgmt_buffers/mprj_dat_o_user[16]
+ mgmt_buffers/mprj_dat_o_user[17] mgmt_buffers/mprj_dat_o_user[18] mgmt_buffers/mprj_dat_o_user[19]
+ mgmt_buffers/mprj_dat_o_user[1] mgmt_buffers/mprj_dat_o_user[20] mgmt_buffers/mprj_dat_o_user[21]
+ mgmt_buffers/mprj_dat_o_user[22] mgmt_buffers/mprj_dat_o_user[23] mgmt_buffers/mprj_dat_o_user[24]
+ mgmt_buffers/mprj_dat_o_user[25] mgmt_buffers/mprj_dat_o_user[26] mgmt_buffers/mprj_dat_o_user[27]
+ mgmt_buffers/mprj_dat_o_user[28] mgmt_buffers/mprj_dat_o_user[29] mgmt_buffers/mprj_dat_o_user[2]
+ mgmt_buffers/mprj_dat_o_user[30] mgmt_buffers/mprj_dat_o_user[31] mgmt_buffers/mprj_dat_o_user[3]
+ mgmt_buffers/mprj_dat_o_user[4] mgmt_buffers/mprj_dat_o_user[5] mgmt_buffers/mprj_dat_o_user[6]
+ mgmt_buffers/mprj_dat_o_user[7] mgmt_buffers/mprj_dat_o_user[8] mgmt_buffers/mprj_dat_o_user[9]
+ soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] mgmt_buffers/mprj_sel_o_user[0]
+ mgmt_buffers/mprj_sel_o_user[1] mgmt_buffers/mprj_sel_o_user[2] mgmt_buffers/mprj_sel_o_user[3]
+ soc/mprj_stb_o mgmt_buffers/mprj_stb_o_user soc/mprj_we_o mgmt_buffers/mprj_we_o_user
+ soc/mprj_vcc_pwrgood soc/mprj_vdd_pwrgood soc/mprj2_vcc_pwrgood soc/mprj2_vdd_pwrgood
+ mgmt_buffers/user_clock mgmt_buffers/user_clock2 mgmt_buffers/user_reset mgmt_buffers/user_resetn
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 mprj/vccd2 mprj/vssd2 mprj/vdda1 mprj/vdda2
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/m1_25_11# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/m1_25_11# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# soc/m2_572_856# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/m3_38_51# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/m1_25_11# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/m3_38_51# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/vss por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/m1_25_11# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/m1_25_11#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/m1_25_11# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/m1_25_11#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# soc/m2_572_856# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# mgmt_protect
Xrstb_level rstb_level/A soc/resetb vddio por/vss soc/VPWR rstb_level/LVGND por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/m1_25_11# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/m1_25_11# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/m1_25_11#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36# por/li_35_36#
+ por/li_35_36# sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped
Xgpio_control_in\[27\] soc/mgmt_in_data[27] gpio_control_in\[27\]/one soc/mgmt_in_data[27]
+ gpio_control_in\[27\]/one padframe/mprj_io_analog_en[27] padframe/mprj_io_analog_pol[27]
+ padframe/mprj_io_analog_sel[27] padframe/mprj_io_dm[81] padframe/mprj_io_dm[82]
+ padframe/mprj_io_dm[83] padframe/mprj_io_holdover[27] padframe/mprj_io_ib_mode_sel[27]
+ padframe/mprj_io_in[27] padframe/mprj_io_inp_dis[27] padframe/mprj_io_out[27] padframe/mprj_io_oeb[27]
+ padframe/mprj_io_slow_sel[27] padframe/mprj_io_vtrip_sel[27] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[27\]/serial_data_in gpio_control_in\[28\]/serial_data_in
+ gpio_control_in\[27\]/user_gpio_in gpio_control_in\[27\]/user_gpio_oeb gpio_control_in\[27\]/user_gpio_out
+ gpio_control_in\[27\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[2\] soc/mgmt_in_data[2] gpio_control_in\[2\]/one soc/mgmt_in_data[2]
+ gpio_control_in\[2\]/one padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2]
+ padframe/mprj_io_analog_sel[2] padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8]
+ padframe/mprj_io_holdover[2] padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_in[2]
+ padframe/mprj_io_inp_dis[2] padframe/mprj_io_out[2] padframe/mprj_io_oeb[2] padframe/mprj_io_slow_sel[2]
+ padframe/mprj_io_vtrip_sel[2] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[2\]/serial_data_in gpio_control_in\[3\]/serial_data_in gpio_control_in\[2\]/user_gpio_in
+ gpio_control_in\[2\]/user_gpio_oeb gpio_control_in\[2\]/user_gpio_out gpio_control_in\[2\]/zero
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[32\] soc/mgmt_in_data[32] gpio_control_in\[32\]/one soc/mgmt_in_data[32]
+ gpio_control_in\[32\]/one padframe/mprj_io_analog_en[32] padframe/mprj_io_analog_pol[32]
+ padframe/mprj_io_analog_sel[32] padframe/mprj_io_dm[96] padframe/mprj_io_dm[97]
+ padframe/mprj_io_dm[98] padframe/mprj_io_holdover[32] padframe/mprj_io_ib_mode_sel[32]
+ padframe/mprj_io_in[32] padframe/mprj_io_inp_dis[32] padframe/mprj_io_out[32] padframe/mprj_io_oeb[32]
+ padframe/mprj_io_slow_sel[32] padframe/mprj_io_vtrip_sel[32] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[32\]/serial_data_in gpio_control_in\[33\]/serial_data_in
+ gpio_control_in\[32\]/user_gpio_in gpio_control_in\[32\]/user_gpio_oeb gpio_control_in\[32\]/user_gpio_out
+ gpio_control_in\[32\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[25\] soc/mgmt_in_data[25] gpio_control_in\[25\]/one soc/mgmt_in_data[25]
+ gpio_control_in\[25\]/one padframe/mprj_io_analog_en[25] padframe/mprj_io_analog_pol[25]
+ padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75] padframe/mprj_io_dm[76]
+ padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_in[25] padframe/mprj_io_inp_dis[25] padframe/mprj_io_out[25] padframe/mprj_io_oeb[25]
+ padframe/mprj_io_slow_sel[25] padframe/mprj_io_vtrip_sel[25] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[25\]/serial_data_in gpio_control_in\[26\]/serial_data_in
+ gpio_control_in\[25\]/user_gpio_in gpio_control_in\[25\]/user_gpio_oeb gpio_control_in\[25\]/user_gpio_out
+ gpio_control_in\[25\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[18\] soc/mgmt_in_data[18] gpio_control_in\[18\]/one soc/mgmt_in_data[18]
+ gpio_control_in\[18\]/one padframe/mprj_io_analog_en[18] padframe/mprj_io_analog_pol[18]
+ padframe/mprj_io_analog_sel[18] padframe/mprj_io_dm[54] padframe/mprj_io_dm[55]
+ padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18] padframe/mprj_io_ib_mode_sel[18]
+ padframe/mprj_io_in[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_out[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[18\]/serial_data_in gpio_control_in\[19\]/serial_data_in
+ gpio_control_in\[18\]/user_gpio_in gpio_control_in\[18\]/user_gpio_oeb gpio_control_in\[18\]/user_gpio_out
+ gpio_control_in\[18\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[30\] soc/mgmt_in_data[30] gpio_control_in\[30\]/one soc/mgmt_in_data[30]
+ gpio_control_in\[30\]/one padframe/mprj_io_analog_en[30] padframe/mprj_io_analog_pol[30]
+ padframe/mprj_io_analog_sel[30] padframe/mprj_io_dm[90] padframe/mprj_io_dm[91]
+ padframe/mprj_io_dm[92] padframe/mprj_io_holdover[30] padframe/mprj_io_ib_mode_sel[30]
+ padframe/mprj_io_in[30] padframe/mprj_io_inp_dis[30] padframe/mprj_io_out[30] padframe/mprj_io_oeb[30]
+ padframe/mprj_io_slow_sel[30] padframe/mprj_io_vtrip_sel[30] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[30\]/serial_data_in gpio_control_in\[31\]/serial_data_in
+ gpio_control_in\[30\]/user_gpio_in gpio_control_in\[30\]/user_gpio_oeb gpio_control_in\[30\]/user_gpio_out
+ gpio_control_in\[30\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[23\] soc/mgmt_in_data[23] gpio_control_in\[23\]/one soc/mgmt_in_data[23]
+ gpio_control_in\[23\]/one padframe/mprj_io_analog_en[23] padframe/mprj_io_analog_pol[23]
+ padframe/mprj_io_analog_sel[23] padframe/mprj_io_dm[69] padframe/mprj_io_dm[70]
+ padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23] padframe/mprj_io_ib_mode_sel[23]
+ padframe/mprj_io_in[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_out[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[23\]/serial_data_in gpio_control_in\[24\]/serial_data_in
+ gpio_control_in\[23\]/user_gpio_in gpio_control_in\[23\]/user_gpio_oeb gpio_control_in\[23\]/user_gpio_out
+ gpio_control_in\[23\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[9\] soc/mgmt_in_data[9] gpio_control_in\[9\]/one soc/mgmt_in_data[9]
+ gpio_control_in\[9\]/one padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9]
+ padframe/mprj_io_analog_sel[9] padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29]
+ padframe/mprj_io_holdover[9] padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_in[9]
+ padframe/mprj_io_inp_dis[9] padframe/mprj_io_out[9] padframe/mprj_io_oeb[9] padframe/mprj_io_slow_sel[9]
+ padframe/mprj_io_vtrip_sel[9] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[9\]/serial_data_in gpio_control_in\[9\]/serial_data_out gpio_control_in\[9\]/user_gpio_in
+ gpio_control_in\[9\]/user_gpio_oeb gpio_control_in\[9\]/user_gpio_out gpio_control_in\[9\]/zero
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_bidir\[0\] soc/mgmt_in_data[0] soc/jtag_outenb soc/jtag_out gpio_control_bidir\[0\]/one
+ padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0] padframe/mprj_io_analog_sel[0]
+ padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2] padframe/mprj_io_holdover[0]
+ padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_in[0] padframe/mprj_io_inp_dis[0]
+ padframe/mprj_io_out[0] padframe/mprj_io_oeb[0] padframe/mprj_io_slow_sel[0] padframe/mprj_io_vtrip_sel[0]
+ soc/mprj_io_loader_resetn soc/mprj_io_loader_clock soc/mprj_io_loader_data gpio_control_bidir\[1\]/serial_data_in
+ gpio_control_bidir\[0\]/user_gpio_in gpio_control_bidir\[0\]/user_gpio_oeb gpio_control_bidir\[0\]/user_gpio_out
+ gpio_control_bidir\[0\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[16\] soc/mgmt_in_data[16] gpio_control_in\[16\]/one soc/mgmt_in_data[16]
+ gpio_control_in\[16\]/one padframe/mprj_io_analog_en[16] padframe/mprj_io_analog_pol[16]
+ padframe/mprj_io_analog_sel[16] padframe/mprj_io_dm[48] padframe/mprj_io_dm[49]
+ padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16] padframe/mprj_io_ib_mode_sel[16]
+ padframe/mprj_io_in[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_out[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[16\]/serial_data_in gpio_control_in\[17\]/serial_data_in
+ gpio_control_in\[16\]/user_gpio_in gpio_control_in\[16\]/user_gpio_oeb gpio_control_in\[16\]/user_gpio_out
+ gpio_control_in\[16\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[21\] soc/mgmt_in_data[21] gpio_control_in\[21\]/one soc/mgmt_in_data[21]
+ gpio_control_in\[21\]/one padframe/mprj_io_analog_en[21] padframe/mprj_io_analog_pol[21]
+ padframe/mprj_io_analog_sel[21] padframe/mprj_io_dm[63] padframe/mprj_io_dm[64]
+ padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21] padframe/mprj_io_ib_mode_sel[21]
+ padframe/mprj_io_in[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_out[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[21\]/serial_data_in gpio_control_in\[22\]/serial_data_in
+ gpio_control_in\[21\]/user_gpio_in gpio_control_in\[21\]/user_gpio_oeb gpio_control_in\[21\]/user_gpio_out
+ gpio_control_in\[21\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xmprj mprj/analog_io[0] mprj/analog_io[10] mprj/analog_io[11] mprj/analog_io[12] mprj/analog_io[13]
+ mprj/analog_io[14] mprj/analog_io[15] mprj/analog_io[16] mprj/analog_io[17] mprj/analog_io[18]
+ mprj/analog_io[19] mprj/analog_io[1] mprj/analog_io[20] mprj/analog_io[21] mprj/analog_io[22]
+ mprj/analog_io[23] mprj/analog_io[24] mprj/analog_io[25] mprj/analog_io[26] mprj/analog_io[27]
+ mprj/analog_io[28] mprj/analog_io[29] mprj/analog_io[2] mprj/analog_io[30] mprj/analog_io[3]
+ mprj/analog_io[4] mprj/analog_io[5] mprj/analog_io[6] mprj/analog_io[7] mprj/analog_io[8]
+ mprj/analog_io[9] mprj/io_in[0] mprj/io_in[10] mprj/io_in[11] mprj/io_in[12] mprj/io_in[13]
+ mprj/io_in[14] mprj/io_in[15] mprj/io_in[16] mprj/io_in[17] mprj/io_in[18] mprj/io_in[19]
+ mprj/io_in[1] mprj/io_in[20] mprj/io_in[21] mprj/io_in[22] mprj/io_in[23] mprj/io_in[24]
+ mprj/io_in[25] mprj/io_in[26] mprj/io_in[27] mprj/io_in[28] mprj/io_in[29] mprj/io_in[2]
+ mprj/io_in[30] mprj/io_in[31] mprj/io_in[32] mprj/io_in[33] mprj/io_in[34] mprj/io_in[35]
+ mprj/io_in[36] mprj/io_in[37] mprj/io_in[3] mprj/io_in[4] mprj/io_in[5] mprj/io_in[6]
+ mprj/io_in[7] mprj/io_in[8] mprj/io_in[9] mprj/io_oeb[0] mprj/io_oeb[10] mprj/io_oeb[11]
+ mprj/io_oeb[12] mprj/io_oeb[13] mprj/io_oeb[14] mprj/io_oeb[15] mprj/io_oeb[16]
+ mprj/io_oeb[17] mprj/io_oeb[18] mprj/io_oeb[19] mprj/io_oeb[1] mprj/io_oeb[20] mprj/io_oeb[21]
+ mprj/io_oeb[22] mprj/io_oeb[23] mprj/io_oeb[24] mprj/io_oeb[25] mprj/io_oeb[26]
+ mprj/io_oeb[27] mprj/io_oeb[28] mprj/io_oeb[29] mprj/io_oeb[2] mprj/io_oeb[30] mprj/io_oeb[31]
+ mprj/io_oeb[32] mprj/io_oeb[33] mprj/io_oeb[34] mprj/io_oeb[35] mprj/io_oeb[36]
+ mprj/io_oeb[37] mprj/io_oeb[3] mprj/io_oeb[4] mprj/io_oeb[5] mprj/io_oeb[6] mprj/io_oeb[7]
+ mprj/io_oeb[8] mprj/io_oeb[9] mprj/io_out[0] mprj/io_out[10] mprj/io_out[11] mprj/io_out[12]
+ mprj/io_out[13] mprj/io_out[14] mprj/io_out[15] mprj/io_out[16] mprj/io_out[17]
+ mprj/io_out[18] mprj/io_out[19] mprj/io_out[1] mprj/io_out[20] mprj/io_out[21] mprj/io_out[22]
+ mprj/io_out[23] mprj/io_out[24] mprj/io_out[25] mprj/io_out[26] mprj/io_out[27]
+ mprj/io_out[28] mprj/io_out[29] mprj/io_out[2] mprj/io_out[30] mprj/io_out[31] mprj/io_out[32]
+ mprj/io_out[33] mprj/io_out[34] mprj/io_out[35] mprj/io_out[36] mprj/io_out[37]
+ mprj/io_out[3] mprj/io_out[4] mprj/io_out[5] mprj/io_out[6] mprj/io_out[7] mprj/io_out[8]
+ mprj/io_out[9] mprj/la_data_in[0] mprj/la_data_in[100] mprj/la_data_in[101] mprj/la_data_in[102]
+ mprj/la_data_in[103] mprj/la_data_in[104] mprj/la_data_in[105] mprj/la_data_in[106]
+ mprj/la_data_in[107] mprj/la_data_in[108] mprj/la_data_in[109] mprj/la_data_in[10]
+ mprj/la_data_in[110] mprj/la_data_in[111] mprj/la_data_in[112] mprj/la_data_in[113]
+ mprj/la_data_in[114] mprj/la_data_in[115] mprj/la_data_in[116] mprj/la_data_in[117]
+ mprj/la_data_in[118] mprj/la_data_in[119] mprj/la_data_in[11] mprj/la_data_in[120]
+ mprj/la_data_in[121] mprj/la_data_in[122] mprj/la_data_in[123] mprj/la_data_in[124]
+ mprj/la_data_in[125] mprj/la_data_in[126] mprj/la_data_in[127] mprj/la_data_in[12]
+ mprj/la_data_in[13] mprj/la_data_in[14] mprj/la_data_in[15] mprj/la_data_in[16]
+ mprj/la_data_in[17] mprj/la_data_in[18] mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20]
+ mprj/la_data_in[21] mprj/la_data_in[22] mprj/la_data_in[23] mprj/la_data_in[24]
+ mprj/la_data_in[25] mprj/la_data_in[26] mprj/la_data_in[27] mprj/la_data_in[28]
+ mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30] mprj/la_data_in[31] mprj/la_data_in[32]
+ mprj/la_data_in[33] mprj/la_data_in[34] mprj/la_data_in[35] mprj/la_data_in[36]
+ mprj/la_data_in[37] mprj/la_data_in[38] mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40]
+ mprj/la_data_in[41] mprj/la_data_in[42] mprj/la_data_in[43] mprj/la_data_in[44]
+ mprj/la_data_in[45] mprj/la_data_in[46] mprj/la_data_in[47] mprj/la_data_in[48]
+ mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50] mprj/la_data_in[51] mprj/la_data_in[52]
+ mprj/la_data_in[53] mprj/la_data_in[54] mprj/la_data_in[55] mprj/la_data_in[56]
+ mprj/la_data_in[57] mprj/la_data_in[58] mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60]
+ mprj/la_data_in[61] mprj/la_data_in[62] mprj/la_data_in[63] mprj/la_data_in[64]
+ mprj/la_data_in[65] mprj/la_data_in[66] mprj/la_data_in[67] mprj/la_data_in[68]
+ mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70] mprj/la_data_in[71] mprj/la_data_in[72]
+ mprj/la_data_in[73] mprj/la_data_in[74] mprj/la_data_in[75] mprj/la_data_in[76]
+ mprj/la_data_in[77] mprj/la_data_in[78] mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80]
+ mprj/la_data_in[81] mprj/la_data_in[82] mprj/la_data_in[83] mprj/la_data_in[84]
+ mprj/la_data_in[85] mprj/la_data_in[86] mprj/la_data_in[87] mprj/la_data_in[88]
+ mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90] mprj/la_data_in[91] mprj/la_data_in[92]
+ mprj/la_data_in[93] mprj/la_data_in[94] mprj/la_data_in[95] mprj/la_data_in[96]
+ mprj/la_data_in[97] mprj/la_data_in[98] mprj/la_data_in[99] mprj/la_data_in[9] mprj/la_data_out[0]
+ mprj/la_data_out[100] mprj/la_data_out[101] mprj/la_data_out[102] mprj/la_data_out[103]
+ mprj/la_data_out[104] mprj/la_data_out[105] mprj/la_data_out[106] mprj/la_data_out[107]
+ mprj/la_data_out[108] mprj/la_data_out[109] mprj/la_data_out[10] mprj/la_data_out[110]
+ mprj/la_data_out[111] mprj/la_data_out[112] mprj/la_data_out[113] mprj/la_data_out[114]
+ mprj/la_data_out[115] mprj/la_data_out[116] mprj/la_data_out[117] mprj/la_data_out[118]
+ mprj/la_data_out[119] mprj/la_data_out[11] mprj/la_data_out[120] mprj/la_data_out[121]
+ mprj/la_data_out[122] mprj/la_data_out[123] mprj/la_data_out[124] mprj/la_data_out[125]
+ mprj/la_data_out[126] mprj/la_data_out[127] mprj/la_data_out[12] mprj/la_data_out[13]
+ mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16] mprj/la_data_out[17]
+ mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1] mprj/la_data_out[20]
+ mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23] mprj/la_data_out[24]
+ mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27] mprj/la_data_out[28]
+ mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30] mprj/la_data_out[31]
+ mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34] mprj/la_data_out[35]
+ mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38] mprj/la_data_out[39]
+ mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41] mprj/la_data_out[42]
+ mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45] mprj/la_data_out[46]
+ mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49] mprj/la_data_out[4]
+ mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52] mprj/la_data_out[53]
+ mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56] mprj/la_data_out[57]
+ mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5] mprj/la_data_out[60]
+ mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63] mprj/la_data_out[64]
+ mprj/la_data_out[65] mprj/la_data_out[66] mprj/la_data_out[67] mprj/la_data_out[68]
+ mprj/la_data_out[69] mprj/la_data_out[6] mprj/la_data_out[70] mprj/la_data_out[71]
+ mprj/la_data_out[72] mprj/la_data_out[73] mprj/la_data_out[74] mprj/la_data_out[75]
+ mprj/la_data_out[76] mprj/la_data_out[77] mprj/la_data_out[78] mprj/la_data_out[79]
+ mprj/la_data_out[7] mprj/la_data_out[80] mprj/la_data_out[81] mprj/la_data_out[82]
+ mprj/la_data_out[83] mprj/la_data_out[84] mprj/la_data_out[85] mprj/la_data_out[86]
+ mprj/la_data_out[87] mprj/la_data_out[88] mprj/la_data_out[89] mprj/la_data_out[8]
+ mprj/la_data_out[90] mprj/la_data_out[91] mprj/la_data_out[92] mprj/la_data_out[93]
+ mprj/la_data_out[94] mprj/la_data_out[95] mprj/la_data_out[96] mprj/la_data_out[97]
+ mprj/la_data_out[98] mprj/la_data_out[99] mprj/la_data_out[9] mprj/la_oen[0] mprj/la_oen[100]
+ mprj/la_oen[101] mprj/la_oen[102] mprj/la_oen[103] mprj/la_oen[104] mprj/la_oen[105]
+ mprj/la_oen[106] mprj/la_oen[107] mprj/la_oen[108] mprj/la_oen[109] mprj/la_oen[10]
+ mprj/la_oen[110] mprj/la_oen[111] mprj/la_oen[112] mprj/la_oen[113] mprj/la_oen[114]
+ mprj/la_oen[115] mprj/la_oen[116] mprj/la_oen[117] mprj/la_oen[118] mprj/la_oen[119]
+ mprj/la_oen[11] mprj/la_oen[120] mprj/la_oen[121] mprj/la_oen[122] mprj/la_oen[123]
+ mprj/la_oen[124] mprj/la_oen[125] mprj/la_oen[126] mprj/la_oen[127] mprj/la_oen[12]
+ mprj/la_oen[13] mprj/la_oen[14] mprj/la_oen[15] mprj/la_oen[16] mprj/la_oen[17]
+ mprj/la_oen[18] mprj/la_oen[19] mprj/la_oen[1] mprj/la_oen[20] mprj/la_oen[21] mprj/la_oen[22]
+ mprj/la_oen[23] mprj/la_oen[24] mprj/la_oen[25] mprj/la_oen[26] mprj/la_oen[27]
+ mprj/la_oen[28] mprj/la_oen[29] mprj/la_oen[2] mprj/la_oen[30] mprj/la_oen[31] mprj/la_oen[32]
+ mprj/la_oen[33] mprj/la_oen[34] mprj/la_oen[35] mprj/la_oen[36] mprj/la_oen[37]
+ mprj/la_oen[38] mprj/la_oen[39] mprj/la_oen[3] mprj/la_oen[40] mprj/la_oen[41] mprj/la_oen[42]
+ mprj/la_oen[43] mprj/la_oen[44] mprj/la_oen[45] mprj/la_oen[46] mprj/la_oen[47]
+ mprj/la_oen[48] mprj/la_oen[49] mprj/la_oen[4] mprj/la_oen[50] mprj/la_oen[51] mprj/la_oen[52]
+ mprj/la_oen[53] mprj/la_oen[54] mprj/la_oen[55] mprj/la_oen[56] mprj/la_oen[57]
+ mprj/la_oen[58] mprj/la_oen[59] mprj/la_oen[5] mprj/la_oen[60] mprj/la_oen[61] mprj/la_oen[62]
+ mprj/la_oen[63] mprj/la_oen[64] mprj/la_oen[65] mprj/la_oen[66] mprj/la_oen[67]
+ mprj/la_oen[68] mprj/la_oen[69] mprj/la_oen[6] mprj/la_oen[70] mprj/la_oen[71] mprj/la_oen[72]
+ mprj/la_oen[73] mprj/la_oen[74] mprj/la_oen[75] mprj/la_oen[76] mprj/la_oen[77]
+ mprj/la_oen[78] mprj/la_oen[79] mprj/la_oen[7] mprj/la_oen[80] mprj/la_oen[81] mprj/la_oen[82]
+ mprj/la_oen[83] mprj/la_oen[84] mprj/la_oen[85] mprj/la_oen[86] mprj/la_oen[87]
+ mprj/la_oen[88] mprj/la_oen[89] mprj/la_oen[8] mprj/la_oen[90] mprj/la_oen[91] mprj/la_oen[92]
+ mprj/la_oen[93] mprj/la_oen[94] mprj/la_oen[95] mprj/la_oen[96] mprj/la_oen[97]
+ mprj/la_oen[98] mprj/la_oen[99] mprj/la_oen[9] mprj/user_clock2 mprj/wb_clk_i mprj/wb_rst_i
+ mprj/wbs_ack_o mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11] mprj/wbs_adr_i[12]
+ mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16] mprj/wbs_adr_i[17]
+ mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20] mprj/wbs_adr_i[21]
+ mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25] mprj/wbs_adr_i[26]
+ mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2] mprj/wbs_adr_i[30]
+ mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5] mprj/wbs_adr_i[6]
+ mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] mprj/wbs_cyc_i mprj/wbs_dat_i[0]
+ mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13] mprj/wbs_dat_i[14]
+ mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18] mprj/wbs_dat_i[19]
+ mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22] mprj/wbs_dat_i[23]
+ mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27] mprj/wbs_dat_i[28]
+ mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31] mprj/wbs_dat_i[3]
+ mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7] mprj/wbs_dat_i[8]
+ mprj/wbs_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11] mprj/wbs_dat_o[12]
+ mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16] mprj/wbs_dat_o[17]
+ mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20] mprj/wbs_dat_o[21]
+ mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25] mprj/wbs_dat_o[26]
+ mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2] mprj/wbs_dat_o[30]
+ mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5] mprj/wbs_dat_o[6]
+ mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] mprj/wbs_sel_i[0] mprj/wbs_sel_i[1]
+ mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] mprj/wbs_stb_i mprj/wbs_we_i mprj/vccd1 mprj/vssd1
+ mprj/vccd2 mprj/vssd2 mprj/vdda1 por/vss mprj/vdda2 por/vss user_project_wrapper
Xgpio_control_in\[14\] soc/mgmt_in_data[14] gpio_control_in\[14\]/one soc/mgmt_in_data[14]
+ gpio_control_in\[14\]/one padframe/mprj_io_analog_en[14] padframe/mprj_io_analog_pol[14]
+ padframe/mprj_io_analog_sel[14] padframe/mprj_io_dm[42] padframe/mprj_io_dm[43]
+ padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14] padframe/mprj_io_ib_mode_sel[14]
+ padframe/mprj_io_in[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_out[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[14\]/serial_data_in gpio_control_in\[15\]/serial_data_in
+ gpio_control_in\[14\]/user_gpio_in gpio_control_in\[14\]/user_gpio_oeb gpio_control_in\[14\]/user_gpio_out
+ gpio_control_in\[14\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[7\] soc/mgmt_in_data[7] gpio_control_in\[7\]/one soc/mgmt_in_data[7]
+ gpio_control_in\[7\]/one padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7]
+ padframe/mprj_io_analog_sel[7] padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23]
+ padframe/mprj_io_holdover[7] padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_in[7]
+ padframe/mprj_io_inp_dis[7] padframe/mprj_io_out[7] padframe/mprj_io_oeb[7] padframe/mprj_io_slow_sel[7]
+ padframe/mprj_io_vtrip_sel[7] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[7\]/serial_data_in gpio_control_in\[8\]/serial_data_in gpio_control_in\[7\]/user_gpio_in
+ gpio_control_in\[7\]/user_gpio_oeb gpio_control_in\[7\]/user_gpio_out gpio_control_in\[7\]/zero
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[5\] soc/mgmt_in_data[5] gpio_control_in\[5\]/one soc/mgmt_in_data[5]
+ gpio_control_in\[5\]/one padframe/mprj_io_analog_en[5] padframe/mprj_io_analog_pol[5]
+ padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15] padframe/mprj_io_dm[16] padframe/mprj_io_dm[17]
+ padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5] padframe/mprj_io_in[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_out[5] padframe/mprj_io_oeb[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[5\]/serial_data_in gpio_control_in\[6\]/serial_data_in gpio_control_in\[5\]/user_gpio_in
+ gpio_control_in\[5\]/user_gpio_oeb gpio_control_in\[5\]/user_gpio_out gpio_control_in\[5\]/zero
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[37\] soc/mgmt_in_data[37] gpio_control_in\[37\]/one soc/mgmt_in_data[37]
+ gpio_control_in\[37\]/one padframe/mprj_io_analog_en[37] padframe/mprj_io_analog_pol[37]
+ padframe/mprj_io_analog_sel[37] padframe/mprj_io_dm[111] padframe/mprj_io_dm[112]
+ padframe/mprj_io_dm[113] padframe/mprj_io_holdover[37] padframe/mprj_io_ib_mode_sel[37]
+ padframe/mprj_io_in[37] padframe/mprj_io_inp_dis[37] padframe/mprj_io_out[37] padframe/mprj_io_oeb[37]
+ padframe/mprj_io_slow_sel[37] padframe/mprj_io_vtrip_sel[37] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[37\]/serial_data_in gpio_control_in\[37\]/serial_data_out
+ gpio_control_in\[37\]/user_gpio_in gpio_control_in\[37\]/user_gpio_oeb gpio_control_in\[37\]/user_gpio_out
+ gpio_control_in\[37\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[12\] soc/mgmt_in_data[12] gpio_control_in\[12\]/one soc/mgmt_in_data[12]
+ gpio_control_in\[12\]/one padframe/mprj_io_analog_en[12] padframe/mprj_io_analog_pol[12]
+ padframe/mprj_io_analog_sel[12] padframe/mprj_io_dm[36] padframe/mprj_io_dm[37]
+ padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12] padframe/mprj_io_ib_mode_sel[12]
+ padframe/mprj_io_in[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_out[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[12\]/serial_data_in gpio_control_in\[13\]/serial_data_in
+ gpio_control_in\[12\]/user_gpio_in gpio_control_in\[12\]/user_gpio_oeb gpio_control_in\[12\]/user_gpio_out
+ gpio_control_in\[12\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xstorage soc/mgmt_addr[0] soc/mgmt_addr[1] soc/mgmt_addr[2] soc/mgmt_addr[3] soc/mgmt_addr[4]
+ soc/mgmt_addr[5] soc/mgmt_addr[6] soc/mgmt_addr[7] soc/mgmt_addr_ro[0] soc/mgmt_addr_ro[1]
+ soc/mgmt_addr_ro[2] soc/mgmt_addr_ro[3] soc/mgmt_addr_ro[4] soc/mgmt_addr_ro[5]
+ soc/mgmt_addr_ro[6] soc/mgmt_addr_ro[7] soc/user_clk soc/mgmt_ena[0] soc/mgmt_ena[1]
+ soc/mgmt_ena_ro soc/mgmt_rdata[0] soc/mgmt_rdata[10] soc/mgmt_rdata[11] soc/mgmt_rdata[12]
+ soc/mgmt_rdata[13] soc/mgmt_rdata[14] soc/mgmt_rdata[15] soc/mgmt_rdata[16] soc/mgmt_rdata[17]
+ soc/mgmt_rdata[18] soc/mgmt_rdata[19] soc/mgmt_rdata[1] soc/mgmt_rdata[20] soc/mgmt_rdata[21]
+ soc/mgmt_rdata[22] soc/mgmt_rdata[23] soc/mgmt_rdata[24] soc/mgmt_rdata[25] soc/mgmt_rdata[26]
+ soc/mgmt_rdata[27] soc/mgmt_rdata[28] soc/mgmt_rdata[29] soc/mgmt_rdata[2] soc/mgmt_rdata[30]
+ soc/mgmt_rdata[31] soc/mgmt_rdata[32] soc/mgmt_rdata[33] soc/mgmt_rdata[34] soc/mgmt_rdata[35]
+ soc/mgmt_rdata[36] soc/mgmt_rdata[37] soc/mgmt_rdata[38] soc/mgmt_rdata[39] soc/mgmt_rdata[3]
+ soc/mgmt_rdata[40] soc/mgmt_rdata[41] soc/mgmt_rdata[42] soc/mgmt_rdata[43] soc/mgmt_rdata[44]
+ soc/mgmt_rdata[45] soc/mgmt_rdata[46] soc/mgmt_rdata[47] soc/mgmt_rdata[48] soc/mgmt_rdata[49]
+ soc/mgmt_rdata[4] soc/mgmt_rdata[50] soc/mgmt_rdata[51] soc/mgmt_rdata[52] soc/mgmt_rdata[53]
+ soc/mgmt_rdata[54] soc/mgmt_rdata[55] soc/mgmt_rdata[56] soc/mgmt_rdata[57] soc/mgmt_rdata[58]
+ soc/mgmt_rdata[59] soc/mgmt_rdata[5] soc/mgmt_rdata[60] soc/mgmt_rdata[61] soc/mgmt_rdata[62]
+ soc/mgmt_rdata[63] soc/mgmt_rdata[6] soc/mgmt_rdata[7] soc/mgmt_rdata[8] soc/mgmt_rdata[9]
+ soc/mgmt_rdata_ro[0] soc/mgmt_rdata_ro[10] soc/mgmt_rdata_ro[11] soc/mgmt_rdata_ro[12]
+ soc/mgmt_rdata_ro[13] soc/mgmt_rdata_ro[14] soc/mgmt_rdata_ro[15] soc/mgmt_rdata_ro[16]
+ soc/mgmt_rdata_ro[17] soc/mgmt_rdata_ro[18] soc/mgmt_rdata_ro[19] soc/mgmt_rdata_ro[1]
+ soc/mgmt_rdata_ro[20] soc/mgmt_rdata_ro[21] soc/mgmt_rdata_ro[22] soc/mgmt_rdata_ro[23]
+ soc/mgmt_rdata_ro[24] soc/mgmt_rdata_ro[25] soc/mgmt_rdata_ro[26] soc/mgmt_rdata_ro[27]
+ soc/mgmt_rdata_ro[28] soc/mgmt_rdata_ro[29] soc/mgmt_rdata_ro[2] soc/mgmt_rdata_ro[30]
+ soc/mgmt_rdata_ro[31] soc/mgmt_rdata_ro[3] soc/mgmt_rdata_ro[4] soc/mgmt_rdata_ro[5]
+ soc/mgmt_rdata_ro[6] soc/mgmt_rdata_ro[7] soc/mgmt_rdata_ro[8] soc/mgmt_rdata_ro[9]
+ soc/mgmt_wdata[0] soc/mgmt_wdata[10] soc/mgmt_wdata[11] soc/mgmt_wdata[12] soc/mgmt_wdata[13]
+ soc/mgmt_wdata[14] soc/mgmt_wdata[15] soc/mgmt_wdata[16] soc/mgmt_wdata[17] soc/mgmt_wdata[18]
+ soc/mgmt_wdata[19] soc/mgmt_wdata[1] soc/mgmt_wdata[20] soc/mgmt_wdata[21] soc/mgmt_wdata[22]
+ soc/mgmt_wdata[23] soc/mgmt_wdata[24] soc/mgmt_wdata[25] soc/mgmt_wdata[26] soc/mgmt_wdata[27]
+ soc/mgmt_wdata[28] soc/mgmt_wdata[29] soc/mgmt_wdata[2] soc/mgmt_wdata[30] soc/mgmt_wdata[31]
+ soc/mgmt_wdata[3] soc/mgmt_wdata[4] soc/mgmt_wdata[5] soc/mgmt_wdata[6] soc/mgmt_wdata[7]
+ soc/mgmt_wdata[8] soc/mgmt_wdata[9] soc/mgmt_wen[0] soc/mgmt_wen[1] soc/mgmt_wen_mask[0]
+ soc/mgmt_wen_mask[1] soc/mgmt_wen_mask[2] soc/mgmt_wen_mask[3] soc/mgmt_wen_mask[4]
+ soc/mgmt_wen_mask[5] soc/mgmt_wen_mask[6] soc/mgmt_wen_mask[7] soc/VPWR por/vss
+ storage
Xgpio_control_in\[35\] soc/mgmt_in_data[35] gpio_control_in\[35\]/one soc/mgmt_in_data[35]
+ gpio_control_in\[35\]/one padframe/mprj_io_analog_en[35] padframe/mprj_io_analog_pol[35]
+ padframe/mprj_io_analog_sel[35] padframe/mprj_io_dm[105] padframe/mprj_io_dm[106]
+ padframe/mprj_io_dm[107] padframe/mprj_io_holdover[35] padframe/mprj_io_ib_mode_sel[35]
+ padframe/mprj_io_in[35] padframe/mprj_io_inp_dis[35] padframe/mprj_io_out[35] padframe/mprj_io_oeb[35]
+ padframe/mprj_io_slow_sel[35] padframe/mprj_io_vtrip_sel[35] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[35\]/serial_data_in gpio_control_in\[36\]/serial_data_in
+ gpio_control_in\[35\]/user_gpio_in gpio_control_in\[35\]/user_gpio_oeb gpio_control_in\[35\]/user_gpio_out
+ gpio_control_in\[35\]/zero soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
Xgpio_control_in\[3\] soc/mgmt_in_data[3] gpio_control_in\[3\]/one soc/mgmt_in_data[3]
+ gpio_control_in\[3\]/one padframe/mprj_io_analog_en[3] padframe/mprj_io_analog_pol[3]
+ padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[9] padframe/mprj_io_dm[10] padframe/mprj_io_dm[11]
+ padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3] padframe/mprj_io_in[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_out[3] padframe/mprj_io_oeb[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[3\]/serial_data_in gpio_control_in\[4\]/serial_data_in gpio_control_in\[3\]/user_gpio_in
+ gpio_control_in\[3\]/user_gpio_oeb gpio_control_in\[3\]/user_gpio_out gpio_control_in\[3\]/zero
+ soc/VPWR por/vss mprj/vccd1 mprj/vssd1 gpio_control_block
.ends

