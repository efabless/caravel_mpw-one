VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_io_alt
  CLASS BLOCK ;
  FOREIGN chip_io_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 938.200 32.990 1000.900 95.440 ;
    END
  END clock
  PIN clock_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.635 208.565 936.915 210.965 ;
    END
  END clock_core
  PIN por
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.215 208.565 970.495 210.965 ;
    END
  END por
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1755.200 32.990 1817.900 95.440 ;
    END
  END flash_clk
  PIN flash_clk_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.835 208.565 1809.115 210.965 ;
    END
  END flash_clk_core
  PIN flash_clk_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.215 208.565 1787.495 210.965 ;
    END
  END flash_clk_ieb_core
  PIN flash_clk_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.475 208.565 1824.755 210.965 ;
    END
  END flash_clk_oeb_core
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1481.200 32.990 1543.900 95.440 ;
    END
  END flash_csb
  PIN flash_csb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.835 208.565 1535.115 210.965 ;
    END
  END flash_csb_core
  PIN flash_csb_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.215 208.565 1513.495 210.965 ;
    END
  END flash_csb_ieb_core
  PIN flash_csb_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.475 208.565 1550.755 210.965 ;
    END
  END flash_csb_oeb_core
  PIN flash_io0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2029.200 32.990 2091.900 95.440 ;
    END
  END flash_io0
  PIN flash_io0_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.635 208.565 2027.915 210.965 ;
    END
  END flash_io0_di_core
  PIN flash_io0_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.835 208.565 2083.115 210.965 ;
    END
  END flash_io0_do_core
  PIN flash_io0_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2046.610 209.000 2046.930 209.060 ;
        RECT 2061.790 209.000 2062.110 209.060 ;
        RECT 2076.050 209.000 2076.370 209.060 ;
        RECT 2046.610 208.860 2076.370 209.000 ;
        RECT 2046.610 208.800 2046.930 208.860 ;
        RECT 2061.790 208.800 2062.110 208.860 ;
        RECT 2076.050 208.800 2076.370 208.860 ;
      LAYER via ;
        RECT 2046.640 208.800 2046.900 209.060 ;
        RECT 2061.820 208.800 2062.080 209.060 ;
        RECT 2076.080 208.800 2076.340 209.060 ;
      LAYER met2 ;
        RECT 2046.035 209.170 2046.315 210.965 ;
        RECT 2061.215 209.170 2061.495 210.965 ;
        RECT 2076.855 209.170 2077.135 210.965 ;
        RECT 2046.035 209.090 2046.840 209.170 ;
        RECT 2061.215 209.090 2062.020 209.170 ;
        RECT 2076.140 209.090 2077.135 209.170 ;
        RECT 2046.035 209.030 2046.900 209.090 ;
        RECT 2046.035 208.565 2046.315 209.030 ;
        RECT 2046.640 208.770 2046.900 209.030 ;
        RECT 2061.215 209.030 2062.080 209.090 ;
        RECT 2061.215 208.565 2061.495 209.030 ;
        RECT 2061.820 208.770 2062.080 209.030 ;
        RECT 2076.080 209.030 2077.135 209.090 ;
        RECT 2076.080 208.770 2076.340 209.030 ;
        RECT 2076.855 208.565 2077.135 209.030 ;
    END
  END flash_io0_ieb_core
  PIN flash_io0_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2055.370 221.835 2055.650 222.205 ;
        RECT 2098.610 221.835 2098.890 222.205 ;
        RECT 2055.440 210.965 2055.580 221.835 ;
        RECT 2098.680 210.965 2098.820 221.835 ;
        RECT 2055.235 209.100 2055.580 210.965 ;
        RECT 2098.475 209.100 2098.820 210.965 ;
        RECT 2055.235 208.565 2055.515 209.100 ;
        RECT 2098.475 208.565 2098.755 209.100 ;
      LAYER via2 ;
        RECT 2055.370 221.880 2055.650 222.160 ;
        RECT 2098.610 221.880 2098.890 222.160 ;
      LAYER met3 ;
        RECT 2055.345 222.170 2055.675 222.185 ;
        RECT 2098.585 222.170 2098.915 222.185 ;
        RECT 2055.345 221.870 2098.915 222.170 ;
        RECT 2055.345 221.855 2055.675 221.870 ;
        RECT 2098.585 221.855 2098.915 221.870 ;
    END
  END flash_io0_oeb_core
  PIN flash_io1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2303.200 32.990 2365.900 95.440 ;
    END
  END flash_io1
  PIN flash_io1_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.635 208.565 2301.915 210.965 ;
    END
  END flash_io1_di_core
  PIN flash_io1_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.835 208.565 2357.115 210.965 ;
    END
  END flash_io1_do_core
  PIN flash_io1_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2320.770 209.000 2321.090 209.060 ;
        RECT 2335.950 209.000 2336.270 209.060 ;
        RECT 2350.210 209.000 2350.530 209.060 ;
        RECT 2320.770 208.860 2350.530 209.000 ;
        RECT 2320.770 208.800 2321.090 208.860 ;
        RECT 2335.950 208.800 2336.270 208.860 ;
        RECT 2350.210 208.800 2350.530 208.860 ;
      LAYER via ;
        RECT 2320.800 208.800 2321.060 209.060 ;
        RECT 2335.980 208.800 2336.240 209.060 ;
        RECT 2350.240 208.800 2350.500 209.060 ;
      LAYER met2 ;
        RECT 2320.035 209.170 2320.315 210.965 ;
        RECT 2335.215 209.170 2335.495 210.965 ;
        RECT 2350.855 209.170 2351.135 210.965 ;
        RECT 2320.035 209.090 2321.000 209.170 ;
        RECT 2335.215 209.090 2336.180 209.170 ;
        RECT 2350.300 209.090 2351.135 209.170 ;
        RECT 2320.035 209.030 2321.060 209.090 ;
        RECT 2320.035 208.565 2320.315 209.030 ;
        RECT 2320.800 208.770 2321.060 209.030 ;
        RECT 2335.215 209.030 2336.240 209.090 ;
        RECT 2335.215 208.565 2335.495 209.030 ;
        RECT 2335.980 208.770 2336.240 209.030 ;
        RECT 2350.240 209.030 2351.135 209.090 ;
        RECT 2350.240 208.770 2350.500 209.030 ;
        RECT 2350.855 208.565 2351.135 209.030 ;
    END
  END flash_io1_ieb_core
  PIN flash_io1_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.070 221.835 2329.350 222.205 ;
        RECT 2372.310 221.835 2372.590 222.205 ;
        RECT 2329.140 210.965 2329.280 221.835 ;
        RECT 2372.380 210.965 2372.520 221.835 ;
        RECT 2329.140 209.030 2329.515 210.965 ;
        RECT 2372.380 209.030 2372.755 210.965 ;
        RECT 2329.235 208.565 2329.515 209.030 ;
        RECT 2372.475 208.565 2372.755 209.030 ;
      LAYER via2 ;
        RECT 2329.070 221.880 2329.350 222.160 ;
        RECT 2372.310 221.880 2372.590 222.160 ;
      LAYER met3 ;
        RECT 2329.045 222.170 2329.375 222.185 ;
        RECT 2372.285 222.170 2372.615 222.185 ;
        RECT 2329.045 221.870 2372.615 222.170 ;
        RECT 2329.045 221.855 2329.375 221.870 ;
        RECT 2372.285 221.855 2372.615 221.870 ;
    END
  END flash_io1_oeb_core
  PIN gpio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2577.200 32.990 2639.900 95.440 ;
    END
  END gpio
  PIN gpio_in_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.635 208.565 2575.915 210.965 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.215 208.565 2609.495 210.965 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.235 208.565 2603.515 210.965 ;
    END
  END gpio_mode0_core
  PIN gpio_mode1_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2594.030 221.155 2594.310 221.525 ;
        RECT 2624.850 221.155 2625.130 221.525 ;
        RECT 2594.100 210.965 2594.240 221.155 ;
        RECT 2624.920 210.965 2625.060 221.155 ;
        RECT 2594.035 208.565 2594.315 210.965 ;
        RECT 2624.855 208.565 2625.135 210.965 ;
      LAYER via2 ;
        RECT 2594.030 221.200 2594.310 221.480 ;
        RECT 2624.850 221.200 2625.130 221.480 ;
      LAYER met3 ;
        RECT 2594.005 221.490 2594.335 221.505 ;
        RECT 2624.825 221.490 2625.155 221.505 ;
        RECT 2594.005 221.190 2625.155 221.490 ;
        RECT 2594.005 221.175 2594.335 221.190 ;
        RECT 2624.825 221.175 2625.155 221.190 ;
    END
  END gpio_mode1_core
  PIN gpio_out_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2630.835 208.565 2631.115 210.965 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.475 208.565 2646.755 210.965 ;
    END
  END gpio_outenb_core
  PIN vccd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 350.270 98.100 404.670 ;
    END
  END vccd_pad
  PIN vdda_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3121.110 34.055 3181.950 94.880 ;
    END
  END vdda_pad
  PIN vddio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 558.050 94.880 618.890 ;
    END
  END vddio_pad
  PIN vddio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4356.050 94.880 4416.890 ;
    END
  END vddio_pad2
  PIN vssa_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 401.110 34.055 461.950 94.880 ;
    END
  END vssa_pad
  PIN vssd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1216.330 30.835 1270.730 98.100 ;
    END
  END vssd_pad
  PIN vssio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2852.110 34.055 2912.950 94.880 ;
    END
  END vssio_pad
  PIN vssio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1674.050 5093.120 1734.890 5153.945 ;
    END
  END vssio_pad2
  PIN mprj_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 506.200 3555.010 568.900 ;
    END
  END mprj_io[0]
  PIN mprj_io_analog_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 529.015 3379.435 529.295 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_pol[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 535.455 3379.435 535.735 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 550.635 3379.435 550.915 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_dm[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 532.235 3379.435 532.515 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 523.035 3379.435 523.315 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 553.855 3379.435 554.135 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_holdover[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 557.075 3379.435 557.355 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 572.255 3379.435 572.535 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_inp_dis[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 538.215 3379.435 538.495 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 575.475 3379.435 575.755 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 559.835 3379.435 560.115 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_slow_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 513.835 3379.435 514.115 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 569.035 3379.435 569.315 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 504.635 3379.435 504.915 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in_3v3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 578.235 3379.435 578.515 ;
    END
  END mprj_io_in_3v3[0]
  PIN mprj_gpio_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3433.055 3379.435 3433.335 ;
    END
  END mprj_gpio_analog[3]
  PIN mprj_gpio_noesd[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3442.255 3379.435 3442.535 ;
    END
  END mprj_gpio_noesd[3]
  PIN mprj_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3422.200 3555.010 3484.900 ;
    END
  END mprj_io[10]
  PIN mprj_io_analog_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3445.015 3379.435 3445.295 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_pol[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3451.455 3379.435 3451.735 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3466.635 3379.435 3466.915 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_dm[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3448.235 3379.435 3448.515 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3439.035 3379.435 3439.315 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3469.855 3379.435 3470.135 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_holdover[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3473.075 3379.435 3473.355 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3488.255 3379.435 3488.535 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_inp_dis[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3454.215 3379.435 3454.495 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3491.475 3379.435 3491.755 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3475.835 3379.435 3476.115 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_slow_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3429.835 3379.435 3430.115 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3485.035 3379.435 3485.315 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3420.635 3379.435 3420.915 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in_3v3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3494.235 3379.435 3494.515 ;
    END
  END mprj_io_in_3v3[10]
  PIN mprj_gpio_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3658.055 3379.435 3658.335 ;
    END
  END mprj_gpio_analog[4]
  PIN mprj_gpio_noesd[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3667.255 3379.435 3667.535 ;
    END
  END mprj_gpio_noesd[4]
  PIN mprj_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3647.200 3555.010 3709.900 ;
    END
  END mprj_io[11]
  PIN mprj_io_analog_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3670.015 3379.435 3670.295 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_pol[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3676.455 3379.435 3676.735 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3691.635 3379.435 3691.915 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_dm[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3673.235 3379.435 3673.515 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3664.035 3379.435 3664.315 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3694.855 3379.435 3695.135 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_holdover[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3698.075 3379.435 3698.355 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3713.255 3379.435 3713.535 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_inp_dis[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3679.215 3379.435 3679.495 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3716.475 3379.435 3716.755 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3700.835 3379.435 3701.115 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_slow_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3654.835 3379.435 3655.115 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3710.035 3379.435 3710.315 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3645.635 3379.435 3645.915 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in_3v3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3719.235 3379.435 3719.515 ;
    END
  END mprj_io_in_3v3[11]
  PIN mprj_gpio_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3883.055 3379.435 3883.335 ;
    END
  END mprj_gpio_analog[5]
  PIN mprj_gpio_noesd[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3892.255 3379.435 3892.535 ;
    END
  END mprj_gpio_noesd[5]
  PIN mprj_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3872.200 3555.010 3934.900 ;
    END
  END mprj_io[12]
  PIN mprj_io_analog_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3895.015 3379.435 3895.295 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_pol[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3901.455 3379.435 3901.735 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3916.635 3379.435 3916.915 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_dm[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3898.235 3379.435 3898.515 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3889.035 3379.435 3889.315 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3919.855 3379.435 3920.135 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_holdover[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3923.075 3379.435 3923.355 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3938.255 3379.435 3938.535 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_inp_dis[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3904.215 3379.435 3904.495 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3941.475 3379.435 3941.755 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3925.835 3379.435 3926.115 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_slow_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3879.835 3379.435 3880.115 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3935.035 3379.435 3935.315 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3870.635 3379.435 3870.915 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in_3v3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3944.235 3379.435 3944.515 ;
    END
  END mprj_io_in_3v3[12]
  PIN mprj_gpio_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4329.055 3379.435 4329.335 ;
    END
  END mprj_gpio_analog[6]
  PIN mprj_gpio_noesd[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4338.255 3379.435 4338.535 ;
    END
  END mprj_gpio_noesd[6]
  PIN mprj_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4318.200 3555.010 4380.900 ;
    END
  END mprj_io[13]
  PIN mprj_io_analog_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4341.015 3379.435 4341.295 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_pol[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4347.455 3379.435 4347.735 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4362.635 3379.435 4362.915 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_dm[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4344.235 3379.435 4344.515 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4335.035 3379.435 4335.315 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4365.855 3379.435 4366.135 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_holdover[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4369.075 3379.435 4369.355 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4384.255 3379.435 4384.535 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_inp_dis[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4350.215 3379.435 4350.495 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4387.475 3379.435 4387.755 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4371.835 3379.435 4372.115 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_slow_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4325.835 3379.435 4326.115 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4381.035 3379.435 4381.315 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4316.635 3379.435 4316.915 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in_3v3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4390.235 3379.435 4390.515 ;
    END
  END mprj_io_in_3v3[13]
  PIN mprj_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 732.200 3555.010 794.900 ;
    END
  END mprj_io[1]
  PIN mprj_io_analog_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 755.015 3379.435 755.295 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_pol[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 761.455 3379.435 761.735 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 776.635 3379.435 776.915 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_dm[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 758.235 3379.435 758.515 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 749.035 3379.435 749.315 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 779.855 3379.435 780.135 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_holdover[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 783.075 3379.435 783.355 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 798.255 3379.435 798.535 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_inp_dis[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 764.215 3379.435 764.495 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 801.475 3379.435 801.755 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 785.835 3379.435 786.115 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_slow_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 739.835 3379.435 740.115 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 795.035 3379.435 795.315 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 730.635 3379.435 730.915 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in_3v3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 804.235 3379.435 804.515 ;
    END
  END mprj_io_in_3v3[1]
  PIN mprj_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 957.200 3555.010 1019.900 ;
    END
  END mprj_io[2]
  PIN mprj_io_analog_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 980.015 3379.435 980.295 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_pol[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 986.455 3379.435 986.735 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1001.635 3379.435 1001.915 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_dm[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 983.235 3379.435 983.515 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 974.035 3379.435 974.315 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1004.855 3379.435 1005.135 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_holdover[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1008.075 3379.435 1008.355 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1023.255 3379.435 1023.535 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_inp_dis[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 989.215 3379.435 989.495 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1026.475 3379.435 1026.755 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1010.835 3379.435 1011.115 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_slow_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 964.835 3379.435 965.115 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1020.035 3379.435 1020.315 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 955.635 3379.435 955.915 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in_3v3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1029.235 3379.435 1029.515 ;
    END
  END mprj_io_in_3v3[2]
  PIN mprj_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1183.200 3555.010 1245.900 ;
    END
  END mprj_io[3]
  PIN mprj_io_analog_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1206.015 3379.435 1206.295 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_pol[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1212.455 3379.435 1212.735 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1227.635 3379.435 1227.915 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_dm[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1200.035 3379.435 1200.315 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1230.855 3379.435 1231.135 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1209.235 3379.435 1209.515 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1234.075 3379.435 1234.355 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1249.255 3379.435 1249.535 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_inp_dis[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1215.215 3379.435 1215.495 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1252.475 3379.435 1252.755 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1236.835 3379.435 1237.115 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_slow_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1190.835 3379.435 1191.115 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1246.035 3379.435 1246.315 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1181.635 3379.435 1181.915 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in_3v3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1255.235 3379.435 1255.515 ;
    END
  END mprj_io_in_3v3[3]
  PIN mprj_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1408.200 3555.010 1470.900 ;
    END
  END mprj_io[4]
  PIN mprj_io_analog_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1431.015 3379.435 1431.295 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_pol[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1437.455 3379.435 1437.735 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1452.635 3379.435 1452.915 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_dm[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1434.235 3379.435 1434.515 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1425.035 3379.435 1425.315 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1455.855 3379.435 1456.135 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_holdover[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1459.075 3379.435 1459.355 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1474.255 3379.435 1474.535 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_inp_dis[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1440.215 3379.435 1440.495 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1477.475 3379.435 1477.755 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1461.835 3379.435 1462.115 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_slow_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1415.835 3379.435 1416.115 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1471.035 3379.435 1471.315 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1406.635 3379.435 1406.915 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in_3v3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1480.235 3379.435 1480.515 ;
    END
  END mprj_io_in_3v3[4]
  PIN mprj_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1633.200 3555.010 1695.900 ;
    END
  END mprj_io[5]
  PIN mprj_io_analog_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1656.015 3379.435 1656.295 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_pol[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1662.455 3379.435 1662.735 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1677.635 3379.435 1677.915 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_dm[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1659.235 3379.435 1659.515 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1650.035 3379.435 1650.315 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1680.855 3379.435 1681.135 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_holdover[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1684.075 3379.435 1684.355 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1699.255 3379.435 1699.535 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_inp_dis[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1665.215 3379.435 1665.495 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1702.475 3379.435 1702.755 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1686.835 3379.435 1687.115 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_slow_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1640.835 3379.435 1641.115 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1696.035 3379.435 1696.315 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1631.635 3379.435 1631.915 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in_3v3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1705.235 3379.435 1705.515 ;
    END
  END mprj_io_in_3v3[5]
  PIN mprj_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1859.200 3555.010 1921.900 ;
    END
  END mprj_io[6]
  PIN mprj_io_analog_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1882.015 3379.435 1882.295 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_pol[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1888.455 3379.435 1888.735 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1903.635 3379.435 1903.915 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_dm[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1885.235 3379.435 1885.515 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1876.035 3379.435 1876.315 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1906.855 3379.435 1907.135 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_holdover[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1910.075 3379.435 1910.355 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1925.255 3379.435 1925.535 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_inp_dis[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1891.215 3379.435 1891.495 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1928.475 3379.435 1928.755 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1912.835 3379.435 1913.115 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_slow_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1866.835 3379.435 1867.115 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1922.035 3379.435 1922.315 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1857.635 3379.435 1857.915 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in_3v3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1931.235 3379.435 1931.515 ;
    END
  END mprj_io_in_3v3[6]
  PIN mprj_gpio_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2756.055 3379.435 2756.335 ;
    END
  END mprj_gpio_analog[0]
  PIN mprj_gpio_noesd[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2765.255 3379.435 2765.535 ;
    END
  END mprj_gpio_noesd[0]
  PIN mprj_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2745.200 3555.010 2807.900 ;
    END
  END mprj_io[7]
  PIN mprj_io_analog_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2768.015 3379.435 2768.295 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_pol[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2774.455 3379.435 2774.735 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2789.635 3379.435 2789.915 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_dm[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2771.235 3379.435 2771.515 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2762.035 3379.435 2762.315 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2792.855 3379.435 2793.135 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_holdover[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2796.075 3379.435 2796.355 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2811.255 3379.435 2811.535 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_inp_dis[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2777.215 3379.435 2777.495 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2814.475 3379.435 2814.755 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2798.835 3379.435 2799.115 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_slow_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2752.835 3379.435 2753.115 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2808.035 3379.435 2808.315 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2743.635 3379.435 2743.915 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in_3v3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2817.235 3379.435 2817.515 ;
    END
  END mprj_io_in_3v3[7]
  PIN mprj_gpio_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2982.055 3379.435 2982.335 ;
    END
  END mprj_gpio_analog[1]
  PIN mprj_gpio_noesd[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2991.255 3379.435 2991.535 ;
    END
  END mprj_gpio_noesd[1]
  PIN mprj_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2971.200 3555.010 3033.900 ;
    END
  END mprj_io[8]
  PIN mprj_io_analog_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2994.015 3379.435 2994.295 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_pol[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3000.455 3379.435 3000.735 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3015.635 3379.435 3015.915 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_dm[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2997.235 3379.435 2997.515 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2988.035 3379.435 2988.315 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3018.855 3379.435 3019.135 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_holdover[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3022.075 3379.435 3022.355 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3037.255 3379.435 3037.535 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_inp_dis[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3003.215 3379.435 3003.495 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3040.475 3379.435 3040.755 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3024.835 3379.435 3025.115 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_slow_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2978.835 3379.435 2979.115 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3034.035 3379.435 3034.315 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2969.635 3379.435 2969.915 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in_3v3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3043.235 3379.435 3043.515 ;
    END
  END mprj_io_in_3v3[8]
  PIN mprj_gpio_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3207.055 3379.435 3207.335 ;
    END
  END mprj_gpio_analog[2]
  PIN mprj_gpio_noesd[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3216.255 3379.435 3216.535 ;
    END
  END mprj_gpio_noesd[2]
  PIN mprj_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3196.200 3555.010 3258.900 ;
    END
  END mprj_io[9]
  PIN mprj_io_analog_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3219.015 3379.435 3219.295 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3225.455 3379.435 3225.735 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3240.635 3379.435 3240.915 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3222.235 3379.435 3222.515 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3213.035 3379.435 3213.315 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3243.855 3379.435 3244.135 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_holdover[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3247.075 3379.435 3247.355 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3262.255 3379.435 3262.535 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_inp_dis[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3228.215 3379.435 3228.495 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3265.475 3379.435 3265.755 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3249.835 3379.435 3250.115 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3203.835 3379.435 3204.115 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3259.035 3379.435 3259.315 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN mprj_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3194.635 3379.435 3194.915 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_in_3v3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3268.235 3379.435 3268.515 ;
    END
  END mprj_io_in_3v3[9]
  PIN mprj_gpio_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3984.665 210.965 3984.945 ;
    END
  END mprj_gpio_analog[7]
  PIN mprj_gpio_noesd[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3975.465 210.965 3975.745 ;
    END
  END mprj_gpio_noesd[7]
  PIN mprj_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3933.100 95.440 3995.800 ;
    END
  END mprj_io[25]
  PIN mprj_io_analog_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3972.705 210.965 3972.985 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_pol[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3966.265 210.965 3966.545 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3951.085 210.965 3951.365 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_dm[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3969.485 210.965 3969.765 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3978.685 210.965 3978.965 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3947.865 210.965 3948.145 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_holdover[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3944.645 210.965 3944.925 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3929.465 210.965 3929.745 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_inp_dis[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3963.505 210.965 3963.785 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3926.245 210.965 3926.525 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3941.885 210.965 3942.165 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_slow_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3987.885 210.965 3988.165 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3932.685 210.965 3932.965 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3997.085 210.965 3997.365 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in_3v3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3923.485 210.965 3923.765 ;
    END
  END mprj_io_in_3v3[14]
  PIN mprj_gpio_analog[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1402.665 210.965 1402.945 ;
    END
  END mprj_gpio_analog[17]
  PIN mprj_gpio_noesd[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1393.465 210.965 1393.745 ;
    END
  END mprj_gpio_noesd[17]
  PIN mprj_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1351.100 95.440 1413.800 ;
    END
  END mprj_io[35]
  PIN mprj_io_analog_en[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1390.705 210.965 1390.985 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_pol[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1384.265 210.965 1384.545 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1369.085 210.965 1369.365 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_dm[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1387.485 210.965 1387.765 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1396.685 210.965 1396.965 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1365.865 210.965 1366.145 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_holdover[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1362.645 210.965 1362.925 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1347.465 210.965 1347.745 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_inp_dis[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1381.505 210.965 1381.785 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1344.245 210.965 1344.525 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1359.885 210.965 1360.165 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_slow_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1405.885 210.965 1406.165 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1350.685 210.965 1350.965 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1415.085 210.965 1415.365 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in_3v3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1341.485 210.965 1341.765 ;
    END
  END mprj_io_in_3v3[24]
  PIN mprj_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1135.100 95.440 1197.800 ;
    END
  END mprj_io[36]
  PIN mprj_io_analog_en[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1174.705 210.965 1174.985 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_pol[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1168.265 210.965 1168.545 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1153.085 210.965 1153.365 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_dm[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1171.485 210.965 1171.765 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1180.685 210.965 1180.965 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1149.865 210.965 1150.145 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_holdover[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1146.645 210.965 1146.925 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1131.465 210.965 1131.745 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_inp_dis[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1165.505 210.965 1165.785 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1128.245 210.965 1128.525 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1143.885 210.965 1144.165 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_slow_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1189.885 210.965 1190.165 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1134.685 210.965 1134.965 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1199.085 210.965 1199.365 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in_3v3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1125.485 210.965 1125.765 ;
    END
  END mprj_io_in_3v3[25]
  PIN mprj_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 919.100 95.440 981.800 ;
    END
  END mprj_io[37]
  PIN mprj_io_analog_en[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 958.705 210.965 958.985 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_pol[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 952.265 210.965 952.545 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 937.085 210.965 937.365 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_dm[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 955.485 210.965 955.765 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 964.685 210.965 964.965 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 933.865 210.965 934.145 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_holdover[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 930.645 210.965 930.925 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 915.465 210.965 915.745 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_inp_dis[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 949.505 210.965 949.785 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 912.245 210.965 912.525 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 927.885 210.965 928.165 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_slow_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 973.885 210.965 974.165 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 918.685 210.965 918.965 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 983.085 210.965 983.365 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in_3v3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 909.485 210.965 909.765 ;
    END
  END mprj_io_in_3v3[26]
  PIN mprj_gpio_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3768.665 210.965 3768.945 ;
    END
  END mprj_gpio_analog[8]
  PIN mprj_gpio_noesd[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3759.465 210.965 3759.745 ;
    END
  END mprj_gpio_noesd[8]
  PIN mprj_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3717.100 95.440 3779.800 ;
    END
  END mprj_io[26]
  PIN mprj_io_analog_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3756.705 210.965 3756.985 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_pol[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3750.265 210.965 3750.545 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3735.085 210.965 3735.365 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_dm[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3753.485 210.965 3753.765 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3762.685 210.965 3762.965 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3731.865 210.965 3732.145 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_holdover[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3728.645 210.965 3728.925 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3713.465 210.965 3713.745 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_inp_dis[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3747.505 210.965 3747.785 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3710.245 210.965 3710.525 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3725.885 210.965 3726.165 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_slow_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3771.885 210.965 3772.165 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3716.685 210.965 3716.965 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3781.085 210.965 3781.365 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in_3v3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3707.485 210.965 3707.765 ;
    END
  END mprj_io_in_3v3[15]
  PIN mprj_gpio_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3552.665 210.965 3552.945 ;
    END
  END mprj_gpio_analog[9]
  PIN mprj_gpio_noesd[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3543.465 210.965 3543.745 ;
    END
  END mprj_gpio_noesd[9]
  PIN mprj_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3501.100 95.440 3563.800 ;
    END
  END mprj_io[27]
  PIN mprj_io_analog_en[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3540.705 210.965 3540.985 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_pol[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3534.265 210.965 3534.545 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3519.085 210.965 3519.365 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_dm[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3537.485 210.965 3537.765 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3546.685 210.965 3546.965 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3515.865 210.965 3516.145 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_holdover[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3512.645 210.965 3512.925 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3497.465 210.965 3497.745 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_inp_dis[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3531.505 210.965 3531.785 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3494.245 210.965 3494.525 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3509.885 210.965 3510.165 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_slow_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3555.885 210.965 3556.165 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3500.685 210.965 3500.965 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3565.085 210.965 3565.365 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in_3v3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3491.485 210.965 3491.765 ;
    END
  END mprj_io_in_3v3[16]
  PIN mprj_gpio_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3336.665 210.965 3336.945 ;
    END
  END mprj_gpio_analog[10]
  PIN mprj_gpio_noesd[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3327.465 210.965 3327.745 ;
    END
  END mprj_gpio_noesd[10]
  PIN mprj_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3285.100 95.440 3347.800 ;
    END
  END mprj_io[28]
  PIN mprj_io_analog_en[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3324.705 210.965 3324.985 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_pol[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3318.265 210.965 3318.545 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3303.085 210.965 3303.365 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_dm[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3321.485 210.965 3321.765 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3330.685 210.965 3330.965 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3299.865 210.965 3300.145 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_holdover[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3296.645 210.965 3296.925 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3281.465 210.965 3281.745 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_inp_dis[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3315.505 210.965 3315.785 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3278.245 210.965 3278.525 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3293.885 210.965 3294.165 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_slow_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3339.885 210.965 3340.165 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3284.685 210.965 3284.965 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3349.085 210.965 3349.365 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in_3v3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3275.485 210.965 3275.765 ;
    END
  END mprj_io_in_3v3[17]
  PIN mprj_gpio_analog[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3120.665 210.965 3120.945 ;
    END
  END mprj_gpio_analog[11]
  PIN mprj_gpio_noesd[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3111.465 210.965 3111.745 ;
    END
  END mprj_gpio_noesd[11]
  PIN mprj_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3069.100 95.440 3131.800 ;
    END
  END mprj_io[29]
  PIN mprj_io_analog_en[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3108.705 210.965 3108.985 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_pol[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3102.265 210.965 3102.545 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3087.085 210.965 3087.365 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_dm[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3105.485 210.965 3105.765 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3114.685 210.965 3114.965 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3083.865 210.965 3084.145 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_holdover[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3080.645 210.965 3080.925 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3065.465 210.965 3065.745 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_inp_dis[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3099.505 210.965 3099.785 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3062.245 210.965 3062.525 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3077.885 210.965 3078.165 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_slow_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3123.885 210.965 3124.165 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3068.685 210.965 3068.965 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3133.085 210.965 3133.365 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in_3v3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3059.485 210.965 3059.765 ;
    END
  END mprj_io_in_3v3[18]
  PIN mprj_gpio_analog[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2904.665 210.965 2904.945 ;
    END
  END mprj_gpio_analog[12]
  PIN mprj_gpio_noesd[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2895.465 210.965 2895.745 ;
    END
  END mprj_gpio_noesd[12]
  PIN mprj_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2853.100 95.440 2915.800 ;
    END
  END mprj_io[30]
  PIN mprj_io_analog_en[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2892.705 210.965 2892.985 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_pol[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2886.265 210.965 2886.545 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2871.085 210.965 2871.365 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_dm[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2889.485 210.965 2889.765 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2898.685 210.965 2898.965 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2867.865 210.965 2868.145 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_holdover[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2864.645 210.965 2864.925 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2849.465 210.965 2849.745 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_inp_dis[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2883.505 210.965 2883.785 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2846.245 210.965 2846.525 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2861.885 210.965 2862.165 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_slow_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2907.885 210.965 2908.165 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2852.685 210.965 2852.965 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2917.085 210.965 2917.365 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in_3v3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2843.485 210.965 2843.765 ;
    END
  END mprj_io_in_3v3[19]
  PIN mprj_gpio_analog[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2688.665 210.965 2688.945 ;
    END
  END mprj_gpio_analog[13]
  PIN mprj_gpio_noesd[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2679.465 210.965 2679.745 ;
    END
  END mprj_gpio_noesd[13]
  PIN mprj_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2637.100 95.440 2699.800 ;
    END
  END mprj_io[31]
  PIN mprj_io_analog_en[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2676.705 210.965 2676.985 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_pol[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2670.265 210.965 2670.545 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2655.085 210.965 2655.365 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_dm[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2673.485 210.965 2673.765 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2682.685 210.965 2682.965 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2651.865 210.965 2652.145 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_holdover[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2648.645 210.965 2648.925 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2633.465 210.965 2633.745 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_inp_dis[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2667.505 210.965 2667.785 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2630.245 210.965 2630.525 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2645.885 210.965 2646.165 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_slow_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2691.885 210.965 2692.165 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2636.685 210.965 2636.965 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2701.085 210.965 2701.365 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in_3v3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2627.485 210.965 2627.765 ;
    END
  END mprj_io_in_3v3[20]
  PIN mprj_gpio_analog[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2050.665 210.965 2050.945 ;
    END
  END mprj_gpio_analog[14]
  PIN mprj_gpio_noesd[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2041.465 210.965 2041.745 ;
    END
  END mprj_gpio_noesd[14]
  PIN mprj_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1999.100 95.440 2061.800 ;
    END
  END mprj_io[32]
  PIN mprj_io_analog_en[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2038.705 210.965 2038.985 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_pol[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2032.265 210.965 2032.545 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2017.085 210.965 2017.365 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_dm[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2035.485 210.965 2035.765 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2044.685 210.965 2044.965 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2013.865 210.965 2014.145 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_holdover[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2010.645 210.965 2010.925 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1995.465 210.965 1995.745 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_inp_dis[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2029.505 210.965 2029.785 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1992.245 210.965 1992.525 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2007.885 210.965 2008.165 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_slow_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2053.885 210.965 2054.165 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1998.685 210.965 1998.965 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2063.085 210.965 2063.365 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in_3v3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1989.485 210.965 1989.765 ;
    END
  END mprj_io_in_3v3[21]
  PIN mprj_gpio_analog[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1834.665 210.965 1834.945 ;
    END
  END mprj_gpio_analog[15]
  PIN mprj_gpio_noesd[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1825.465 210.965 1825.745 ;
    END
  END mprj_gpio_noesd[15]
  PIN mprj_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1783.100 95.440 1845.800 ;
    END
  END mprj_io[33]
  PIN mprj_io_analog_en[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1822.705 210.965 1822.985 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_pol[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1816.265 210.965 1816.545 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1801.085 210.965 1801.365 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_dm[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1819.485 210.965 1819.765 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1828.685 210.965 1828.965 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1797.865 210.965 1798.145 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_holdover[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1794.645 210.965 1794.925 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1779.465 210.965 1779.745 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_inp_dis[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1813.505 210.965 1813.785 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1776.245 210.965 1776.525 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1791.885 210.965 1792.165 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_slow_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1837.885 210.965 1838.165 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1782.685 210.965 1782.965 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1847.085 210.965 1847.365 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in_3v3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1773.485 210.965 1773.765 ;
    END
  END mprj_io_in_3v3[22]
  PIN mprj_gpio_analog[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1618.665 210.965 1618.945 ;
    END
  END mprj_gpio_analog[16]
  PIN mprj_gpio_noesd[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1609.465 210.965 1609.745 ;
    END
  END mprj_gpio_noesd[16]
  PIN mprj_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1567.100 95.440 1629.800 ;
    END
  END mprj_io[34]
  PIN mprj_io_analog_en[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1606.705 210.965 1606.985 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_pol[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1600.265 210.965 1600.545 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1585.085 210.965 1585.365 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_dm[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1603.485 210.965 1603.765 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1612.685 210.965 1612.965 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1581.865 210.965 1582.145 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_holdover[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1578.645 210.965 1578.925 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1563.465 210.965 1563.745 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_inp_dis[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1597.505 210.965 1597.785 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1560.245 210.965 1560.525 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1575.885 210.965 1576.165 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_slow_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1621.885 210.965 1622.165 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1566.685 210.965 1566.965 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1631.085 210.965 1631.365 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in_3v3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1557.485 210.965 1557.765 ;
    END
  END mprj_io_in_3v3[23]
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3368.650 4354.280 3368.970 4354.340 ;
        RECT 3376.930 4354.280 3377.250 4354.340 ;
        RECT 3368.650 4354.140 3377.250 4354.280 ;
        RECT 3368.650 4354.080 3368.970 4354.140 ;
        RECT 3376.930 4354.080 3377.250 4354.140 ;
        RECT 211.210 3936.420 211.530 3936.480 ;
        RECT 212.130 3936.420 212.450 3936.480 ;
        RECT 211.210 3936.280 212.450 3936.420 ;
        RECT 211.210 3936.220 211.530 3936.280 ;
        RECT 212.130 3936.220 212.450 3936.280 ;
        RECT 3368.650 3929.960 3368.970 3930.020 ;
        RECT 3376.010 3929.960 3376.330 3930.020 ;
        RECT 3376.930 3929.960 3377.250 3930.020 ;
        RECT 3368.650 3929.820 3377.250 3929.960 ;
        RECT 3368.650 3929.760 3368.970 3929.820 ;
        RECT 3376.010 3929.760 3376.330 3929.820 ;
        RECT 3376.930 3929.760 3377.250 3929.820 ;
        RECT 3368.650 3908.200 3368.970 3908.260 ;
        RECT 3376.010 3908.200 3376.330 3908.260 ;
        RECT 3376.930 3908.200 3377.250 3908.260 ;
        RECT 3368.650 3908.060 3377.250 3908.200 ;
        RECT 3368.650 3908.000 3368.970 3908.060 ;
        RECT 3376.010 3908.000 3376.330 3908.060 ;
        RECT 3376.930 3908.000 3377.250 3908.060 ;
        RECT 3368.650 3704.880 3368.970 3704.940 ;
        RECT 3376.010 3704.880 3376.330 3704.940 ;
        RECT 3376.930 3704.880 3377.250 3704.940 ;
        RECT 3368.650 3704.740 3377.250 3704.880 ;
        RECT 3368.650 3704.680 3368.970 3704.740 ;
        RECT 3376.010 3704.680 3376.330 3704.740 ;
        RECT 3376.930 3704.680 3377.250 3704.740 ;
        RECT 3368.650 3685.160 3368.970 3685.220 ;
        RECT 3376.010 3685.160 3376.330 3685.220 ;
        RECT 3376.930 3685.160 3377.250 3685.220 ;
        RECT 3368.650 3685.020 3377.250 3685.160 ;
        RECT 3368.650 3684.960 3368.970 3685.020 ;
        RECT 3376.010 3684.960 3376.330 3685.020 ;
        RECT 3376.930 3684.960 3377.250 3685.020 ;
        RECT 3368.650 3479.800 3368.970 3479.860 ;
        RECT 3376.010 3479.800 3376.330 3479.860 ;
        RECT 3376.930 3479.800 3377.250 3479.860 ;
        RECT 3368.650 3479.660 3377.250 3479.800 ;
        RECT 3368.650 3479.600 3368.970 3479.660 ;
        RECT 3376.010 3479.600 3376.330 3479.660 ;
        RECT 3376.930 3479.600 3377.250 3479.660 ;
        RECT 3368.650 3460.420 3368.970 3460.480 ;
        RECT 3376.010 3460.420 3376.330 3460.480 ;
        RECT 3376.930 3460.420 3377.250 3460.480 ;
        RECT 3368.650 3460.280 3377.250 3460.420 ;
        RECT 3368.650 3460.220 3368.970 3460.280 ;
        RECT 3376.010 3460.220 3376.330 3460.280 ;
        RECT 3376.930 3460.220 3377.250 3460.280 ;
        RECT 3368.650 3255.740 3368.970 3255.800 ;
        RECT 3376.930 3255.740 3377.250 3255.800 ;
        RECT 3368.650 3255.600 3377.250 3255.740 ;
        RECT 3368.650 3255.540 3368.970 3255.600 ;
        RECT 3376.930 3255.540 3377.250 3255.600 ;
        RECT 3368.650 3232.280 3368.970 3232.340 ;
        RECT 3376.930 3232.280 3377.250 3232.340 ;
        RECT 3368.650 3232.140 3377.250 3232.280 ;
        RECT 3368.650 3232.080 3368.970 3232.140 ;
        RECT 3376.930 3232.080 3377.250 3232.140 ;
        RECT 3368.650 3028.960 3368.970 3029.020 ;
        RECT 3376.010 3028.960 3376.330 3029.020 ;
        RECT 3376.930 3028.960 3377.250 3029.020 ;
        RECT 3368.650 3028.820 3377.250 3028.960 ;
        RECT 3368.650 3028.760 3368.970 3028.820 ;
        RECT 3376.010 3028.760 3376.330 3028.820 ;
        RECT 3376.930 3028.760 3377.250 3028.820 ;
        RECT 3368.650 3009.240 3368.970 3009.300 ;
        RECT 3376.010 3009.240 3376.330 3009.300 ;
        RECT 3376.930 3009.240 3377.250 3009.300 ;
        RECT 3368.650 3009.100 3377.250 3009.240 ;
        RECT 3368.650 3009.040 3368.970 3009.100 ;
        RECT 3376.010 3009.040 3376.330 3009.100 ;
        RECT 3376.930 3009.040 3377.250 3009.100 ;
        RECT 3368.650 2805.580 3368.970 2805.640 ;
        RECT 3376.010 2805.580 3376.330 2805.640 ;
        RECT 3368.650 2805.440 3376.330 2805.580 ;
        RECT 3368.650 2805.380 3368.970 2805.440 ;
        RECT 3376.010 2805.380 3376.330 2805.440 ;
        RECT 3368.190 2783.140 3368.510 2783.200 ;
        RECT 3376.010 2783.140 3376.330 2783.200 ;
        RECT 3376.930 2783.140 3377.250 2783.200 ;
        RECT 3368.190 2783.000 3377.250 2783.140 ;
        RECT 3368.190 2782.940 3368.510 2783.000 ;
        RECT 3376.010 2782.940 3376.330 2783.000 ;
        RECT 3376.930 2782.940 3377.250 2783.000 ;
        RECT 3368.190 1921.580 3368.510 1921.640 ;
        RECT 3376.930 1921.580 3377.250 1921.640 ;
        RECT 3368.190 1921.440 3377.250 1921.580 ;
        RECT 3368.190 1921.380 3368.510 1921.440 ;
        RECT 3376.930 1921.380 3377.250 1921.440 ;
        RECT 3368.190 1895.400 3368.510 1895.460 ;
        RECT 3376.930 1895.400 3377.250 1895.460 ;
        RECT 3368.190 1895.260 3377.250 1895.400 ;
        RECT 3368.190 1895.200 3368.510 1895.260 ;
        RECT 3376.930 1895.200 3377.250 1895.260 ;
        RECT 3368.190 1694.120 3368.510 1694.180 ;
        RECT 3376.930 1694.120 3377.250 1694.180 ;
        RECT 3368.190 1693.980 3377.250 1694.120 ;
        RECT 3368.190 1693.920 3368.510 1693.980 ;
        RECT 3376.930 1693.920 3377.250 1693.980 ;
        RECT 3369.110 1671.340 3369.430 1671.400 ;
        RECT 3376.930 1671.340 3377.250 1671.400 ;
        RECT 3369.110 1671.200 3377.250 1671.340 ;
        RECT 3369.110 1671.140 3369.430 1671.200 ;
        RECT 3376.930 1671.140 3377.250 1671.200 ;
        RECT 3369.110 1473.460 3369.430 1473.520 ;
        RECT 3376.470 1473.460 3376.790 1473.520 ;
        RECT 3369.110 1473.320 3376.790 1473.460 ;
        RECT 3369.110 1473.260 3369.430 1473.320 ;
        RECT 3376.470 1473.260 3376.790 1473.320 ;
        RECT 3368.190 1444.220 3368.510 1444.280 ;
        RECT 3376.930 1444.220 3377.250 1444.280 ;
        RECT 3368.190 1444.080 3377.250 1444.220 ;
        RECT 3368.190 1444.020 3368.510 1444.080 ;
        RECT 3376.930 1444.020 3377.250 1444.080 ;
        RECT 3368.190 1245.660 3368.510 1245.720 ;
        RECT 3376.930 1245.660 3377.250 1245.720 ;
        RECT 3368.190 1245.520 3377.250 1245.660 ;
        RECT 3368.190 1245.460 3368.510 1245.520 ;
        RECT 3376.930 1245.460 3377.250 1245.520 ;
        RECT 3369.110 1219.140 3369.430 1219.200 ;
        RECT 3376.930 1219.140 3377.250 1219.200 ;
        RECT 3369.110 1219.000 3377.250 1219.140 ;
        RECT 3369.110 1218.940 3369.430 1219.000 ;
        RECT 3376.930 1218.940 3377.250 1219.000 ;
        RECT 3369.110 1017.520 3369.430 1017.580 ;
        RECT 3376.470 1017.520 3376.790 1017.580 ;
        RECT 3369.110 1017.380 3376.790 1017.520 ;
        RECT 3369.110 1017.320 3369.430 1017.380 ;
        RECT 3376.470 1017.320 3376.790 1017.380 ;
        RECT 3368.650 995.420 3368.970 995.480 ;
        RECT 3376.930 995.420 3377.250 995.480 ;
        RECT 3368.650 995.280 3377.250 995.420 ;
        RECT 3368.650 995.220 3368.970 995.280 ;
        RECT 3376.930 995.220 3377.250 995.280 ;
        RECT 208.910 945.780 209.230 945.840 ;
        RECT 212.130 945.780 212.450 945.840 ;
        RECT 208.910 945.640 212.450 945.780 ;
        RECT 208.910 945.580 209.230 945.640 ;
        RECT 212.130 945.580 212.450 945.640 ;
        RECT 3368.650 793.120 3368.970 793.180 ;
        RECT 3376.930 793.120 3377.250 793.180 ;
        RECT 3368.650 792.980 3377.250 793.120 ;
        RECT 3368.650 792.920 3368.970 792.980 ;
        RECT 3376.930 792.920 3377.250 792.980 ;
        RECT 3368.190 770.680 3368.510 770.740 ;
        RECT 3376.470 770.680 3376.790 770.740 ;
        RECT 3368.190 770.540 3376.790 770.680 ;
        RECT 3368.190 770.480 3368.510 770.540 ;
        RECT 3376.470 770.480 3376.790 770.540 ;
        RECT 3368.190 568.720 3368.510 568.780 ;
        RECT 3376.930 568.720 3377.250 568.780 ;
        RECT 3368.190 568.580 3377.250 568.720 ;
        RECT 3368.190 568.520 3368.510 568.580 ;
        RECT 3376.930 568.520 3377.250 568.580 ;
        RECT 3368.190 542.200 3368.510 542.260 ;
        RECT 3376.930 542.200 3377.250 542.260 ;
        RECT 3368.190 542.060 3377.250 542.200 ;
        RECT 3368.190 542.000 3368.510 542.060 ;
        RECT 3376.930 542.000 3377.250 542.060 ;
        RECT 3368.190 234.840 3368.510 234.900 ;
        RECT 2637.340 234.700 3368.510 234.840 ;
        RECT 2637.340 234.560 2637.480 234.700 ;
        RECT 3368.190 234.640 3368.510 234.700 ;
        RECT 262.270 234.500 262.590 234.560 ;
        RECT 717.670 234.500 717.990 234.560 ;
        RECT 262.270 234.360 717.990 234.500 ;
        RECT 262.270 234.300 262.590 234.360 ;
        RECT 717.670 234.300 717.990 234.360 ;
        RECT 2637.250 234.300 2637.570 234.560 ;
        RECT 2341.470 221.920 2341.790 221.980 ;
        RECT 2363.090 221.920 2363.410 221.980 ;
        RECT 2089.480 221.780 2387.470 221.920 ;
        RECT 1793.610 221.580 1793.930 221.640 ;
        RECT 1815.230 221.580 1815.550 221.640 ;
        RECT 1749.540 221.440 1816.840 221.580 ;
        RECT 1519.450 221.240 1519.770 221.300 ;
        RECT 1541.070 221.240 1541.390 221.300 ;
        RECT 1749.540 221.240 1749.680 221.440 ;
        RECT 1793.610 221.380 1793.930 221.440 ;
        RECT 1815.230 221.380 1815.550 221.440 ;
        RECT 1034.930 221.100 1749.680 221.240 ;
        RECT 1816.700 221.240 1816.840 221.440 ;
        RECT 2089.480 221.300 2089.620 221.780 ;
        RECT 2341.470 221.720 2341.790 221.780 ;
        RECT 2363.090 221.720 2363.410 221.780 ;
        RECT 2387.330 221.580 2387.470 221.780 ;
        RECT 2387.330 221.440 2615.860 221.580 ;
        RECT 2067.770 221.240 2068.090 221.300 ;
        RECT 2089.390 221.240 2089.710 221.300 ;
        RECT 1816.700 221.100 2089.710 221.240 ;
        RECT 717.670 220.900 717.990 220.960 ;
        RECT 725.490 220.900 725.810 220.960 ;
        RECT 976.650 220.900 976.970 220.960 ;
        RECT 998.270 220.900 998.590 220.960 ;
        RECT 1034.930 220.900 1035.070 221.100 ;
        RECT 1519.450 221.040 1519.770 221.100 ;
        RECT 1541.070 221.040 1541.390 221.100 ;
        RECT 2067.770 221.040 2068.090 221.100 ;
        RECT 2089.390 221.040 2089.710 221.100 ;
        RECT 2615.720 220.960 2615.860 221.440 ;
        RECT 717.670 220.760 1035.070 220.900 ;
        RECT 2615.630 220.900 2615.950 220.960 ;
        RECT 2637.250 220.900 2637.570 220.960 ;
        RECT 2615.630 220.760 2637.570 220.900 ;
        RECT 717.670 220.700 717.990 220.760 ;
        RECT 725.490 220.700 725.810 220.760 ;
        RECT 976.650 220.700 976.970 220.760 ;
        RECT 998.270 220.700 998.590 220.760 ;
        RECT 2615.630 220.700 2615.950 220.760 ;
        RECT 2637.250 220.700 2637.570 220.760 ;
      LAYER via ;
        RECT 3368.680 4354.080 3368.940 4354.340 ;
        RECT 3376.960 4354.080 3377.220 4354.340 ;
        RECT 211.240 3936.220 211.500 3936.480 ;
        RECT 212.160 3936.220 212.420 3936.480 ;
        RECT 3368.680 3929.760 3368.940 3930.020 ;
        RECT 3376.040 3929.760 3376.300 3930.020 ;
        RECT 3376.960 3929.760 3377.220 3930.020 ;
        RECT 3368.680 3908.000 3368.940 3908.260 ;
        RECT 3376.040 3908.000 3376.300 3908.260 ;
        RECT 3376.960 3908.000 3377.220 3908.260 ;
        RECT 3368.680 3704.680 3368.940 3704.940 ;
        RECT 3376.040 3704.680 3376.300 3704.940 ;
        RECT 3376.960 3704.680 3377.220 3704.940 ;
        RECT 3368.680 3684.960 3368.940 3685.220 ;
        RECT 3376.040 3684.960 3376.300 3685.220 ;
        RECT 3376.960 3684.960 3377.220 3685.220 ;
        RECT 3368.680 3479.600 3368.940 3479.860 ;
        RECT 3376.040 3479.600 3376.300 3479.860 ;
        RECT 3376.960 3479.600 3377.220 3479.860 ;
        RECT 3368.680 3460.220 3368.940 3460.480 ;
        RECT 3376.040 3460.220 3376.300 3460.480 ;
        RECT 3376.960 3460.220 3377.220 3460.480 ;
        RECT 3368.680 3255.540 3368.940 3255.800 ;
        RECT 3376.960 3255.540 3377.220 3255.800 ;
        RECT 3368.680 3232.080 3368.940 3232.340 ;
        RECT 3376.960 3232.080 3377.220 3232.340 ;
        RECT 3368.680 3028.760 3368.940 3029.020 ;
        RECT 3376.040 3028.760 3376.300 3029.020 ;
        RECT 3376.960 3028.760 3377.220 3029.020 ;
        RECT 3368.680 3009.040 3368.940 3009.300 ;
        RECT 3376.040 3009.040 3376.300 3009.300 ;
        RECT 3376.960 3009.040 3377.220 3009.300 ;
        RECT 3368.680 2805.380 3368.940 2805.640 ;
        RECT 3376.040 2805.380 3376.300 2805.640 ;
        RECT 3368.220 2782.940 3368.480 2783.200 ;
        RECT 3376.040 2782.940 3376.300 2783.200 ;
        RECT 3376.960 2782.940 3377.220 2783.200 ;
        RECT 3368.220 1921.380 3368.480 1921.640 ;
        RECT 3376.960 1921.380 3377.220 1921.640 ;
        RECT 3368.220 1895.200 3368.480 1895.460 ;
        RECT 3376.960 1895.200 3377.220 1895.460 ;
        RECT 3368.220 1693.920 3368.480 1694.180 ;
        RECT 3376.960 1693.920 3377.220 1694.180 ;
        RECT 3369.140 1671.140 3369.400 1671.400 ;
        RECT 3376.960 1671.140 3377.220 1671.400 ;
        RECT 3369.140 1473.260 3369.400 1473.520 ;
        RECT 3376.500 1473.260 3376.760 1473.520 ;
        RECT 3368.220 1444.020 3368.480 1444.280 ;
        RECT 3376.960 1444.020 3377.220 1444.280 ;
        RECT 3368.220 1245.460 3368.480 1245.720 ;
        RECT 3376.960 1245.460 3377.220 1245.720 ;
        RECT 3369.140 1218.940 3369.400 1219.200 ;
        RECT 3376.960 1218.940 3377.220 1219.200 ;
        RECT 3369.140 1017.320 3369.400 1017.580 ;
        RECT 3376.500 1017.320 3376.760 1017.580 ;
        RECT 3368.680 995.220 3368.940 995.480 ;
        RECT 3376.960 995.220 3377.220 995.480 ;
        RECT 208.940 945.580 209.200 945.840 ;
        RECT 212.160 945.580 212.420 945.840 ;
        RECT 3368.680 792.920 3368.940 793.180 ;
        RECT 3376.960 792.920 3377.220 793.180 ;
        RECT 3368.220 770.480 3368.480 770.740 ;
        RECT 3376.500 770.480 3376.760 770.740 ;
        RECT 3368.220 568.520 3368.480 568.780 ;
        RECT 3376.960 568.520 3377.220 568.780 ;
        RECT 3368.220 542.000 3368.480 542.260 ;
        RECT 3376.960 542.000 3377.220 542.260 ;
        RECT 3368.220 234.640 3368.480 234.900 ;
        RECT 262.300 234.300 262.560 234.560 ;
        RECT 717.700 234.300 717.960 234.560 ;
        RECT 2637.280 234.300 2637.540 234.560 ;
        RECT 717.700 220.700 717.960 220.960 ;
        RECT 725.520 220.700 725.780 220.960 ;
        RECT 976.680 220.700 976.940 220.960 ;
        RECT 998.300 220.700 998.560 220.960 ;
        RECT 1519.480 221.040 1519.740 221.300 ;
        RECT 1541.100 221.040 1541.360 221.300 ;
        RECT 1793.640 221.380 1793.900 221.640 ;
        RECT 1815.260 221.380 1815.520 221.640 ;
        RECT 2341.500 221.720 2341.760 221.980 ;
        RECT 2363.120 221.720 2363.380 221.980 ;
        RECT 2067.800 221.040 2068.060 221.300 ;
        RECT 2089.420 221.040 2089.680 221.300 ;
        RECT 2615.660 220.700 2615.920 220.960 ;
        RECT 2637.280 220.700 2637.540 220.960 ;
      LAYER met2 ;
        RECT 3377.035 4378.485 3379.435 4378.555 ;
        RECT 3376.560 4378.345 3379.435 4378.485 ;
        RECT 3376.560 4356.865 3376.700 4378.345 ;
        RECT 3377.035 4378.275 3379.435 4378.345 ;
        RECT 3377.035 4356.865 3379.435 4356.935 ;
        RECT 3376.560 4356.725 3379.435 4356.865 ;
        RECT 3377.020 4356.655 3379.435 4356.725 ;
        RECT 3377.020 4354.370 3377.160 4356.655 ;
        RECT 3368.680 4354.050 3368.940 4354.370 ;
        RECT 3376.960 4354.050 3377.220 4354.370 ;
        RECT 208.565 3957.330 210.965 3957.345 ;
        RECT 208.565 3957.190 211.440 3957.330 ;
        RECT 208.565 3957.065 210.965 3957.190 ;
        RECT 211.300 3936.510 211.440 3957.190 ;
        RECT 211.240 3936.250 211.500 3936.510 ;
        RECT 209.460 3936.190 211.500 3936.250 ;
        RECT 212.160 3936.190 212.420 3936.510 ;
        RECT 209.460 3936.110 211.440 3936.190 ;
        RECT 209.460 3935.725 209.600 3936.110 ;
        RECT 208.565 3935.445 210.965 3935.725 ;
        RECT 208.610 3935.430 209.600 3935.445 ;
        RECT 208.565 3741.065 210.965 3741.345 ;
        RECT 209.460 3739.870 209.600 3741.065 ;
        RECT 212.220 3739.870 212.360 3936.190 ;
        RECT 3368.740 3930.050 3368.880 4354.050 ;
        RECT 3377.035 3932.415 3379.435 3932.555 ;
        RECT 3377.020 3932.275 3379.435 3932.415 ;
        RECT 3377.020 3930.050 3377.160 3932.275 ;
        RECT 3368.680 3929.730 3368.940 3930.050 ;
        RECT 3376.040 3929.730 3376.300 3930.050 ;
        RECT 3376.960 3929.730 3377.220 3930.050 ;
        RECT 3376.100 3908.290 3376.240 3929.730 ;
        RECT 3377.035 3910.795 3379.435 3910.935 ;
        RECT 3377.020 3910.655 3379.435 3910.795 ;
        RECT 3377.020 3908.290 3377.160 3910.655 ;
        RECT 3368.680 3907.970 3368.940 3908.290 ;
        RECT 3376.040 3907.970 3376.300 3908.290 ;
        RECT 3376.960 3907.970 3377.220 3908.290 ;
        RECT 209.460 3739.730 212.360 3739.870 ;
        RECT 208.565 3719.445 210.965 3719.725 ;
        RECT 209.000 3718.650 209.140 3719.445 ;
        RECT 211.300 3718.650 211.440 3739.730 ;
        RECT 209.000 3718.510 211.440 3718.650 ;
        RECT 211.300 3643.270 211.440 3718.510 ;
        RECT 3368.740 3704.970 3368.880 3907.970 ;
        RECT 3377.035 3707.415 3379.435 3707.555 ;
        RECT 3377.020 3707.275 3379.435 3707.415 ;
        RECT 3377.020 3704.970 3377.160 3707.275 ;
        RECT 3368.680 3704.650 3368.940 3704.970 ;
        RECT 3376.040 3704.650 3376.300 3704.970 ;
        RECT 3376.960 3704.650 3377.220 3704.970 ;
        RECT 3376.100 3685.250 3376.240 3704.650 ;
        RECT 3377.035 3685.795 3379.435 3685.935 ;
        RECT 3377.020 3685.655 3379.435 3685.795 ;
        RECT 3377.020 3685.250 3377.160 3685.655 ;
        RECT 3368.680 3684.930 3368.940 3685.250 ;
        RECT 3376.040 3684.930 3376.300 3685.250 ;
        RECT 3376.960 3684.930 3377.220 3685.250 ;
        RECT 211.300 3643.130 211.900 3643.270 ;
        RECT 208.565 3525.065 210.965 3525.345 ;
        RECT 209.460 3524.850 209.600 3525.065 ;
        RECT 211.760 3524.850 211.900 3643.130 ;
        RECT 209.460 3524.710 211.900 3524.850 ;
        RECT 208.610 3503.725 209.600 3503.770 ;
        RECT 208.565 3503.445 210.965 3503.725 ;
        RECT 209.460 3503.090 209.600 3503.445 ;
        RECT 211.300 3503.090 211.440 3524.710 ;
        RECT 209.460 3502.950 211.440 3503.090 ;
        RECT 211.300 3450.070 211.440 3502.950 ;
        RECT 3368.740 3479.890 3368.880 3684.930 ;
        RECT 3377.035 3482.415 3379.435 3482.555 ;
        RECT 3377.020 3482.275 3379.435 3482.415 ;
        RECT 3377.020 3479.890 3377.160 3482.275 ;
        RECT 3368.680 3479.570 3368.940 3479.890 ;
        RECT 3376.040 3479.570 3376.300 3479.890 ;
        RECT 3376.960 3479.570 3377.220 3479.890 ;
        RECT 3376.100 3460.510 3376.240 3479.570 ;
        RECT 3377.035 3460.860 3379.435 3460.935 ;
        RECT 3377.020 3460.655 3379.435 3460.860 ;
        RECT 3377.020 3460.510 3377.160 3460.655 ;
        RECT 3368.680 3460.190 3368.940 3460.510 ;
        RECT 3376.040 3460.190 3376.300 3460.510 ;
        RECT 3376.960 3460.190 3377.220 3460.510 ;
        RECT 211.300 3449.930 211.900 3450.070 ;
        RECT 211.760 3309.970 211.900 3449.930 ;
        RECT 209.000 3309.830 211.900 3309.970 ;
        RECT 209.000 3309.345 209.140 3309.830 ;
        RECT 208.565 3309.065 210.965 3309.345 ;
        RECT 211.300 3288.210 211.440 3309.830 ;
        RECT 209.460 3288.070 211.440 3288.210 ;
        RECT 209.460 3287.725 209.600 3288.070 ;
        RECT 208.565 3287.445 210.965 3287.725 ;
        RECT 208.610 3287.390 209.600 3287.445 ;
        RECT 211.300 3256.870 211.440 3288.070 ;
        RECT 211.300 3256.730 211.900 3256.870 ;
        RECT 211.760 3093.730 211.900 3256.730 ;
        RECT 3368.740 3255.830 3368.880 3460.190 ;
        RECT 3377.035 3256.415 3379.435 3256.555 ;
        RECT 3377.020 3256.275 3379.435 3256.415 ;
        RECT 3377.020 3255.830 3377.160 3256.275 ;
        RECT 3368.680 3255.510 3368.940 3255.830 ;
        RECT 3376.960 3255.510 3377.220 3255.830 ;
        RECT 3368.740 3232.370 3368.880 3255.510 ;
        RECT 3377.035 3234.795 3379.435 3234.935 ;
        RECT 3377.020 3234.655 3379.435 3234.795 ;
        RECT 3377.020 3232.370 3377.160 3234.655 ;
        RECT 3368.680 3232.050 3368.940 3232.370 ;
        RECT 3376.960 3232.050 3377.220 3232.370 ;
        RECT 209.000 3093.590 211.900 3093.730 ;
        RECT 209.000 3093.345 209.140 3093.590 ;
        RECT 208.565 3093.065 210.965 3093.345 ;
        RECT 208.565 3071.655 210.965 3071.725 ;
        RECT 211.300 3071.655 211.440 3093.590 ;
        RECT 208.565 3071.515 211.440 3071.655 ;
        RECT 208.565 3071.445 210.965 3071.515 ;
        RECT 211.300 3063.670 211.440 3071.515 ;
        RECT 211.300 3063.530 211.900 3063.670 ;
        RECT 208.565 2877.275 210.965 2877.345 ;
        RECT 211.760 2877.275 211.900 3063.530 ;
        RECT 3368.740 3029.050 3368.880 3232.050 ;
        RECT 3377.035 3031.415 3379.435 3031.555 ;
        RECT 3377.020 3031.275 3379.435 3031.415 ;
        RECT 3377.020 3029.050 3377.160 3031.275 ;
        RECT 3368.680 3028.730 3368.940 3029.050 ;
        RECT 3376.040 3028.730 3376.300 3029.050 ;
        RECT 3376.960 3028.730 3377.220 3029.050 ;
        RECT 3376.100 3009.330 3376.240 3028.730 ;
        RECT 3377.035 3009.795 3379.435 3009.935 ;
        RECT 3377.020 3009.655 3379.435 3009.795 ;
        RECT 3377.020 3009.330 3377.160 3009.655 ;
        RECT 3368.680 3009.010 3368.940 3009.330 ;
        RECT 3376.040 3009.010 3376.300 3009.330 ;
        RECT 3376.960 3009.010 3377.220 3009.330 ;
        RECT 208.565 2877.135 211.900 2877.275 ;
        RECT 208.565 2877.065 210.965 2877.135 ;
        RECT 211.300 2856.410 211.440 2877.135 ;
        RECT 209.000 2856.270 211.900 2856.410 ;
        RECT 209.000 2855.730 209.140 2856.270 ;
        RECT 208.610 2855.725 209.140 2855.730 ;
        RECT 208.565 2855.445 210.965 2855.725 ;
        RECT 208.565 2661.065 210.965 2661.345 ;
        RECT 209.460 2660.570 209.600 2661.065 ;
        RECT 211.760 2660.570 211.900 2856.270 ;
        RECT 3368.740 2805.670 3368.880 3009.010 ;
        RECT 3376.100 2805.670 3376.240 2805.825 ;
        RECT 3368.680 2805.350 3368.940 2805.670 ;
        RECT 3376.040 2805.410 3376.300 2805.670 ;
        RECT 3377.035 2805.410 3379.435 2805.555 ;
        RECT 3376.040 2805.350 3379.435 2805.410 ;
        RECT 3376.100 2805.275 3379.435 2805.350 ;
        RECT 3376.100 2805.270 3377.090 2805.275 ;
        RECT 3376.100 2783.230 3376.240 2805.270 ;
        RECT 3377.035 2783.795 3379.435 2783.935 ;
        RECT 3377.020 2783.655 3379.435 2783.795 ;
        RECT 3377.020 2783.230 3377.160 2783.655 ;
        RECT 3368.220 2782.910 3368.480 2783.230 ;
        RECT 3376.040 2782.910 3376.300 2783.230 ;
        RECT 3376.960 2782.910 3377.220 2783.230 ;
        RECT 209.460 2660.430 211.900 2660.570 ;
        RECT 208.565 2639.585 210.965 2639.725 ;
        RECT 208.540 2639.490 210.965 2639.585 ;
        RECT 211.300 2639.490 211.440 2660.430 ;
        RECT 208.540 2639.350 211.440 2639.490 ;
        RECT 211.300 2097.670 211.440 2639.350 ;
        RECT 211.300 2097.530 211.900 2097.670 ;
        RECT 211.760 2026.130 211.900 2097.530 ;
        RECT 209.000 2025.990 211.900 2026.130 ;
        RECT 209.000 2023.410 209.140 2025.990 ;
        RECT 208.610 2023.345 209.140 2023.410 ;
        RECT 208.565 2023.065 210.965 2023.345 ;
        RECT 208.565 2001.650 210.965 2001.725 ;
        RECT 211.300 2001.650 211.440 2025.990 ;
        RECT 208.565 2001.510 211.440 2001.650 ;
        RECT 208.565 2001.445 210.965 2001.510 ;
        RECT 208.565 1807.170 210.965 1807.345 ;
        RECT 211.300 1807.170 211.440 2001.510 ;
        RECT 3368.280 1921.670 3368.420 2782.910 ;
        RECT 3368.220 1921.350 3368.480 1921.670 ;
        RECT 3376.960 1921.350 3377.220 1921.670 ;
        RECT 3377.020 1920.050 3377.160 1921.350 ;
        RECT 3376.560 1919.910 3377.160 1920.050 ;
        RECT 3376.560 1897.865 3376.700 1919.910 ;
        RECT 3377.020 1919.555 3377.160 1919.910 ;
        RECT 3377.020 1919.300 3379.435 1919.555 ;
        RECT 3377.035 1919.275 3379.435 1919.300 ;
        RECT 3377.035 1897.865 3379.435 1897.935 ;
        RECT 3376.560 1897.725 3379.435 1897.865 ;
        RECT 3377.020 1897.655 3379.435 1897.725 ;
        RECT 3377.020 1895.490 3377.160 1897.655 ;
        RECT 3368.220 1895.170 3368.480 1895.490 ;
        RECT 3376.960 1895.170 3377.220 1895.490 ;
        RECT 208.565 1807.065 211.440 1807.170 ;
        RECT 208.610 1807.030 211.440 1807.065 ;
        RECT 208.565 1785.445 210.965 1785.725 ;
        RECT 209.920 1783.370 210.060 1785.445 ;
        RECT 211.300 1783.370 211.440 1807.030 ;
        RECT 209.920 1783.230 211.440 1783.370 ;
        RECT 211.300 1663.010 211.440 1783.230 ;
        RECT 3368.280 1694.210 3368.420 1895.170 ;
        RECT 3368.220 1693.890 3368.480 1694.210 ;
        RECT 3376.960 1693.890 3377.220 1694.210 ;
        RECT 3377.020 1693.555 3377.160 1693.890 ;
        RECT 3377.020 1693.275 3379.435 1693.555 ;
        RECT 3377.020 1690.890 3377.160 1693.275 ;
        RECT 3376.560 1690.750 3377.160 1690.890 ;
        RECT 3376.560 1671.850 3376.700 1690.750 ;
        RECT 3377.035 1671.850 3379.435 1671.935 ;
        RECT 3376.560 1671.710 3379.435 1671.850 ;
        RECT 3377.020 1671.655 3379.435 1671.710 ;
        RECT 3377.020 1671.430 3377.160 1671.655 ;
        RECT 3369.140 1671.110 3369.400 1671.430 ;
        RECT 3376.960 1671.110 3377.220 1671.430 ;
        RECT 211.300 1662.870 211.900 1663.010 ;
        RECT 208.565 1591.275 210.965 1591.345 ;
        RECT 211.760 1591.275 211.900 1662.870 ;
        RECT 208.565 1591.135 211.900 1591.275 ;
        RECT 208.565 1591.065 210.965 1591.135 ;
        RECT 208.565 1569.445 210.965 1569.725 ;
        RECT 209.000 1569.170 209.140 1569.445 ;
        RECT 211.300 1569.170 211.440 1591.135 ;
        RECT 209.000 1569.030 211.440 1569.170 ;
        RECT 211.300 1518.070 211.440 1569.030 ;
        RECT 211.300 1517.930 211.900 1518.070 ;
        RECT 211.760 1376.050 211.900 1517.930 ;
        RECT 3369.200 1473.550 3369.340 1671.110 ;
        RECT 3369.140 1473.230 3369.400 1473.550 ;
        RECT 3376.500 1473.230 3376.760 1473.550 ;
        RECT 3376.560 1468.530 3376.700 1473.230 ;
        RECT 3377.035 1468.530 3379.435 1468.555 ;
        RECT 3376.560 1468.390 3379.435 1468.530 ;
        RECT 3376.560 1446.770 3376.700 1468.390 ;
        RECT 3377.035 1468.275 3379.435 1468.390 ;
        RECT 3377.035 1446.770 3379.435 1446.935 ;
        RECT 3376.560 1446.655 3379.435 1446.770 ;
        RECT 3376.560 1446.630 3377.160 1446.655 ;
        RECT 3377.020 1444.310 3377.160 1446.630 ;
        RECT 3368.220 1443.990 3368.480 1444.310 ;
        RECT 3376.960 1443.990 3377.220 1444.310 ;
        RECT 209.000 1375.910 211.900 1376.050 ;
        RECT 209.000 1375.370 209.140 1375.910 ;
        RECT 208.610 1375.345 209.140 1375.370 ;
        RECT 208.565 1375.065 210.965 1375.345 ;
        RECT 211.300 1354.290 211.440 1375.910 ;
        RECT 209.460 1354.150 211.440 1354.290 ;
        RECT 209.460 1353.725 209.600 1354.150 ;
        RECT 208.565 1353.445 210.965 1353.725 ;
        RECT 211.300 1324.870 211.440 1354.150 ;
        RECT 211.300 1324.730 211.900 1324.870 ;
        RECT 208.565 1159.275 210.965 1159.345 ;
        RECT 211.760 1159.275 211.900 1324.730 ;
        RECT 3368.280 1245.750 3368.420 1443.990 ;
        RECT 3368.220 1245.430 3368.480 1245.750 ;
        RECT 3376.960 1245.430 3377.220 1245.750 ;
        RECT 3377.020 1243.555 3377.160 1245.430 ;
        RECT 3377.020 1243.450 3379.435 1243.555 ;
        RECT 3376.560 1243.310 3379.435 1243.450 ;
        RECT 3376.560 1221.865 3376.700 1243.310 ;
        RECT 3377.035 1243.275 3379.435 1243.310 ;
        RECT 3377.035 1221.865 3379.435 1221.935 ;
        RECT 3376.560 1221.725 3379.435 1221.865 ;
        RECT 3377.020 1221.655 3379.435 1221.725 ;
        RECT 3377.020 1219.230 3377.160 1221.655 ;
        RECT 3369.140 1218.910 3369.400 1219.230 ;
        RECT 3376.960 1218.910 3377.220 1219.230 ;
        RECT 208.565 1159.135 211.900 1159.275 ;
        RECT 208.565 1159.065 210.965 1159.135 ;
        RECT 211.300 1138.050 211.440 1159.135 ;
        RECT 209.000 1137.910 211.900 1138.050 ;
        RECT 209.000 1137.725 209.140 1137.910 ;
        RECT 208.565 1137.445 210.965 1137.725 ;
        RECT 211.760 987.770 211.900 1137.910 ;
        RECT 3369.200 1017.610 3369.340 1218.910 ;
        RECT 3376.560 1017.610 3376.700 1017.900 ;
        RECT 3369.140 1017.290 3369.400 1017.610 ;
        RECT 3376.500 1017.485 3376.760 1017.610 ;
        RECT 3377.035 1017.485 3379.435 1017.555 ;
        RECT 3376.500 1017.345 3379.435 1017.485 ;
        RECT 3376.500 1017.290 3376.760 1017.345 ;
        RECT 3376.560 995.930 3376.700 1017.290 ;
        RECT 3377.035 1017.275 3379.435 1017.345 ;
        RECT 3377.035 995.930 3379.435 995.935 ;
        RECT 3376.560 995.790 3379.435 995.930 ;
        RECT 3377.020 995.655 3379.435 995.790 ;
        RECT 3377.020 995.510 3377.160 995.655 ;
        RECT 3368.680 995.190 3368.940 995.510 ;
        RECT 3376.960 995.190 3377.220 995.510 ;
        RECT 211.760 987.630 212.360 987.770 ;
        RECT 212.220 945.870 212.360 987.630 ;
        RECT 208.940 945.550 209.200 945.870 ;
        RECT 212.160 945.550 212.420 945.870 ;
        RECT 209.000 943.345 209.140 945.550 ;
        RECT 208.565 943.065 210.965 943.345 ;
        RECT 212.220 940.170 212.360 945.550 ;
        RECT 211.300 940.030 212.360 940.170 ;
        RECT 208.565 921.655 210.965 921.725 ;
        RECT 211.300 921.655 211.440 940.030 ;
        RECT 208.565 921.515 211.900 921.655 ;
        RECT 208.565 921.445 210.965 921.515 ;
        RECT 211.760 235.125 211.900 921.515 ;
        RECT 3368.740 793.210 3368.880 995.190 ;
        RECT 3368.680 792.890 3368.940 793.210 ;
        RECT 3376.960 792.890 3377.220 793.210 ;
        RECT 3377.020 792.610 3377.160 792.890 ;
        RECT 3376.560 792.555 3377.160 792.610 ;
        RECT 3376.560 792.470 3379.435 792.555 ;
        RECT 3376.560 770.850 3376.700 792.470 ;
        RECT 3377.035 792.275 3379.435 792.470 ;
        RECT 3377.035 770.850 3379.435 770.935 ;
        RECT 3376.560 770.770 3379.435 770.850 ;
        RECT 3368.220 770.450 3368.480 770.770 ;
        RECT 3376.500 770.710 3379.435 770.770 ;
        RECT 3376.500 770.450 3376.760 770.710 ;
        RECT 3377.035 770.655 3379.435 770.710 ;
        RECT 3368.280 568.810 3368.420 770.450 ;
        RECT 3376.560 770.295 3376.700 770.450 ;
        RECT 3368.220 568.490 3368.480 568.810 ;
        RECT 3376.960 568.490 3377.220 568.810 ;
        RECT 3377.020 566.555 3377.160 568.490 ;
        RECT 3377.020 566.485 3379.435 566.555 ;
        RECT 3376.560 566.345 3379.435 566.485 ;
        RECT 3376.560 544.865 3376.700 566.345 ;
        RECT 3377.035 566.275 3379.435 566.345 ;
        RECT 3377.035 544.865 3379.435 544.935 ;
        RECT 3376.560 544.725 3379.435 544.865 ;
        RECT 3377.020 544.655 3379.435 544.725 ;
        RECT 3377.020 542.290 3377.160 544.655 ;
        RECT 3368.220 541.970 3368.480 542.290 ;
        RECT 3376.960 541.970 3377.220 542.290 ;
        RECT 211.690 234.755 211.970 235.125 ;
        RECT 3368.280 234.930 3368.420 541.970 ;
        RECT 3368.220 234.610 3368.480 234.930 ;
        RECT 262.300 234.445 262.560 234.590 ;
        RECT 262.290 234.075 262.570 234.445 ;
        RECT 717.700 234.270 717.960 234.590 ;
        RECT 2637.280 234.270 2637.540 234.590 ;
        RECT 717.760 220.990 717.900 234.270 ;
        RECT 2341.500 221.690 2341.760 222.010 ;
        RECT 2363.120 221.690 2363.380 222.010 ;
        RECT 1793.640 221.350 1793.900 221.670 ;
        RECT 1815.260 221.350 1815.520 221.670 ;
        RECT 1519.480 221.010 1519.740 221.330 ;
        RECT 1541.100 221.010 1541.360 221.330 ;
        RECT 717.700 220.670 717.960 220.990 ;
        RECT 725.520 220.670 725.780 220.990 ;
        RECT 976.680 220.670 976.940 220.990 ;
        RECT 998.300 220.670 998.560 220.990 ;
        RECT 725.580 201.010 725.720 220.670 ;
        RECT 976.740 210.965 976.880 220.670 ;
        RECT 998.360 210.965 998.500 220.670 ;
        RECT 1519.540 210.965 1519.680 221.010 ;
        RECT 1541.160 210.965 1541.300 221.010 ;
        RECT 1793.700 210.965 1793.840 221.350 ;
        RECT 1815.320 210.965 1815.460 221.350 ;
        RECT 2067.800 221.010 2068.060 221.330 ;
        RECT 2089.420 221.010 2089.680 221.330 ;
        RECT 2067.860 210.965 2068.000 221.010 ;
        RECT 2089.480 210.965 2089.620 221.010 ;
        RECT 976.655 208.565 976.935 210.965 ;
        RECT 998.275 208.565 998.555 210.965 ;
        RECT 1519.540 209.030 1519.935 210.965 ;
        RECT 1541.160 209.030 1541.555 210.965 ;
        RECT 1519.655 208.565 1519.935 209.030 ;
        RECT 1541.275 208.565 1541.555 209.030 ;
        RECT 1793.655 208.565 1793.935 210.965 ;
        RECT 1815.275 208.565 1815.555 210.965 ;
        RECT 2067.655 209.100 2068.000 210.965 ;
        RECT 2089.275 209.100 2089.620 210.965 ;
        RECT 2341.560 210.965 2341.700 221.690 ;
        RECT 2363.180 210.965 2363.320 221.690 ;
        RECT 2637.340 220.990 2637.480 234.270 ;
        RECT 2615.660 220.670 2615.920 220.990 ;
        RECT 2637.280 220.670 2637.540 220.990 ;
        RECT 2615.720 210.965 2615.860 220.670 ;
        RECT 2637.340 210.965 2637.480 220.670 ;
        RECT 2067.655 208.565 2067.935 209.100 ;
        RECT 2089.275 208.565 2089.555 209.100 ;
        RECT 2341.560 209.030 2341.935 210.965 ;
        RECT 2363.180 209.030 2363.555 210.965 ;
        RECT 2341.655 208.565 2341.935 209.030 ;
        RECT 2363.275 208.565 2363.555 209.030 ;
        RECT 2615.655 208.565 2615.935 210.965 ;
        RECT 2637.275 208.565 2637.555 210.965 ;
        RECT 725.515 200.870 725.720 201.010 ;
        RECT 725.515 200.000 725.655 200.870 ;
        RECT 725.455 198.530 725.715 200.000 ;
      LAYER via2 ;
        RECT 211.690 234.800 211.970 235.080 ;
        RECT 262.290 234.120 262.570 234.400 ;
      LAYER met3 ;
        RECT 211.665 235.090 211.995 235.105 ;
        RECT 211.665 234.790 224.170 235.090 ;
        RECT 211.665 234.775 211.995 234.790 ;
        RECT 223.870 234.410 224.170 234.790 ;
        RECT 262.265 234.410 262.595 234.425 ;
        RECT 223.870 234.110 262.595 234.410 ;
        RECT 262.265 234.095 262.595 234.110 ;
    END
  END porb_h
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 683.565 35.715 720.750 91.545 ;
    END
  END resetb
  PIN resetb_core_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 708.335 190.155 709.065 200.000 ;
        RECT 708.335 189.855 709.365 190.155 ;
        RECT 708.335 189.555 709.100 189.855 ;
        RECT 709.365 189.555 709.830 189.855 ;
        RECT 708.335 189.090 709.830 189.555 ;
        RECT 709.100 185.230 709.830 189.090 ;
    END
  END resetb_core_h
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 468.035 181.615 663.965 185.065 ;
    END
  END vdda
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 143.265 964.910 143.595 ;
    END
  END vssa
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 158.370 664.270 158.415 ;
        RECT 467.730 153.810 664.345 158.370 ;
        RECT 467.730 153.765 664.270 153.810 ;
    END
  END vssd
  PIN mprj_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3154.720 4988.000 3179.720 5070.350 ;
    END
  END mprj_analog[1]
  PIN mprj_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3137.050 5093.120 3197.890 5153.945 ;
    END
  END mprj_io[15]
  PIN mprj_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2645.720 4988.000 2670.720 5070.350 ;
    END
  END mprj_analog[2]
  PIN mprj_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2628.050 5093.120 2688.890 5153.945 ;
    END
  END mprj_io[16]
  PIN mprj_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2388.720 4988.000 2413.720 5070.350 ;
    END
  END mprj_analog[3]
  PIN mprj_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2371.050 5093.120 2431.890 5153.945 ;
    END
  END mprj_io[17]
  PIN mprj_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1943.720 4988.000 1968.720 5070.350 ;
    END
  END mprj_analog[4]
  PIN mprj_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1926.050 5093.120 1986.890 5153.945 ;
    END
  END mprj_io[18]
  PIN mprj_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3388.000 4716.000 3403.685 4787.610 ;
    END
  END mprj_analog[0]
  PIN mprj_clamp_high[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3388.000 4763.710 3413.660 4787.610 ;
    END
  END mprj_clamp_high[0]
  PIN mprj_clamp_low[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3388.000 4813.605 3390.055 4837.505 ;
    END
  END mprj_clamp_low[0]
  PIN mprj_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4770.110 3553.945 4830.950 ;
    END
  END mprj_io[14]
  PIN vccd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 4548.330 3557.165 4602.730 ;
    END
  END vccd1_pad
  PIN vdda1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4099.110 3553.945 4159.950 ;
    END
  END vdda1_pad
  PIN vdda1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2526.110 3553.945 2586.950 ;
    END
  END vdda1_pad2
  PIN vssa1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2885.050 5093.120 2945.890 5153.945 ;
    END
  END vssa1_pad
  PIN vssa1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2085.110 3553.945 2145.950 ;
    END
  END vssa1_pad2
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3396.885 2151.730 3401.535 2300.270 ;
    END
  END vccd1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3402.935 2152.035 3406.385 2299.965 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3444.405 2151.730 3444.735 2771.910 ;
    END
  END vssa1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3390.000 2349.500 3429.600 2373.500 ;
    END
  END vssd1
  PIN vssd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 2309.330 3557.165 2363.730 ;
    END
  END vssd1_pad
  PIN mprj_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 919.720 4988.000 944.720 5070.350 ;
    END
  END mprj_analog[7]
  PIN mprj_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 902.050 5093.120 962.890 5153.945 ;
    END
  END mprj_io[21]
  PIN mprj_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 662.720 4988.000 687.720 5070.350 ;
    END
  END mprj_analog[8]
  PIN mprj_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 645.050 5093.120 705.890 5153.945 ;
    END
  END mprj_io[22]
  PIN mprj_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 405.720 4988.000 430.720 5070.350 ;
    END
  END mprj_analog[9]
  PIN mprj_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 388.050 5093.120 448.890 5153.945 ;
    END
  END mprj_io[23]
  PIN mprj_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.650 4795.720 200.000 4820.720 ;
    END
  END mprj_analog[10]
  PIN mprj_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4778.050 94.880 4838.890 ;
    END
  END mprj_io[24]
  PIN mprj_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1460.390 4988.000 1532.000 5003.685 ;
    END
  END mprj_analog[5]
  PIN mprj_clamp_high[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.390 4988.000 1484.290 5013.660 ;
    END
  END mprj_clamp_high[1]
  PIN mprj_clamp_low[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.495 4988.000 1434.395 4990.055 ;
    END
  END mprj_clamp_low[1]
  PIN mprj_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1417.050 5093.120 1477.890 5153.945 ;
    END
  END mprj_io[19]
  PIN mprj_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1202.390 4988.000 1274.000 5003.685 ;
    END
  END mprj_analog[6]
  PIN mprj_clamp_high[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 4988.000 1226.290 5013.660 ;
    END
  END mprj_clamp_high[2]
  PIN mprj_clamp_low[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.495 4988.000 1176.395 4990.055 ;
    END
  END mprj_clamp_low[2]
  PIN mprj_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1159.050 5093.120 1219.890 5153.945 ;
    END
  END mprj_io[20]
  PIN vccd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 4570.270 98.100 4624.670 ;
    END
  END vccd2_pad
  PIN vdda2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 2422.050 94.880 2482.890 ;
    END
  END vdda2_pad
  PIN vssa2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4145.050 94.880 4205.890 ;
    END
  END vssa2_pad
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 192.515 2277.730 197.965 2416.270 ;
    END
  END vccd
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 186.465 2277.730 191.115 2416.270 ;
    END
  END vccd2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 181.615 2278.035 185.065 2415.965 ;
    END
  END vdda2
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 164.665 2277.730 168.115 2416.270 ;
    END
  END vddio
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.265 2035.090 143.595 2628.610 ;
    END
  END vssa2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.400 2204.500 198.000 2228.500 ;
    END
  END vssd2
  PIN vssd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 2214.270 98.100 2268.670 ;
    END
  END vssd2_pad
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.035 2279.000 24.215 2280.465 ;
        RECT 0.000 2277.730 24.215 2279.000 ;
    END
  END vssio
  OBS
      LAYER pwell ;
        RECT 1155.495 4988.935 1163.285 5011.790 ;
      LAYER nwell ;
        RECT 1163.860 4988.685 1222.965 4990.205 ;
      LAYER pwell ;
        RECT 1413.495 4988.935 1421.285 5011.790 ;
      LAYER nwell ;
        RECT 1421.860 4988.685 1480.965 4990.205 ;
        RECT 1678.860 4988.685 1737.965 4990.205 ;
        RECT 2889.860 4988.685 2948.965 4990.205 ;
      LAYER pwell ;
        RECT 3388.935 4826.715 3411.790 4834.505 ;
      LAYER nwell ;
        RECT 3388.685 4767.035 3390.205 4826.140 ;
        RECT 197.795 4360.860 199.315 4419.965 ;
        RECT 3393.665 4388.890 3397.325 4392.415 ;
        RECT 3444.590 4391.285 3469.235 4392.715 ;
        RECT 3476.485 4392.120 3480.400 4392.415 ;
      LAYER pwell ;
        RECT 176.210 4352.495 199.065 4360.285 ;
      LAYER nwell ;
        RECT 3407.155 4327.170 3411.080 4387.420 ;
        RECT 3444.590 4368.485 3446.020 4391.285 ;
        RECT 3448.180 4388.190 3450.340 4391.285 ;
        RECT 3448.180 4381.540 3449.020 4388.190 ;
        RECT 3448.770 4378.465 3449.020 4381.540 ;
        RECT 3467.805 4367.185 3469.235 4391.285 ;
        RECT 3473.580 4389.205 3480.400 4392.120 ;
        RECT 3473.580 4387.470 3479.820 4389.205 ;
        RECT 3474.660 4386.025 3479.820 4387.470 ;
      LAYER pwell ;
        RECT 3480.935 4386.785 3518.355 4392.215 ;
      LAYER nwell ;
        RECT 3474.660 4383.580 3476.280 4386.025 ;
        RECT 3474.660 4383.505 3475.740 4383.580 ;
      LAYER pwell ;
        RECT 3480.935 4382.700 3484.255 4386.785 ;
        RECT 3482.955 4352.615 3484.255 4382.700 ;
        RECT 3489.965 4386.265 3518.355 4386.785 ;
        RECT 3489.965 4352.615 3491.550 4386.265 ;
        RECT 3482.955 4346.160 3485.985 4352.615 ;
        RECT 3482.955 4345.410 3483.260 4346.160 ;
      LAYER nwell ;
        RECT 3422.265 4333.725 3424.055 4343.085 ;
        RECT 3420.410 4327.170 3424.055 4333.725 ;
        RECT 3407.155 4311.550 3413.345 4327.170 ;
        RECT 3417.785 4311.550 3424.055 4327.170 ;
        RECT 3460.595 4329.350 3461.265 4345.060 ;
        RECT 3438.620 4312.875 3440.050 4321.665 ;
        RECT 3453.195 4312.875 3454.045 4321.665 ;
        RECT 3460.595 4312.875 3461.775 4329.350 ;
        RECT 3438.620 4312.760 3461.775 4312.875 ;
        RECT 3471.165 4312.760 3472.345 4345.060 ;
        RECT 3482.245 4329.350 3483.165 4345.060 ;
        RECT 3481.735 4312.760 3483.165 4329.350 ;
        RECT 3438.620 4311.330 3483.165 4312.760 ;
      LAYER pwell ;
        RECT 3483.975 4315.230 3485.985 4346.160 ;
        RECT 3488.820 4339.120 3491.550 4352.615 ;
        RECT 3487.520 4315.230 3491.550 4339.120 ;
        RECT 3483.975 4314.135 3491.550 4315.230 ;
        RECT 3513.135 4351.755 3518.355 4386.265 ;
        RECT 3513.135 4325.090 3517.315 4351.755 ;
      LAYER nwell ;
        RECT 3518.665 4345.960 3528.380 4392.415 ;
      LAYER pwell ;
        RECT 3513.135 4314.135 3518.355 4325.090 ;
        RECT 3483.975 4311.710 3518.355 4314.135 ;
      LAYER nwell ;
        RECT 3518.665 4311.560 3528.385 4345.960 ;
      LAYER pwell ;
        RECT 3528.685 4311.710 3532.565 4392.290 ;
      LAYER nwell ;
        RECT 3532.880 4385.615 3566.975 4392.415 ;
        RECT 3532.880 4313.370 3534.690 4385.615 ;
        RECT 3556.515 4384.485 3566.975 4385.615 ;
        RECT 3556.515 4325.030 3558.475 4384.485 ;
        RECT 3561.545 4325.030 3566.975 4384.485 ;
        RECT 3556.515 4313.370 3566.975 4325.030 ;
        RECT 3532.880 4311.565 3566.975 4313.370 ;
        RECT 3532.880 4311.560 3558.230 4311.565 ;
        RECT 197.795 4149.860 199.315 4208.965 ;
      LAYER pwell ;
        RECT 3388.935 4155.715 3411.790 4163.505 ;
      LAYER nwell ;
        RECT 3388.685 4096.035 3390.205 4155.140 ;
        RECT 29.770 4002.435 55.120 4002.440 ;
        RECT 21.025 4000.630 55.120 4002.435 ;
        RECT 21.025 3988.970 31.485 4000.630 ;
        RECT 21.025 3929.515 26.455 3988.970 ;
        RECT 29.525 3929.515 31.485 3988.970 ;
        RECT 21.025 3928.385 31.485 3929.515 ;
        RECT 53.310 3928.385 55.120 4000.630 ;
        RECT 21.025 3921.585 55.120 3928.385 ;
      LAYER pwell ;
        RECT 55.435 3921.710 59.315 4002.290 ;
      LAYER nwell ;
        RECT 59.615 3968.040 69.335 4002.440 ;
      LAYER pwell ;
        RECT 69.645 3999.865 104.025 4002.290 ;
        RECT 69.645 3988.910 74.865 3999.865 ;
      LAYER nwell ;
        RECT 59.620 3921.585 69.335 3968.040 ;
      LAYER pwell ;
        RECT 70.685 3962.245 74.865 3988.910 ;
        RECT 69.645 3927.735 74.865 3962.245 ;
        RECT 96.450 3998.770 104.025 3999.865 ;
        RECT 96.450 3974.880 100.480 3998.770 ;
        RECT 96.450 3961.385 99.180 3974.880 ;
        RECT 102.015 3967.840 104.025 3998.770 ;
      LAYER nwell ;
        RECT 104.835 4001.240 149.380 4002.670 ;
        RECT 104.835 3984.650 106.265 4001.240 ;
        RECT 104.835 3968.940 105.755 3984.650 ;
        RECT 115.655 3968.940 116.835 4001.240 ;
        RECT 126.225 4001.125 149.380 4001.240 ;
        RECT 126.225 3984.650 127.405 4001.125 ;
        RECT 133.955 3992.335 134.805 4001.125 ;
        RECT 147.950 3992.335 149.380 4001.125 ;
        RECT 126.735 3968.940 127.405 3984.650 ;
        RECT 163.945 3986.830 170.215 4002.450 ;
        RECT 174.655 3986.830 180.845 4002.450 ;
        RECT 163.945 3980.275 167.590 3986.830 ;
        RECT 163.945 3970.915 165.735 3980.275 ;
      LAYER pwell ;
        RECT 104.740 3967.840 105.045 3968.590 ;
        RECT 102.015 3961.385 105.045 3967.840 ;
        RECT 96.450 3927.735 98.035 3961.385 ;
        RECT 69.645 3927.215 98.035 3927.735 ;
        RECT 103.745 3931.300 105.045 3961.385 ;
        RECT 103.745 3927.215 107.065 3931.300 ;
      LAYER nwell ;
        RECT 112.260 3930.420 113.340 3930.495 ;
        RECT 111.720 3927.975 113.340 3930.420 ;
      LAYER pwell ;
        RECT 69.645 3921.785 107.065 3927.215 ;
      LAYER nwell ;
        RECT 108.180 3926.530 113.340 3927.975 ;
        RECT 108.180 3924.795 114.420 3926.530 ;
        RECT 107.600 3921.880 114.420 3924.795 ;
        RECT 118.765 3922.715 120.195 3946.815 ;
        RECT 138.980 3932.460 139.230 3935.535 ;
        RECT 138.980 3925.810 139.820 3932.460 ;
        RECT 137.660 3922.715 139.820 3925.810 ;
        RECT 141.980 3922.715 143.410 3945.515 ;
        RECT 176.920 3926.580 180.845 3986.830 ;
        RECT 3393.665 3942.890 3397.325 3946.415 ;
        RECT 3444.590 3945.285 3469.235 3946.715 ;
        RECT 3476.485 3946.120 3480.400 3946.415 ;
        RECT 107.600 3921.585 111.515 3921.880 ;
        RECT 118.765 3921.285 143.410 3922.715 ;
        RECT 190.675 3921.585 194.335 3925.110 ;
        RECT 3407.155 3881.170 3411.080 3941.420 ;
        RECT 3444.590 3922.485 3446.020 3945.285 ;
        RECT 3448.180 3942.190 3450.340 3945.285 ;
        RECT 3448.180 3935.540 3449.020 3942.190 ;
        RECT 3448.770 3932.465 3449.020 3935.540 ;
        RECT 3467.805 3921.185 3469.235 3945.285 ;
        RECT 3473.580 3943.205 3480.400 3946.120 ;
        RECT 3473.580 3941.470 3479.820 3943.205 ;
        RECT 3474.660 3940.025 3479.820 3941.470 ;
      LAYER pwell ;
        RECT 3480.935 3940.785 3518.355 3946.215 ;
      LAYER nwell ;
        RECT 3474.660 3937.580 3476.280 3940.025 ;
        RECT 3474.660 3937.505 3475.740 3937.580 ;
      LAYER pwell ;
        RECT 3480.935 3936.700 3484.255 3940.785 ;
        RECT 3482.955 3906.615 3484.255 3936.700 ;
        RECT 3489.965 3940.265 3518.355 3940.785 ;
        RECT 3489.965 3906.615 3491.550 3940.265 ;
        RECT 3482.955 3900.160 3485.985 3906.615 ;
        RECT 3482.955 3899.410 3483.260 3900.160 ;
      LAYER nwell ;
        RECT 3422.265 3887.725 3424.055 3897.085 ;
        RECT 3420.410 3881.170 3424.055 3887.725 ;
        RECT 3407.155 3865.550 3413.345 3881.170 ;
        RECT 3417.785 3865.550 3424.055 3881.170 ;
        RECT 3460.595 3883.350 3461.265 3899.060 ;
        RECT 3438.620 3866.875 3440.050 3875.665 ;
        RECT 3453.195 3866.875 3454.045 3875.665 ;
        RECT 3460.595 3866.875 3461.775 3883.350 ;
        RECT 3438.620 3866.760 3461.775 3866.875 ;
        RECT 3471.165 3866.760 3472.345 3899.060 ;
        RECT 3482.245 3883.350 3483.165 3899.060 ;
        RECT 3481.735 3866.760 3483.165 3883.350 ;
        RECT 3438.620 3865.330 3483.165 3866.760 ;
      LAYER pwell ;
        RECT 3483.975 3869.230 3485.985 3900.160 ;
        RECT 3488.820 3893.120 3491.550 3906.615 ;
        RECT 3487.520 3869.230 3491.550 3893.120 ;
        RECT 3483.975 3868.135 3491.550 3869.230 ;
        RECT 3513.135 3905.755 3518.355 3940.265 ;
        RECT 3513.135 3879.090 3517.315 3905.755 ;
      LAYER nwell ;
        RECT 3518.665 3899.960 3528.380 3946.415 ;
      LAYER pwell ;
        RECT 3513.135 3868.135 3518.355 3879.090 ;
        RECT 3483.975 3865.710 3518.355 3868.135 ;
      LAYER nwell ;
        RECT 3518.665 3865.560 3528.385 3899.960 ;
      LAYER pwell ;
        RECT 3528.685 3865.710 3532.565 3946.290 ;
      LAYER nwell ;
        RECT 3532.880 3939.615 3566.975 3946.415 ;
        RECT 3532.880 3867.370 3534.690 3939.615 ;
        RECT 3556.515 3938.485 3566.975 3939.615 ;
        RECT 3556.515 3879.030 3558.475 3938.485 ;
        RECT 3561.545 3879.030 3566.975 3938.485 ;
        RECT 3556.515 3867.370 3566.975 3879.030 ;
        RECT 3532.880 3865.565 3566.975 3867.370 ;
        RECT 3532.880 3865.560 3558.230 3865.565 ;
        RECT 29.770 3786.435 55.120 3786.440 ;
        RECT 21.025 3784.630 55.120 3786.435 ;
        RECT 21.025 3772.970 31.485 3784.630 ;
        RECT 21.025 3713.515 26.455 3772.970 ;
        RECT 29.525 3713.515 31.485 3772.970 ;
        RECT 21.025 3712.385 31.485 3713.515 ;
        RECT 53.310 3712.385 55.120 3784.630 ;
        RECT 21.025 3705.585 55.120 3712.385 ;
      LAYER pwell ;
        RECT 55.435 3705.710 59.315 3786.290 ;
      LAYER nwell ;
        RECT 59.615 3752.040 69.335 3786.440 ;
      LAYER pwell ;
        RECT 69.645 3783.865 104.025 3786.290 ;
        RECT 69.645 3772.910 74.865 3783.865 ;
      LAYER nwell ;
        RECT 59.620 3705.585 69.335 3752.040 ;
      LAYER pwell ;
        RECT 70.685 3746.245 74.865 3772.910 ;
        RECT 69.645 3711.735 74.865 3746.245 ;
        RECT 96.450 3782.770 104.025 3783.865 ;
        RECT 96.450 3758.880 100.480 3782.770 ;
        RECT 96.450 3745.385 99.180 3758.880 ;
        RECT 102.015 3751.840 104.025 3782.770 ;
      LAYER nwell ;
        RECT 104.835 3785.240 149.380 3786.670 ;
        RECT 104.835 3768.650 106.265 3785.240 ;
        RECT 104.835 3752.940 105.755 3768.650 ;
        RECT 115.655 3752.940 116.835 3785.240 ;
        RECT 126.225 3785.125 149.380 3785.240 ;
        RECT 126.225 3768.650 127.405 3785.125 ;
        RECT 133.955 3776.335 134.805 3785.125 ;
        RECT 147.950 3776.335 149.380 3785.125 ;
        RECT 126.735 3752.940 127.405 3768.650 ;
        RECT 163.945 3770.830 170.215 3786.450 ;
        RECT 174.655 3770.830 180.845 3786.450 ;
        RECT 163.945 3764.275 167.590 3770.830 ;
        RECT 163.945 3754.915 165.735 3764.275 ;
      LAYER pwell ;
        RECT 104.740 3751.840 105.045 3752.590 ;
        RECT 102.015 3745.385 105.045 3751.840 ;
        RECT 96.450 3711.735 98.035 3745.385 ;
        RECT 69.645 3711.215 98.035 3711.735 ;
        RECT 103.745 3715.300 105.045 3745.385 ;
        RECT 103.745 3711.215 107.065 3715.300 ;
      LAYER nwell ;
        RECT 112.260 3714.420 113.340 3714.495 ;
        RECT 111.720 3711.975 113.340 3714.420 ;
      LAYER pwell ;
        RECT 69.645 3705.785 107.065 3711.215 ;
      LAYER nwell ;
        RECT 108.180 3710.530 113.340 3711.975 ;
        RECT 108.180 3708.795 114.420 3710.530 ;
        RECT 107.600 3705.880 114.420 3708.795 ;
        RECT 118.765 3706.715 120.195 3730.815 ;
        RECT 138.980 3716.460 139.230 3719.535 ;
        RECT 138.980 3709.810 139.820 3716.460 ;
        RECT 137.660 3706.715 139.820 3709.810 ;
        RECT 141.980 3706.715 143.410 3729.515 ;
        RECT 176.920 3710.580 180.845 3770.830 ;
        RECT 3393.665 3717.890 3397.325 3721.415 ;
        RECT 3444.590 3720.285 3469.235 3721.715 ;
        RECT 3476.485 3721.120 3480.400 3721.415 ;
        RECT 107.600 3705.585 111.515 3705.880 ;
        RECT 118.765 3705.285 143.410 3706.715 ;
        RECT 190.675 3705.585 194.335 3709.110 ;
        RECT 3407.155 3656.170 3411.080 3716.420 ;
        RECT 3444.590 3697.485 3446.020 3720.285 ;
        RECT 3448.180 3717.190 3450.340 3720.285 ;
        RECT 3448.180 3710.540 3449.020 3717.190 ;
        RECT 3448.770 3707.465 3449.020 3710.540 ;
        RECT 3467.805 3696.185 3469.235 3720.285 ;
        RECT 3473.580 3718.205 3480.400 3721.120 ;
        RECT 3473.580 3716.470 3479.820 3718.205 ;
        RECT 3474.660 3715.025 3479.820 3716.470 ;
      LAYER pwell ;
        RECT 3480.935 3715.785 3518.355 3721.215 ;
      LAYER nwell ;
        RECT 3474.660 3712.580 3476.280 3715.025 ;
        RECT 3474.660 3712.505 3475.740 3712.580 ;
      LAYER pwell ;
        RECT 3480.935 3711.700 3484.255 3715.785 ;
        RECT 3482.955 3681.615 3484.255 3711.700 ;
        RECT 3489.965 3715.265 3518.355 3715.785 ;
        RECT 3489.965 3681.615 3491.550 3715.265 ;
        RECT 3482.955 3675.160 3485.985 3681.615 ;
        RECT 3482.955 3674.410 3483.260 3675.160 ;
      LAYER nwell ;
        RECT 3422.265 3662.725 3424.055 3672.085 ;
        RECT 3420.410 3656.170 3424.055 3662.725 ;
        RECT 3407.155 3640.550 3413.345 3656.170 ;
        RECT 3417.785 3640.550 3424.055 3656.170 ;
        RECT 3460.595 3658.350 3461.265 3674.060 ;
        RECT 3438.620 3641.875 3440.050 3650.665 ;
        RECT 3453.195 3641.875 3454.045 3650.665 ;
        RECT 3460.595 3641.875 3461.775 3658.350 ;
        RECT 3438.620 3641.760 3461.775 3641.875 ;
        RECT 3471.165 3641.760 3472.345 3674.060 ;
        RECT 3482.245 3658.350 3483.165 3674.060 ;
        RECT 3481.735 3641.760 3483.165 3658.350 ;
        RECT 3438.620 3640.330 3483.165 3641.760 ;
      LAYER pwell ;
        RECT 3483.975 3644.230 3485.985 3675.160 ;
        RECT 3488.820 3668.120 3491.550 3681.615 ;
        RECT 3487.520 3644.230 3491.550 3668.120 ;
        RECT 3483.975 3643.135 3491.550 3644.230 ;
        RECT 3513.135 3680.755 3518.355 3715.265 ;
        RECT 3513.135 3654.090 3517.315 3680.755 ;
      LAYER nwell ;
        RECT 3518.665 3674.960 3528.380 3721.415 ;
      LAYER pwell ;
        RECT 3513.135 3643.135 3518.355 3654.090 ;
        RECT 3483.975 3640.710 3518.355 3643.135 ;
      LAYER nwell ;
        RECT 3518.665 3640.560 3528.385 3674.960 ;
      LAYER pwell ;
        RECT 3528.685 3640.710 3532.565 3721.290 ;
      LAYER nwell ;
        RECT 3532.880 3714.615 3566.975 3721.415 ;
        RECT 3532.880 3642.370 3534.690 3714.615 ;
        RECT 3556.515 3713.485 3566.975 3714.615 ;
        RECT 3556.515 3654.030 3558.475 3713.485 ;
        RECT 3561.545 3654.030 3566.975 3713.485 ;
        RECT 3556.515 3642.370 3566.975 3654.030 ;
        RECT 3532.880 3640.565 3566.975 3642.370 ;
        RECT 3532.880 3640.560 3558.230 3640.565 ;
        RECT 29.770 3570.435 55.120 3570.440 ;
        RECT 21.025 3568.630 55.120 3570.435 ;
        RECT 21.025 3556.970 31.485 3568.630 ;
        RECT 21.025 3497.515 26.455 3556.970 ;
        RECT 29.525 3497.515 31.485 3556.970 ;
        RECT 21.025 3496.385 31.485 3497.515 ;
        RECT 53.310 3496.385 55.120 3568.630 ;
        RECT 21.025 3489.585 55.120 3496.385 ;
      LAYER pwell ;
        RECT 55.435 3489.710 59.315 3570.290 ;
      LAYER nwell ;
        RECT 59.615 3536.040 69.335 3570.440 ;
      LAYER pwell ;
        RECT 69.645 3567.865 104.025 3570.290 ;
        RECT 69.645 3556.910 74.865 3567.865 ;
      LAYER nwell ;
        RECT 59.620 3489.585 69.335 3536.040 ;
      LAYER pwell ;
        RECT 70.685 3530.245 74.865 3556.910 ;
        RECT 69.645 3495.735 74.865 3530.245 ;
        RECT 96.450 3566.770 104.025 3567.865 ;
        RECT 96.450 3542.880 100.480 3566.770 ;
        RECT 96.450 3529.385 99.180 3542.880 ;
        RECT 102.015 3535.840 104.025 3566.770 ;
      LAYER nwell ;
        RECT 104.835 3569.240 149.380 3570.670 ;
        RECT 104.835 3552.650 106.265 3569.240 ;
        RECT 104.835 3536.940 105.755 3552.650 ;
        RECT 115.655 3536.940 116.835 3569.240 ;
        RECT 126.225 3569.125 149.380 3569.240 ;
        RECT 126.225 3552.650 127.405 3569.125 ;
        RECT 133.955 3560.335 134.805 3569.125 ;
        RECT 147.950 3560.335 149.380 3569.125 ;
        RECT 126.735 3536.940 127.405 3552.650 ;
        RECT 163.945 3554.830 170.215 3570.450 ;
        RECT 174.655 3554.830 180.845 3570.450 ;
        RECT 163.945 3548.275 167.590 3554.830 ;
        RECT 163.945 3538.915 165.735 3548.275 ;
      LAYER pwell ;
        RECT 104.740 3535.840 105.045 3536.590 ;
        RECT 102.015 3529.385 105.045 3535.840 ;
        RECT 96.450 3495.735 98.035 3529.385 ;
        RECT 69.645 3495.215 98.035 3495.735 ;
        RECT 103.745 3499.300 105.045 3529.385 ;
        RECT 103.745 3495.215 107.065 3499.300 ;
      LAYER nwell ;
        RECT 112.260 3498.420 113.340 3498.495 ;
        RECT 111.720 3495.975 113.340 3498.420 ;
      LAYER pwell ;
        RECT 69.645 3489.785 107.065 3495.215 ;
      LAYER nwell ;
        RECT 108.180 3494.530 113.340 3495.975 ;
        RECT 108.180 3492.795 114.420 3494.530 ;
        RECT 107.600 3489.880 114.420 3492.795 ;
        RECT 118.765 3490.715 120.195 3514.815 ;
        RECT 138.980 3500.460 139.230 3503.535 ;
        RECT 138.980 3493.810 139.820 3500.460 ;
        RECT 137.660 3490.715 139.820 3493.810 ;
        RECT 141.980 3490.715 143.410 3513.515 ;
        RECT 176.920 3494.580 180.845 3554.830 ;
        RECT 107.600 3489.585 111.515 3489.880 ;
        RECT 118.765 3489.285 143.410 3490.715 ;
        RECT 190.675 3489.585 194.335 3493.110 ;
        RECT 3393.665 3492.890 3397.325 3496.415 ;
        RECT 3444.590 3495.285 3469.235 3496.715 ;
        RECT 3476.485 3496.120 3480.400 3496.415 ;
        RECT 3407.155 3431.170 3411.080 3491.420 ;
        RECT 3444.590 3472.485 3446.020 3495.285 ;
        RECT 3448.180 3492.190 3450.340 3495.285 ;
        RECT 3448.180 3485.540 3449.020 3492.190 ;
        RECT 3448.770 3482.465 3449.020 3485.540 ;
        RECT 3467.805 3471.185 3469.235 3495.285 ;
        RECT 3473.580 3493.205 3480.400 3496.120 ;
        RECT 3473.580 3491.470 3479.820 3493.205 ;
        RECT 3474.660 3490.025 3479.820 3491.470 ;
      LAYER pwell ;
        RECT 3480.935 3490.785 3518.355 3496.215 ;
      LAYER nwell ;
        RECT 3474.660 3487.580 3476.280 3490.025 ;
        RECT 3474.660 3487.505 3475.740 3487.580 ;
      LAYER pwell ;
        RECT 3480.935 3486.700 3484.255 3490.785 ;
        RECT 3482.955 3456.615 3484.255 3486.700 ;
        RECT 3489.965 3490.265 3518.355 3490.785 ;
        RECT 3489.965 3456.615 3491.550 3490.265 ;
        RECT 3482.955 3450.160 3485.985 3456.615 ;
        RECT 3482.955 3449.410 3483.260 3450.160 ;
      LAYER nwell ;
        RECT 3422.265 3437.725 3424.055 3447.085 ;
        RECT 3420.410 3431.170 3424.055 3437.725 ;
        RECT 3407.155 3415.550 3413.345 3431.170 ;
        RECT 3417.785 3415.550 3424.055 3431.170 ;
        RECT 3460.595 3433.350 3461.265 3449.060 ;
        RECT 3438.620 3416.875 3440.050 3425.665 ;
        RECT 3453.195 3416.875 3454.045 3425.665 ;
        RECT 3460.595 3416.875 3461.775 3433.350 ;
        RECT 3438.620 3416.760 3461.775 3416.875 ;
        RECT 3471.165 3416.760 3472.345 3449.060 ;
        RECT 3482.245 3433.350 3483.165 3449.060 ;
        RECT 3481.735 3416.760 3483.165 3433.350 ;
        RECT 3438.620 3415.330 3483.165 3416.760 ;
      LAYER pwell ;
        RECT 3483.975 3419.230 3485.985 3450.160 ;
        RECT 3488.820 3443.120 3491.550 3456.615 ;
        RECT 3487.520 3419.230 3491.550 3443.120 ;
        RECT 3483.975 3418.135 3491.550 3419.230 ;
        RECT 3513.135 3455.755 3518.355 3490.265 ;
        RECT 3513.135 3429.090 3517.315 3455.755 ;
      LAYER nwell ;
        RECT 3518.665 3449.960 3528.380 3496.415 ;
      LAYER pwell ;
        RECT 3513.135 3418.135 3518.355 3429.090 ;
        RECT 3483.975 3415.710 3518.355 3418.135 ;
      LAYER nwell ;
        RECT 3518.665 3415.560 3528.385 3449.960 ;
      LAYER pwell ;
        RECT 3528.685 3415.710 3532.565 3496.290 ;
      LAYER nwell ;
        RECT 3532.880 3489.615 3566.975 3496.415 ;
        RECT 3532.880 3417.370 3534.690 3489.615 ;
        RECT 3556.515 3488.485 3566.975 3489.615 ;
        RECT 3556.515 3429.030 3558.475 3488.485 ;
        RECT 3561.545 3429.030 3566.975 3488.485 ;
        RECT 3556.515 3417.370 3566.975 3429.030 ;
        RECT 3532.880 3415.565 3566.975 3417.370 ;
        RECT 3532.880 3415.560 3558.230 3415.565 ;
        RECT 29.770 3354.435 55.120 3354.440 ;
        RECT 21.025 3352.630 55.120 3354.435 ;
        RECT 21.025 3340.970 31.485 3352.630 ;
        RECT 21.025 3281.515 26.455 3340.970 ;
        RECT 29.525 3281.515 31.485 3340.970 ;
        RECT 21.025 3280.385 31.485 3281.515 ;
        RECT 53.310 3280.385 55.120 3352.630 ;
        RECT 21.025 3273.585 55.120 3280.385 ;
      LAYER pwell ;
        RECT 55.435 3273.710 59.315 3354.290 ;
      LAYER nwell ;
        RECT 59.615 3320.040 69.335 3354.440 ;
      LAYER pwell ;
        RECT 69.645 3351.865 104.025 3354.290 ;
        RECT 69.645 3340.910 74.865 3351.865 ;
      LAYER nwell ;
        RECT 59.620 3273.585 69.335 3320.040 ;
      LAYER pwell ;
        RECT 70.685 3314.245 74.865 3340.910 ;
        RECT 69.645 3279.735 74.865 3314.245 ;
        RECT 96.450 3350.770 104.025 3351.865 ;
        RECT 96.450 3326.880 100.480 3350.770 ;
        RECT 96.450 3313.385 99.180 3326.880 ;
        RECT 102.015 3319.840 104.025 3350.770 ;
      LAYER nwell ;
        RECT 104.835 3353.240 149.380 3354.670 ;
        RECT 104.835 3336.650 106.265 3353.240 ;
        RECT 104.835 3320.940 105.755 3336.650 ;
        RECT 115.655 3320.940 116.835 3353.240 ;
        RECT 126.225 3353.125 149.380 3353.240 ;
        RECT 126.225 3336.650 127.405 3353.125 ;
        RECT 133.955 3344.335 134.805 3353.125 ;
        RECT 147.950 3344.335 149.380 3353.125 ;
        RECT 126.735 3320.940 127.405 3336.650 ;
        RECT 163.945 3338.830 170.215 3354.450 ;
        RECT 174.655 3338.830 180.845 3354.450 ;
        RECT 163.945 3332.275 167.590 3338.830 ;
        RECT 163.945 3322.915 165.735 3332.275 ;
      LAYER pwell ;
        RECT 104.740 3319.840 105.045 3320.590 ;
        RECT 102.015 3313.385 105.045 3319.840 ;
        RECT 96.450 3279.735 98.035 3313.385 ;
        RECT 69.645 3279.215 98.035 3279.735 ;
        RECT 103.745 3283.300 105.045 3313.385 ;
        RECT 103.745 3279.215 107.065 3283.300 ;
      LAYER nwell ;
        RECT 112.260 3282.420 113.340 3282.495 ;
        RECT 111.720 3279.975 113.340 3282.420 ;
      LAYER pwell ;
        RECT 69.645 3273.785 107.065 3279.215 ;
      LAYER nwell ;
        RECT 108.180 3278.530 113.340 3279.975 ;
        RECT 108.180 3276.795 114.420 3278.530 ;
        RECT 107.600 3273.880 114.420 3276.795 ;
        RECT 118.765 3274.715 120.195 3298.815 ;
        RECT 138.980 3284.460 139.230 3287.535 ;
        RECT 138.980 3277.810 139.820 3284.460 ;
        RECT 137.660 3274.715 139.820 3277.810 ;
        RECT 141.980 3274.715 143.410 3297.515 ;
        RECT 176.920 3278.580 180.845 3338.830 ;
        RECT 107.600 3273.585 111.515 3273.880 ;
        RECT 118.765 3273.285 143.410 3274.715 ;
        RECT 190.675 3273.585 194.335 3277.110 ;
        RECT 3393.665 3266.890 3397.325 3270.415 ;
        RECT 3444.590 3269.285 3469.235 3270.715 ;
        RECT 3476.485 3270.120 3480.400 3270.415 ;
        RECT 3407.155 3205.170 3411.080 3265.420 ;
        RECT 3444.590 3246.485 3446.020 3269.285 ;
        RECT 3448.180 3266.190 3450.340 3269.285 ;
        RECT 3448.180 3259.540 3449.020 3266.190 ;
        RECT 3448.770 3256.465 3449.020 3259.540 ;
        RECT 3467.805 3245.185 3469.235 3269.285 ;
        RECT 3473.580 3267.205 3480.400 3270.120 ;
        RECT 3473.580 3265.470 3479.820 3267.205 ;
        RECT 3474.660 3264.025 3479.820 3265.470 ;
      LAYER pwell ;
        RECT 3480.935 3264.785 3518.355 3270.215 ;
      LAYER nwell ;
        RECT 3474.660 3261.580 3476.280 3264.025 ;
        RECT 3474.660 3261.505 3475.740 3261.580 ;
      LAYER pwell ;
        RECT 3480.935 3260.700 3484.255 3264.785 ;
        RECT 3482.955 3230.615 3484.255 3260.700 ;
        RECT 3489.965 3264.265 3518.355 3264.785 ;
        RECT 3489.965 3230.615 3491.550 3264.265 ;
        RECT 3482.955 3224.160 3485.985 3230.615 ;
        RECT 3482.955 3223.410 3483.260 3224.160 ;
      LAYER nwell ;
        RECT 3422.265 3211.725 3424.055 3221.085 ;
        RECT 3420.410 3205.170 3424.055 3211.725 ;
        RECT 3407.155 3189.550 3413.345 3205.170 ;
        RECT 3417.785 3189.550 3424.055 3205.170 ;
        RECT 3460.595 3207.350 3461.265 3223.060 ;
        RECT 3438.620 3190.875 3440.050 3199.665 ;
        RECT 3453.195 3190.875 3454.045 3199.665 ;
        RECT 3460.595 3190.875 3461.775 3207.350 ;
        RECT 3438.620 3190.760 3461.775 3190.875 ;
        RECT 3471.165 3190.760 3472.345 3223.060 ;
        RECT 3482.245 3207.350 3483.165 3223.060 ;
        RECT 3481.735 3190.760 3483.165 3207.350 ;
        RECT 3438.620 3189.330 3483.165 3190.760 ;
      LAYER pwell ;
        RECT 3483.975 3193.230 3485.985 3224.160 ;
        RECT 3488.820 3217.120 3491.550 3230.615 ;
        RECT 3487.520 3193.230 3491.550 3217.120 ;
        RECT 3483.975 3192.135 3491.550 3193.230 ;
        RECT 3513.135 3229.755 3518.355 3264.265 ;
        RECT 3513.135 3203.090 3517.315 3229.755 ;
      LAYER nwell ;
        RECT 3518.665 3223.960 3528.380 3270.415 ;
      LAYER pwell ;
        RECT 3513.135 3192.135 3518.355 3203.090 ;
        RECT 3483.975 3189.710 3518.355 3192.135 ;
      LAYER nwell ;
        RECT 3518.665 3189.560 3528.385 3223.960 ;
      LAYER pwell ;
        RECT 3528.685 3189.710 3532.565 3270.290 ;
      LAYER nwell ;
        RECT 3532.880 3263.615 3566.975 3270.415 ;
        RECT 3532.880 3191.370 3534.690 3263.615 ;
        RECT 3556.515 3262.485 3566.975 3263.615 ;
        RECT 3556.515 3203.030 3558.475 3262.485 ;
        RECT 3561.545 3203.030 3566.975 3262.485 ;
        RECT 3556.515 3191.370 3566.975 3203.030 ;
        RECT 3532.880 3189.565 3566.975 3191.370 ;
        RECT 3532.880 3189.560 3558.230 3189.565 ;
        RECT 29.770 3138.435 55.120 3138.440 ;
        RECT 21.025 3136.630 55.120 3138.435 ;
        RECT 21.025 3124.970 31.485 3136.630 ;
        RECT 21.025 3065.515 26.455 3124.970 ;
        RECT 29.525 3065.515 31.485 3124.970 ;
        RECT 21.025 3064.385 31.485 3065.515 ;
        RECT 53.310 3064.385 55.120 3136.630 ;
        RECT 21.025 3057.585 55.120 3064.385 ;
      LAYER pwell ;
        RECT 55.435 3057.710 59.315 3138.290 ;
      LAYER nwell ;
        RECT 59.615 3104.040 69.335 3138.440 ;
      LAYER pwell ;
        RECT 69.645 3135.865 104.025 3138.290 ;
        RECT 69.645 3124.910 74.865 3135.865 ;
      LAYER nwell ;
        RECT 59.620 3057.585 69.335 3104.040 ;
      LAYER pwell ;
        RECT 70.685 3098.245 74.865 3124.910 ;
        RECT 69.645 3063.735 74.865 3098.245 ;
        RECT 96.450 3134.770 104.025 3135.865 ;
        RECT 96.450 3110.880 100.480 3134.770 ;
        RECT 96.450 3097.385 99.180 3110.880 ;
        RECT 102.015 3103.840 104.025 3134.770 ;
      LAYER nwell ;
        RECT 104.835 3137.240 149.380 3138.670 ;
        RECT 104.835 3120.650 106.265 3137.240 ;
        RECT 104.835 3104.940 105.755 3120.650 ;
        RECT 115.655 3104.940 116.835 3137.240 ;
        RECT 126.225 3137.125 149.380 3137.240 ;
        RECT 126.225 3120.650 127.405 3137.125 ;
        RECT 133.955 3128.335 134.805 3137.125 ;
        RECT 147.950 3128.335 149.380 3137.125 ;
        RECT 126.735 3104.940 127.405 3120.650 ;
        RECT 163.945 3122.830 170.215 3138.450 ;
        RECT 174.655 3122.830 180.845 3138.450 ;
        RECT 163.945 3116.275 167.590 3122.830 ;
        RECT 163.945 3106.915 165.735 3116.275 ;
      LAYER pwell ;
        RECT 104.740 3103.840 105.045 3104.590 ;
        RECT 102.015 3097.385 105.045 3103.840 ;
        RECT 96.450 3063.735 98.035 3097.385 ;
        RECT 69.645 3063.215 98.035 3063.735 ;
        RECT 103.745 3067.300 105.045 3097.385 ;
        RECT 103.745 3063.215 107.065 3067.300 ;
      LAYER nwell ;
        RECT 112.260 3066.420 113.340 3066.495 ;
        RECT 111.720 3063.975 113.340 3066.420 ;
      LAYER pwell ;
        RECT 69.645 3057.785 107.065 3063.215 ;
      LAYER nwell ;
        RECT 108.180 3062.530 113.340 3063.975 ;
        RECT 108.180 3060.795 114.420 3062.530 ;
        RECT 107.600 3057.880 114.420 3060.795 ;
        RECT 118.765 3058.715 120.195 3082.815 ;
        RECT 138.980 3068.460 139.230 3071.535 ;
        RECT 138.980 3061.810 139.820 3068.460 ;
        RECT 137.660 3058.715 139.820 3061.810 ;
        RECT 141.980 3058.715 143.410 3081.515 ;
        RECT 176.920 3062.580 180.845 3122.830 ;
        RECT 107.600 3057.585 111.515 3057.880 ;
        RECT 118.765 3057.285 143.410 3058.715 ;
        RECT 190.675 3057.585 194.335 3061.110 ;
        RECT 3393.665 3041.890 3397.325 3045.415 ;
        RECT 3444.590 3044.285 3469.235 3045.715 ;
        RECT 3476.485 3045.120 3480.400 3045.415 ;
        RECT 3407.155 2980.170 3411.080 3040.420 ;
        RECT 3444.590 3021.485 3446.020 3044.285 ;
        RECT 3448.180 3041.190 3450.340 3044.285 ;
        RECT 3448.180 3034.540 3449.020 3041.190 ;
        RECT 3448.770 3031.465 3449.020 3034.540 ;
        RECT 3467.805 3020.185 3469.235 3044.285 ;
        RECT 3473.580 3042.205 3480.400 3045.120 ;
        RECT 3473.580 3040.470 3479.820 3042.205 ;
        RECT 3474.660 3039.025 3479.820 3040.470 ;
      LAYER pwell ;
        RECT 3480.935 3039.785 3518.355 3045.215 ;
      LAYER nwell ;
        RECT 3474.660 3036.580 3476.280 3039.025 ;
        RECT 3474.660 3036.505 3475.740 3036.580 ;
      LAYER pwell ;
        RECT 3480.935 3035.700 3484.255 3039.785 ;
        RECT 3482.955 3005.615 3484.255 3035.700 ;
        RECT 3489.965 3039.265 3518.355 3039.785 ;
        RECT 3489.965 3005.615 3491.550 3039.265 ;
        RECT 3482.955 2999.160 3485.985 3005.615 ;
        RECT 3482.955 2998.410 3483.260 2999.160 ;
      LAYER nwell ;
        RECT 3422.265 2986.725 3424.055 2996.085 ;
        RECT 3420.410 2980.170 3424.055 2986.725 ;
        RECT 3407.155 2964.550 3413.345 2980.170 ;
        RECT 3417.785 2964.550 3424.055 2980.170 ;
        RECT 3460.595 2982.350 3461.265 2998.060 ;
        RECT 3438.620 2965.875 3440.050 2974.665 ;
        RECT 3453.195 2965.875 3454.045 2974.665 ;
        RECT 3460.595 2965.875 3461.775 2982.350 ;
        RECT 3438.620 2965.760 3461.775 2965.875 ;
        RECT 3471.165 2965.760 3472.345 2998.060 ;
        RECT 3482.245 2982.350 3483.165 2998.060 ;
        RECT 3481.735 2965.760 3483.165 2982.350 ;
        RECT 3438.620 2964.330 3483.165 2965.760 ;
      LAYER pwell ;
        RECT 3483.975 2968.230 3485.985 2999.160 ;
        RECT 3488.820 2992.120 3491.550 3005.615 ;
        RECT 3487.520 2968.230 3491.550 2992.120 ;
        RECT 3483.975 2967.135 3491.550 2968.230 ;
        RECT 3513.135 3004.755 3518.355 3039.265 ;
        RECT 3513.135 2978.090 3517.315 3004.755 ;
      LAYER nwell ;
        RECT 3518.665 2998.960 3528.380 3045.415 ;
      LAYER pwell ;
        RECT 3513.135 2967.135 3518.355 2978.090 ;
        RECT 3483.975 2964.710 3518.355 2967.135 ;
      LAYER nwell ;
        RECT 3518.665 2964.560 3528.385 2998.960 ;
      LAYER pwell ;
        RECT 3528.685 2964.710 3532.565 3045.290 ;
      LAYER nwell ;
        RECT 3532.880 3038.615 3566.975 3045.415 ;
        RECT 3532.880 2966.370 3534.690 3038.615 ;
        RECT 3556.515 3037.485 3566.975 3038.615 ;
        RECT 3556.515 2978.030 3558.475 3037.485 ;
        RECT 3561.545 2978.030 3566.975 3037.485 ;
        RECT 3556.515 2966.370 3566.975 2978.030 ;
        RECT 3532.880 2964.565 3566.975 2966.370 ;
        RECT 3532.880 2964.560 3558.230 2964.565 ;
        RECT 29.770 2922.435 55.120 2922.440 ;
        RECT 21.025 2920.630 55.120 2922.435 ;
        RECT 21.025 2908.970 31.485 2920.630 ;
        RECT 21.025 2849.515 26.455 2908.970 ;
        RECT 29.525 2849.515 31.485 2908.970 ;
        RECT 21.025 2848.385 31.485 2849.515 ;
        RECT 53.310 2848.385 55.120 2920.630 ;
        RECT 21.025 2841.585 55.120 2848.385 ;
      LAYER pwell ;
        RECT 55.435 2841.710 59.315 2922.290 ;
      LAYER nwell ;
        RECT 59.615 2888.040 69.335 2922.440 ;
      LAYER pwell ;
        RECT 69.645 2919.865 104.025 2922.290 ;
        RECT 69.645 2908.910 74.865 2919.865 ;
      LAYER nwell ;
        RECT 59.620 2841.585 69.335 2888.040 ;
      LAYER pwell ;
        RECT 70.685 2882.245 74.865 2908.910 ;
        RECT 69.645 2847.735 74.865 2882.245 ;
        RECT 96.450 2918.770 104.025 2919.865 ;
        RECT 96.450 2894.880 100.480 2918.770 ;
        RECT 96.450 2881.385 99.180 2894.880 ;
        RECT 102.015 2887.840 104.025 2918.770 ;
      LAYER nwell ;
        RECT 104.835 2921.240 149.380 2922.670 ;
        RECT 104.835 2904.650 106.265 2921.240 ;
        RECT 104.835 2888.940 105.755 2904.650 ;
        RECT 115.655 2888.940 116.835 2921.240 ;
        RECT 126.225 2921.125 149.380 2921.240 ;
        RECT 126.225 2904.650 127.405 2921.125 ;
        RECT 133.955 2912.335 134.805 2921.125 ;
        RECT 147.950 2912.335 149.380 2921.125 ;
        RECT 126.735 2888.940 127.405 2904.650 ;
        RECT 163.945 2906.830 170.215 2922.450 ;
        RECT 174.655 2906.830 180.845 2922.450 ;
        RECT 163.945 2900.275 167.590 2906.830 ;
        RECT 163.945 2890.915 165.735 2900.275 ;
      LAYER pwell ;
        RECT 104.740 2887.840 105.045 2888.590 ;
        RECT 102.015 2881.385 105.045 2887.840 ;
        RECT 96.450 2847.735 98.035 2881.385 ;
        RECT 69.645 2847.215 98.035 2847.735 ;
        RECT 103.745 2851.300 105.045 2881.385 ;
        RECT 103.745 2847.215 107.065 2851.300 ;
      LAYER nwell ;
        RECT 112.260 2850.420 113.340 2850.495 ;
        RECT 111.720 2847.975 113.340 2850.420 ;
      LAYER pwell ;
        RECT 69.645 2841.785 107.065 2847.215 ;
      LAYER nwell ;
        RECT 108.180 2846.530 113.340 2847.975 ;
        RECT 108.180 2844.795 114.420 2846.530 ;
        RECT 107.600 2841.880 114.420 2844.795 ;
        RECT 118.765 2842.715 120.195 2866.815 ;
        RECT 138.980 2852.460 139.230 2855.535 ;
        RECT 138.980 2845.810 139.820 2852.460 ;
        RECT 137.660 2842.715 139.820 2845.810 ;
        RECT 141.980 2842.715 143.410 2865.515 ;
        RECT 176.920 2846.580 180.845 2906.830 ;
        RECT 107.600 2841.585 111.515 2841.880 ;
        RECT 118.765 2841.285 143.410 2842.715 ;
        RECT 190.675 2841.585 194.335 2845.110 ;
        RECT 3393.665 2815.890 3397.325 2819.415 ;
        RECT 3444.590 2818.285 3469.235 2819.715 ;
        RECT 3476.485 2819.120 3480.400 2819.415 ;
        RECT 3407.155 2754.170 3411.080 2814.420 ;
        RECT 3444.590 2795.485 3446.020 2818.285 ;
        RECT 3448.180 2815.190 3450.340 2818.285 ;
        RECT 3448.180 2808.540 3449.020 2815.190 ;
        RECT 3448.770 2805.465 3449.020 2808.540 ;
        RECT 3467.805 2794.185 3469.235 2818.285 ;
        RECT 3473.580 2816.205 3480.400 2819.120 ;
        RECT 3473.580 2814.470 3479.820 2816.205 ;
        RECT 3474.660 2813.025 3479.820 2814.470 ;
      LAYER pwell ;
        RECT 3480.935 2813.785 3518.355 2819.215 ;
      LAYER nwell ;
        RECT 3474.660 2810.580 3476.280 2813.025 ;
        RECT 3474.660 2810.505 3475.740 2810.580 ;
      LAYER pwell ;
        RECT 3480.935 2809.700 3484.255 2813.785 ;
        RECT 3482.955 2779.615 3484.255 2809.700 ;
        RECT 3489.965 2813.265 3518.355 2813.785 ;
        RECT 3489.965 2779.615 3491.550 2813.265 ;
        RECT 3482.955 2773.160 3485.985 2779.615 ;
        RECT 3482.955 2772.410 3483.260 2773.160 ;
      LAYER nwell ;
        RECT 3422.265 2760.725 3424.055 2770.085 ;
        RECT 3420.410 2754.170 3424.055 2760.725 ;
        RECT 3407.155 2738.550 3413.345 2754.170 ;
        RECT 3417.785 2738.550 3424.055 2754.170 ;
        RECT 3460.595 2756.350 3461.265 2772.060 ;
        RECT 3438.620 2739.875 3440.050 2748.665 ;
        RECT 3453.195 2739.875 3454.045 2748.665 ;
        RECT 3460.595 2739.875 3461.775 2756.350 ;
        RECT 3438.620 2739.760 3461.775 2739.875 ;
        RECT 3471.165 2739.760 3472.345 2772.060 ;
        RECT 3482.245 2756.350 3483.165 2772.060 ;
        RECT 3481.735 2739.760 3483.165 2756.350 ;
        RECT 3438.620 2738.330 3483.165 2739.760 ;
      LAYER pwell ;
        RECT 3483.975 2742.230 3485.985 2773.160 ;
        RECT 3488.820 2766.120 3491.550 2779.615 ;
        RECT 3487.520 2742.230 3491.550 2766.120 ;
        RECT 3483.975 2741.135 3491.550 2742.230 ;
        RECT 3513.135 2778.755 3518.355 2813.265 ;
        RECT 3513.135 2752.090 3517.315 2778.755 ;
      LAYER nwell ;
        RECT 3518.665 2772.960 3528.380 2819.415 ;
      LAYER pwell ;
        RECT 3513.135 2741.135 3518.355 2752.090 ;
        RECT 3483.975 2738.710 3518.355 2741.135 ;
      LAYER nwell ;
        RECT 3518.665 2738.560 3528.385 2772.960 ;
      LAYER pwell ;
        RECT 3528.685 2738.710 3532.565 2819.290 ;
      LAYER nwell ;
        RECT 3532.880 2812.615 3566.975 2819.415 ;
        RECT 3532.880 2740.370 3534.690 2812.615 ;
        RECT 3556.515 2811.485 3566.975 2812.615 ;
        RECT 3556.515 2752.030 3558.475 2811.485 ;
        RECT 3561.545 2752.030 3566.975 2811.485 ;
        RECT 3556.515 2740.370 3566.975 2752.030 ;
        RECT 3532.880 2738.565 3566.975 2740.370 ;
        RECT 3532.880 2738.560 3558.230 2738.565 ;
        RECT 29.770 2706.435 55.120 2706.440 ;
        RECT 21.025 2704.630 55.120 2706.435 ;
        RECT 21.025 2692.970 31.485 2704.630 ;
        RECT 21.025 2633.515 26.455 2692.970 ;
        RECT 29.525 2633.515 31.485 2692.970 ;
        RECT 21.025 2632.385 31.485 2633.515 ;
        RECT 53.310 2632.385 55.120 2704.630 ;
        RECT 21.025 2625.585 55.120 2632.385 ;
      LAYER pwell ;
        RECT 55.435 2625.710 59.315 2706.290 ;
      LAYER nwell ;
        RECT 59.615 2672.040 69.335 2706.440 ;
      LAYER pwell ;
        RECT 69.645 2703.865 104.025 2706.290 ;
        RECT 69.645 2692.910 74.865 2703.865 ;
      LAYER nwell ;
        RECT 59.620 2625.585 69.335 2672.040 ;
      LAYER pwell ;
        RECT 70.685 2666.245 74.865 2692.910 ;
        RECT 69.645 2631.735 74.865 2666.245 ;
        RECT 96.450 2702.770 104.025 2703.865 ;
        RECT 96.450 2678.880 100.480 2702.770 ;
        RECT 96.450 2665.385 99.180 2678.880 ;
        RECT 102.015 2671.840 104.025 2702.770 ;
      LAYER nwell ;
        RECT 104.835 2705.240 149.380 2706.670 ;
        RECT 104.835 2688.650 106.265 2705.240 ;
        RECT 104.835 2672.940 105.755 2688.650 ;
        RECT 115.655 2672.940 116.835 2705.240 ;
        RECT 126.225 2705.125 149.380 2705.240 ;
        RECT 126.225 2688.650 127.405 2705.125 ;
        RECT 133.955 2696.335 134.805 2705.125 ;
        RECT 147.950 2696.335 149.380 2705.125 ;
        RECT 126.735 2672.940 127.405 2688.650 ;
        RECT 163.945 2690.830 170.215 2706.450 ;
        RECT 174.655 2690.830 180.845 2706.450 ;
        RECT 163.945 2684.275 167.590 2690.830 ;
        RECT 163.945 2674.915 165.735 2684.275 ;
      LAYER pwell ;
        RECT 104.740 2671.840 105.045 2672.590 ;
        RECT 102.015 2665.385 105.045 2671.840 ;
        RECT 96.450 2631.735 98.035 2665.385 ;
        RECT 69.645 2631.215 98.035 2631.735 ;
        RECT 103.745 2635.300 105.045 2665.385 ;
        RECT 103.745 2631.215 107.065 2635.300 ;
      LAYER nwell ;
        RECT 112.260 2634.420 113.340 2634.495 ;
        RECT 111.720 2631.975 113.340 2634.420 ;
      LAYER pwell ;
        RECT 69.645 2625.785 107.065 2631.215 ;
      LAYER nwell ;
        RECT 108.180 2630.530 113.340 2631.975 ;
        RECT 108.180 2628.795 114.420 2630.530 ;
        RECT 107.600 2625.880 114.420 2628.795 ;
        RECT 118.765 2626.715 120.195 2650.815 ;
        RECT 138.980 2636.460 139.230 2639.535 ;
        RECT 138.980 2629.810 139.820 2636.460 ;
        RECT 137.660 2626.715 139.820 2629.810 ;
        RECT 141.980 2626.715 143.410 2649.515 ;
        RECT 176.920 2630.580 180.845 2690.830 ;
        RECT 107.600 2625.585 111.515 2625.880 ;
        RECT 118.765 2625.285 143.410 2626.715 ;
        RECT 190.675 2625.585 194.335 2629.110 ;
      LAYER pwell ;
        RECT 3388.935 2582.715 3411.790 2590.505 ;
      LAYER nwell ;
        RECT 3388.685 2523.035 3390.205 2582.140 ;
        RECT 197.795 2426.860 199.315 2485.965 ;
      LAYER pwell ;
        RECT 176.210 2418.495 199.065 2426.285 ;
      LAYER nwell ;
        RECT 3388.685 2082.035 3390.205 2141.140 ;
        RECT 29.770 2068.435 55.120 2068.440 ;
        RECT 21.025 2066.630 55.120 2068.435 ;
        RECT 21.025 2054.970 31.485 2066.630 ;
        RECT 21.025 1995.515 26.455 2054.970 ;
        RECT 29.525 1995.515 31.485 2054.970 ;
        RECT 21.025 1994.385 31.485 1995.515 ;
        RECT 53.310 1994.385 55.120 2066.630 ;
        RECT 21.025 1987.585 55.120 1994.385 ;
      LAYER pwell ;
        RECT 55.435 1987.710 59.315 2068.290 ;
      LAYER nwell ;
        RECT 59.615 2034.040 69.335 2068.440 ;
      LAYER pwell ;
        RECT 69.645 2065.865 104.025 2068.290 ;
        RECT 69.645 2054.910 74.865 2065.865 ;
      LAYER nwell ;
        RECT 59.620 1987.585 69.335 2034.040 ;
      LAYER pwell ;
        RECT 70.685 2028.245 74.865 2054.910 ;
        RECT 69.645 1993.735 74.865 2028.245 ;
        RECT 96.450 2064.770 104.025 2065.865 ;
        RECT 96.450 2040.880 100.480 2064.770 ;
        RECT 96.450 2027.385 99.180 2040.880 ;
        RECT 102.015 2033.840 104.025 2064.770 ;
      LAYER nwell ;
        RECT 104.835 2067.240 149.380 2068.670 ;
        RECT 104.835 2050.650 106.265 2067.240 ;
        RECT 104.835 2034.940 105.755 2050.650 ;
        RECT 115.655 2034.940 116.835 2067.240 ;
        RECT 126.225 2067.125 149.380 2067.240 ;
        RECT 126.225 2050.650 127.405 2067.125 ;
        RECT 133.955 2058.335 134.805 2067.125 ;
        RECT 147.950 2058.335 149.380 2067.125 ;
        RECT 126.735 2034.940 127.405 2050.650 ;
        RECT 163.945 2052.830 170.215 2068.450 ;
        RECT 174.655 2052.830 180.845 2068.450 ;
        RECT 163.945 2046.275 167.590 2052.830 ;
        RECT 163.945 2036.915 165.735 2046.275 ;
      LAYER pwell ;
        RECT 104.740 2033.840 105.045 2034.590 ;
        RECT 102.015 2027.385 105.045 2033.840 ;
        RECT 96.450 1993.735 98.035 2027.385 ;
        RECT 69.645 1993.215 98.035 1993.735 ;
        RECT 103.745 1997.300 105.045 2027.385 ;
        RECT 103.745 1993.215 107.065 1997.300 ;
      LAYER nwell ;
        RECT 112.260 1996.420 113.340 1996.495 ;
        RECT 111.720 1993.975 113.340 1996.420 ;
      LAYER pwell ;
        RECT 69.645 1987.785 107.065 1993.215 ;
      LAYER nwell ;
        RECT 108.180 1992.530 113.340 1993.975 ;
        RECT 108.180 1990.795 114.420 1992.530 ;
        RECT 107.600 1987.880 114.420 1990.795 ;
        RECT 118.765 1988.715 120.195 2012.815 ;
        RECT 138.980 1998.460 139.230 2001.535 ;
        RECT 138.980 1991.810 139.820 1998.460 ;
        RECT 137.660 1988.715 139.820 1991.810 ;
        RECT 141.980 1988.715 143.410 2011.515 ;
        RECT 176.920 1992.580 180.845 2052.830 ;
        RECT 107.600 1987.585 111.515 1987.880 ;
        RECT 118.765 1987.285 143.410 1988.715 ;
        RECT 190.675 1987.585 194.335 1991.110 ;
        RECT 3393.665 1929.890 3397.325 1933.415 ;
        RECT 3444.590 1932.285 3469.235 1933.715 ;
        RECT 3476.485 1933.120 3480.400 1933.415 ;
        RECT 3407.155 1868.170 3411.080 1928.420 ;
        RECT 3444.590 1909.485 3446.020 1932.285 ;
        RECT 3448.180 1929.190 3450.340 1932.285 ;
        RECT 3448.180 1922.540 3449.020 1929.190 ;
        RECT 3448.770 1919.465 3449.020 1922.540 ;
        RECT 3467.805 1908.185 3469.235 1932.285 ;
        RECT 3473.580 1930.205 3480.400 1933.120 ;
        RECT 3473.580 1928.470 3479.820 1930.205 ;
        RECT 3474.660 1927.025 3479.820 1928.470 ;
      LAYER pwell ;
        RECT 3480.935 1927.785 3518.355 1933.215 ;
      LAYER nwell ;
        RECT 3474.660 1924.580 3476.280 1927.025 ;
        RECT 3474.660 1924.505 3475.740 1924.580 ;
      LAYER pwell ;
        RECT 3480.935 1923.700 3484.255 1927.785 ;
        RECT 3482.955 1893.615 3484.255 1923.700 ;
        RECT 3489.965 1927.265 3518.355 1927.785 ;
        RECT 3489.965 1893.615 3491.550 1927.265 ;
        RECT 3482.955 1887.160 3485.985 1893.615 ;
        RECT 3482.955 1886.410 3483.260 1887.160 ;
      LAYER nwell ;
        RECT 3422.265 1874.725 3424.055 1884.085 ;
        RECT 3420.410 1868.170 3424.055 1874.725 ;
        RECT 29.770 1852.435 55.120 1852.440 ;
        RECT 21.025 1850.630 55.120 1852.435 ;
        RECT 21.025 1838.970 31.485 1850.630 ;
        RECT 21.025 1779.515 26.455 1838.970 ;
        RECT 29.525 1779.515 31.485 1838.970 ;
        RECT 21.025 1778.385 31.485 1779.515 ;
        RECT 53.310 1778.385 55.120 1850.630 ;
        RECT 21.025 1771.585 55.120 1778.385 ;
      LAYER pwell ;
        RECT 55.435 1771.710 59.315 1852.290 ;
      LAYER nwell ;
        RECT 59.615 1818.040 69.335 1852.440 ;
      LAYER pwell ;
        RECT 69.645 1849.865 104.025 1852.290 ;
        RECT 69.645 1838.910 74.865 1849.865 ;
      LAYER nwell ;
        RECT 59.620 1771.585 69.335 1818.040 ;
      LAYER pwell ;
        RECT 70.685 1812.245 74.865 1838.910 ;
        RECT 69.645 1777.735 74.865 1812.245 ;
        RECT 96.450 1848.770 104.025 1849.865 ;
        RECT 96.450 1824.880 100.480 1848.770 ;
        RECT 96.450 1811.385 99.180 1824.880 ;
        RECT 102.015 1817.840 104.025 1848.770 ;
      LAYER nwell ;
        RECT 104.835 1851.240 149.380 1852.670 ;
        RECT 3407.155 1852.550 3413.345 1868.170 ;
        RECT 3417.785 1852.550 3424.055 1868.170 ;
        RECT 3460.595 1870.350 3461.265 1886.060 ;
        RECT 3438.620 1853.875 3440.050 1862.665 ;
        RECT 3453.195 1853.875 3454.045 1862.665 ;
        RECT 3460.595 1853.875 3461.775 1870.350 ;
        RECT 3438.620 1853.760 3461.775 1853.875 ;
        RECT 3471.165 1853.760 3472.345 1886.060 ;
        RECT 3482.245 1870.350 3483.165 1886.060 ;
        RECT 3481.735 1853.760 3483.165 1870.350 ;
        RECT 104.835 1834.650 106.265 1851.240 ;
        RECT 104.835 1818.940 105.755 1834.650 ;
        RECT 115.655 1818.940 116.835 1851.240 ;
        RECT 126.225 1851.125 149.380 1851.240 ;
        RECT 126.225 1834.650 127.405 1851.125 ;
        RECT 133.955 1842.335 134.805 1851.125 ;
        RECT 147.950 1842.335 149.380 1851.125 ;
        RECT 126.735 1818.940 127.405 1834.650 ;
        RECT 163.945 1836.830 170.215 1852.450 ;
        RECT 174.655 1836.830 180.845 1852.450 ;
        RECT 3438.620 1852.330 3483.165 1853.760 ;
      LAYER pwell ;
        RECT 3483.975 1856.230 3485.985 1887.160 ;
        RECT 3488.820 1880.120 3491.550 1893.615 ;
        RECT 3487.520 1856.230 3491.550 1880.120 ;
        RECT 3483.975 1855.135 3491.550 1856.230 ;
        RECT 3513.135 1892.755 3518.355 1927.265 ;
        RECT 3513.135 1866.090 3517.315 1892.755 ;
      LAYER nwell ;
        RECT 3518.665 1886.960 3528.380 1933.415 ;
      LAYER pwell ;
        RECT 3513.135 1855.135 3518.355 1866.090 ;
        RECT 3483.975 1852.710 3518.355 1855.135 ;
      LAYER nwell ;
        RECT 3518.665 1852.560 3528.385 1886.960 ;
      LAYER pwell ;
        RECT 3528.685 1852.710 3532.565 1933.290 ;
      LAYER nwell ;
        RECT 3532.880 1926.615 3566.975 1933.415 ;
        RECT 3532.880 1854.370 3534.690 1926.615 ;
        RECT 3556.515 1925.485 3566.975 1926.615 ;
        RECT 3556.515 1866.030 3558.475 1925.485 ;
        RECT 3561.545 1866.030 3566.975 1925.485 ;
        RECT 3556.515 1854.370 3566.975 1866.030 ;
        RECT 3532.880 1852.565 3566.975 1854.370 ;
        RECT 3532.880 1852.560 3558.230 1852.565 ;
        RECT 163.945 1830.275 167.590 1836.830 ;
        RECT 163.945 1820.915 165.735 1830.275 ;
      LAYER pwell ;
        RECT 104.740 1817.840 105.045 1818.590 ;
        RECT 102.015 1811.385 105.045 1817.840 ;
        RECT 96.450 1777.735 98.035 1811.385 ;
        RECT 69.645 1777.215 98.035 1777.735 ;
        RECT 103.745 1781.300 105.045 1811.385 ;
        RECT 103.745 1777.215 107.065 1781.300 ;
      LAYER nwell ;
        RECT 112.260 1780.420 113.340 1780.495 ;
        RECT 111.720 1777.975 113.340 1780.420 ;
      LAYER pwell ;
        RECT 69.645 1771.785 107.065 1777.215 ;
      LAYER nwell ;
        RECT 108.180 1776.530 113.340 1777.975 ;
        RECT 108.180 1774.795 114.420 1776.530 ;
        RECT 107.600 1771.880 114.420 1774.795 ;
        RECT 118.765 1772.715 120.195 1796.815 ;
        RECT 138.980 1782.460 139.230 1785.535 ;
        RECT 138.980 1775.810 139.820 1782.460 ;
        RECT 137.660 1772.715 139.820 1775.810 ;
        RECT 141.980 1772.715 143.410 1795.515 ;
        RECT 176.920 1776.580 180.845 1836.830 ;
        RECT 107.600 1771.585 111.515 1771.880 ;
        RECT 118.765 1771.285 143.410 1772.715 ;
        RECT 190.675 1771.585 194.335 1775.110 ;
        RECT 3393.665 1703.890 3397.325 1707.415 ;
        RECT 3444.590 1706.285 3469.235 1707.715 ;
        RECT 3476.485 1707.120 3480.400 1707.415 ;
        RECT 3407.155 1642.170 3411.080 1702.420 ;
        RECT 3444.590 1683.485 3446.020 1706.285 ;
        RECT 3448.180 1703.190 3450.340 1706.285 ;
        RECT 3448.180 1696.540 3449.020 1703.190 ;
        RECT 3448.770 1693.465 3449.020 1696.540 ;
        RECT 3467.805 1682.185 3469.235 1706.285 ;
        RECT 3473.580 1704.205 3480.400 1707.120 ;
        RECT 3473.580 1702.470 3479.820 1704.205 ;
        RECT 3474.660 1701.025 3479.820 1702.470 ;
      LAYER pwell ;
        RECT 3480.935 1701.785 3518.355 1707.215 ;
      LAYER nwell ;
        RECT 3474.660 1698.580 3476.280 1701.025 ;
        RECT 3474.660 1698.505 3475.740 1698.580 ;
      LAYER pwell ;
        RECT 3480.935 1697.700 3484.255 1701.785 ;
        RECT 3482.955 1667.615 3484.255 1697.700 ;
        RECT 3489.965 1701.265 3518.355 1701.785 ;
        RECT 3489.965 1667.615 3491.550 1701.265 ;
        RECT 3482.955 1661.160 3485.985 1667.615 ;
        RECT 3482.955 1660.410 3483.260 1661.160 ;
      LAYER nwell ;
        RECT 3422.265 1648.725 3424.055 1658.085 ;
        RECT 3420.410 1642.170 3424.055 1648.725 ;
        RECT 29.770 1636.435 55.120 1636.440 ;
        RECT 21.025 1634.630 55.120 1636.435 ;
        RECT 21.025 1622.970 31.485 1634.630 ;
        RECT 21.025 1563.515 26.455 1622.970 ;
        RECT 29.525 1563.515 31.485 1622.970 ;
        RECT 21.025 1562.385 31.485 1563.515 ;
        RECT 53.310 1562.385 55.120 1634.630 ;
        RECT 21.025 1555.585 55.120 1562.385 ;
      LAYER pwell ;
        RECT 55.435 1555.710 59.315 1636.290 ;
      LAYER nwell ;
        RECT 59.615 1602.040 69.335 1636.440 ;
      LAYER pwell ;
        RECT 69.645 1633.865 104.025 1636.290 ;
        RECT 69.645 1622.910 74.865 1633.865 ;
      LAYER nwell ;
        RECT 59.620 1555.585 69.335 1602.040 ;
      LAYER pwell ;
        RECT 70.685 1596.245 74.865 1622.910 ;
        RECT 69.645 1561.735 74.865 1596.245 ;
        RECT 96.450 1632.770 104.025 1633.865 ;
        RECT 96.450 1608.880 100.480 1632.770 ;
        RECT 96.450 1595.385 99.180 1608.880 ;
        RECT 102.015 1601.840 104.025 1632.770 ;
      LAYER nwell ;
        RECT 104.835 1635.240 149.380 1636.670 ;
        RECT 104.835 1618.650 106.265 1635.240 ;
        RECT 104.835 1602.940 105.755 1618.650 ;
        RECT 115.655 1602.940 116.835 1635.240 ;
        RECT 126.225 1635.125 149.380 1635.240 ;
        RECT 126.225 1618.650 127.405 1635.125 ;
        RECT 133.955 1626.335 134.805 1635.125 ;
        RECT 147.950 1626.335 149.380 1635.125 ;
        RECT 126.735 1602.940 127.405 1618.650 ;
        RECT 163.945 1620.830 170.215 1636.450 ;
        RECT 174.655 1620.830 180.845 1636.450 ;
        RECT 3407.155 1626.550 3413.345 1642.170 ;
        RECT 3417.785 1626.550 3424.055 1642.170 ;
        RECT 3460.595 1644.350 3461.265 1660.060 ;
        RECT 3438.620 1627.875 3440.050 1636.665 ;
        RECT 3453.195 1627.875 3454.045 1636.665 ;
        RECT 3460.595 1627.875 3461.775 1644.350 ;
        RECT 3438.620 1627.760 3461.775 1627.875 ;
        RECT 3471.165 1627.760 3472.345 1660.060 ;
        RECT 3482.245 1644.350 3483.165 1660.060 ;
        RECT 3481.735 1627.760 3483.165 1644.350 ;
        RECT 3438.620 1626.330 3483.165 1627.760 ;
      LAYER pwell ;
        RECT 3483.975 1630.230 3485.985 1661.160 ;
        RECT 3488.820 1654.120 3491.550 1667.615 ;
        RECT 3487.520 1630.230 3491.550 1654.120 ;
        RECT 3483.975 1629.135 3491.550 1630.230 ;
        RECT 3513.135 1666.755 3518.355 1701.265 ;
        RECT 3513.135 1640.090 3517.315 1666.755 ;
      LAYER nwell ;
        RECT 3518.665 1660.960 3528.380 1707.415 ;
      LAYER pwell ;
        RECT 3513.135 1629.135 3518.355 1640.090 ;
        RECT 3483.975 1626.710 3518.355 1629.135 ;
      LAYER nwell ;
        RECT 3518.665 1626.560 3528.385 1660.960 ;
      LAYER pwell ;
        RECT 3528.685 1626.710 3532.565 1707.290 ;
      LAYER nwell ;
        RECT 3532.880 1700.615 3566.975 1707.415 ;
        RECT 3532.880 1628.370 3534.690 1700.615 ;
        RECT 3556.515 1699.485 3566.975 1700.615 ;
        RECT 3556.515 1640.030 3558.475 1699.485 ;
        RECT 3561.545 1640.030 3566.975 1699.485 ;
        RECT 3556.515 1628.370 3566.975 1640.030 ;
        RECT 3532.880 1626.565 3566.975 1628.370 ;
        RECT 3532.880 1626.560 3558.230 1626.565 ;
        RECT 163.945 1614.275 167.590 1620.830 ;
        RECT 163.945 1604.915 165.735 1614.275 ;
      LAYER pwell ;
        RECT 104.740 1601.840 105.045 1602.590 ;
        RECT 102.015 1595.385 105.045 1601.840 ;
        RECT 96.450 1561.735 98.035 1595.385 ;
        RECT 69.645 1561.215 98.035 1561.735 ;
        RECT 103.745 1565.300 105.045 1595.385 ;
        RECT 103.745 1561.215 107.065 1565.300 ;
      LAYER nwell ;
        RECT 112.260 1564.420 113.340 1564.495 ;
        RECT 111.720 1561.975 113.340 1564.420 ;
      LAYER pwell ;
        RECT 69.645 1555.785 107.065 1561.215 ;
      LAYER nwell ;
        RECT 108.180 1560.530 113.340 1561.975 ;
        RECT 108.180 1558.795 114.420 1560.530 ;
        RECT 107.600 1555.880 114.420 1558.795 ;
        RECT 118.765 1556.715 120.195 1580.815 ;
        RECT 138.980 1566.460 139.230 1569.535 ;
        RECT 138.980 1559.810 139.820 1566.460 ;
        RECT 137.660 1556.715 139.820 1559.810 ;
        RECT 141.980 1556.715 143.410 1579.515 ;
        RECT 176.920 1560.580 180.845 1620.830 ;
        RECT 107.600 1555.585 111.515 1555.880 ;
        RECT 118.765 1555.285 143.410 1556.715 ;
        RECT 190.675 1555.585 194.335 1559.110 ;
        RECT 3393.665 1478.890 3397.325 1482.415 ;
        RECT 3444.590 1481.285 3469.235 1482.715 ;
        RECT 3476.485 1482.120 3480.400 1482.415 ;
        RECT 29.770 1420.435 55.120 1420.440 ;
        RECT 21.025 1418.630 55.120 1420.435 ;
        RECT 21.025 1406.970 31.485 1418.630 ;
        RECT 21.025 1347.515 26.455 1406.970 ;
        RECT 29.525 1347.515 31.485 1406.970 ;
        RECT 21.025 1346.385 31.485 1347.515 ;
        RECT 53.310 1346.385 55.120 1418.630 ;
        RECT 21.025 1339.585 55.120 1346.385 ;
      LAYER pwell ;
        RECT 55.435 1339.710 59.315 1420.290 ;
      LAYER nwell ;
        RECT 59.615 1386.040 69.335 1420.440 ;
      LAYER pwell ;
        RECT 69.645 1417.865 104.025 1420.290 ;
        RECT 69.645 1406.910 74.865 1417.865 ;
      LAYER nwell ;
        RECT 59.620 1339.585 69.335 1386.040 ;
      LAYER pwell ;
        RECT 70.685 1380.245 74.865 1406.910 ;
        RECT 69.645 1345.735 74.865 1380.245 ;
        RECT 96.450 1416.770 104.025 1417.865 ;
        RECT 96.450 1392.880 100.480 1416.770 ;
        RECT 96.450 1379.385 99.180 1392.880 ;
        RECT 102.015 1385.840 104.025 1416.770 ;
      LAYER nwell ;
        RECT 104.835 1419.240 149.380 1420.670 ;
        RECT 104.835 1402.650 106.265 1419.240 ;
        RECT 104.835 1386.940 105.755 1402.650 ;
        RECT 115.655 1386.940 116.835 1419.240 ;
        RECT 126.225 1419.125 149.380 1419.240 ;
        RECT 126.225 1402.650 127.405 1419.125 ;
        RECT 133.955 1410.335 134.805 1419.125 ;
        RECT 147.950 1410.335 149.380 1419.125 ;
        RECT 126.735 1386.940 127.405 1402.650 ;
        RECT 163.945 1404.830 170.215 1420.450 ;
        RECT 174.655 1404.830 180.845 1420.450 ;
        RECT 163.945 1398.275 167.590 1404.830 ;
        RECT 163.945 1388.915 165.735 1398.275 ;
      LAYER pwell ;
        RECT 104.740 1385.840 105.045 1386.590 ;
        RECT 102.015 1379.385 105.045 1385.840 ;
        RECT 96.450 1345.735 98.035 1379.385 ;
        RECT 69.645 1345.215 98.035 1345.735 ;
        RECT 103.745 1349.300 105.045 1379.385 ;
        RECT 103.745 1345.215 107.065 1349.300 ;
      LAYER nwell ;
        RECT 112.260 1348.420 113.340 1348.495 ;
        RECT 111.720 1345.975 113.340 1348.420 ;
      LAYER pwell ;
        RECT 69.645 1339.785 107.065 1345.215 ;
      LAYER nwell ;
        RECT 108.180 1344.530 113.340 1345.975 ;
        RECT 108.180 1342.795 114.420 1344.530 ;
        RECT 107.600 1339.880 114.420 1342.795 ;
        RECT 118.765 1340.715 120.195 1364.815 ;
        RECT 138.980 1350.460 139.230 1353.535 ;
        RECT 138.980 1343.810 139.820 1350.460 ;
        RECT 137.660 1340.715 139.820 1343.810 ;
        RECT 141.980 1340.715 143.410 1363.515 ;
        RECT 176.920 1344.580 180.845 1404.830 ;
        RECT 3407.155 1417.170 3411.080 1477.420 ;
        RECT 3444.590 1458.485 3446.020 1481.285 ;
        RECT 3448.180 1478.190 3450.340 1481.285 ;
        RECT 3448.180 1471.540 3449.020 1478.190 ;
        RECT 3448.770 1468.465 3449.020 1471.540 ;
        RECT 3467.805 1457.185 3469.235 1481.285 ;
        RECT 3473.580 1479.205 3480.400 1482.120 ;
        RECT 3473.580 1477.470 3479.820 1479.205 ;
        RECT 3474.660 1476.025 3479.820 1477.470 ;
      LAYER pwell ;
        RECT 3480.935 1476.785 3518.355 1482.215 ;
      LAYER nwell ;
        RECT 3474.660 1473.580 3476.280 1476.025 ;
        RECT 3474.660 1473.505 3475.740 1473.580 ;
      LAYER pwell ;
        RECT 3480.935 1472.700 3484.255 1476.785 ;
        RECT 3482.955 1442.615 3484.255 1472.700 ;
        RECT 3489.965 1476.265 3518.355 1476.785 ;
        RECT 3489.965 1442.615 3491.550 1476.265 ;
        RECT 3482.955 1436.160 3485.985 1442.615 ;
        RECT 3482.955 1435.410 3483.260 1436.160 ;
      LAYER nwell ;
        RECT 3422.265 1423.725 3424.055 1433.085 ;
        RECT 3420.410 1417.170 3424.055 1423.725 ;
        RECT 3407.155 1401.550 3413.345 1417.170 ;
        RECT 3417.785 1401.550 3424.055 1417.170 ;
        RECT 3460.595 1419.350 3461.265 1435.060 ;
        RECT 3438.620 1402.875 3440.050 1411.665 ;
        RECT 3453.195 1402.875 3454.045 1411.665 ;
        RECT 3460.595 1402.875 3461.775 1419.350 ;
        RECT 3438.620 1402.760 3461.775 1402.875 ;
        RECT 3471.165 1402.760 3472.345 1435.060 ;
        RECT 3482.245 1419.350 3483.165 1435.060 ;
        RECT 3481.735 1402.760 3483.165 1419.350 ;
        RECT 3438.620 1401.330 3483.165 1402.760 ;
      LAYER pwell ;
        RECT 3483.975 1405.230 3485.985 1436.160 ;
        RECT 3488.820 1429.120 3491.550 1442.615 ;
        RECT 3487.520 1405.230 3491.550 1429.120 ;
        RECT 3483.975 1404.135 3491.550 1405.230 ;
        RECT 3513.135 1441.755 3518.355 1476.265 ;
        RECT 3513.135 1415.090 3517.315 1441.755 ;
      LAYER nwell ;
        RECT 3518.665 1435.960 3528.380 1482.415 ;
      LAYER pwell ;
        RECT 3513.135 1404.135 3518.355 1415.090 ;
        RECT 3483.975 1401.710 3518.355 1404.135 ;
      LAYER nwell ;
        RECT 3518.665 1401.560 3528.385 1435.960 ;
      LAYER pwell ;
        RECT 3528.685 1401.710 3532.565 1482.290 ;
      LAYER nwell ;
        RECT 3532.880 1475.615 3566.975 1482.415 ;
        RECT 3532.880 1403.370 3534.690 1475.615 ;
        RECT 3556.515 1474.485 3566.975 1475.615 ;
        RECT 3556.515 1415.030 3558.475 1474.485 ;
        RECT 3561.545 1415.030 3566.975 1474.485 ;
        RECT 3556.515 1403.370 3566.975 1415.030 ;
        RECT 3532.880 1401.565 3566.975 1403.370 ;
        RECT 3532.880 1401.560 3558.230 1401.565 ;
        RECT 107.600 1339.585 111.515 1339.880 ;
        RECT 118.765 1339.285 143.410 1340.715 ;
        RECT 190.675 1339.585 194.335 1343.110 ;
        RECT 3393.665 1253.890 3397.325 1257.415 ;
        RECT 3444.590 1256.285 3469.235 1257.715 ;
        RECT 3476.485 1257.120 3480.400 1257.415 ;
        RECT 29.770 1204.435 55.120 1204.440 ;
        RECT 21.025 1202.630 55.120 1204.435 ;
        RECT 21.025 1190.970 31.485 1202.630 ;
        RECT 21.025 1131.515 26.455 1190.970 ;
        RECT 29.525 1131.515 31.485 1190.970 ;
        RECT 21.025 1130.385 31.485 1131.515 ;
        RECT 53.310 1130.385 55.120 1202.630 ;
        RECT 21.025 1123.585 55.120 1130.385 ;
      LAYER pwell ;
        RECT 55.435 1123.710 59.315 1204.290 ;
      LAYER nwell ;
        RECT 59.615 1170.040 69.335 1204.440 ;
      LAYER pwell ;
        RECT 69.645 1201.865 104.025 1204.290 ;
        RECT 69.645 1190.910 74.865 1201.865 ;
      LAYER nwell ;
        RECT 59.620 1123.585 69.335 1170.040 ;
      LAYER pwell ;
        RECT 70.685 1164.245 74.865 1190.910 ;
        RECT 69.645 1129.735 74.865 1164.245 ;
        RECT 96.450 1200.770 104.025 1201.865 ;
        RECT 96.450 1176.880 100.480 1200.770 ;
        RECT 96.450 1163.385 99.180 1176.880 ;
        RECT 102.015 1169.840 104.025 1200.770 ;
      LAYER nwell ;
        RECT 104.835 1203.240 149.380 1204.670 ;
        RECT 104.835 1186.650 106.265 1203.240 ;
        RECT 104.835 1170.940 105.755 1186.650 ;
        RECT 115.655 1170.940 116.835 1203.240 ;
        RECT 126.225 1203.125 149.380 1203.240 ;
        RECT 126.225 1186.650 127.405 1203.125 ;
        RECT 133.955 1194.335 134.805 1203.125 ;
        RECT 147.950 1194.335 149.380 1203.125 ;
        RECT 126.735 1170.940 127.405 1186.650 ;
        RECT 163.945 1188.830 170.215 1204.450 ;
        RECT 174.655 1188.830 180.845 1204.450 ;
        RECT 163.945 1182.275 167.590 1188.830 ;
        RECT 163.945 1172.915 165.735 1182.275 ;
      LAYER pwell ;
        RECT 104.740 1169.840 105.045 1170.590 ;
        RECT 102.015 1163.385 105.045 1169.840 ;
        RECT 96.450 1129.735 98.035 1163.385 ;
        RECT 69.645 1129.215 98.035 1129.735 ;
        RECT 103.745 1133.300 105.045 1163.385 ;
        RECT 103.745 1129.215 107.065 1133.300 ;
      LAYER nwell ;
        RECT 112.260 1132.420 113.340 1132.495 ;
        RECT 111.720 1129.975 113.340 1132.420 ;
      LAYER pwell ;
        RECT 69.645 1123.785 107.065 1129.215 ;
      LAYER nwell ;
        RECT 108.180 1128.530 113.340 1129.975 ;
        RECT 108.180 1126.795 114.420 1128.530 ;
        RECT 107.600 1123.880 114.420 1126.795 ;
        RECT 118.765 1124.715 120.195 1148.815 ;
        RECT 138.980 1134.460 139.230 1137.535 ;
        RECT 138.980 1127.810 139.820 1134.460 ;
        RECT 137.660 1124.715 139.820 1127.810 ;
        RECT 141.980 1124.715 143.410 1147.515 ;
        RECT 176.920 1128.580 180.845 1188.830 ;
        RECT 3407.155 1192.170 3411.080 1252.420 ;
        RECT 3444.590 1233.485 3446.020 1256.285 ;
        RECT 3448.180 1253.190 3450.340 1256.285 ;
        RECT 3448.180 1246.540 3449.020 1253.190 ;
        RECT 3448.770 1243.465 3449.020 1246.540 ;
        RECT 3467.805 1232.185 3469.235 1256.285 ;
        RECT 3473.580 1254.205 3480.400 1257.120 ;
        RECT 3473.580 1252.470 3479.820 1254.205 ;
        RECT 3474.660 1251.025 3479.820 1252.470 ;
      LAYER pwell ;
        RECT 3480.935 1251.785 3518.355 1257.215 ;
      LAYER nwell ;
        RECT 3474.660 1248.580 3476.280 1251.025 ;
        RECT 3474.660 1248.505 3475.740 1248.580 ;
      LAYER pwell ;
        RECT 3480.935 1247.700 3484.255 1251.785 ;
        RECT 3482.955 1217.615 3484.255 1247.700 ;
        RECT 3489.965 1251.265 3518.355 1251.785 ;
        RECT 3489.965 1217.615 3491.550 1251.265 ;
        RECT 3482.955 1211.160 3485.985 1217.615 ;
        RECT 3482.955 1210.410 3483.260 1211.160 ;
      LAYER nwell ;
        RECT 3422.265 1198.725 3424.055 1208.085 ;
        RECT 3420.410 1192.170 3424.055 1198.725 ;
        RECT 3407.155 1176.550 3413.345 1192.170 ;
        RECT 3417.785 1176.550 3424.055 1192.170 ;
        RECT 3460.595 1194.350 3461.265 1210.060 ;
        RECT 3438.620 1177.875 3440.050 1186.665 ;
        RECT 3453.195 1177.875 3454.045 1186.665 ;
        RECT 3460.595 1177.875 3461.775 1194.350 ;
        RECT 3438.620 1177.760 3461.775 1177.875 ;
        RECT 3471.165 1177.760 3472.345 1210.060 ;
        RECT 3482.245 1194.350 3483.165 1210.060 ;
        RECT 3481.735 1177.760 3483.165 1194.350 ;
        RECT 3438.620 1176.330 3483.165 1177.760 ;
      LAYER pwell ;
        RECT 3483.975 1180.230 3485.985 1211.160 ;
        RECT 3488.820 1204.120 3491.550 1217.615 ;
        RECT 3487.520 1180.230 3491.550 1204.120 ;
        RECT 3483.975 1179.135 3491.550 1180.230 ;
        RECT 3513.135 1216.755 3518.355 1251.265 ;
        RECT 3513.135 1190.090 3517.315 1216.755 ;
      LAYER nwell ;
        RECT 3518.665 1210.960 3528.380 1257.415 ;
      LAYER pwell ;
        RECT 3513.135 1179.135 3518.355 1190.090 ;
        RECT 3483.975 1176.710 3518.355 1179.135 ;
      LAYER nwell ;
        RECT 3518.665 1176.560 3528.385 1210.960 ;
      LAYER pwell ;
        RECT 3528.685 1176.710 3532.565 1257.290 ;
      LAYER nwell ;
        RECT 3532.880 1250.615 3566.975 1257.415 ;
        RECT 3532.880 1178.370 3534.690 1250.615 ;
        RECT 3556.515 1249.485 3566.975 1250.615 ;
        RECT 3556.515 1190.030 3558.475 1249.485 ;
        RECT 3561.545 1190.030 3566.975 1249.485 ;
        RECT 3556.515 1178.370 3566.975 1190.030 ;
        RECT 3532.880 1176.565 3566.975 1178.370 ;
        RECT 3532.880 1176.560 3558.230 1176.565 ;
        RECT 107.600 1123.585 111.515 1123.880 ;
        RECT 118.765 1123.285 143.410 1124.715 ;
        RECT 190.675 1123.585 194.335 1127.110 ;
        RECT 3393.665 1027.890 3397.325 1031.415 ;
        RECT 3444.590 1030.285 3469.235 1031.715 ;
        RECT 3476.485 1031.120 3480.400 1031.415 ;
        RECT 29.770 988.435 55.120 988.440 ;
        RECT 21.025 986.630 55.120 988.435 ;
        RECT 21.025 974.970 31.485 986.630 ;
        RECT 21.025 915.515 26.455 974.970 ;
        RECT 29.525 915.515 31.485 974.970 ;
        RECT 21.025 914.385 31.485 915.515 ;
        RECT 53.310 914.385 55.120 986.630 ;
        RECT 21.025 907.585 55.120 914.385 ;
      LAYER pwell ;
        RECT 55.435 907.710 59.315 988.290 ;
      LAYER nwell ;
        RECT 59.615 954.040 69.335 988.440 ;
      LAYER pwell ;
        RECT 69.645 985.865 104.025 988.290 ;
        RECT 69.645 974.910 74.865 985.865 ;
      LAYER nwell ;
        RECT 59.620 907.585 69.335 954.040 ;
      LAYER pwell ;
        RECT 70.685 948.245 74.865 974.910 ;
        RECT 69.645 913.735 74.865 948.245 ;
        RECT 96.450 984.770 104.025 985.865 ;
        RECT 96.450 960.880 100.480 984.770 ;
        RECT 96.450 947.385 99.180 960.880 ;
        RECT 102.015 953.840 104.025 984.770 ;
      LAYER nwell ;
        RECT 104.835 987.240 149.380 988.670 ;
        RECT 104.835 970.650 106.265 987.240 ;
        RECT 104.835 954.940 105.755 970.650 ;
        RECT 115.655 954.940 116.835 987.240 ;
        RECT 126.225 987.125 149.380 987.240 ;
        RECT 126.225 970.650 127.405 987.125 ;
        RECT 133.955 978.335 134.805 987.125 ;
        RECT 147.950 978.335 149.380 987.125 ;
        RECT 126.735 954.940 127.405 970.650 ;
        RECT 163.945 972.830 170.215 988.450 ;
        RECT 174.655 972.830 180.845 988.450 ;
        RECT 163.945 966.275 167.590 972.830 ;
        RECT 163.945 956.915 165.735 966.275 ;
      LAYER pwell ;
        RECT 104.740 953.840 105.045 954.590 ;
        RECT 102.015 947.385 105.045 953.840 ;
        RECT 96.450 913.735 98.035 947.385 ;
        RECT 69.645 913.215 98.035 913.735 ;
        RECT 103.745 917.300 105.045 947.385 ;
        RECT 103.745 913.215 107.065 917.300 ;
      LAYER nwell ;
        RECT 112.260 916.420 113.340 916.495 ;
        RECT 111.720 913.975 113.340 916.420 ;
      LAYER pwell ;
        RECT 69.645 907.785 107.065 913.215 ;
      LAYER nwell ;
        RECT 108.180 912.530 113.340 913.975 ;
        RECT 108.180 910.795 114.420 912.530 ;
        RECT 107.600 907.880 114.420 910.795 ;
        RECT 118.765 908.715 120.195 932.815 ;
        RECT 138.980 918.460 139.230 921.535 ;
        RECT 138.980 911.810 139.820 918.460 ;
        RECT 137.660 908.715 139.820 911.810 ;
        RECT 141.980 908.715 143.410 931.515 ;
        RECT 176.920 912.580 180.845 972.830 ;
        RECT 3407.155 966.170 3411.080 1026.420 ;
        RECT 3444.590 1007.485 3446.020 1030.285 ;
        RECT 3448.180 1027.190 3450.340 1030.285 ;
        RECT 3448.180 1020.540 3449.020 1027.190 ;
        RECT 3448.770 1017.465 3449.020 1020.540 ;
        RECT 3467.805 1006.185 3469.235 1030.285 ;
        RECT 3473.580 1028.205 3480.400 1031.120 ;
        RECT 3473.580 1026.470 3479.820 1028.205 ;
        RECT 3474.660 1025.025 3479.820 1026.470 ;
      LAYER pwell ;
        RECT 3480.935 1025.785 3518.355 1031.215 ;
      LAYER nwell ;
        RECT 3474.660 1022.580 3476.280 1025.025 ;
        RECT 3474.660 1022.505 3475.740 1022.580 ;
      LAYER pwell ;
        RECT 3480.935 1021.700 3484.255 1025.785 ;
        RECT 3482.955 991.615 3484.255 1021.700 ;
        RECT 3489.965 1025.265 3518.355 1025.785 ;
        RECT 3489.965 991.615 3491.550 1025.265 ;
        RECT 3482.955 985.160 3485.985 991.615 ;
        RECT 3482.955 984.410 3483.260 985.160 ;
      LAYER nwell ;
        RECT 3422.265 972.725 3424.055 982.085 ;
        RECT 3420.410 966.170 3424.055 972.725 ;
        RECT 3407.155 950.550 3413.345 966.170 ;
        RECT 3417.785 950.550 3424.055 966.170 ;
        RECT 3460.595 968.350 3461.265 984.060 ;
        RECT 3438.620 951.875 3440.050 960.665 ;
        RECT 3453.195 951.875 3454.045 960.665 ;
        RECT 3460.595 951.875 3461.775 968.350 ;
        RECT 3438.620 951.760 3461.775 951.875 ;
        RECT 3471.165 951.760 3472.345 984.060 ;
        RECT 3482.245 968.350 3483.165 984.060 ;
        RECT 3481.735 951.760 3483.165 968.350 ;
        RECT 3438.620 950.330 3483.165 951.760 ;
      LAYER pwell ;
        RECT 3483.975 954.230 3485.985 985.160 ;
        RECT 3488.820 978.120 3491.550 991.615 ;
        RECT 3487.520 954.230 3491.550 978.120 ;
        RECT 3483.975 953.135 3491.550 954.230 ;
        RECT 3513.135 990.755 3518.355 1025.265 ;
        RECT 3513.135 964.090 3517.315 990.755 ;
      LAYER nwell ;
        RECT 3518.665 984.960 3528.380 1031.415 ;
      LAYER pwell ;
        RECT 3513.135 953.135 3518.355 964.090 ;
        RECT 3483.975 950.710 3518.355 953.135 ;
      LAYER nwell ;
        RECT 3518.665 950.560 3528.385 984.960 ;
      LAYER pwell ;
        RECT 3528.685 950.710 3532.565 1031.290 ;
      LAYER nwell ;
        RECT 3532.880 1024.615 3566.975 1031.415 ;
        RECT 3532.880 952.370 3534.690 1024.615 ;
        RECT 3556.515 1023.485 3566.975 1024.615 ;
        RECT 3556.515 964.030 3558.475 1023.485 ;
        RECT 3561.545 964.030 3566.975 1023.485 ;
        RECT 3556.515 952.370 3566.975 964.030 ;
        RECT 3532.880 950.565 3566.975 952.370 ;
        RECT 3532.880 950.560 3558.230 950.565 ;
        RECT 107.600 907.585 111.515 907.880 ;
        RECT 118.765 907.285 143.410 908.715 ;
        RECT 190.675 907.585 194.335 911.110 ;
        RECT 3393.665 802.890 3397.325 806.415 ;
        RECT 3444.590 805.285 3469.235 806.715 ;
        RECT 3476.485 806.120 3480.400 806.415 ;
        RECT 3407.155 741.170 3411.080 801.420 ;
        RECT 3444.590 782.485 3446.020 805.285 ;
        RECT 3448.180 802.190 3450.340 805.285 ;
        RECT 3448.180 795.540 3449.020 802.190 ;
        RECT 3448.770 792.465 3449.020 795.540 ;
        RECT 3467.805 781.185 3469.235 805.285 ;
        RECT 3473.580 803.205 3480.400 806.120 ;
        RECT 3473.580 801.470 3479.820 803.205 ;
        RECT 3474.660 800.025 3479.820 801.470 ;
      LAYER pwell ;
        RECT 3480.935 800.785 3518.355 806.215 ;
      LAYER nwell ;
        RECT 3474.660 797.580 3476.280 800.025 ;
        RECT 3474.660 797.505 3475.740 797.580 ;
      LAYER pwell ;
        RECT 3480.935 796.700 3484.255 800.785 ;
        RECT 3482.955 766.615 3484.255 796.700 ;
        RECT 3489.965 800.265 3518.355 800.785 ;
        RECT 3489.965 766.615 3491.550 800.265 ;
        RECT 3482.955 760.160 3485.985 766.615 ;
        RECT 3482.955 759.410 3483.260 760.160 ;
      LAYER nwell ;
        RECT 3422.265 747.725 3424.055 757.085 ;
        RECT 3420.410 741.170 3424.055 747.725 ;
        RECT 3407.155 725.550 3413.345 741.170 ;
        RECT 3417.785 725.550 3424.055 741.170 ;
        RECT 3460.595 743.350 3461.265 759.060 ;
        RECT 3438.620 726.875 3440.050 735.665 ;
        RECT 3453.195 726.875 3454.045 735.665 ;
        RECT 3460.595 726.875 3461.775 743.350 ;
        RECT 3438.620 726.760 3461.775 726.875 ;
        RECT 3471.165 726.760 3472.345 759.060 ;
        RECT 3482.245 743.350 3483.165 759.060 ;
        RECT 3481.735 726.760 3483.165 743.350 ;
        RECT 3438.620 725.330 3483.165 726.760 ;
      LAYER pwell ;
        RECT 3483.975 729.230 3485.985 760.160 ;
        RECT 3488.820 753.120 3491.550 766.615 ;
        RECT 3487.520 729.230 3491.550 753.120 ;
        RECT 3483.975 728.135 3491.550 729.230 ;
        RECT 3513.135 765.755 3518.355 800.265 ;
        RECT 3513.135 739.090 3517.315 765.755 ;
      LAYER nwell ;
        RECT 3518.665 759.960 3528.380 806.415 ;
      LAYER pwell ;
        RECT 3513.135 728.135 3518.355 739.090 ;
        RECT 3483.975 725.710 3518.355 728.135 ;
      LAYER nwell ;
        RECT 3518.665 725.560 3528.385 759.960 ;
      LAYER pwell ;
        RECT 3528.685 725.710 3532.565 806.290 ;
      LAYER nwell ;
        RECT 3532.880 799.615 3566.975 806.415 ;
        RECT 3532.880 727.370 3534.690 799.615 ;
        RECT 3556.515 798.485 3566.975 799.615 ;
        RECT 3556.515 739.030 3558.475 798.485 ;
        RECT 3561.545 739.030 3566.975 798.485 ;
        RECT 3556.515 727.370 3566.975 739.030 ;
        RECT 3532.880 725.565 3566.975 727.370 ;
        RECT 3532.880 725.560 3558.230 725.565 ;
        RECT 197.795 562.860 199.315 621.965 ;
        RECT 3393.665 576.890 3397.325 580.415 ;
        RECT 3444.590 579.285 3469.235 580.715 ;
        RECT 3476.485 580.120 3480.400 580.415 ;
      LAYER pwell ;
        RECT 176.210 554.495 199.065 562.285 ;
      LAYER nwell ;
        RECT 3407.155 515.170 3411.080 575.420 ;
        RECT 3444.590 556.485 3446.020 579.285 ;
        RECT 3448.180 576.190 3450.340 579.285 ;
        RECT 3448.180 569.540 3449.020 576.190 ;
        RECT 3448.770 566.465 3449.020 569.540 ;
        RECT 3467.805 555.185 3469.235 579.285 ;
        RECT 3473.580 577.205 3480.400 580.120 ;
        RECT 3473.580 575.470 3479.820 577.205 ;
        RECT 3474.660 574.025 3479.820 575.470 ;
      LAYER pwell ;
        RECT 3480.935 574.785 3518.355 580.215 ;
      LAYER nwell ;
        RECT 3474.660 571.580 3476.280 574.025 ;
        RECT 3474.660 571.505 3475.740 571.580 ;
      LAYER pwell ;
        RECT 3480.935 570.700 3484.255 574.785 ;
        RECT 3482.955 540.615 3484.255 570.700 ;
        RECT 3489.965 574.265 3518.355 574.785 ;
        RECT 3489.965 540.615 3491.550 574.265 ;
        RECT 3482.955 534.160 3485.985 540.615 ;
        RECT 3482.955 533.410 3483.260 534.160 ;
      LAYER nwell ;
        RECT 3422.265 521.725 3424.055 531.085 ;
        RECT 3420.410 515.170 3424.055 521.725 ;
        RECT 3407.155 499.550 3413.345 515.170 ;
        RECT 3417.785 499.550 3424.055 515.170 ;
        RECT 3460.595 517.350 3461.265 533.060 ;
        RECT 3438.620 500.875 3440.050 509.665 ;
        RECT 3453.195 500.875 3454.045 509.665 ;
        RECT 3460.595 500.875 3461.775 517.350 ;
        RECT 3438.620 500.760 3461.775 500.875 ;
        RECT 3471.165 500.760 3472.345 533.060 ;
        RECT 3482.245 517.350 3483.165 533.060 ;
        RECT 3481.735 500.760 3483.165 517.350 ;
        RECT 3438.620 499.330 3483.165 500.760 ;
      LAYER pwell ;
        RECT 3483.975 503.230 3485.985 534.160 ;
        RECT 3488.820 527.120 3491.550 540.615 ;
        RECT 3487.520 503.230 3491.550 527.120 ;
        RECT 3483.975 502.135 3491.550 503.230 ;
        RECT 3513.135 539.755 3518.355 574.265 ;
        RECT 3513.135 513.090 3517.315 539.755 ;
      LAYER nwell ;
        RECT 3518.665 533.960 3528.380 580.415 ;
      LAYER pwell ;
        RECT 3513.135 502.135 3518.355 513.090 ;
        RECT 3483.975 499.710 3518.355 502.135 ;
      LAYER nwell ;
        RECT 3518.665 499.560 3528.385 533.960 ;
      LAYER pwell ;
        RECT 3528.685 499.710 3532.565 580.290 ;
      LAYER nwell ;
        RECT 3532.880 573.615 3566.975 580.415 ;
        RECT 3532.880 501.370 3534.690 573.615 ;
        RECT 3556.515 572.485 3566.975 573.615 ;
        RECT 3556.515 513.030 3558.475 572.485 ;
        RECT 3561.545 513.030 3566.975 572.485 ;
        RECT 3556.515 501.370 3566.975 513.030 ;
        RECT 3532.880 499.565 3566.975 501.370 ;
        RECT 3532.880 499.560 3558.230 499.565 ;
        RECT 398.035 197.795 457.140 199.315 ;
        RECT 2849.035 197.795 2908.140 199.315 ;
        RECT 3118.035 197.795 3177.140 199.315 ;
        RECT 1008.890 190.675 1012.415 194.335 ;
        RECT 1551.890 190.675 1555.415 194.335 ;
        RECT 1825.890 190.675 1829.415 194.335 ;
        RECT 2099.890 190.675 2103.415 194.335 ;
        RECT 2373.890 190.675 2377.415 194.335 ;
        RECT 2647.890 190.675 2651.415 194.335 ;
        RECT 931.550 176.920 1007.420 180.845 ;
        RECT 1474.550 176.920 1550.420 180.845 ;
        RECT 1748.550 176.920 1824.420 180.845 ;
        RECT 2022.550 176.920 2098.420 180.845 ;
        RECT 2296.550 176.920 2372.420 180.845 ;
        RECT 2570.550 176.920 2646.420 180.845 ;
        RECT 931.550 174.655 947.170 176.920 ;
        RECT 1474.550 174.655 1490.170 176.920 ;
        RECT 1748.550 174.655 1764.170 176.920 ;
        RECT 2022.550 174.655 2038.170 176.920 ;
        RECT 2296.550 174.655 2312.170 176.920 ;
        RECT 2570.550 174.655 2586.170 176.920 ;
      LAYER pwell ;
        RECT 3177.715 176.210 3185.505 199.065 ;
      LAYER nwell ;
        RECT 931.550 167.590 947.170 170.215 ;
        RECT 1474.550 167.590 1490.170 170.215 ;
        RECT 1748.550 167.590 1764.170 170.215 ;
        RECT 2022.550 167.590 2038.170 170.215 ;
        RECT 2296.550 167.590 2312.170 170.215 ;
        RECT 2570.550 167.590 2586.170 170.215 ;
        RECT 931.550 165.735 953.725 167.590 ;
        RECT 1474.550 165.735 1496.725 167.590 ;
        RECT 1748.550 165.735 1770.725 167.590 ;
        RECT 2022.550 165.735 2044.725 167.590 ;
        RECT 2296.550 165.735 2318.725 167.590 ;
        RECT 2570.550 165.735 2592.725 167.590 ;
        RECT 931.550 163.945 963.085 165.735 ;
        RECT 1474.550 163.945 1506.085 165.735 ;
        RECT 1748.550 163.945 1780.085 165.735 ;
        RECT 2022.550 163.945 2054.085 165.735 ;
        RECT 2296.550 163.945 2328.085 165.735 ;
        RECT 2570.550 163.945 2602.085 165.735 ;
        RECT 931.330 147.950 941.665 149.380 ;
        RECT 1474.330 147.950 1484.665 149.380 ;
        RECT 1748.330 147.950 1758.665 149.380 ;
        RECT 2022.330 147.950 2032.665 149.380 ;
        RECT 2296.330 147.950 2306.665 149.380 ;
        RECT 2570.330 147.950 2580.665 149.380 ;
        RECT 931.330 134.805 932.875 147.950 ;
        RECT 988.485 141.980 1012.715 143.410 ;
        RECT 1011.285 139.820 1012.715 141.980 ;
        RECT 1001.540 139.230 1012.715 139.820 ;
        RECT 998.465 138.980 1012.715 139.230 ;
        RECT 1008.190 137.660 1012.715 138.980 ;
        RECT 931.330 133.955 941.665 134.805 ;
        RECT 931.330 127.405 932.875 133.955 ;
        RECT 931.330 126.735 965.060 127.405 ;
        RECT 931.330 126.225 949.350 126.735 ;
        RECT 931.330 116.835 932.760 126.225 ;
        RECT 1011.285 120.195 1012.715 137.660 ;
        RECT 987.185 118.765 1012.715 120.195 ;
        RECT 1474.330 134.805 1475.875 147.950 ;
        RECT 1531.485 141.980 1555.715 143.410 ;
        RECT 1554.285 139.820 1555.715 141.980 ;
        RECT 1544.540 139.230 1555.715 139.820 ;
        RECT 1541.465 138.980 1555.715 139.230 ;
        RECT 1551.190 137.660 1555.715 138.980 ;
        RECT 1474.330 133.955 1484.665 134.805 ;
        RECT 1474.330 127.405 1475.875 133.955 ;
        RECT 1474.330 126.735 1508.060 127.405 ;
        RECT 1474.330 126.225 1492.350 126.735 ;
        RECT 1474.330 116.835 1475.760 126.225 ;
        RECT 1554.285 120.195 1555.715 137.660 ;
        RECT 1530.185 118.765 1555.715 120.195 ;
        RECT 1748.330 134.805 1749.875 147.950 ;
        RECT 1805.485 141.980 1829.715 143.410 ;
        RECT 1828.285 139.820 1829.715 141.980 ;
        RECT 1818.540 139.230 1829.715 139.820 ;
        RECT 1815.465 138.980 1829.715 139.230 ;
        RECT 1825.190 137.660 1829.715 138.980 ;
        RECT 1748.330 133.955 1758.665 134.805 ;
        RECT 1748.330 127.405 1749.875 133.955 ;
        RECT 1748.330 126.735 1782.060 127.405 ;
        RECT 1748.330 126.225 1766.350 126.735 ;
        RECT 1748.330 116.835 1749.760 126.225 ;
        RECT 1828.285 120.195 1829.715 137.660 ;
        RECT 1804.185 118.765 1829.715 120.195 ;
        RECT 2022.330 134.805 2023.875 147.950 ;
        RECT 2079.485 141.980 2103.715 143.410 ;
        RECT 2102.285 139.820 2103.715 141.980 ;
        RECT 2092.540 139.230 2103.715 139.820 ;
        RECT 2089.465 138.980 2103.715 139.230 ;
        RECT 2099.190 137.660 2103.715 138.980 ;
        RECT 2022.330 133.955 2032.665 134.805 ;
        RECT 2022.330 127.405 2023.875 133.955 ;
        RECT 2022.330 126.735 2056.060 127.405 ;
        RECT 2022.330 126.225 2040.350 126.735 ;
        RECT 2022.330 116.835 2023.760 126.225 ;
        RECT 2102.285 120.195 2103.715 137.660 ;
        RECT 2078.185 118.765 2103.715 120.195 ;
        RECT 2296.330 134.805 2297.875 147.950 ;
        RECT 2353.485 141.980 2377.715 143.410 ;
        RECT 2376.285 139.820 2377.715 141.980 ;
        RECT 2366.540 139.230 2377.715 139.820 ;
        RECT 2363.465 138.980 2377.715 139.230 ;
        RECT 2373.190 137.660 2377.715 138.980 ;
        RECT 2296.330 133.955 2306.665 134.805 ;
        RECT 2296.330 127.405 2297.875 133.955 ;
        RECT 2296.330 126.735 2330.060 127.405 ;
        RECT 2296.330 126.225 2314.350 126.735 ;
        RECT 2296.330 116.835 2297.760 126.225 ;
        RECT 2376.285 120.195 2377.715 137.660 ;
        RECT 2352.185 118.765 2377.715 120.195 ;
        RECT 2570.330 134.805 2571.875 147.950 ;
        RECT 2627.485 141.980 2651.715 143.410 ;
        RECT 2650.285 139.820 2651.715 141.980 ;
        RECT 2640.540 139.230 2651.715 139.820 ;
        RECT 2637.465 138.980 2651.715 139.230 ;
        RECT 2647.190 137.660 2651.715 138.980 ;
        RECT 2570.330 133.955 2580.665 134.805 ;
        RECT 2570.330 127.405 2571.875 133.955 ;
        RECT 2570.330 126.735 2604.060 127.405 ;
        RECT 2570.330 126.225 2588.350 126.735 ;
        RECT 2570.330 116.835 2571.760 126.225 ;
        RECT 2650.285 120.195 2651.715 137.660 ;
        RECT 2626.185 118.765 2651.715 120.195 ;
        RECT 931.330 115.655 965.060 116.835 ;
        RECT 1474.330 115.655 1508.060 116.835 ;
        RECT 1748.330 115.655 1782.060 116.835 ;
        RECT 2022.330 115.655 2056.060 116.835 ;
        RECT 2296.330 115.655 2330.060 116.835 ;
        RECT 2570.330 115.655 2604.060 116.835 ;
        RECT 931.330 106.265 932.760 115.655 ;
        RECT 1007.470 113.340 1012.120 114.420 ;
        RECT 1003.505 112.260 1012.120 113.340 ;
        RECT 1003.580 111.720 1012.120 112.260 ;
        RECT 1006.025 111.515 1012.120 111.720 ;
        RECT 1006.025 108.180 1012.415 111.515 ;
        RECT 1009.205 107.600 1012.415 108.180 ;
        RECT 931.330 105.755 949.350 106.265 ;
        RECT 931.330 104.835 965.060 105.755 ;
      LAYER pwell ;
        RECT 1002.700 105.045 1012.215 107.065 ;
        RECT 965.410 104.740 1012.215 105.045 ;
      LAYER nwell ;
        RECT 1474.330 106.265 1475.760 115.655 ;
        RECT 1550.470 113.340 1555.120 114.420 ;
        RECT 1546.505 112.260 1555.120 113.340 ;
        RECT 1546.580 111.720 1555.120 112.260 ;
        RECT 1549.025 111.515 1555.120 111.720 ;
        RECT 1549.025 108.180 1555.415 111.515 ;
        RECT 1552.205 107.600 1555.415 108.180 ;
        RECT 1474.330 105.755 1492.350 106.265 ;
        RECT 1474.330 104.835 1508.060 105.755 ;
      LAYER pwell ;
        RECT 1545.700 105.045 1555.215 107.065 ;
        RECT 1508.410 104.740 1555.215 105.045 ;
      LAYER nwell ;
        RECT 1748.330 106.265 1749.760 115.655 ;
        RECT 1824.470 113.340 1829.120 114.420 ;
        RECT 1820.505 112.260 1829.120 113.340 ;
        RECT 1820.580 111.720 1829.120 112.260 ;
        RECT 1823.025 111.515 1829.120 111.720 ;
        RECT 1823.025 108.180 1829.415 111.515 ;
        RECT 1826.205 107.600 1829.415 108.180 ;
        RECT 1748.330 105.755 1766.350 106.265 ;
        RECT 1748.330 104.835 1782.060 105.755 ;
      LAYER pwell ;
        RECT 1819.700 105.045 1829.215 107.065 ;
        RECT 1782.410 104.740 1829.215 105.045 ;
      LAYER nwell ;
        RECT 2022.330 106.265 2023.760 115.655 ;
        RECT 2098.470 113.340 2103.120 114.420 ;
        RECT 2094.505 112.260 2103.120 113.340 ;
        RECT 2094.580 111.720 2103.120 112.260 ;
        RECT 2097.025 111.515 2103.120 111.720 ;
        RECT 2097.025 108.180 2103.415 111.515 ;
        RECT 2100.205 107.600 2103.415 108.180 ;
        RECT 2022.330 105.755 2040.350 106.265 ;
        RECT 2022.330 104.835 2056.060 105.755 ;
      LAYER pwell ;
        RECT 2093.700 105.045 2103.215 107.065 ;
        RECT 2056.410 104.740 2103.215 105.045 ;
      LAYER nwell ;
        RECT 2296.330 106.265 2297.760 115.655 ;
        RECT 2372.470 113.340 2377.120 114.420 ;
        RECT 2368.505 112.260 2377.120 113.340 ;
        RECT 2368.580 111.720 2377.120 112.260 ;
        RECT 2371.025 111.515 2377.120 111.720 ;
        RECT 2371.025 108.180 2377.415 111.515 ;
        RECT 2374.205 107.600 2377.415 108.180 ;
        RECT 2296.330 105.755 2314.350 106.265 ;
        RECT 2296.330 104.835 2330.060 105.755 ;
      LAYER pwell ;
        RECT 2367.700 105.045 2377.215 107.065 ;
        RECT 2330.410 104.740 2377.215 105.045 ;
      LAYER nwell ;
        RECT 2570.330 106.265 2571.760 115.655 ;
        RECT 2646.470 113.340 2651.120 114.420 ;
        RECT 2642.505 112.260 2651.120 113.340 ;
        RECT 2642.580 111.720 2651.120 112.260 ;
        RECT 2645.025 111.515 2651.120 111.720 ;
        RECT 2645.025 108.180 2651.415 111.515 ;
        RECT 2648.205 107.600 2651.415 108.180 ;
        RECT 2570.330 105.755 2588.350 106.265 ;
        RECT 2570.330 104.835 2604.060 105.755 ;
      LAYER pwell ;
        RECT 2641.700 105.045 2651.215 107.065 ;
        RECT 2604.410 104.740 2651.215 105.045 ;
        RECT 966.160 104.025 1012.215 104.740 ;
        RECT 1509.160 104.025 1555.215 104.740 ;
        RECT 1783.160 104.025 1829.215 104.740 ;
        RECT 2057.160 104.025 2103.215 104.740 ;
        RECT 2331.160 104.025 2377.215 104.740 ;
        RECT 2605.160 104.025 2651.215 104.740 ;
        RECT 931.710 103.745 1012.215 104.025 ;
        RECT 679.530 103.265 738.130 103.270 ;
        RECT 662.870 102.005 738.130 103.265 ;
        RECT 662.870 100.770 666.070 102.005 ;
        RECT 679.530 100.770 738.130 102.005 ;
        RECT 662.870 97.475 738.130 100.770 ;
        RECT 662.870 75.865 664.440 97.475 ;
        RECT 736.565 75.865 738.130 97.475 ;
        RECT 662.870 70.685 738.130 75.865 ;
        RECT 662.870 69.645 676.090 70.685 ;
        RECT 696.250 69.645 738.130 70.685 ;
        RECT 931.710 102.015 972.615 103.745 ;
        RECT 931.710 100.480 935.230 102.015 ;
        RECT 931.710 99.180 959.120 100.480 ;
        RECT 931.710 98.035 972.615 99.180 ;
        RECT 1006.785 98.035 1012.215 103.745 ;
        RECT 931.710 96.450 1012.215 98.035 ;
        RECT 931.710 74.865 934.135 96.450 ;
        RECT 1006.265 74.865 1012.215 96.450 ;
        RECT 931.710 70.685 1012.215 74.865 ;
        RECT 931.710 69.645 945.090 70.685 ;
        RECT 971.755 69.645 1012.215 70.685 ;
        RECT 1474.710 103.745 1555.215 104.025 ;
        RECT 1474.710 102.015 1515.615 103.745 ;
        RECT 1474.710 100.480 1478.230 102.015 ;
        RECT 1474.710 99.180 1502.120 100.480 ;
        RECT 1474.710 98.035 1515.615 99.180 ;
        RECT 1549.785 98.035 1555.215 103.745 ;
        RECT 1474.710 96.450 1555.215 98.035 ;
        RECT 1474.710 74.865 1477.135 96.450 ;
        RECT 1549.265 74.865 1555.215 96.450 ;
        RECT 1474.710 70.685 1555.215 74.865 ;
        RECT 1474.710 69.645 1488.090 70.685 ;
        RECT 1514.755 69.645 1555.215 70.685 ;
        RECT 1748.710 103.745 1829.215 104.025 ;
        RECT 1748.710 102.015 1789.615 103.745 ;
        RECT 1748.710 100.480 1752.230 102.015 ;
        RECT 1748.710 99.180 1776.120 100.480 ;
        RECT 1748.710 98.035 1789.615 99.180 ;
        RECT 1823.785 98.035 1829.215 103.745 ;
        RECT 1748.710 96.450 1829.215 98.035 ;
        RECT 1748.710 74.865 1751.135 96.450 ;
        RECT 1823.265 74.865 1829.215 96.450 ;
        RECT 1748.710 70.685 1829.215 74.865 ;
        RECT 1748.710 69.645 1762.090 70.685 ;
        RECT 1788.755 69.645 1829.215 70.685 ;
        RECT 2022.710 103.745 2103.215 104.025 ;
        RECT 2022.710 102.015 2063.615 103.745 ;
        RECT 2022.710 100.480 2026.230 102.015 ;
        RECT 2022.710 99.180 2050.120 100.480 ;
        RECT 2022.710 98.035 2063.615 99.180 ;
        RECT 2097.785 98.035 2103.215 103.745 ;
        RECT 2022.710 96.450 2103.215 98.035 ;
        RECT 2022.710 74.865 2025.135 96.450 ;
        RECT 2097.265 74.865 2103.215 96.450 ;
        RECT 2022.710 70.685 2103.215 74.865 ;
        RECT 2022.710 69.645 2036.090 70.685 ;
        RECT 2062.755 69.645 2103.215 70.685 ;
        RECT 2296.710 103.745 2377.215 104.025 ;
        RECT 2296.710 102.015 2337.615 103.745 ;
        RECT 2296.710 100.480 2300.230 102.015 ;
        RECT 2296.710 99.180 2324.120 100.480 ;
        RECT 2296.710 98.035 2337.615 99.180 ;
        RECT 2371.785 98.035 2377.215 103.745 ;
        RECT 2296.710 96.450 2377.215 98.035 ;
        RECT 2296.710 74.865 2299.135 96.450 ;
        RECT 2371.265 74.865 2377.215 96.450 ;
        RECT 2296.710 70.685 2377.215 74.865 ;
        RECT 2296.710 69.645 2310.090 70.685 ;
        RECT 2336.755 69.645 2377.215 70.685 ;
        RECT 2570.710 103.745 2651.215 104.025 ;
        RECT 2570.710 102.015 2611.615 103.745 ;
        RECT 2570.710 100.480 2574.230 102.015 ;
        RECT 2570.710 99.180 2598.120 100.480 ;
        RECT 2570.710 98.035 2611.615 99.180 ;
        RECT 2645.785 98.035 2651.215 103.745 ;
        RECT 2570.710 96.450 2651.215 98.035 ;
        RECT 2570.710 74.865 2573.135 96.450 ;
        RECT 2645.265 74.865 2651.215 96.450 ;
        RECT 2570.710 70.685 2651.215 74.865 ;
        RECT 2570.710 69.645 2584.090 70.685 ;
        RECT 2610.755 69.645 2651.215 70.685 ;
      LAYER nwell ;
        RECT 662.670 59.620 738.330 69.335 ;
        RECT 931.560 59.620 1012.415 69.335 ;
        RECT 1474.560 59.620 1555.415 69.335 ;
        RECT 1748.560 59.620 1829.415 69.335 ;
        RECT 2022.560 59.620 2103.415 69.335 ;
        RECT 2296.560 59.620 2377.415 69.335 ;
        RECT 2570.560 59.620 2651.415 69.335 ;
        RECT 931.560 59.615 965.960 59.620 ;
        RECT 1474.560 59.615 1508.960 59.620 ;
        RECT 1748.560 59.615 1782.960 59.620 ;
        RECT 2022.560 59.615 2056.960 59.620 ;
        RECT 2296.560 59.615 2330.960 59.620 ;
        RECT 2570.560 59.615 2604.960 59.620 ;
      LAYER pwell ;
        RECT 662.710 55.435 738.290 59.315 ;
        RECT 931.710 55.435 1012.290 59.315 ;
        RECT 1474.710 55.435 1555.290 59.315 ;
        RECT 1748.710 55.435 1829.290 59.315 ;
        RECT 2022.710 55.435 2103.290 59.315 ;
        RECT 2296.710 55.435 2377.290 59.315 ;
        RECT 2570.710 55.435 2651.290 59.315 ;
      LAYER nwell ;
        RECT 662.380 53.310 738.515 55.120 ;
        RECT 662.380 31.485 664.905 53.310 ;
        RECT 736.325 31.485 738.515 53.310 ;
        RECT 662.380 29.790 738.515 31.485 ;
        RECT 931.560 53.310 1012.415 55.120 ;
        RECT 931.560 31.485 933.370 53.310 ;
        RECT 1005.615 31.485 1012.415 53.310 ;
        RECT 931.560 29.770 1012.415 31.485 ;
        RECT 1474.560 53.310 1555.415 55.120 ;
        RECT 1474.560 31.485 1476.370 53.310 ;
        RECT 1548.615 31.485 1555.415 53.310 ;
        RECT 1474.560 29.770 1555.415 31.485 ;
        RECT 1748.560 53.310 1829.415 55.120 ;
        RECT 1748.560 31.485 1750.370 53.310 ;
        RECT 1822.615 31.485 1829.415 53.310 ;
        RECT 1748.560 29.770 1829.415 31.485 ;
        RECT 2022.560 53.310 2103.415 55.120 ;
        RECT 2022.560 31.485 2024.370 53.310 ;
        RECT 2096.615 31.485 2103.415 53.310 ;
        RECT 2022.560 29.770 2103.415 31.485 ;
        RECT 2296.560 53.310 2377.415 55.120 ;
        RECT 2296.560 31.485 2298.370 53.310 ;
        RECT 2370.615 31.485 2377.415 53.310 ;
        RECT 2296.560 29.770 2377.415 31.485 ;
        RECT 2570.560 53.310 2651.415 55.120 ;
        RECT 2570.560 31.485 2572.370 53.310 ;
        RECT 2644.615 31.485 2651.415 53.310 ;
        RECT 2570.560 29.770 2651.415 31.485 ;
        RECT 931.565 29.525 1012.415 29.770 ;
        RECT 931.565 26.455 945.030 29.525 ;
        RECT 1004.485 26.455 1012.415 29.525 ;
        RECT 931.565 21.025 1012.415 26.455 ;
        RECT 1474.565 29.525 1555.415 29.770 ;
        RECT 1474.565 26.455 1488.030 29.525 ;
        RECT 1547.485 26.455 1555.415 29.525 ;
        RECT 1474.565 21.025 1555.415 26.455 ;
        RECT 1748.565 29.525 1829.415 29.770 ;
        RECT 1748.565 26.455 1762.030 29.525 ;
        RECT 1821.485 26.455 1829.415 29.525 ;
        RECT 1748.565 21.025 1829.415 26.455 ;
        RECT 2022.565 29.525 2103.415 29.770 ;
        RECT 2022.565 26.455 2036.030 29.525 ;
        RECT 2095.485 26.455 2103.415 29.525 ;
        RECT 2022.565 21.025 2103.415 26.455 ;
        RECT 2296.565 29.525 2377.415 29.770 ;
        RECT 2296.565 26.455 2310.030 29.525 ;
        RECT 2369.485 26.455 2377.415 29.525 ;
        RECT 2296.565 21.025 2377.415 26.455 ;
        RECT 2570.565 29.525 2651.415 29.770 ;
        RECT 2570.565 26.455 2584.030 29.525 ;
        RECT 2643.485 26.455 2651.415 29.525 ;
        RECT 2570.565 21.025 2651.415 26.455 ;
      LAYER li1 ;
        RECT 383.905 5036.265 453.045 5169.100 ;
        RECT 640.905 5036.265 710.045 5169.100 ;
        RECT 897.905 5036.265 967.045 5169.100 ;
        RECT 1152.610 4990.035 1224.855 5187.695 ;
        RECT 1410.610 4990.035 1482.855 5187.695 ;
        RECT 1668.070 4990.035 1739.775 5187.695 ;
        RECT 1921.905 5036.265 1991.045 5169.100 ;
        RECT 2366.905 5036.265 2436.045 5169.100 ;
        RECT 2623.905 5036.265 2693.045 5169.100 ;
        RECT 2879.070 4990.035 2950.775 5187.695 ;
        RECT 3132.905 5036.265 3202.045 5169.100 ;
        RECT 1152.610 4989.065 1163.155 4990.035 ;
        RECT 1164.035 4989.920 1165.045 4990.035 ;
        RECT 1221.730 4989.920 1222.680 4990.035 ;
        RECT 1164.035 4988.970 1222.680 4989.920 ;
        RECT 1410.610 4989.065 1421.155 4990.035 ;
        RECT 1422.035 4989.920 1423.045 4990.035 ;
        RECT 1479.730 4989.920 1480.680 4990.035 ;
        RECT 1422.035 4988.970 1480.680 4989.920 ;
        RECT 1679.065 4989.890 1680.045 4990.035 ;
        RECT 1736.760 4989.890 1737.650 4990.035 ;
        RECT 1679.065 4989.000 1737.650 4989.890 ;
        RECT 2890.065 4989.890 2891.045 4990.035 ;
        RECT 2947.760 4989.890 2948.650 4990.035 ;
        RECT 2890.065 4989.000 2948.650 4989.890 ;
        RECT 18.900 4773.905 151.735 4843.045 ;
        RECT 3389.065 4826.845 3587.695 4837.390 ;
        RECT 3390.035 4825.965 3587.695 4826.845 ;
        RECT 3388.970 4824.955 3587.695 4825.965 ;
        RECT 3388.970 4768.270 3389.920 4824.955 ;
        RECT 3390.035 4768.270 3587.695 4824.955 ;
        RECT 3388.970 4767.320 3587.695 4768.270 ;
        RECT 3390.035 4765.145 3587.695 4767.320 ;
        RECT 0.220 4560.240 196.980 4634.755 ;
        RECT 3391.020 4538.245 3587.780 4612.760 ;
        RECT 0.305 4419.680 197.965 4421.855 ;
        RECT 0.305 4418.730 199.030 4419.680 ;
        RECT 0.305 4362.045 197.965 4418.730 ;
        RECT 198.080 4362.045 199.030 4418.730 ;
        RECT 3483.895 4392.085 3518.220 4392.115 ;
        RECT 3519.275 4392.085 3528.150 4392.115 ;
        RECT 3393.995 4392.000 3396.995 4392.085 ;
        RECT 3445.220 4392.000 3468.605 4392.085 ;
        RECT 3476.815 4392.000 3480.070 4392.085 ;
        RECT 3481.065 4392.000 3518.225 4392.085 ;
        RECT 3518.995 4392.000 3528.150 4392.085 ;
        RECT 3528.815 4392.000 3532.435 4392.160 ;
        RECT 3533.155 4392.085 3558.090 4392.115 ;
        RECT 3533.155 4392.000 3566.645 4392.085 ;
        RECT 0.305 4361.035 199.030 4362.045 ;
        RECT 0.305 4360.155 197.965 4361.035 ;
        RECT 0.305 4349.610 198.935 4360.155 ;
        RECT 3388.230 4312.000 3587.705 4392.000 ;
        RECT 3407.485 4311.880 3413.015 4312.000 ;
        RECT 3418.115 4311.880 3423.725 4312.000 ;
        RECT 3439.250 4311.915 3482.580 4312.000 ;
        RECT 3484.105 4311.840 3518.225 4312.000 ;
        RECT 3518.995 4311.915 3528.055 4312.000 ;
        RECT 3528.815 4311.840 3532.435 4312.000 ;
        RECT 3533.215 4311.895 3566.645 4312.000 ;
        RECT 0.305 4208.650 197.965 4210.775 ;
        RECT 0.305 4207.760 199.000 4208.650 ;
        RECT 0.305 4151.045 197.965 4207.760 ;
        RECT 198.110 4151.045 199.000 4207.760 ;
        RECT 3389.065 4155.845 3587.695 4166.390 ;
        RECT 3390.035 4154.965 3587.695 4155.845 ;
        RECT 0.305 4150.065 199.000 4151.045 ;
        RECT 3388.970 4153.955 3587.695 4154.965 ;
        RECT 0.305 4139.070 197.965 4150.065 ;
        RECT 3388.970 4097.270 3389.920 4153.955 ;
        RECT 3390.035 4097.270 3587.695 4153.955 ;
        RECT 3388.970 4096.320 3587.695 4097.270 ;
        RECT 3390.035 4094.145 3587.695 4096.320 ;
        RECT 21.355 4002.000 54.785 4002.105 ;
        RECT 55.565 4002.000 59.185 4002.160 ;
        RECT 59.945 4002.000 69.005 4002.085 ;
        RECT 69.775 4002.000 103.895 4002.160 ;
        RECT 105.420 4002.000 148.750 4002.085 ;
        RECT 164.275 4002.000 169.885 4002.120 ;
        RECT 174.985 4002.000 180.515 4002.120 ;
        RECT 0.295 3922.000 199.770 4002.000 ;
        RECT 3483.895 3946.085 3518.220 3946.115 ;
        RECT 3519.275 3946.085 3528.150 3946.115 ;
        RECT 3393.995 3946.000 3396.995 3946.085 ;
        RECT 3445.220 3946.000 3468.605 3946.085 ;
        RECT 3476.815 3946.000 3480.070 3946.085 ;
        RECT 3481.065 3946.000 3518.225 3946.085 ;
        RECT 3518.995 3946.000 3528.150 3946.085 ;
        RECT 3528.815 3946.000 3532.435 3946.160 ;
        RECT 3533.155 3946.085 3558.090 3946.115 ;
        RECT 3533.155 3946.000 3566.645 3946.085 ;
        RECT 21.355 3921.915 54.845 3922.000 ;
        RECT 29.910 3921.885 54.845 3921.915 ;
        RECT 55.565 3921.840 59.185 3922.000 ;
        RECT 59.850 3921.915 69.005 3922.000 ;
        RECT 69.775 3921.915 106.935 3922.000 ;
        RECT 107.930 3921.915 111.185 3922.000 ;
        RECT 119.395 3921.915 142.780 3922.000 ;
        RECT 191.005 3921.915 194.005 3922.000 ;
        RECT 59.850 3921.885 68.725 3921.915 ;
        RECT 69.780 3921.885 104.105 3921.915 ;
        RECT 3388.230 3866.000 3587.705 3946.000 ;
        RECT 3407.485 3865.880 3413.015 3866.000 ;
        RECT 3418.115 3865.880 3423.725 3866.000 ;
        RECT 3439.250 3865.915 3482.580 3866.000 ;
        RECT 3484.105 3865.840 3518.225 3866.000 ;
        RECT 3518.995 3865.915 3528.055 3866.000 ;
        RECT 3528.815 3865.840 3532.435 3866.000 ;
        RECT 3533.215 3865.895 3566.645 3866.000 ;
        RECT 21.355 3786.000 54.785 3786.105 ;
        RECT 55.565 3786.000 59.185 3786.160 ;
        RECT 59.945 3786.000 69.005 3786.085 ;
        RECT 69.775 3786.000 103.895 3786.160 ;
        RECT 105.420 3786.000 148.750 3786.085 ;
        RECT 164.275 3786.000 169.885 3786.120 ;
        RECT 174.985 3786.000 180.515 3786.120 ;
        RECT 0.295 3706.000 199.770 3786.000 ;
        RECT 3483.895 3721.085 3518.220 3721.115 ;
        RECT 3519.275 3721.085 3528.150 3721.115 ;
        RECT 3393.995 3721.000 3396.995 3721.085 ;
        RECT 3445.220 3721.000 3468.605 3721.085 ;
        RECT 3476.815 3721.000 3480.070 3721.085 ;
        RECT 3481.065 3721.000 3518.225 3721.085 ;
        RECT 3518.995 3721.000 3528.150 3721.085 ;
        RECT 3528.815 3721.000 3532.435 3721.160 ;
        RECT 3533.155 3721.085 3558.090 3721.115 ;
        RECT 3533.155 3721.000 3566.645 3721.085 ;
        RECT 21.355 3705.915 54.845 3706.000 ;
        RECT 29.910 3705.885 54.845 3705.915 ;
        RECT 55.565 3705.840 59.185 3706.000 ;
        RECT 59.850 3705.915 69.005 3706.000 ;
        RECT 69.775 3705.915 106.935 3706.000 ;
        RECT 107.930 3705.915 111.185 3706.000 ;
        RECT 119.395 3705.915 142.780 3706.000 ;
        RECT 191.005 3705.915 194.005 3706.000 ;
        RECT 59.850 3705.885 68.725 3705.915 ;
        RECT 69.780 3705.885 104.105 3705.915 ;
        RECT 3388.230 3641.000 3587.705 3721.000 ;
        RECT 3407.485 3640.880 3413.015 3641.000 ;
        RECT 3418.115 3640.880 3423.725 3641.000 ;
        RECT 3439.250 3640.915 3482.580 3641.000 ;
        RECT 3484.105 3640.840 3518.225 3641.000 ;
        RECT 3518.995 3640.915 3528.055 3641.000 ;
        RECT 3528.815 3640.840 3532.435 3641.000 ;
        RECT 3533.215 3640.895 3566.645 3641.000 ;
        RECT 21.355 3570.000 54.785 3570.105 ;
        RECT 55.565 3570.000 59.185 3570.160 ;
        RECT 59.945 3570.000 69.005 3570.085 ;
        RECT 69.775 3570.000 103.895 3570.160 ;
        RECT 105.420 3570.000 148.750 3570.085 ;
        RECT 164.275 3570.000 169.885 3570.120 ;
        RECT 174.985 3570.000 180.515 3570.120 ;
        RECT 0.295 3490.000 199.770 3570.000 ;
        RECT 3483.895 3496.085 3518.220 3496.115 ;
        RECT 3519.275 3496.085 3528.150 3496.115 ;
        RECT 3393.995 3496.000 3396.995 3496.085 ;
        RECT 3445.220 3496.000 3468.605 3496.085 ;
        RECT 3476.815 3496.000 3480.070 3496.085 ;
        RECT 3481.065 3496.000 3518.225 3496.085 ;
        RECT 3518.995 3496.000 3528.150 3496.085 ;
        RECT 3528.815 3496.000 3532.435 3496.160 ;
        RECT 3533.155 3496.085 3558.090 3496.115 ;
        RECT 3533.155 3496.000 3566.645 3496.085 ;
        RECT 21.355 3489.915 54.845 3490.000 ;
        RECT 29.910 3489.885 54.845 3489.915 ;
        RECT 55.565 3489.840 59.185 3490.000 ;
        RECT 59.850 3489.915 69.005 3490.000 ;
        RECT 69.775 3489.915 106.935 3490.000 ;
        RECT 107.930 3489.915 111.185 3490.000 ;
        RECT 119.395 3489.915 142.780 3490.000 ;
        RECT 191.005 3489.915 194.005 3490.000 ;
        RECT 59.850 3489.885 68.725 3489.915 ;
        RECT 69.780 3489.885 104.105 3489.915 ;
        RECT 3388.230 3416.000 3587.705 3496.000 ;
        RECT 3407.485 3415.880 3413.015 3416.000 ;
        RECT 3418.115 3415.880 3423.725 3416.000 ;
        RECT 3439.250 3415.915 3482.580 3416.000 ;
        RECT 3484.105 3415.840 3518.225 3416.000 ;
        RECT 3518.995 3415.915 3528.055 3416.000 ;
        RECT 3528.815 3415.840 3532.435 3416.000 ;
        RECT 3533.215 3415.895 3566.645 3416.000 ;
        RECT 21.355 3354.000 54.785 3354.105 ;
        RECT 55.565 3354.000 59.185 3354.160 ;
        RECT 59.945 3354.000 69.005 3354.085 ;
        RECT 69.775 3354.000 103.895 3354.160 ;
        RECT 105.420 3354.000 148.750 3354.085 ;
        RECT 164.275 3354.000 169.885 3354.120 ;
        RECT 174.985 3354.000 180.515 3354.120 ;
        RECT 0.295 3274.000 199.770 3354.000 ;
        RECT 21.355 3273.915 54.845 3274.000 ;
        RECT 29.910 3273.885 54.845 3273.915 ;
        RECT 55.565 3273.840 59.185 3274.000 ;
        RECT 59.850 3273.915 69.005 3274.000 ;
        RECT 69.775 3273.915 106.935 3274.000 ;
        RECT 107.930 3273.915 111.185 3274.000 ;
        RECT 119.395 3273.915 142.780 3274.000 ;
        RECT 191.005 3273.915 194.005 3274.000 ;
        RECT 59.850 3273.885 68.725 3273.915 ;
        RECT 69.780 3273.885 104.105 3273.915 ;
        RECT 3483.895 3270.085 3518.220 3270.115 ;
        RECT 3519.275 3270.085 3528.150 3270.115 ;
        RECT 3393.995 3270.000 3396.995 3270.085 ;
        RECT 3445.220 3270.000 3468.605 3270.085 ;
        RECT 3476.815 3270.000 3480.070 3270.085 ;
        RECT 3481.065 3270.000 3518.225 3270.085 ;
        RECT 3518.995 3270.000 3528.150 3270.085 ;
        RECT 3528.815 3270.000 3532.435 3270.160 ;
        RECT 3533.155 3270.085 3558.090 3270.115 ;
        RECT 3533.155 3270.000 3566.645 3270.085 ;
        RECT 3388.230 3190.000 3587.705 3270.000 ;
        RECT 3407.485 3189.880 3413.015 3190.000 ;
        RECT 3418.115 3189.880 3423.725 3190.000 ;
        RECT 3439.250 3189.915 3482.580 3190.000 ;
        RECT 3484.105 3189.840 3518.225 3190.000 ;
        RECT 3518.995 3189.915 3528.055 3190.000 ;
        RECT 3528.815 3189.840 3532.435 3190.000 ;
        RECT 3533.215 3189.895 3566.645 3190.000 ;
        RECT 21.355 3138.000 54.785 3138.105 ;
        RECT 55.565 3138.000 59.185 3138.160 ;
        RECT 59.945 3138.000 69.005 3138.085 ;
        RECT 69.775 3138.000 103.895 3138.160 ;
        RECT 105.420 3138.000 148.750 3138.085 ;
        RECT 164.275 3138.000 169.885 3138.120 ;
        RECT 174.985 3138.000 180.515 3138.120 ;
        RECT 0.295 3058.000 199.770 3138.000 ;
        RECT 21.355 3057.915 54.845 3058.000 ;
        RECT 29.910 3057.885 54.845 3057.915 ;
        RECT 55.565 3057.840 59.185 3058.000 ;
        RECT 59.850 3057.915 69.005 3058.000 ;
        RECT 69.775 3057.915 106.935 3058.000 ;
        RECT 107.930 3057.915 111.185 3058.000 ;
        RECT 119.395 3057.915 142.780 3058.000 ;
        RECT 191.005 3057.915 194.005 3058.000 ;
        RECT 59.850 3057.885 68.725 3057.915 ;
        RECT 69.780 3057.885 104.105 3057.915 ;
        RECT 3483.895 3045.085 3518.220 3045.115 ;
        RECT 3519.275 3045.085 3528.150 3045.115 ;
        RECT 3393.995 3045.000 3396.995 3045.085 ;
        RECT 3445.220 3045.000 3468.605 3045.085 ;
        RECT 3476.815 3045.000 3480.070 3045.085 ;
        RECT 3481.065 3045.000 3518.225 3045.085 ;
        RECT 3518.995 3045.000 3528.150 3045.085 ;
        RECT 3528.815 3045.000 3532.435 3045.160 ;
        RECT 3533.155 3045.085 3558.090 3045.115 ;
        RECT 3533.155 3045.000 3566.645 3045.085 ;
        RECT 3388.230 2965.000 3587.705 3045.000 ;
        RECT 3407.485 2964.880 3413.015 2965.000 ;
        RECT 3418.115 2964.880 3423.725 2965.000 ;
        RECT 3439.250 2964.915 3482.580 2965.000 ;
        RECT 3484.105 2964.840 3518.225 2965.000 ;
        RECT 3518.995 2964.915 3528.055 2965.000 ;
        RECT 3528.815 2964.840 3532.435 2965.000 ;
        RECT 3533.215 2964.895 3566.645 2965.000 ;
        RECT 21.355 2922.000 54.785 2922.105 ;
        RECT 55.565 2922.000 59.185 2922.160 ;
        RECT 59.945 2922.000 69.005 2922.085 ;
        RECT 69.775 2922.000 103.895 2922.160 ;
        RECT 105.420 2922.000 148.750 2922.085 ;
        RECT 164.275 2922.000 169.885 2922.120 ;
        RECT 174.985 2922.000 180.515 2922.120 ;
        RECT 0.295 2842.000 199.770 2922.000 ;
        RECT 21.355 2841.915 54.845 2842.000 ;
        RECT 29.910 2841.885 54.845 2841.915 ;
        RECT 55.565 2841.840 59.185 2842.000 ;
        RECT 59.850 2841.915 69.005 2842.000 ;
        RECT 69.775 2841.915 106.935 2842.000 ;
        RECT 107.930 2841.915 111.185 2842.000 ;
        RECT 119.395 2841.915 142.780 2842.000 ;
        RECT 191.005 2841.915 194.005 2842.000 ;
        RECT 59.850 2841.885 68.725 2841.915 ;
        RECT 69.780 2841.885 104.105 2841.915 ;
        RECT 3483.895 2819.085 3518.220 2819.115 ;
        RECT 3519.275 2819.085 3528.150 2819.115 ;
        RECT 3393.995 2819.000 3396.995 2819.085 ;
        RECT 3445.220 2819.000 3468.605 2819.085 ;
        RECT 3476.815 2819.000 3480.070 2819.085 ;
        RECT 3481.065 2819.000 3518.225 2819.085 ;
        RECT 3518.995 2819.000 3528.150 2819.085 ;
        RECT 3528.815 2819.000 3532.435 2819.160 ;
        RECT 3533.155 2819.085 3558.090 2819.115 ;
        RECT 3533.155 2819.000 3566.645 2819.085 ;
        RECT 3388.230 2739.000 3587.705 2819.000 ;
        RECT 3407.485 2738.880 3413.015 2739.000 ;
        RECT 3418.115 2738.880 3423.725 2739.000 ;
        RECT 3439.250 2738.915 3482.580 2739.000 ;
        RECT 3484.105 2738.840 3518.225 2739.000 ;
        RECT 3518.995 2738.915 3528.055 2739.000 ;
        RECT 3528.815 2738.840 3532.435 2739.000 ;
        RECT 3533.215 2738.895 3566.645 2739.000 ;
        RECT 21.355 2706.000 54.785 2706.105 ;
        RECT 55.565 2706.000 59.185 2706.160 ;
        RECT 59.945 2706.000 69.005 2706.085 ;
        RECT 69.775 2706.000 103.895 2706.160 ;
        RECT 105.420 2706.000 148.750 2706.085 ;
        RECT 164.275 2706.000 169.885 2706.120 ;
        RECT 174.985 2706.000 180.515 2706.120 ;
        RECT 0.295 2626.000 199.770 2706.000 ;
        RECT 21.355 2625.915 54.845 2626.000 ;
        RECT 29.910 2625.885 54.845 2625.915 ;
        RECT 55.565 2625.840 59.185 2626.000 ;
        RECT 59.850 2625.915 69.005 2626.000 ;
        RECT 69.775 2625.915 106.935 2626.000 ;
        RECT 107.930 2625.915 111.185 2626.000 ;
        RECT 119.395 2625.915 142.780 2626.000 ;
        RECT 191.005 2625.915 194.005 2626.000 ;
        RECT 59.850 2625.885 68.725 2625.915 ;
        RECT 69.780 2625.885 104.105 2625.915 ;
        RECT 3389.065 2582.845 3587.695 2593.390 ;
        RECT 3390.035 2581.965 3587.695 2582.845 ;
        RECT 3388.970 2580.955 3587.695 2581.965 ;
        RECT 3388.970 2524.270 3389.920 2580.955 ;
        RECT 3390.035 2524.270 3587.695 2580.955 ;
        RECT 3388.970 2523.320 3587.695 2524.270 ;
        RECT 3390.035 2521.145 3587.695 2523.320 ;
        RECT 0.305 2485.680 197.965 2487.855 ;
        RECT 0.305 2484.730 199.030 2485.680 ;
        RECT 0.305 2428.045 197.965 2484.730 ;
        RECT 198.080 2428.045 199.030 2484.730 ;
        RECT 0.305 2427.035 199.030 2428.045 ;
        RECT 0.305 2426.155 197.965 2427.035 ;
        RECT 0.305 2415.610 198.935 2426.155 ;
        RECT 3391.020 2299.245 3587.780 2373.760 ;
        RECT 0.220 2204.240 196.980 2278.755 ;
        RECT 3390.035 2140.935 3587.695 2151.930 ;
        RECT 3389.000 2139.955 3587.695 2140.935 ;
        RECT 3389.000 2083.240 3389.890 2139.955 ;
        RECT 3390.035 2083.240 3587.695 2139.955 ;
        RECT 3389.000 2082.350 3587.695 2083.240 ;
        RECT 3390.035 2080.225 3587.695 2082.350 ;
        RECT 21.355 2068.000 54.785 2068.105 ;
        RECT 55.565 2068.000 59.185 2068.160 ;
        RECT 59.945 2068.000 69.005 2068.085 ;
        RECT 69.775 2068.000 103.895 2068.160 ;
        RECT 105.420 2068.000 148.750 2068.085 ;
        RECT 164.275 2068.000 169.885 2068.120 ;
        RECT 174.985 2068.000 180.515 2068.120 ;
        RECT 0.295 1988.000 199.770 2068.000 ;
        RECT 21.355 1987.915 54.845 1988.000 ;
        RECT 29.910 1987.885 54.845 1987.915 ;
        RECT 55.565 1987.840 59.185 1988.000 ;
        RECT 59.850 1987.915 69.005 1988.000 ;
        RECT 69.775 1987.915 106.935 1988.000 ;
        RECT 107.930 1987.915 111.185 1988.000 ;
        RECT 119.395 1987.915 142.780 1988.000 ;
        RECT 191.005 1987.915 194.005 1988.000 ;
        RECT 59.850 1987.885 68.725 1987.915 ;
        RECT 69.780 1987.885 104.105 1987.915 ;
        RECT 3483.895 1933.085 3518.220 1933.115 ;
        RECT 3519.275 1933.085 3528.150 1933.115 ;
        RECT 3393.995 1933.000 3396.995 1933.085 ;
        RECT 3445.220 1933.000 3468.605 1933.085 ;
        RECT 3476.815 1933.000 3480.070 1933.085 ;
        RECT 3481.065 1933.000 3518.225 1933.085 ;
        RECT 3518.995 1933.000 3528.150 1933.085 ;
        RECT 3528.815 1933.000 3532.435 1933.160 ;
        RECT 3533.155 1933.085 3558.090 1933.115 ;
        RECT 3533.155 1933.000 3566.645 1933.085 ;
        RECT 3388.230 1853.000 3587.705 1933.000 ;
        RECT 3407.485 1852.880 3413.015 1853.000 ;
        RECT 3418.115 1852.880 3423.725 1853.000 ;
        RECT 3439.250 1852.915 3482.580 1853.000 ;
        RECT 3484.105 1852.840 3518.225 1853.000 ;
        RECT 3518.995 1852.915 3528.055 1853.000 ;
        RECT 3528.815 1852.840 3532.435 1853.000 ;
        RECT 3533.215 1852.895 3566.645 1853.000 ;
        RECT 21.355 1852.000 54.785 1852.105 ;
        RECT 55.565 1852.000 59.185 1852.160 ;
        RECT 59.945 1852.000 69.005 1852.085 ;
        RECT 69.775 1852.000 103.895 1852.160 ;
        RECT 105.420 1852.000 148.750 1852.085 ;
        RECT 164.275 1852.000 169.885 1852.120 ;
        RECT 174.985 1852.000 180.515 1852.120 ;
        RECT 0.295 1772.000 199.770 1852.000 ;
        RECT 21.355 1771.915 54.845 1772.000 ;
        RECT 29.910 1771.885 54.845 1771.915 ;
        RECT 55.565 1771.840 59.185 1772.000 ;
        RECT 59.850 1771.915 69.005 1772.000 ;
        RECT 69.775 1771.915 106.935 1772.000 ;
        RECT 107.930 1771.915 111.185 1772.000 ;
        RECT 119.395 1771.915 142.780 1772.000 ;
        RECT 191.005 1771.915 194.005 1772.000 ;
        RECT 59.850 1771.885 68.725 1771.915 ;
        RECT 69.780 1771.885 104.105 1771.915 ;
        RECT 3483.895 1707.085 3518.220 1707.115 ;
        RECT 3519.275 1707.085 3528.150 1707.115 ;
        RECT 3393.995 1707.000 3396.995 1707.085 ;
        RECT 3445.220 1707.000 3468.605 1707.085 ;
        RECT 3476.815 1707.000 3480.070 1707.085 ;
        RECT 3481.065 1707.000 3518.225 1707.085 ;
        RECT 3518.995 1707.000 3528.150 1707.085 ;
        RECT 3528.815 1707.000 3532.435 1707.160 ;
        RECT 3533.155 1707.085 3558.090 1707.115 ;
        RECT 3533.155 1707.000 3566.645 1707.085 ;
        RECT 21.355 1636.000 54.785 1636.105 ;
        RECT 55.565 1636.000 59.185 1636.160 ;
        RECT 59.945 1636.000 69.005 1636.085 ;
        RECT 69.775 1636.000 103.895 1636.160 ;
        RECT 105.420 1636.000 148.750 1636.085 ;
        RECT 164.275 1636.000 169.885 1636.120 ;
        RECT 174.985 1636.000 180.515 1636.120 ;
        RECT 0.295 1556.000 199.770 1636.000 ;
        RECT 3388.230 1627.000 3587.705 1707.000 ;
        RECT 3407.485 1626.880 3413.015 1627.000 ;
        RECT 3418.115 1626.880 3423.725 1627.000 ;
        RECT 3439.250 1626.915 3482.580 1627.000 ;
        RECT 3484.105 1626.840 3518.225 1627.000 ;
        RECT 3518.995 1626.915 3528.055 1627.000 ;
        RECT 3528.815 1626.840 3532.435 1627.000 ;
        RECT 3533.215 1626.895 3566.645 1627.000 ;
        RECT 21.355 1555.915 54.845 1556.000 ;
        RECT 29.910 1555.885 54.845 1555.915 ;
        RECT 55.565 1555.840 59.185 1556.000 ;
        RECT 59.850 1555.915 69.005 1556.000 ;
        RECT 69.775 1555.915 106.935 1556.000 ;
        RECT 107.930 1555.915 111.185 1556.000 ;
        RECT 119.395 1555.915 142.780 1556.000 ;
        RECT 191.005 1555.915 194.005 1556.000 ;
        RECT 59.850 1555.885 68.725 1555.915 ;
        RECT 69.780 1555.885 104.105 1555.915 ;
        RECT 3483.895 1482.085 3518.220 1482.115 ;
        RECT 3519.275 1482.085 3528.150 1482.115 ;
        RECT 3393.995 1482.000 3396.995 1482.085 ;
        RECT 3445.220 1482.000 3468.605 1482.085 ;
        RECT 3476.815 1482.000 3480.070 1482.085 ;
        RECT 3481.065 1482.000 3518.225 1482.085 ;
        RECT 3518.995 1482.000 3528.150 1482.085 ;
        RECT 3528.815 1482.000 3532.435 1482.160 ;
        RECT 3533.155 1482.085 3558.090 1482.115 ;
        RECT 3533.155 1482.000 3566.645 1482.085 ;
        RECT 21.355 1420.000 54.785 1420.105 ;
        RECT 55.565 1420.000 59.185 1420.160 ;
        RECT 59.945 1420.000 69.005 1420.085 ;
        RECT 69.775 1420.000 103.895 1420.160 ;
        RECT 105.420 1420.000 148.750 1420.085 ;
        RECT 164.275 1420.000 169.885 1420.120 ;
        RECT 174.985 1420.000 180.515 1420.120 ;
        RECT 0.295 1340.000 199.770 1420.000 ;
        RECT 3388.230 1402.000 3587.705 1482.000 ;
        RECT 3407.485 1401.880 3413.015 1402.000 ;
        RECT 3418.115 1401.880 3423.725 1402.000 ;
        RECT 3439.250 1401.915 3482.580 1402.000 ;
        RECT 3484.105 1401.840 3518.225 1402.000 ;
        RECT 3518.995 1401.915 3528.055 1402.000 ;
        RECT 3528.815 1401.840 3532.435 1402.000 ;
        RECT 3533.215 1401.895 3566.645 1402.000 ;
        RECT 21.355 1339.915 54.845 1340.000 ;
        RECT 29.910 1339.885 54.845 1339.915 ;
        RECT 55.565 1339.840 59.185 1340.000 ;
        RECT 59.850 1339.915 69.005 1340.000 ;
        RECT 69.775 1339.915 106.935 1340.000 ;
        RECT 107.930 1339.915 111.185 1340.000 ;
        RECT 119.395 1339.915 142.780 1340.000 ;
        RECT 191.005 1339.915 194.005 1340.000 ;
        RECT 59.850 1339.885 68.725 1339.915 ;
        RECT 69.780 1339.885 104.105 1339.915 ;
        RECT 3483.895 1257.085 3518.220 1257.115 ;
        RECT 3519.275 1257.085 3528.150 1257.115 ;
        RECT 3393.995 1257.000 3396.995 1257.085 ;
        RECT 3445.220 1257.000 3468.605 1257.085 ;
        RECT 3476.815 1257.000 3480.070 1257.085 ;
        RECT 3481.065 1257.000 3518.225 1257.085 ;
        RECT 3518.995 1257.000 3528.150 1257.085 ;
        RECT 3528.815 1257.000 3532.435 1257.160 ;
        RECT 3533.155 1257.085 3558.090 1257.115 ;
        RECT 3533.155 1257.000 3566.645 1257.085 ;
        RECT 21.355 1204.000 54.785 1204.105 ;
        RECT 55.565 1204.000 59.185 1204.160 ;
        RECT 59.945 1204.000 69.005 1204.085 ;
        RECT 69.775 1204.000 103.895 1204.160 ;
        RECT 105.420 1204.000 148.750 1204.085 ;
        RECT 164.275 1204.000 169.885 1204.120 ;
        RECT 174.985 1204.000 180.515 1204.120 ;
        RECT 0.295 1124.000 199.770 1204.000 ;
        RECT 3388.230 1177.000 3587.705 1257.000 ;
        RECT 3407.485 1176.880 3413.015 1177.000 ;
        RECT 3418.115 1176.880 3423.725 1177.000 ;
        RECT 3439.250 1176.915 3482.580 1177.000 ;
        RECT 3484.105 1176.840 3518.225 1177.000 ;
        RECT 3518.995 1176.915 3528.055 1177.000 ;
        RECT 3528.815 1176.840 3532.435 1177.000 ;
        RECT 3533.215 1176.895 3566.645 1177.000 ;
        RECT 21.355 1123.915 54.845 1124.000 ;
        RECT 29.910 1123.885 54.845 1123.915 ;
        RECT 55.565 1123.840 59.185 1124.000 ;
        RECT 59.850 1123.915 69.005 1124.000 ;
        RECT 69.775 1123.915 106.935 1124.000 ;
        RECT 107.930 1123.915 111.185 1124.000 ;
        RECT 119.395 1123.915 142.780 1124.000 ;
        RECT 191.005 1123.915 194.005 1124.000 ;
        RECT 59.850 1123.885 68.725 1123.915 ;
        RECT 69.780 1123.885 104.105 1123.915 ;
        RECT 3483.895 1031.085 3518.220 1031.115 ;
        RECT 3519.275 1031.085 3528.150 1031.115 ;
        RECT 3393.995 1031.000 3396.995 1031.085 ;
        RECT 3445.220 1031.000 3468.605 1031.085 ;
        RECT 3476.815 1031.000 3480.070 1031.085 ;
        RECT 3481.065 1031.000 3518.225 1031.085 ;
        RECT 3518.995 1031.000 3528.150 1031.085 ;
        RECT 3528.815 1031.000 3532.435 1031.160 ;
        RECT 3533.155 1031.085 3558.090 1031.115 ;
        RECT 3533.155 1031.000 3566.645 1031.085 ;
        RECT 21.355 988.000 54.785 988.105 ;
        RECT 55.565 988.000 59.185 988.160 ;
        RECT 59.945 988.000 69.005 988.085 ;
        RECT 69.775 988.000 103.895 988.160 ;
        RECT 105.420 988.000 148.750 988.085 ;
        RECT 164.275 988.000 169.885 988.120 ;
        RECT 174.985 988.000 180.515 988.120 ;
        RECT 0.295 908.000 199.770 988.000 ;
        RECT 3388.230 951.000 3587.705 1031.000 ;
        RECT 3407.485 950.880 3413.015 951.000 ;
        RECT 3418.115 950.880 3423.725 951.000 ;
        RECT 3439.250 950.915 3482.580 951.000 ;
        RECT 3484.105 950.840 3518.225 951.000 ;
        RECT 3518.995 950.915 3528.055 951.000 ;
        RECT 3528.815 950.840 3532.435 951.000 ;
        RECT 3533.215 950.895 3566.645 951.000 ;
        RECT 21.355 907.915 54.845 908.000 ;
        RECT 29.910 907.885 54.845 907.915 ;
        RECT 55.565 907.840 59.185 908.000 ;
        RECT 59.850 907.915 69.005 908.000 ;
        RECT 69.775 907.915 106.935 908.000 ;
        RECT 107.930 907.915 111.185 908.000 ;
        RECT 119.395 907.915 142.780 908.000 ;
        RECT 191.005 907.915 194.005 908.000 ;
        RECT 59.850 907.885 68.725 907.915 ;
        RECT 69.780 907.885 104.105 907.915 ;
        RECT 3483.895 806.085 3518.220 806.115 ;
        RECT 3519.275 806.085 3528.150 806.115 ;
        RECT 3393.995 806.000 3396.995 806.085 ;
        RECT 3445.220 806.000 3468.605 806.085 ;
        RECT 3476.815 806.000 3480.070 806.085 ;
        RECT 3481.065 806.000 3518.225 806.085 ;
        RECT 3518.995 806.000 3528.150 806.085 ;
        RECT 3528.815 806.000 3532.435 806.160 ;
        RECT 3533.155 806.085 3558.090 806.115 ;
        RECT 3533.155 806.000 3566.645 806.085 ;
        RECT 3388.230 726.000 3587.705 806.000 ;
        RECT 3407.485 725.880 3413.015 726.000 ;
        RECT 3418.115 725.880 3423.725 726.000 ;
        RECT 3439.250 725.915 3482.580 726.000 ;
        RECT 3484.105 725.840 3518.225 726.000 ;
        RECT 3518.995 725.915 3528.055 726.000 ;
        RECT 3528.815 725.840 3532.435 726.000 ;
        RECT 3533.215 725.895 3566.645 726.000 ;
        RECT 0.305 621.680 197.965 623.855 ;
        RECT 0.305 620.730 199.030 621.680 ;
        RECT 0.305 564.045 197.965 620.730 ;
        RECT 198.080 564.045 199.030 620.730 ;
        RECT 3483.895 580.085 3518.220 580.115 ;
        RECT 3519.275 580.085 3528.150 580.115 ;
        RECT 3393.995 580.000 3396.995 580.085 ;
        RECT 3445.220 580.000 3468.605 580.085 ;
        RECT 3476.815 580.000 3480.070 580.085 ;
        RECT 3481.065 580.000 3518.225 580.085 ;
        RECT 3518.995 580.000 3528.150 580.085 ;
        RECT 3528.815 580.000 3532.435 580.160 ;
        RECT 3533.155 580.085 3558.090 580.115 ;
        RECT 3533.155 580.000 3566.645 580.085 ;
        RECT 0.305 563.035 199.030 564.045 ;
        RECT 0.305 562.155 197.965 563.035 ;
        RECT 0.305 551.610 198.935 562.155 ;
        RECT 3388.230 500.000 3587.705 580.000 ;
        RECT 3407.485 499.880 3413.015 500.000 ;
        RECT 3418.115 499.880 3423.725 500.000 ;
        RECT 3439.250 499.915 3482.580 500.000 ;
        RECT 3484.105 499.840 3518.225 500.000 ;
        RECT 3518.995 499.915 3528.055 500.000 ;
        RECT 3528.815 499.840 3532.435 500.000 ;
        RECT 3533.215 499.895 3566.645 500.000 ;
        RECT 0.220 340.240 196.980 414.755 ;
        RECT 398.350 198.110 456.935 199.000 ;
        RECT 398.350 197.965 399.240 198.110 ;
        RECT 455.955 197.965 456.935 198.110 ;
        RECT 396.225 0.305 467.930 197.965 ;
        RECT 663.000 98.605 738.000 199.815 ;
        RECT 932.000 194.005 1012.000 199.770 ;
        RECT 932.000 191.005 1012.085 194.005 ;
        RECT 932.000 180.515 1012.000 191.005 ;
        RECT 931.880 174.985 1012.000 180.515 ;
        RECT 932.000 169.885 1012.000 174.985 ;
        RECT 931.880 164.275 1012.000 169.885 ;
        RECT 932.000 148.750 1012.000 164.275 ;
        RECT 931.915 142.780 1012.000 148.750 ;
        RECT 931.915 119.395 1012.085 142.780 ;
        RECT 931.915 111.185 1012.000 119.395 ;
        RECT 931.915 107.930 1012.085 111.185 ;
        RECT 931.915 106.935 1012.000 107.930 ;
        RECT 931.915 105.420 1012.085 106.935 ;
        RECT 932.000 104.105 1012.085 105.420 ;
        RECT 932.000 103.895 1012.115 104.105 ;
        RECT 663.000 69.775 738.265 98.605 ;
        RECT 931.840 69.780 1012.115 103.895 ;
        RECT 931.840 69.775 1012.085 69.780 ;
        RECT 663.000 59.185 738.000 69.775 ;
        RECT 932.000 69.005 1012.000 69.775 ;
        RECT 931.915 68.725 1012.085 69.005 ;
        RECT 931.915 59.945 1012.115 68.725 ;
        RECT 932.000 59.850 1012.115 59.945 ;
        RECT 932.000 59.185 1012.000 59.850 ;
        RECT 662.840 55.565 738.160 59.185 ;
        RECT 931.840 55.565 1012.160 59.185 ;
        RECT 663.000 0.780 738.000 55.565 ;
        RECT 932.000 54.845 1012.000 55.565 ;
        RECT 932.000 54.785 1012.115 54.845 ;
        RECT 931.895 29.910 1012.115 54.785 ;
        RECT 931.895 21.355 1012.085 29.910 ;
        RECT 932.000 0.295 1012.000 21.355 ;
        RECT 1206.245 0.220 1280.760 196.980 ;
        RECT 1475.000 194.005 1555.000 199.770 ;
        RECT 1749.000 194.005 1829.000 199.770 ;
        RECT 2023.000 194.005 2103.000 199.770 ;
        RECT 2297.000 194.005 2377.000 199.770 ;
        RECT 2571.000 194.005 2651.000 199.770 ;
        RECT 2849.350 198.110 2907.935 199.000 ;
        RECT 2849.350 197.965 2850.240 198.110 ;
        RECT 2906.955 197.965 2907.935 198.110 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.270 198.080 ;
        RECT 3175.955 197.965 3176.965 198.080 ;
        RECT 3177.845 197.965 3188.390 198.935 ;
        RECT 1475.000 191.005 1555.085 194.005 ;
        RECT 1749.000 191.005 1829.085 194.005 ;
        RECT 2023.000 191.005 2103.085 194.005 ;
        RECT 2297.000 191.005 2377.085 194.005 ;
        RECT 2571.000 191.005 2651.085 194.005 ;
        RECT 1475.000 180.515 1555.000 191.005 ;
        RECT 1749.000 180.515 1829.000 191.005 ;
        RECT 2023.000 180.515 2103.000 191.005 ;
        RECT 2297.000 180.515 2377.000 191.005 ;
        RECT 2571.000 180.515 2651.000 191.005 ;
        RECT 1474.880 174.985 1555.000 180.515 ;
        RECT 1748.880 174.985 1829.000 180.515 ;
        RECT 2022.880 174.985 2103.000 180.515 ;
        RECT 2296.880 174.985 2377.000 180.515 ;
        RECT 2570.880 174.985 2651.000 180.515 ;
        RECT 1475.000 169.885 1555.000 174.985 ;
        RECT 1749.000 169.885 1829.000 174.985 ;
        RECT 2023.000 169.885 2103.000 174.985 ;
        RECT 2297.000 169.885 2377.000 174.985 ;
        RECT 2571.000 169.885 2651.000 174.985 ;
        RECT 1474.880 164.275 1555.000 169.885 ;
        RECT 1748.880 164.275 1829.000 169.885 ;
        RECT 2022.880 164.275 2103.000 169.885 ;
        RECT 2296.880 164.275 2377.000 169.885 ;
        RECT 2570.880 164.275 2651.000 169.885 ;
        RECT 1475.000 148.750 1555.000 164.275 ;
        RECT 1749.000 148.750 1829.000 164.275 ;
        RECT 2023.000 148.750 2103.000 164.275 ;
        RECT 2297.000 148.750 2377.000 164.275 ;
        RECT 2571.000 148.750 2651.000 164.275 ;
        RECT 1474.915 142.780 1555.000 148.750 ;
        RECT 1748.915 142.780 1829.000 148.750 ;
        RECT 2022.915 142.780 2103.000 148.750 ;
        RECT 2296.915 142.780 2377.000 148.750 ;
        RECT 2570.915 142.780 2651.000 148.750 ;
        RECT 1474.915 119.395 1555.085 142.780 ;
        RECT 1748.915 119.395 1829.085 142.780 ;
        RECT 2022.915 119.395 2103.085 142.780 ;
        RECT 2296.915 119.395 2377.085 142.780 ;
        RECT 2570.915 119.395 2651.085 142.780 ;
        RECT 1474.915 111.185 1555.000 119.395 ;
        RECT 1748.915 111.185 1829.000 119.395 ;
        RECT 2022.915 111.185 2103.000 119.395 ;
        RECT 2296.915 111.185 2377.000 119.395 ;
        RECT 2570.915 111.185 2651.000 119.395 ;
        RECT 1474.915 107.930 1555.085 111.185 ;
        RECT 1748.915 107.930 1829.085 111.185 ;
        RECT 2022.915 107.930 2103.085 111.185 ;
        RECT 2296.915 107.930 2377.085 111.185 ;
        RECT 2570.915 107.930 2651.085 111.185 ;
        RECT 1474.915 106.935 1555.000 107.930 ;
        RECT 1748.915 106.935 1829.000 107.930 ;
        RECT 2022.915 106.935 2103.000 107.930 ;
        RECT 2296.915 106.935 2377.000 107.930 ;
        RECT 2570.915 106.935 2651.000 107.930 ;
        RECT 1474.915 105.420 1555.085 106.935 ;
        RECT 1748.915 105.420 1829.085 106.935 ;
        RECT 2022.915 105.420 2103.085 106.935 ;
        RECT 2296.915 105.420 2377.085 106.935 ;
        RECT 2570.915 105.420 2651.085 106.935 ;
        RECT 1475.000 104.105 1555.085 105.420 ;
        RECT 1749.000 104.105 1829.085 105.420 ;
        RECT 2023.000 104.105 2103.085 105.420 ;
        RECT 2297.000 104.105 2377.085 105.420 ;
        RECT 2571.000 104.105 2651.085 105.420 ;
        RECT 1475.000 103.895 1555.115 104.105 ;
        RECT 1749.000 103.895 1829.115 104.105 ;
        RECT 2023.000 103.895 2103.115 104.105 ;
        RECT 2297.000 103.895 2377.115 104.105 ;
        RECT 2571.000 103.895 2651.115 104.105 ;
        RECT 1474.840 69.780 1555.115 103.895 ;
        RECT 1748.840 69.780 1829.115 103.895 ;
        RECT 2022.840 69.780 2103.115 103.895 ;
        RECT 2296.840 69.780 2377.115 103.895 ;
        RECT 2570.840 69.780 2651.115 103.895 ;
        RECT 1474.840 69.775 1555.085 69.780 ;
        RECT 1748.840 69.775 1829.085 69.780 ;
        RECT 2022.840 69.775 2103.085 69.780 ;
        RECT 2296.840 69.775 2377.085 69.780 ;
        RECT 2570.840 69.775 2651.085 69.780 ;
        RECT 1475.000 69.005 1555.000 69.775 ;
        RECT 1749.000 69.005 1829.000 69.775 ;
        RECT 2023.000 69.005 2103.000 69.775 ;
        RECT 2297.000 69.005 2377.000 69.775 ;
        RECT 2571.000 69.005 2651.000 69.775 ;
        RECT 1474.915 68.725 1555.085 69.005 ;
        RECT 1748.915 68.725 1829.085 69.005 ;
        RECT 2022.915 68.725 2103.085 69.005 ;
        RECT 2296.915 68.725 2377.085 69.005 ;
        RECT 2570.915 68.725 2651.085 69.005 ;
        RECT 1474.915 59.945 1555.115 68.725 ;
        RECT 1748.915 59.945 1829.115 68.725 ;
        RECT 2022.915 59.945 2103.115 68.725 ;
        RECT 2296.915 59.945 2377.115 68.725 ;
        RECT 2570.915 59.945 2651.115 68.725 ;
        RECT 1475.000 59.850 1555.115 59.945 ;
        RECT 1749.000 59.850 1829.115 59.945 ;
        RECT 2023.000 59.850 2103.115 59.945 ;
        RECT 2297.000 59.850 2377.115 59.945 ;
        RECT 2571.000 59.850 2651.115 59.945 ;
        RECT 1475.000 59.185 1555.000 59.850 ;
        RECT 1749.000 59.185 1829.000 59.850 ;
        RECT 2023.000 59.185 2103.000 59.850 ;
        RECT 2297.000 59.185 2377.000 59.850 ;
        RECT 2571.000 59.185 2651.000 59.850 ;
        RECT 1474.840 55.565 1555.160 59.185 ;
        RECT 1748.840 55.565 1829.160 59.185 ;
        RECT 2022.840 55.565 2103.160 59.185 ;
        RECT 2296.840 55.565 2377.160 59.185 ;
        RECT 2570.840 55.565 2651.160 59.185 ;
        RECT 1475.000 54.845 1555.000 55.565 ;
        RECT 1749.000 54.845 1829.000 55.565 ;
        RECT 2023.000 54.845 2103.000 55.565 ;
        RECT 2297.000 54.845 2377.000 55.565 ;
        RECT 2571.000 54.845 2651.000 55.565 ;
        RECT 1475.000 54.785 1555.115 54.845 ;
        RECT 1749.000 54.785 1829.115 54.845 ;
        RECT 2023.000 54.785 2103.115 54.845 ;
        RECT 2297.000 54.785 2377.115 54.845 ;
        RECT 2571.000 54.785 2651.115 54.845 ;
        RECT 1474.895 29.910 1555.115 54.785 ;
        RECT 1748.895 29.910 1829.115 54.785 ;
        RECT 2022.895 29.910 2103.115 54.785 ;
        RECT 2296.895 29.910 2377.115 54.785 ;
        RECT 2570.895 29.910 2651.115 54.785 ;
        RECT 1474.895 21.355 1555.085 29.910 ;
        RECT 1748.895 21.355 1829.085 29.910 ;
        RECT 2022.895 21.355 2103.085 29.910 ;
        RECT 2296.895 21.355 2377.085 29.910 ;
        RECT 2570.895 21.355 2651.085 29.910 ;
        RECT 1475.000 0.295 1555.000 21.355 ;
        RECT 1749.000 0.295 1829.000 21.355 ;
        RECT 2023.000 0.295 2103.000 21.355 ;
        RECT 2297.000 0.295 2377.000 21.355 ;
        RECT 2571.000 0.295 2651.000 21.355 ;
        RECT 2847.225 0.305 2918.930 197.965 ;
        RECT 3116.145 0.305 3188.390 197.965 ;
      LAYER met1 ;
        RECT 385.250 5034.255 451.440 5036.855 ;
        RECT 642.250 5034.255 708.440 5036.855 ;
        RECT 899.250 5034.255 965.440 5036.855 ;
        RECT 1152.185 4990.035 1224.915 5187.725 ;
        RECT 1410.185 4990.035 1482.915 5187.725 ;
        RECT 1667.185 4990.035 1740.620 5187.725 ;
        RECT 1923.250 5034.255 1989.440 5036.855 ;
        RECT 2368.250 5034.255 2434.440 5036.855 ;
        RECT 2625.250 5034.255 2691.440 5036.855 ;
        RECT 2878.185 4990.035 2951.620 5187.725 ;
        RECT 3134.250 5034.255 3200.440 5036.855 ;
        RECT 1155.625 4989.130 1160.855 4990.035 ;
        RECT 1164.035 4989.920 1165.350 4990.035 ;
        POLYGON 1165.350 4990.035 1165.465 4989.920 1165.350 4989.920 ;
        POLYGON 1221.540 4990.035 1221.540 4989.920 1221.425 4989.920 ;
        RECT 1221.540 4989.920 1222.680 4990.035 ;
        RECT 1164.035 4988.970 1222.680 4989.920 ;
        RECT 1413.625 4989.130 1418.855 4990.035 ;
        RECT 1422.035 4989.920 1423.350 4990.035 ;
        POLYGON 1423.350 4990.035 1423.465 4989.920 1423.350 4989.920 ;
        POLYGON 1479.540 4990.035 1479.540 4989.920 1479.425 4989.920 ;
        RECT 1479.540 4989.920 1480.680 4990.035 ;
        RECT 1422.035 4988.970 1480.680 4989.920 ;
        RECT 1679.035 4989.920 1680.350 4990.035 ;
        POLYGON 1680.350 4990.035 1680.465 4989.920 1680.350 4989.920 ;
        POLYGON 1736.540 4990.035 1736.540 4989.920 1736.425 4989.920 ;
        RECT 1736.540 4989.920 1737.680 4990.035 ;
        RECT 1679.035 4988.970 1737.680 4989.920 ;
        RECT 2890.035 4989.920 2891.350 4990.035 ;
        POLYGON 2891.350 4990.035 2891.465 4989.920 2891.350 4989.920 ;
        POLYGON 2947.540 4990.035 2947.540 4989.920 2947.425 4989.920 ;
        RECT 2947.540 4989.920 2948.680 4990.035 ;
        RECT 2890.035 4988.970 2948.680 4989.920 ;
      LAYER met1 ;
        RECT 2925.210 4981.920 2925.530 4981.980 ;
        RECT 3373.710 4981.920 3374.030 4981.980 ;
        RECT 2925.210 4981.780 3374.030 4981.920 ;
        RECT 2925.210 4981.720 2925.530 4981.780 ;
        RECT 3373.710 4981.720 3374.030 4981.780 ;
        RECT 1780.270 4954.380 1780.590 4954.440 ;
        RECT 3367.730 4954.380 3368.050 4954.440 ;
        RECT 1780.270 4954.240 3368.050 4954.380 ;
        RECT 1780.270 4954.180 1780.590 4954.240 ;
        RECT 3367.730 4954.180 3368.050 4954.240 ;
        RECT 211.210 4950.980 211.530 4951.040 ;
        RECT 211.210 4950.840 262.270 4950.980 ;
        RECT 211.210 4950.780 211.530 4950.840 ;
        RECT 224.550 4950.440 224.870 4950.700 ;
        RECT 262.130 4950.640 262.270 4950.840 ;
        RECT 1718.170 4950.640 1718.490 4950.700 ;
        RECT 1780.270 4950.640 1780.590 4950.700 ;
        RECT 262.130 4950.500 1780.590 4950.640 ;
        RECT 1718.170 4950.440 1718.490 4950.500 ;
        RECT 1780.270 4950.440 1780.590 4950.500 ;
        RECT 224.640 4950.300 224.780 4950.440 ;
        RECT 3367.270 4950.300 3367.590 4950.360 ;
        RECT 224.640 4950.160 3367.590 4950.300 ;
        RECT 3367.270 4950.100 3367.590 4950.160 ;
      LAYER met1 ;
        RECT 151.145 4775.250 153.745 4841.440 ;
        RECT 3390.035 4834.375 3587.725 4837.815 ;
        RECT 3389.130 4829.145 3587.725 4834.375 ;
        RECT 3390.035 4825.965 3587.725 4829.145 ;
        RECT 3388.970 4824.650 3587.725 4825.965 ;
        RECT 3388.970 4768.460 3389.920 4824.650 ;
        POLYGON 3389.920 4824.650 3390.035 4824.650 3389.920 4824.535 ;
        POLYGON 3389.920 4768.575 3390.035 4768.460 3389.920 4768.460 ;
        RECT 3390.035 4768.460 3587.725 4824.650 ;
        RECT 3388.970 4767.320 3587.725 4768.460 ;
        RECT 3390.035 4765.085 3587.725 4767.320 ;
        RECT 122.615 4641.935 204.885 4645.935 ;
        POLYGON 204.885 4645.935 208.885 4641.935 204.885 4641.935 ;
        RECT 122.615 4636.200 208.885 4641.935 ;
        RECT 0.160 4616.565 197.965 4635.000 ;
        RECT 198.780 4616.565 208.885 4636.200 ;
        RECT 0.160 4580.925 208.885 4616.565 ;
        RECT 3390.035 4596.345 3587.840 4612.880 ;
        RECT 3390.000 4592.075 3587.840 4596.345 ;
        RECT 0.160 4576.655 198.000 4580.925 ;
        RECT 0.160 4560.120 197.965 4576.655 ;
        RECT 3379.115 4556.435 3587.840 4592.075 ;
        RECT 3379.115 4536.800 3389.220 4556.435 ;
        RECT 3390.035 4538.000 3587.840 4556.435 ;
        RECT 3379.115 4531.065 3465.385 4536.800 ;
        POLYGON 3379.115 4531.065 3383.115 4531.065 3383.115 4527.065 ;
        RECT 3383.115 4527.065 3465.385 4531.065 ;
        RECT 0.275 4419.680 197.965 4421.915 ;
        RECT 0.275 4418.540 199.030 4419.680 ;
        RECT 0.275 4362.350 197.965 4418.540 ;
        POLYGON 197.965 4418.540 198.080 4418.540 198.080 4418.425 ;
        POLYGON 198.080 4362.465 198.080 4362.350 197.965 4362.350 ;
        RECT 198.080 4362.350 199.030 4418.540 ;
        RECT 3445.190 4392.000 3468.635 4392.115 ;
        RECT 3477.750 4392.000 3479.480 4392.145 ;
        RECT 3483.895 4392.000 3518.220 4392.115 ;
        RECT 3519.275 4392.000 3558.090 4392.115 ;
      LAYER met1 ;
        RECT 3367.730 4372.640 3368.050 4372.700 ;
        RECT 3376.930 4372.640 3377.250 4372.700 ;
        RECT 3367.730 4372.500 3377.250 4372.640 ;
        RECT 3367.730 4372.440 3368.050 4372.500 ;
        RECT 3376.930 4372.440 3377.250 4372.500 ;
      LAYER met1 ;
        RECT 0.275 4361.035 199.030 4362.350 ;
      LAYER met1 ;
        RECT 3367.270 4362.100 3367.590 4362.160 ;
        RECT 3368.190 4362.100 3368.510 4362.160 ;
        RECT 3376.930 4362.100 3377.250 4362.160 ;
        RECT 3367.270 4361.960 3377.250 4362.100 ;
        RECT 3367.270 4361.900 3367.590 4361.960 ;
        RECT 3368.190 4361.900 3368.510 4361.960 ;
        RECT 3376.930 4361.900 3377.250 4361.960 ;
      LAYER met1 ;
        RECT 0.275 4357.855 197.965 4361.035 ;
        RECT 0.275 4352.625 198.870 4357.855 ;
        RECT 0.275 4349.185 197.965 4352.625 ;
      LAYER met1 ;
        RECT 3369.110 4350.880 3369.430 4350.940 ;
        RECT 3376.930 4350.880 3377.250 4350.940 ;
        RECT 3369.110 4350.740 3377.250 4350.880 ;
        RECT 3369.110 4350.680 3369.430 4350.740 ;
        RECT 3376.930 4350.680 3377.250 4350.740 ;
        RECT 3367.270 4321.300 3367.590 4321.360 ;
        RECT 3376.930 4321.300 3377.250 4321.360 ;
        RECT 3367.270 4321.160 3377.250 4321.300 ;
        RECT 3367.270 4321.100 3367.590 4321.160 ;
        RECT 3376.930 4321.100 3377.250 4321.160 ;
        RECT 3369.110 4316.200 3369.430 4316.260 ;
        RECT 3376.930 4316.200 3377.250 4316.260 ;
        RECT 3369.110 4316.060 3377.250 4316.200 ;
        RECT 3369.110 4316.000 3369.430 4316.060 ;
        RECT 3376.930 4316.000 3377.250 4316.060 ;
      LAYER met1 ;
        RECT 3381.155 4312.000 3588.000 4392.000 ;
        RECT 3407.485 4311.885 3413.015 4312.000 ;
        RECT 3418.120 4311.885 3423.725 4312.000 ;
        RECT 3439.220 4311.940 3482.580 4312.000 ;
        RECT 3439.220 4311.885 3460.930 4311.940 ;
        POLYGON 3460.930 4311.940 3460.985 4311.940 3460.930 4311.885 ;
        RECT 3483.895 4311.855 3518.220 4312.000 ;
        RECT 3519.275 4311.855 3558.090 4312.000 ;
        RECT 3566.900 4311.980 3568.975 4312.000 ;
        RECT 0.275 4208.680 197.965 4211.620 ;
        RECT 0.275 4207.540 199.030 4208.680 ;
        RECT 0.275 4151.350 197.965 4207.540 ;
        POLYGON 197.965 4207.540 198.080 4207.540 198.080 4207.425 ;
        POLYGON 198.080 4151.465 198.080 4151.350 197.965 4151.350 ;
        RECT 198.080 4151.350 199.030 4207.540 ;
        RECT 3390.035 4163.375 3587.725 4166.815 ;
        RECT 3389.130 4158.145 3587.725 4163.375 ;
        RECT 3390.035 4154.965 3587.725 4158.145 ;
        RECT 0.275 4150.035 199.030 4151.350 ;
        RECT 3388.970 4153.650 3587.725 4154.965 ;
        RECT 0.275 4138.185 197.965 4150.035 ;
        RECT 3388.970 4097.460 3389.920 4153.650 ;
        POLYGON 3389.920 4153.650 3390.035 4153.650 3389.920 4153.535 ;
        POLYGON 3389.920 4097.575 3390.035 4097.460 3389.920 4097.460 ;
        RECT 3390.035 4097.460 3587.725 4153.650 ;
        RECT 3388.970 4096.320 3587.725 4097.460 ;
        RECT 3390.035 4094.085 3587.725 4096.320 ;
      LAYER met1 ;
        RECT 3376.470 4091.800 3376.790 4091.860 ;
        RECT 3387.970 4091.800 3388.290 4091.860 ;
        RECT 3376.470 4091.660 3388.290 4091.800 ;
        RECT 3376.470 4091.600 3376.790 4091.660 ;
        RECT 3387.970 4091.600 3388.290 4091.660 ;
      LAYER met1 ;
        RECT 19.025 4002.000 21.100 4002.020 ;
        RECT 29.910 4002.000 68.725 4002.145 ;
        RECT 69.780 4002.000 104.105 4002.145 ;
        POLYGON 127.070 4002.115 127.070 4002.060 127.015 4002.060 ;
        RECT 127.070 4002.060 148.780 4002.115 ;
        RECT 105.420 4002.000 148.780 4002.060 ;
        RECT 164.275 4002.000 169.880 4002.115 ;
        RECT 174.985 4002.000 180.515 4002.115 ;
        RECT 0.000 3922.000 206.845 4002.000 ;
      LAYER met1 ;
        RECT 208.910 3988.780 209.230 3988.840 ;
        RECT 213.050 3988.780 213.370 3988.840 ;
        RECT 208.910 3988.640 213.370 3988.780 ;
        RECT 208.910 3988.580 209.230 3988.640 ;
        RECT 213.050 3988.580 213.370 3988.640 ;
        RECT 208.910 3956.820 209.230 3956.880 ;
        RECT 212.130 3956.820 212.450 3956.880 ;
        RECT 208.910 3956.680 212.450 3956.820 ;
        RECT 208.910 3956.620 209.230 3956.680 ;
        RECT 212.130 3956.620 212.450 3956.680 ;
      LAYER met1 ;
        RECT 3445.190 3946.000 3468.635 3946.115 ;
        RECT 3477.750 3946.000 3479.480 3946.145 ;
        RECT 3483.895 3946.000 3518.220 3946.115 ;
        RECT 3519.275 3946.000 3558.090 3946.115 ;
      LAYER met1 ;
        RECT 208.910 3941.520 209.230 3941.580 ;
        RECT 211.670 3941.520 211.990 3941.580 ;
        RECT 208.910 3941.380 211.990 3941.520 ;
        RECT 208.910 3941.320 209.230 3941.380 ;
        RECT 211.670 3941.320 211.990 3941.380 ;
        RECT 208.910 3936.220 209.230 3936.480 ;
        RECT 209.000 3935.400 209.140 3936.220 ;
        RECT 211.210 3935.400 211.530 3935.460 ;
        RECT 209.000 3935.260 211.530 3935.400 ;
        RECT 211.210 3935.200 211.530 3935.260 ;
        RECT 211.670 3935.060 211.990 3935.120 ;
        RECT 212.590 3935.060 212.910 3935.120 ;
        RECT 211.670 3934.920 212.910 3935.060 ;
        RECT 211.670 3934.860 211.990 3934.920 ;
        RECT 212.590 3934.860 212.910 3934.920 ;
        RECT 3367.730 3928.600 3368.050 3928.660 ;
        RECT 3376.930 3928.600 3377.250 3928.660 ;
        RECT 3367.730 3928.460 3377.250 3928.600 ;
        RECT 3367.730 3928.400 3368.050 3928.460 ;
        RECT 3376.930 3928.400 3377.250 3928.460 ;
      LAYER met1 ;
        RECT 29.910 3921.885 68.725 3922.000 ;
        RECT 69.780 3921.885 104.105 3922.000 ;
        RECT 108.520 3921.855 110.250 3922.000 ;
        RECT 119.365 3921.885 142.810 3922.000 ;
      LAYER met1 ;
        RECT 3368.190 3911.600 3368.510 3911.660 ;
        RECT 3376.930 3911.600 3377.250 3911.660 ;
        RECT 3368.190 3911.460 3377.250 3911.600 ;
        RECT 3368.190 3911.400 3368.510 3911.460 ;
        RECT 3376.930 3911.400 3377.250 3911.460 ;
        RECT 3376.010 3905.140 3376.330 3905.200 ;
        RECT 3376.930 3905.140 3377.250 3905.200 ;
        RECT 3376.010 3905.000 3377.250 3905.140 ;
        RECT 3376.010 3904.940 3376.330 3905.000 ;
        RECT 3376.930 3904.940 3377.250 3905.000 ;
        RECT 3367.270 3879.300 3367.590 3879.360 ;
        RECT 3376.930 3879.300 3377.250 3879.360 ;
        RECT 3367.270 3879.160 3377.250 3879.300 ;
        RECT 3367.270 3879.100 3367.590 3879.160 ;
        RECT 3376.930 3879.100 3377.250 3879.160 ;
      LAYER met1 ;
        RECT 3381.155 3866.000 3588.000 3946.000 ;
        RECT 3407.485 3865.885 3413.015 3866.000 ;
        RECT 3418.120 3865.885 3423.725 3866.000 ;
        RECT 3439.220 3865.940 3482.580 3866.000 ;
        RECT 3439.220 3865.885 3460.930 3865.940 ;
        POLYGON 3460.930 3865.940 3460.985 3865.940 3460.930 3865.885 ;
        RECT 3483.895 3865.855 3518.220 3866.000 ;
        RECT 3519.275 3865.855 3558.090 3866.000 ;
        RECT 3566.900 3865.980 3568.975 3866.000 ;
      LAYER met1 ;
        RECT 211.210 3788.180 211.530 3788.240 ;
        RECT 213.970 3788.180 214.290 3788.240 ;
        RECT 211.210 3788.040 214.290 3788.180 ;
        RECT 211.210 3787.980 211.530 3788.040 ;
        RECT 213.970 3787.980 214.290 3788.040 ;
        RECT 211.670 3787.840 211.990 3787.900 ;
        RECT 213.510 3787.840 213.830 3787.900 ;
        RECT 211.670 3787.700 213.830 3787.840 ;
        RECT 211.670 3787.640 211.990 3787.700 ;
        RECT 213.510 3787.640 213.830 3787.700 ;
      LAYER met1 ;
        RECT 19.025 3786.000 21.100 3786.020 ;
        RECT 29.910 3786.000 68.725 3786.145 ;
        RECT 69.780 3786.000 104.105 3786.145 ;
        POLYGON 127.070 3786.115 127.070 3786.060 127.015 3786.060 ;
        RECT 127.070 3786.060 148.780 3786.115 ;
        RECT 105.420 3786.000 148.780 3786.060 ;
        RECT 164.275 3786.000 169.880 3786.115 ;
        RECT 174.985 3786.000 180.515 3786.115 ;
        RECT 0.000 3706.000 206.845 3786.000 ;
      LAYER met1 ;
        RECT 208.910 3777.300 209.230 3777.360 ;
        RECT 213.050 3777.300 213.370 3777.360 ;
        RECT 208.910 3777.160 213.370 3777.300 ;
        RECT 208.910 3777.100 209.230 3777.160 ;
        RECT 213.050 3777.100 213.370 3777.160 ;
        RECT 208.910 3738.540 209.230 3738.600 ;
        RECT 213.510 3738.540 213.830 3738.600 ;
        RECT 208.910 3738.400 213.830 3738.540 ;
        RECT 208.910 3738.340 209.230 3738.400 ;
        RECT 213.510 3738.340 213.830 3738.400 ;
      LAYER met1 ;
        RECT 3445.190 3721.000 3468.635 3721.115 ;
        RECT 3477.750 3721.000 3479.480 3721.145 ;
        RECT 3483.895 3721.000 3518.220 3721.115 ;
        RECT 3519.275 3721.000 3558.090 3721.115 ;
      LAYER met1 ;
        RECT 208.910 3720.180 209.230 3720.240 ;
        RECT 213.970 3720.180 214.290 3720.240 ;
        RECT 208.910 3720.040 214.290 3720.180 ;
        RECT 208.910 3719.980 209.230 3720.040 ;
        RECT 213.970 3719.980 214.290 3720.040 ;
      LAYER met1 ;
        RECT 29.910 3705.885 68.725 3706.000 ;
        RECT 69.780 3705.885 104.105 3706.000 ;
        RECT 108.520 3705.855 110.250 3706.000 ;
        RECT 119.365 3705.885 142.810 3706.000 ;
      LAYER met1 ;
        RECT 3367.730 3701.820 3368.050 3701.880 ;
        RECT 3369.110 3701.820 3369.430 3701.880 ;
        RECT 3376.930 3701.820 3377.250 3701.880 ;
        RECT 3367.730 3701.680 3377.250 3701.820 ;
        RECT 3367.730 3701.620 3368.050 3701.680 ;
        RECT 3369.110 3701.620 3369.430 3701.680 ;
        RECT 3376.930 3701.620 3377.250 3701.680 ;
        RECT 3368.190 3690.600 3368.510 3690.660 ;
        RECT 3376.930 3690.600 3377.250 3690.660 ;
        RECT 3368.190 3690.460 3377.250 3690.600 ;
        RECT 3368.190 3690.400 3368.510 3690.460 ;
        RECT 3376.930 3690.400 3377.250 3690.460 ;
        RECT 3367.270 3654.560 3367.590 3654.620 ;
        RECT 3370.030 3654.560 3370.350 3654.620 ;
        RECT 3376.930 3654.560 3377.250 3654.620 ;
        RECT 3367.270 3654.420 3377.250 3654.560 ;
        RECT 3367.270 3654.360 3367.590 3654.420 ;
        RECT 3370.030 3654.360 3370.350 3654.420 ;
        RECT 3376.930 3654.360 3377.250 3654.420 ;
      LAYER met1 ;
        RECT 3381.155 3641.000 3588.000 3721.000 ;
        RECT 3407.485 3640.885 3413.015 3641.000 ;
        RECT 3418.120 3640.885 3423.725 3641.000 ;
        RECT 3439.220 3640.940 3482.580 3641.000 ;
        RECT 3439.220 3640.885 3460.930 3640.940 ;
        POLYGON 3460.930 3640.940 3460.985 3640.940 3460.930 3640.885 ;
        RECT 3483.895 3640.855 3518.220 3641.000 ;
        RECT 3519.275 3640.855 3558.090 3641.000 ;
        RECT 3566.900 3640.980 3568.975 3641.000 ;
        RECT 19.025 3570.000 21.100 3570.020 ;
        RECT 29.910 3570.000 68.725 3570.145 ;
        RECT 69.780 3570.000 104.105 3570.145 ;
        POLYGON 127.070 3570.115 127.070 3570.060 127.015 3570.060 ;
        RECT 127.070 3570.060 148.780 3570.115 ;
        RECT 105.420 3570.000 148.780 3570.060 ;
        RECT 164.275 3570.000 169.880 3570.115 ;
        RECT 174.985 3570.000 180.515 3570.115 ;
        RECT 0.000 3490.000 206.845 3570.000 ;
      LAYER met1 ;
        RECT 208.910 3561.400 209.230 3561.460 ;
        RECT 213.050 3561.400 213.370 3561.460 ;
        RECT 208.910 3561.260 213.370 3561.400 ;
        RECT 208.910 3561.200 209.230 3561.260 ;
        RECT 213.050 3561.200 213.370 3561.260 ;
        RECT 208.910 3519.920 209.230 3519.980 ;
        RECT 212.130 3519.920 212.450 3519.980 ;
        RECT 213.510 3519.920 213.830 3519.980 ;
        RECT 208.910 3519.780 213.830 3519.920 ;
        RECT 208.910 3519.720 209.230 3519.780 ;
        RECT 212.130 3519.720 212.450 3519.780 ;
        RECT 213.510 3519.720 213.830 3519.780 ;
        RECT 208.910 3504.280 209.230 3504.340 ;
        RECT 213.050 3504.280 213.370 3504.340 ;
        RECT 208.910 3504.140 213.370 3504.280 ;
        RECT 208.910 3504.080 209.230 3504.140 ;
        RECT 213.050 3504.080 213.370 3504.140 ;
      LAYER met1 ;
        RECT 3445.190 3496.000 3468.635 3496.115 ;
        RECT 3477.750 3496.000 3479.480 3496.145 ;
        RECT 3483.895 3496.000 3518.220 3496.115 ;
        RECT 3519.275 3496.000 3558.090 3496.115 ;
        RECT 29.910 3489.885 68.725 3490.000 ;
        RECT 69.780 3489.885 104.105 3490.000 ;
        RECT 108.520 3489.855 110.250 3490.000 ;
        RECT 119.365 3489.885 142.810 3490.000 ;
      LAYER met1 ;
        RECT 3367.270 3476.740 3367.590 3476.800 ;
        RECT 3369.110 3476.740 3369.430 3476.800 ;
        RECT 3376.930 3476.740 3377.250 3476.800 ;
        RECT 3367.270 3476.600 3377.250 3476.740 ;
        RECT 3367.270 3476.540 3367.590 3476.600 ;
        RECT 3369.110 3476.540 3369.430 3476.600 ;
        RECT 3376.930 3476.540 3377.250 3476.600 ;
        RECT 3369.570 3461.440 3369.890 3461.500 ;
        RECT 3376.930 3461.440 3377.250 3461.500 ;
        RECT 3369.570 3461.300 3377.250 3461.440 ;
        RECT 3369.570 3461.240 3369.890 3461.300 ;
        RECT 3376.930 3461.240 3377.250 3461.300 ;
        RECT 3367.730 3426.080 3368.050 3426.140 ;
        RECT 3370.030 3426.080 3370.350 3426.140 ;
        RECT 3376.930 3426.080 3377.250 3426.140 ;
        RECT 3367.730 3425.940 3377.250 3426.080 ;
        RECT 3367.730 3425.880 3368.050 3425.940 ;
        RECT 3370.030 3425.880 3370.350 3425.940 ;
        RECT 3376.930 3425.880 3377.250 3425.940 ;
      LAYER met1 ;
        RECT 3381.155 3416.000 3588.000 3496.000 ;
        RECT 3407.485 3415.885 3413.015 3416.000 ;
        RECT 3418.120 3415.885 3423.725 3416.000 ;
        RECT 3439.220 3415.940 3482.580 3416.000 ;
        RECT 3439.220 3415.885 3460.930 3415.940 ;
        POLYGON 3460.930 3415.940 3460.985 3415.940 3460.930 3415.885 ;
        RECT 3483.895 3415.855 3518.220 3416.000 ;
        RECT 3519.275 3415.855 3558.090 3416.000 ;
        RECT 3566.900 3415.980 3568.975 3416.000 ;
        RECT 19.025 3354.000 21.100 3354.020 ;
        RECT 29.910 3354.000 68.725 3354.145 ;
        RECT 69.780 3354.000 104.105 3354.145 ;
        POLYGON 127.070 3354.115 127.070 3354.060 127.015 3354.060 ;
        RECT 127.070 3354.060 148.780 3354.115 ;
        RECT 105.420 3354.000 148.780 3354.060 ;
        RECT 164.275 3354.000 169.880 3354.115 ;
        RECT 174.985 3354.000 180.515 3354.115 ;
        RECT 0.000 3274.000 206.845 3354.000 ;
      LAYER met1 ;
        RECT 208.910 3340.740 209.230 3340.800 ;
        RECT 212.590 3340.740 212.910 3340.800 ;
        RECT 208.910 3340.600 212.910 3340.740 ;
        RECT 208.910 3340.540 209.230 3340.600 ;
        RECT 212.590 3340.540 212.910 3340.600 ;
        RECT 208.910 3305.380 209.230 3305.440 ;
        RECT 212.130 3305.380 212.450 3305.440 ;
        RECT 208.910 3305.240 212.450 3305.380 ;
        RECT 208.910 3305.180 209.230 3305.240 ;
        RECT 212.130 3305.180 212.450 3305.240 ;
        RECT 208.910 3293.480 209.230 3293.540 ;
        RECT 213.050 3293.480 213.370 3293.540 ;
        RECT 208.910 3293.340 213.370 3293.480 ;
        RECT 208.910 3293.280 209.230 3293.340 ;
        RECT 213.050 3293.280 213.370 3293.340 ;
      LAYER met1 ;
        RECT 29.910 3273.885 68.725 3274.000 ;
        RECT 69.780 3273.885 104.105 3274.000 ;
        RECT 108.520 3273.855 110.250 3274.000 ;
        RECT 119.365 3273.885 142.810 3274.000 ;
        RECT 3445.190 3270.000 3468.635 3270.115 ;
        RECT 3477.750 3270.000 3479.480 3270.145 ;
        RECT 3483.895 3270.000 3518.220 3270.115 ;
        RECT 3519.275 3270.000 3558.090 3270.115 ;
      LAYER met1 ;
        RECT 3367.270 3252.680 3367.590 3252.740 ;
        RECT 3376.930 3252.680 3377.250 3252.740 ;
        RECT 3367.270 3252.540 3377.250 3252.680 ;
        RECT 3367.270 3252.480 3367.590 3252.540 ;
        RECT 3376.930 3252.480 3377.250 3252.540 ;
        RECT 3367.270 3236.020 3367.590 3236.080 ;
        RECT 3368.190 3236.020 3368.510 3236.080 ;
        RECT 3367.270 3235.880 3368.510 3236.020 ;
        RECT 3367.270 3235.820 3367.590 3235.880 ;
        RECT 3368.190 3235.820 3368.510 3235.880 ;
        RECT 3367.270 3235.340 3367.590 3235.400 ;
        RECT 3369.570 3235.340 3369.890 3235.400 ;
        RECT 3376.930 3235.340 3377.250 3235.400 ;
        RECT 3367.270 3235.200 3377.250 3235.340 ;
        RECT 3367.270 3235.140 3367.590 3235.200 ;
        RECT 3369.570 3235.140 3369.890 3235.200 ;
        RECT 3376.930 3235.140 3377.250 3235.200 ;
        RECT 3376.010 3228.880 3376.330 3228.940 ;
        RECT 3376.930 3228.880 3377.250 3228.940 ;
        RECT 3376.010 3228.740 3377.250 3228.880 ;
        RECT 3376.010 3228.680 3376.330 3228.740 ;
        RECT 3376.930 3228.680 3377.250 3228.740 ;
        RECT 3367.730 3203.380 3368.050 3203.440 ;
        RECT 3376.930 3203.380 3377.250 3203.440 ;
        RECT 3367.730 3203.240 3377.250 3203.380 ;
        RECT 3367.730 3203.180 3368.050 3203.240 ;
        RECT 3376.930 3203.180 3377.250 3203.240 ;
      LAYER met1 ;
        RECT 3381.155 3190.000 3588.000 3270.000 ;
        RECT 3407.485 3189.885 3413.015 3190.000 ;
        RECT 3418.120 3189.885 3423.725 3190.000 ;
        RECT 3439.220 3189.940 3482.580 3190.000 ;
        RECT 3439.220 3189.885 3460.930 3189.940 ;
        POLYGON 3460.930 3189.940 3460.985 3189.940 3460.930 3189.885 ;
        RECT 3483.895 3189.855 3518.220 3190.000 ;
        RECT 3519.275 3189.855 3558.090 3190.000 ;
        RECT 3566.900 3189.980 3568.975 3190.000 ;
        RECT 19.025 3138.000 21.100 3138.020 ;
        RECT 29.910 3138.000 68.725 3138.145 ;
        RECT 69.780 3138.000 104.105 3138.145 ;
        POLYGON 127.070 3138.115 127.070 3138.060 127.015 3138.060 ;
        RECT 127.070 3138.060 148.780 3138.115 ;
        RECT 105.420 3138.000 148.780 3138.060 ;
        RECT 164.275 3138.000 169.880 3138.115 ;
        RECT 174.985 3138.000 180.515 3138.115 ;
        RECT 0.000 3058.000 206.845 3138.000 ;
      LAYER met1 ;
        RECT 208.910 3124.840 209.230 3124.900 ;
        RECT 212.590 3124.840 212.910 3124.900 ;
        RECT 208.910 3124.700 212.910 3124.840 ;
        RECT 208.910 3124.640 209.230 3124.700 ;
        RECT 212.590 3124.640 212.910 3124.700 ;
        RECT 208.910 3092.540 209.230 3092.600 ;
        RECT 212.130 3092.540 212.450 3092.600 ;
        RECT 208.910 3092.400 212.450 3092.540 ;
        RECT 208.910 3092.340 209.230 3092.400 ;
        RECT 212.130 3092.340 212.450 3092.400 ;
        RECT 208.910 3077.580 209.230 3077.640 ;
        RECT 213.050 3077.580 213.370 3077.640 ;
        RECT 208.910 3077.440 213.370 3077.580 ;
        RECT 208.910 3077.380 209.230 3077.440 ;
        RECT 213.050 3077.380 213.370 3077.440 ;
      LAYER met1 ;
        RECT 29.910 3057.885 68.725 3058.000 ;
        RECT 69.780 3057.885 104.105 3058.000 ;
        RECT 108.520 3057.855 110.250 3058.000 ;
        RECT 119.365 3057.885 142.810 3058.000 ;
        RECT 3445.190 3045.000 3468.635 3045.115 ;
        RECT 3477.750 3045.000 3479.480 3045.145 ;
        RECT 3483.895 3045.000 3518.220 3045.115 ;
        RECT 3519.275 3045.000 3558.090 3045.115 ;
      LAYER met1 ;
        RECT 3368.190 3025.560 3368.510 3025.620 ;
        RECT 3376.930 3025.560 3377.250 3025.620 ;
        RECT 3368.190 3025.420 3377.250 3025.560 ;
        RECT 3368.190 3025.360 3368.510 3025.420 ;
        RECT 3376.930 3025.360 3377.250 3025.420 ;
        RECT 212.590 3015.840 212.910 3016.100 ;
        RECT 212.680 3015.080 212.820 3015.840 ;
        RECT 212.590 3014.820 212.910 3015.080 ;
        RECT 3367.270 3014.680 3367.590 3014.740 ;
        RECT 3376.930 3014.680 3377.250 3014.740 ;
        RECT 3367.270 3014.540 3377.250 3014.680 ;
        RECT 3367.270 3014.480 3367.590 3014.540 ;
        RECT 3376.930 3014.480 3377.250 3014.540 ;
        RECT 3367.730 2975.240 3368.050 2975.300 ;
        RECT 3376.930 2975.240 3377.250 2975.300 ;
        RECT 3367.730 2975.100 3377.250 2975.240 ;
        RECT 3367.730 2975.040 3368.050 2975.100 ;
        RECT 3376.930 2975.040 3377.250 2975.100 ;
      LAYER met1 ;
        RECT 3381.155 2965.000 3588.000 3045.000 ;
        RECT 3407.485 2964.885 3413.015 2965.000 ;
        RECT 3418.120 2964.885 3423.725 2965.000 ;
        RECT 3439.220 2964.940 3482.580 2965.000 ;
        RECT 3439.220 2964.885 3460.930 2964.940 ;
        POLYGON 3460.930 2964.940 3460.985 2964.940 3460.930 2964.885 ;
        RECT 3483.895 2964.855 3518.220 2965.000 ;
        RECT 3519.275 2964.855 3558.090 2965.000 ;
        RECT 3566.900 2964.980 3568.975 2965.000 ;
        RECT 19.025 2922.000 21.100 2922.020 ;
        RECT 29.910 2922.000 68.725 2922.145 ;
        RECT 69.780 2922.000 104.105 2922.145 ;
        POLYGON 127.070 2922.115 127.070 2922.060 127.015 2922.060 ;
        RECT 127.070 2922.060 148.780 2922.115 ;
        RECT 105.420 2922.000 148.780 2922.060 ;
        RECT 164.275 2922.000 169.880 2922.115 ;
        RECT 174.985 2922.000 180.515 2922.115 ;
        RECT 0.000 2842.000 206.845 2922.000 ;
      LAYER met1 ;
        RECT 208.910 2908.600 209.230 2908.660 ;
        RECT 212.130 2908.600 212.450 2908.660 ;
        RECT 208.910 2908.460 212.450 2908.600 ;
        RECT 208.910 2908.400 209.230 2908.460 ;
        RECT 212.130 2908.400 212.450 2908.460 ;
        RECT 208.910 2876.300 209.230 2876.360 ;
        RECT 213.510 2876.300 213.830 2876.360 ;
        RECT 208.910 2876.160 213.830 2876.300 ;
        RECT 208.910 2876.100 209.230 2876.160 ;
        RECT 213.510 2876.100 213.830 2876.160 ;
        RECT 208.910 2861.340 209.230 2861.400 ;
        RECT 212.590 2861.340 212.910 2861.400 ;
        RECT 213.970 2861.340 214.290 2861.400 ;
        RECT 208.910 2861.200 214.290 2861.340 ;
        RECT 208.910 2861.140 209.230 2861.200 ;
        RECT 212.590 2861.140 212.910 2861.200 ;
        RECT 213.970 2861.140 214.290 2861.200 ;
        RECT 211.210 2855.900 211.530 2855.960 ;
        RECT 212.130 2855.900 212.450 2855.960 ;
        RECT 211.210 2855.760 212.450 2855.900 ;
        RECT 211.210 2855.700 211.530 2855.760 ;
        RECT 212.130 2855.700 212.450 2855.760 ;
      LAYER met1 ;
        RECT 29.910 2841.885 68.725 2842.000 ;
        RECT 69.780 2841.885 104.105 2842.000 ;
        RECT 108.520 2841.855 110.250 2842.000 ;
        RECT 119.365 2841.885 142.810 2842.000 ;
        RECT 3445.190 2819.000 3468.635 2819.115 ;
        RECT 3477.750 2819.000 3479.480 2819.145 ;
        RECT 3483.895 2819.000 3518.220 2819.115 ;
        RECT 3519.275 2819.000 3558.090 2819.115 ;
      LAYER met1 ;
        RECT 3368.190 2804.900 3368.510 2804.960 ;
        RECT 3376.930 2804.900 3377.250 2804.960 ;
        RECT 3368.190 2804.760 3377.250 2804.900 ;
        RECT 3368.190 2804.700 3368.510 2804.760 ;
        RECT 3376.930 2804.700 3377.250 2804.760 ;
        RECT 3367.270 2789.260 3367.590 2789.320 ;
        RECT 3376.930 2789.260 3377.250 2789.320 ;
        RECT 3367.270 2789.120 3377.250 2789.260 ;
        RECT 3367.270 2789.060 3367.590 2789.120 ;
        RECT 3376.930 2789.060 3377.250 2789.120 ;
        RECT 3376.010 2778.040 3376.330 2778.100 ;
        RECT 3376.930 2778.040 3377.250 2778.100 ;
        RECT 3376.010 2777.900 3377.250 2778.040 ;
        RECT 3376.010 2777.840 3376.330 2777.900 ;
        RECT 3376.930 2777.840 3377.250 2777.900 ;
        RECT 3367.730 2752.540 3368.050 2752.600 ;
        RECT 3376.930 2752.540 3377.250 2752.600 ;
        RECT 3367.730 2752.400 3377.250 2752.540 ;
        RECT 3367.730 2752.340 3368.050 2752.400 ;
        RECT 3376.930 2752.340 3377.250 2752.400 ;
      LAYER met1 ;
        RECT 3381.155 2739.000 3588.000 2819.000 ;
        RECT 3407.485 2738.885 3413.015 2739.000 ;
        RECT 3418.120 2738.885 3423.725 2739.000 ;
        RECT 3439.220 2738.940 3482.580 2739.000 ;
        RECT 3439.220 2738.885 3460.930 2738.940 ;
        POLYGON 3460.930 2738.940 3460.985 2738.940 3460.930 2738.885 ;
        RECT 3483.895 2738.855 3518.220 2739.000 ;
        RECT 3519.275 2738.855 3558.090 2739.000 ;
        RECT 3566.900 2738.980 3568.975 2739.000 ;
      LAYER met1 ;
        RECT 211.210 2715.480 211.530 2715.540 ;
        RECT 212.130 2715.480 212.450 2715.540 ;
        RECT 211.210 2715.340 212.450 2715.480 ;
        RECT 211.210 2715.280 211.530 2715.340 ;
        RECT 212.130 2715.280 212.450 2715.340 ;
      LAYER met1 ;
        RECT 19.025 2706.000 21.100 2706.020 ;
        RECT 29.910 2706.000 68.725 2706.145 ;
        RECT 69.780 2706.000 104.105 2706.145 ;
        POLYGON 127.070 2706.115 127.070 2706.060 127.015 2706.060 ;
        RECT 127.070 2706.060 148.780 2706.115 ;
        RECT 105.420 2706.000 148.780 2706.060 ;
        RECT 164.275 2706.000 169.880 2706.115 ;
        RECT 174.985 2706.000 180.515 2706.115 ;
        RECT 0.000 2626.000 206.845 2706.000 ;
      LAYER met1 ;
        RECT 208.910 2697.460 209.230 2697.520 ;
        RECT 212.130 2697.460 212.450 2697.520 ;
        RECT 213.970 2697.460 214.290 2697.520 ;
        RECT 208.910 2697.320 214.290 2697.460 ;
        RECT 208.910 2697.260 209.230 2697.320 ;
        RECT 212.130 2697.260 212.450 2697.320 ;
        RECT 213.970 2697.260 214.290 2697.320 ;
        RECT 208.910 2655.980 209.230 2656.040 ;
        RECT 212.130 2655.980 212.450 2656.040 ;
        RECT 208.910 2655.840 212.450 2655.980 ;
        RECT 208.910 2655.780 209.230 2655.840 ;
        RECT 212.130 2655.780 212.450 2655.840 ;
        RECT 208.910 2640.340 209.230 2640.400 ;
        RECT 211.670 2640.340 211.990 2640.400 ;
        RECT 213.510 2640.340 213.830 2640.400 ;
        RECT 208.910 2640.200 213.830 2640.340 ;
        RECT 208.910 2640.140 209.230 2640.200 ;
        RECT 211.670 2640.140 211.990 2640.200 ;
        RECT 213.510 2640.140 213.830 2640.200 ;
      LAYER met1 ;
        RECT 29.910 2625.885 68.725 2626.000 ;
        RECT 69.780 2625.885 104.105 2626.000 ;
        RECT 108.520 2625.855 110.250 2626.000 ;
        RECT 119.365 2625.885 142.810 2626.000 ;
        RECT 3390.035 2590.375 3587.725 2593.815 ;
        RECT 3389.130 2585.145 3587.725 2590.375 ;
        RECT 3390.035 2581.965 3587.725 2585.145 ;
        RECT 3388.970 2580.650 3587.725 2581.965 ;
      LAYER met1 ;
        RECT 3376.470 2568.940 3376.790 2569.000 ;
        RECT 3388.430 2568.940 3388.750 2569.000 ;
        RECT 3376.470 2568.800 3388.750 2568.940 ;
        RECT 3376.470 2568.740 3376.790 2568.800 ;
        RECT 3388.430 2568.740 3388.750 2568.800 ;
      LAYER met1 ;
        RECT 3388.970 2524.460 3389.920 2580.650 ;
        POLYGON 3389.920 2580.650 3390.035 2580.650 3389.920 2580.535 ;
        POLYGON 3389.920 2524.575 3390.035 2524.460 3389.920 2524.460 ;
        RECT 3390.035 2524.460 3587.725 2580.650 ;
        RECT 3388.970 2523.320 3587.725 2524.460 ;
        RECT 3390.035 2521.085 3587.725 2523.320 ;
        RECT 0.275 2485.680 197.965 2487.915 ;
        RECT 0.275 2484.540 199.030 2485.680 ;
        RECT 0.275 2428.350 197.965 2484.540 ;
        POLYGON 197.965 2484.540 198.080 2484.540 198.080 2484.425 ;
        POLYGON 198.080 2428.465 198.080 2428.350 197.965 2428.350 ;
        RECT 198.080 2428.350 199.030 2484.540 ;
        RECT 0.275 2427.035 199.030 2428.350 ;
        RECT 0.275 2423.855 197.965 2427.035 ;
        RECT 0.275 2418.625 198.870 2423.855 ;
        RECT 0.275 2415.185 197.965 2418.625 ;
        RECT 3390.035 2357.345 3587.840 2373.880 ;
        RECT 3390.000 2353.075 3587.840 2357.345 ;
        RECT 3379.115 2317.435 3587.840 2353.075 ;
        RECT 3379.115 2297.800 3389.220 2317.435 ;
        RECT 3390.035 2299.000 3587.840 2317.435 ;
        RECT 3379.115 2292.065 3465.385 2297.800 ;
        POLYGON 3379.115 2292.065 3381.245 2292.065 3381.245 2289.935 ;
        RECT 3381.245 2289.935 3465.385 2292.065 ;
        RECT 122.615 2285.935 204.885 2289.935 ;
        POLYGON 204.885 2289.935 208.885 2285.935 204.885 2285.935 ;
        POLYGON 3381.245 2289.935 3383.115 2289.935 3383.115 2288.065 ;
        RECT 3383.115 2288.065 3465.385 2289.935 ;
        RECT 122.615 2280.200 208.885 2285.935 ;
        RECT 0.160 2260.565 197.965 2279.000 ;
        RECT 198.780 2260.565 208.885 2280.200 ;
        RECT 0.160 2224.925 208.885 2260.565 ;
        RECT 0.160 2220.655 198.000 2224.925 ;
        RECT 0.160 2204.120 197.965 2220.655 ;
        RECT 3390.035 2140.965 3587.725 2152.815 ;
        RECT 3388.970 2139.650 3587.725 2140.965 ;
      LAYER met1 ;
        RECT 3373.710 2139.180 3374.030 2139.240 ;
        RECT 3387.510 2139.180 3387.830 2139.240 ;
        RECT 3373.710 2139.040 3387.830 2139.180 ;
        RECT 3373.710 2138.980 3374.030 2139.040 ;
        RECT 3387.510 2138.980 3387.830 2139.040 ;
      LAYER met1 ;
        RECT 3388.970 2083.460 3389.920 2139.650 ;
        POLYGON 3389.920 2139.650 3390.035 2139.650 3389.920 2139.535 ;
        POLYGON 3389.920 2083.575 3390.035 2083.460 3389.920 2083.460 ;
        RECT 3390.035 2083.460 3587.725 2139.650 ;
        RECT 3388.970 2082.320 3587.725 2083.460 ;
        RECT 3390.035 2079.380 3587.725 2082.320 ;
        RECT 19.025 2068.000 21.100 2068.020 ;
        RECT 29.910 2068.000 68.725 2068.145 ;
        RECT 69.780 2068.000 104.105 2068.145 ;
        POLYGON 127.070 2068.115 127.070 2068.060 127.015 2068.060 ;
        RECT 127.070 2068.060 148.780 2068.115 ;
        RECT 105.420 2068.000 148.780 2068.060 ;
        RECT 164.275 2068.000 169.880 2068.115 ;
        RECT 174.985 2068.000 180.515 2068.115 ;
        RECT 0.000 1988.000 206.845 2068.000 ;
      LAYER met1 ;
        RECT 208.910 2054.860 209.230 2054.920 ;
        RECT 212.590 2054.860 212.910 2054.920 ;
        RECT 213.970 2054.860 214.290 2054.920 ;
        RECT 208.910 2054.720 214.290 2054.860 ;
        RECT 208.910 2054.660 209.230 2054.720 ;
        RECT 212.590 2054.660 212.910 2054.720 ;
        RECT 213.970 2054.660 214.290 2054.720 ;
        RECT 208.910 2022.560 209.230 2022.620 ;
        RECT 212.130 2022.560 212.450 2022.620 ;
        RECT 213.050 2022.560 213.370 2022.620 ;
        RECT 208.910 2022.420 213.370 2022.560 ;
        RECT 208.910 2022.360 209.230 2022.420 ;
        RECT 212.130 2022.360 212.450 2022.420 ;
        RECT 213.050 2022.360 213.370 2022.420 ;
        RECT 208.910 2004.200 209.230 2004.260 ;
        RECT 213.510 2004.200 213.830 2004.260 ;
        RECT 208.910 2004.060 213.830 2004.200 ;
        RECT 208.910 2004.000 209.230 2004.060 ;
        RECT 213.510 2004.000 213.830 2004.060 ;
      LAYER met1 ;
        RECT 29.910 1987.885 68.725 1988.000 ;
        RECT 69.780 1987.885 104.105 1988.000 ;
        RECT 108.520 1987.855 110.250 1988.000 ;
        RECT 119.365 1987.885 142.810 1988.000 ;
        RECT 3445.190 1933.000 3468.635 1933.115 ;
        RECT 3477.750 1933.000 3479.480 1933.145 ;
        RECT 3483.895 1933.000 3518.220 1933.115 ;
        RECT 3519.275 1933.000 3558.090 1933.115 ;
      LAYER met1 ;
        RECT 3367.730 1913.760 3368.050 1913.820 ;
        RECT 3376.930 1913.760 3377.250 1913.820 ;
        RECT 3367.730 1913.620 3377.250 1913.760 ;
        RECT 3367.730 1913.560 3368.050 1913.620 ;
        RECT 3376.930 1913.560 3377.250 1913.620 ;
        RECT 3368.650 1898.460 3368.970 1898.520 ;
        RECT 3376.930 1898.460 3377.250 1898.520 ;
        RECT 3368.650 1898.320 3377.250 1898.460 ;
        RECT 3368.650 1898.260 3368.970 1898.320 ;
        RECT 3376.930 1898.260 3377.250 1898.320 ;
        RECT 3367.270 1861.740 3367.590 1861.800 ;
        RECT 3369.570 1861.740 3369.890 1861.800 ;
        RECT 3376.930 1861.740 3377.250 1861.800 ;
        RECT 3367.270 1861.600 3377.250 1861.740 ;
        RECT 3367.270 1861.540 3367.590 1861.600 ;
        RECT 3369.570 1861.540 3369.890 1861.600 ;
        RECT 3376.930 1861.540 3377.250 1861.600 ;
      LAYER met1 ;
        RECT 3381.155 1853.000 3588.000 1933.000 ;
        RECT 3407.485 1852.885 3413.015 1853.000 ;
        RECT 3418.120 1852.885 3423.725 1853.000 ;
        RECT 3439.220 1852.940 3482.580 1853.000 ;
        RECT 3439.220 1852.885 3460.930 1852.940 ;
        POLYGON 3460.930 1852.940 3460.985 1852.940 3460.930 1852.885 ;
        RECT 3483.895 1852.855 3518.220 1853.000 ;
        RECT 3519.275 1852.855 3558.090 1853.000 ;
        RECT 3566.900 1852.980 3568.975 1853.000 ;
        RECT 19.025 1852.000 21.100 1852.020 ;
        RECT 29.910 1852.000 68.725 1852.145 ;
        RECT 69.780 1852.000 104.105 1852.145 ;
        POLYGON 127.070 1852.115 127.070 1852.060 127.015 1852.060 ;
        RECT 127.070 1852.060 148.780 1852.115 ;
        RECT 105.420 1852.000 148.780 1852.060 ;
        RECT 164.275 1852.000 169.880 1852.115 ;
        RECT 174.985 1852.000 180.515 1852.115 ;
        RECT 0.000 1772.000 206.845 1852.000 ;
      LAYER met1 ;
        RECT 208.910 1847.800 209.230 1847.860 ;
        RECT 211.670 1847.800 211.990 1847.860 ;
        RECT 208.910 1847.660 211.990 1847.800 ;
        RECT 208.910 1847.600 209.230 1847.660 ;
        RECT 211.670 1847.600 211.990 1847.660 ;
        RECT 208.910 1843.380 209.230 1843.440 ;
        RECT 212.590 1843.380 212.910 1843.440 ;
        RECT 208.910 1843.240 212.910 1843.380 ;
        RECT 208.910 1843.180 209.230 1843.240 ;
        RECT 212.590 1843.180 212.910 1843.240 ;
        RECT 208.910 1813.120 209.230 1813.180 ;
        RECT 211.670 1813.120 211.990 1813.180 ;
        RECT 208.910 1812.980 211.990 1813.120 ;
        RECT 208.910 1812.920 209.230 1812.980 ;
        RECT 211.670 1812.920 211.990 1812.980 ;
        RECT 208.910 1803.600 209.230 1803.660 ;
        RECT 213.050 1803.600 213.370 1803.660 ;
        RECT 208.910 1803.460 213.370 1803.600 ;
        RECT 208.910 1803.400 209.230 1803.460 ;
        RECT 213.050 1803.400 213.370 1803.460 ;
        RECT 208.910 1786.260 209.230 1786.320 ;
        RECT 212.590 1786.260 212.910 1786.320 ;
        RECT 213.510 1786.260 213.830 1786.320 ;
        RECT 208.910 1786.120 213.830 1786.260 ;
        RECT 208.910 1786.060 209.230 1786.120 ;
        RECT 212.590 1786.060 212.910 1786.120 ;
        RECT 213.510 1786.060 213.830 1786.120 ;
      LAYER met1 ;
        RECT 29.910 1771.885 68.725 1772.000 ;
        RECT 69.780 1771.885 104.105 1772.000 ;
        RECT 108.520 1771.855 110.250 1772.000 ;
        RECT 119.365 1771.885 142.810 1772.000 ;
        RECT 3445.190 1707.000 3468.635 1707.115 ;
        RECT 3477.750 1707.000 3479.480 1707.145 ;
        RECT 3483.895 1707.000 3518.220 1707.115 ;
        RECT 3519.275 1707.000 3558.090 1707.115 ;
      LAYER met1 ;
        RECT 3367.730 1687.660 3368.050 1687.720 ;
        RECT 3376.930 1687.660 3377.250 1687.720 ;
        RECT 3367.730 1687.520 3377.250 1687.660 ;
        RECT 3367.730 1687.460 3368.050 1687.520 ;
        RECT 3376.930 1687.460 3377.250 1687.520 ;
        RECT 3368.650 1672.360 3368.970 1672.420 ;
        RECT 3370.030 1672.360 3370.350 1672.420 ;
        RECT 3376.930 1672.360 3377.250 1672.420 ;
        RECT 3368.650 1672.220 3377.250 1672.360 ;
        RECT 3368.650 1672.160 3368.970 1672.220 ;
        RECT 3370.030 1672.160 3370.350 1672.220 ;
        RECT 3376.930 1672.160 3377.250 1672.220 ;
        RECT 3369.570 1640.400 3369.890 1640.460 ;
        RECT 3376.930 1640.400 3377.250 1640.460 ;
        RECT 3369.570 1640.260 3377.250 1640.400 ;
        RECT 3369.570 1640.200 3369.890 1640.260 ;
        RECT 3376.930 1640.200 3377.250 1640.260 ;
      LAYER met1 ;
        RECT 19.025 1636.000 21.100 1636.020 ;
        RECT 29.910 1636.000 68.725 1636.145 ;
        RECT 69.780 1636.000 104.105 1636.145 ;
        POLYGON 127.070 1636.115 127.070 1636.060 127.015 1636.060 ;
        RECT 127.070 1636.060 148.780 1636.115 ;
        RECT 105.420 1636.000 148.780 1636.060 ;
        RECT 164.275 1636.000 169.880 1636.115 ;
        RECT 174.985 1636.000 180.515 1636.115 ;
        RECT 0.000 1556.000 206.845 1636.000 ;
      LAYER met1 ;
        RECT 208.910 1627.480 209.230 1627.540 ;
        RECT 212.130 1627.480 212.450 1627.540 ;
        RECT 213.970 1627.480 214.290 1627.540 ;
        RECT 208.910 1627.340 214.290 1627.480 ;
        RECT 208.910 1627.280 209.230 1627.340 ;
        RECT 212.130 1627.280 212.450 1627.340 ;
        RECT 213.970 1627.280 214.290 1627.340 ;
      LAYER met1 ;
        RECT 3381.155 1627.000 3588.000 1707.000 ;
        RECT 3407.485 1626.885 3413.015 1627.000 ;
        RECT 3418.120 1626.885 3423.725 1627.000 ;
        RECT 3439.220 1626.940 3482.580 1627.000 ;
        RECT 3439.220 1626.885 3460.930 1626.940 ;
        POLYGON 3460.930 1626.940 3460.985 1626.940 3460.930 1626.885 ;
        RECT 3483.895 1626.855 3518.220 1627.000 ;
        RECT 3519.275 1626.855 3558.090 1627.000 ;
        RECT 3566.900 1626.980 3568.975 1627.000 ;
      LAYER met1 ;
        RECT 208.910 1586.000 209.230 1586.060 ;
        RECT 213.050 1586.000 213.370 1586.060 ;
        RECT 208.910 1585.860 213.370 1586.000 ;
        RECT 208.910 1585.800 209.230 1585.860 ;
        RECT 213.050 1585.800 213.370 1585.860 ;
        RECT 208.910 1570.360 209.230 1570.420 ;
        RECT 212.590 1570.360 212.910 1570.420 ;
        RECT 213.510 1570.360 213.830 1570.420 ;
        RECT 208.910 1570.220 213.830 1570.360 ;
        RECT 208.910 1570.160 209.230 1570.220 ;
        RECT 212.590 1570.160 212.910 1570.220 ;
        RECT 213.510 1570.160 213.830 1570.220 ;
      LAYER met1 ;
        RECT 29.910 1555.885 68.725 1556.000 ;
        RECT 69.780 1555.885 104.105 1556.000 ;
        RECT 108.520 1555.855 110.250 1556.000 ;
        RECT 119.365 1555.885 142.810 1556.000 ;
        RECT 3445.190 1482.000 3468.635 1482.115 ;
        RECT 3477.750 1482.000 3479.480 1482.145 ;
        RECT 3483.895 1482.000 3518.220 1482.115 ;
        RECT 3519.275 1482.000 3558.090 1482.115 ;
      LAYER met1 ;
        RECT 3367.270 1465.980 3367.590 1466.040 ;
        RECT 3376.930 1465.980 3377.250 1466.040 ;
        RECT 3367.270 1465.840 3377.250 1465.980 ;
        RECT 3367.270 1465.780 3367.590 1465.840 ;
        RECT 3376.930 1465.780 3377.250 1465.840 ;
        RECT 3367.730 1447.620 3368.050 1447.680 ;
        RECT 3370.030 1447.620 3370.350 1447.680 ;
        RECT 3376.930 1447.620 3377.250 1447.680 ;
        RECT 3367.730 1447.480 3377.250 1447.620 ;
        RECT 3367.730 1447.420 3368.050 1447.480 ;
        RECT 3370.030 1447.420 3370.350 1447.480 ;
        RECT 3376.930 1447.420 3377.250 1447.480 ;
      LAYER met1 ;
        RECT 19.025 1420.000 21.100 1420.020 ;
        RECT 29.910 1420.000 68.725 1420.145 ;
        RECT 69.780 1420.000 104.105 1420.145 ;
        POLYGON 127.070 1420.115 127.070 1420.060 127.015 1420.060 ;
        RECT 127.070 1420.060 148.780 1420.115 ;
        RECT 105.420 1420.000 148.780 1420.060 ;
        RECT 164.275 1420.000 169.880 1420.115 ;
        RECT 174.985 1420.000 180.515 1420.115 ;
        RECT 0.000 1340.000 206.845 1420.000 ;
      LAYER met1 ;
        RECT 3369.570 1415.320 3369.890 1415.380 ;
        RECT 3376.930 1415.320 3377.250 1415.380 ;
        RECT 3369.570 1415.180 3377.250 1415.320 ;
        RECT 3369.570 1415.120 3369.890 1415.180 ;
        RECT 3376.930 1415.120 3377.250 1415.180 ;
        RECT 208.910 1406.820 209.230 1406.880 ;
        RECT 212.130 1406.820 212.450 1406.880 ;
        RECT 213.970 1406.820 214.290 1406.880 ;
        RECT 208.910 1406.680 214.290 1406.820 ;
        RECT 208.910 1406.620 209.230 1406.680 ;
        RECT 212.130 1406.620 212.450 1406.680 ;
        RECT 213.970 1406.620 214.290 1406.680 ;
      LAYER met1 ;
        RECT 3381.155 1402.000 3588.000 1482.000 ;
        RECT 3407.485 1401.885 3413.015 1402.000 ;
        RECT 3418.120 1401.885 3423.725 1402.000 ;
        RECT 3439.220 1401.940 3482.580 1402.000 ;
        RECT 3439.220 1401.885 3460.930 1401.940 ;
        POLYGON 3460.930 1401.940 3460.985 1401.940 3460.930 1401.885 ;
        RECT 3483.895 1401.855 3518.220 1402.000 ;
        RECT 3519.275 1401.855 3558.090 1402.000 ;
        RECT 3566.900 1401.980 3568.975 1402.000 ;
      LAYER met1 ;
        RECT 208.910 1372.820 209.230 1372.880 ;
        RECT 213.050 1372.820 213.370 1372.880 ;
        RECT 208.910 1372.680 213.370 1372.820 ;
        RECT 208.910 1372.620 209.230 1372.680 ;
        RECT 213.050 1372.620 213.370 1372.680 ;
        RECT 208.910 1359.560 209.230 1359.620 ;
        RECT 213.510 1359.560 213.830 1359.620 ;
        RECT 208.910 1359.420 213.830 1359.560 ;
        RECT 208.910 1359.360 209.230 1359.420 ;
        RECT 213.510 1359.360 213.830 1359.420 ;
      LAYER met1 ;
        RECT 29.910 1339.885 68.725 1340.000 ;
        RECT 69.780 1339.885 104.105 1340.000 ;
        RECT 108.520 1339.855 110.250 1340.000 ;
        RECT 119.365 1339.885 142.810 1340.000 ;
        RECT 3445.190 1257.000 3468.635 1257.115 ;
        RECT 3477.750 1257.000 3479.480 1257.145 ;
        RECT 3483.895 1257.000 3518.220 1257.115 ;
        RECT 3519.275 1257.000 3558.090 1257.115 ;
      LAYER met1 ;
        RECT 3367.270 1242.940 3367.590 1243.000 ;
        RECT 3370.030 1242.940 3370.350 1243.000 ;
        RECT 3376.930 1242.940 3377.250 1243.000 ;
        RECT 3367.270 1242.800 3377.250 1242.940 ;
        RECT 3367.270 1242.740 3367.590 1242.800 ;
        RECT 3370.030 1242.740 3370.350 1242.800 ;
        RECT 3376.930 1242.740 3377.250 1242.800 ;
        RECT 3367.730 1224.580 3368.050 1224.640 ;
        RECT 3376.930 1224.580 3377.250 1224.640 ;
        RECT 3367.730 1224.440 3377.250 1224.580 ;
        RECT 3367.730 1224.380 3368.050 1224.440 ;
        RECT 3376.930 1224.380 3377.250 1224.440 ;
      LAYER met1 ;
        RECT 19.025 1204.000 21.100 1204.020 ;
        RECT 29.910 1204.000 68.725 1204.145 ;
        RECT 69.780 1204.000 104.105 1204.145 ;
        POLYGON 127.070 1204.115 127.070 1204.060 127.015 1204.060 ;
        RECT 127.070 1204.060 148.780 1204.115 ;
        RECT 105.420 1204.000 148.780 1204.060 ;
        RECT 164.275 1204.000 169.880 1204.115 ;
        RECT 174.985 1204.000 180.515 1204.115 ;
        RECT 0.000 1124.000 206.845 1204.000 ;
      LAYER met1 ;
        RECT 208.910 1190.580 209.230 1190.640 ;
        RECT 212.130 1190.580 212.450 1190.640 ;
        RECT 208.910 1190.440 212.450 1190.580 ;
        RECT 208.910 1190.380 209.230 1190.440 ;
        RECT 212.130 1190.380 212.450 1190.440 ;
        RECT 3369.570 1188.540 3369.890 1188.600 ;
        RECT 3376.930 1188.540 3377.250 1188.600 ;
        RECT 3369.570 1188.400 3377.250 1188.540 ;
        RECT 3369.570 1188.340 3369.890 1188.400 ;
        RECT 3376.930 1188.340 3377.250 1188.400 ;
      LAYER met1 ;
        RECT 3381.155 1177.000 3588.000 1257.000 ;
        RECT 3407.485 1176.885 3413.015 1177.000 ;
        RECT 3418.120 1176.885 3423.725 1177.000 ;
        RECT 3439.220 1176.940 3482.580 1177.000 ;
        RECT 3439.220 1176.885 3460.930 1176.940 ;
        POLYGON 3460.930 1176.940 3460.985 1176.940 3460.930 1176.885 ;
        RECT 3483.895 1176.855 3518.220 1177.000 ;
        RECT 3519.275 1176.855 3558.090 1177.000 ;
        RECT 3566.900 1176.980 3568.975 1177.000 ;
      LAYER met1 ;
        RECT 208.910 1158.620 209.230 1158.680 ;
        RECT 212.590 1158.620 212.910 1158.680 ;
        RECT 208.910 1158.480 212.910 1158.620 ;
        RECT 208.910 1158.420 209.230 1158.480 ;
        RECT 212.590 1158.420 212.910 1158.480 ;
        RECT 208.910 1143.320 209.230 1143.380 ;
        RECT 213.050 1143.320 213.370 1143.380 ;
        RECT 208.910 1143.180 213.370 1143.320 ;
        RECT 208.910 1143.120 209.230 1143.180 ;
        RECT 213.050 1143.120 213.370 1143.180 ;
        RECT 211.210 1137.540 211.530 1137.600 ;
        RECT 212.590 1137.540 212.910 1137.600 ;
        RECT 211.210 1137.400 212.910 1137.540 ;
        RECT 211.210 1137.340 211.530 1137.400 ;
        RECT 212.590 1137.340 212.910 1137.400 ;
      LAYER met1 ;
        RECT 29.910 1123.885 68.725 1124.000 ;
        RECT 69.780 1123.885 104.105 1124.000 ;
        RECT 108.520 1123.855 110.250 1124.000 ;
        RECT 119.365 1123.885 142.810 1124.000 ;
        RECT 3445.190 1031.000 3468.635 1031.115 ;
        RECT 3477.750 1031.000 3479.480 1031.145 ;
        RECT 3483.895 1031.000 3518.220 1031.115 ;
        RECT 3519.275 1031.000 3558.090 1031.115 ;
      LAYER met1 ;
        RECT 3370.030 1011.740 3370.350 1011.800 ;
        RECT 3376.930 1011.740 3377.250 1011.800 ;
        RECT 3370.030 1011.600 3377.250 1011.740 ;
        RECT 3370.030 1011.540 3370.350 1011.600 ;
        RECT 3376.930 1011.540 3377.250 1011.600 ;
        RECT 3367.730 996.440 3368.050 996.500 ;
        RECT 3376.930 996.440 3377.250 996.500 ;
        RECT 3367.730 996.300 3377.250 996.440 ;
        RECT 3367.730 996.240 3368.050 996.300 ;
        RECT 3376.930 996.240 3377.250 996.300 ;
      LAYER met1 ;
        RECT 19.025 988.000 21.100 988.020 ;
        RECT 29.910 988.000 68.725 988.145 ;
        RECT 69.780 988.000 104.105 988.145 ;
        POLYGON 127.070 988.115 127.070 988.060 127.015 988.060 ;
        RECT 127.070 988.060 148.780 988.115 ;
        RECT 105.420 988.000 148.780 988.060 ;
        RECT 164.275 988.000 169.880 988.115 ;
        RECT 174.985 988.000 180.515 988.115 ;
        RECT 0.000 908.000 206.845 988.000 ;
      LAYER met1 ;
        RECT 208.910 979.440 209.230 979.500 ;
        RECT 212.590 979.440 212.910 979.500 ;
        RECT 208.910 979.300 212.910 979.440 ;
        RECT 208.910 979.240 209.230 979.300 ;
        RECT 212.590 979.240 212.910 979.300 ;
        RECT 3369.570 959.720 3369.890 959.780 ;
        RECT 3376.930 959.720 3377.250 959.780 ;
        RECT 3369.570 959.580 3377.250 959.720 ;
        RECT 3369.570 959.520 3369.890 959.580 ;
        RECT 3376.930 959.520 3377.250 959.580 ;
      LAYER met1 ;
        RECT 3381.155 951.000 3588.000 1031.000 ;
        RECT 3407.485 950.885 3413.015 951.000 ;
        RECT 3418.120 950.885 3423.725 951.000 ;
        RECT 3439.220 950.940 3482.580 951.000 ;
        RECT 3439.220 950.885 3460.930 950.940 ;
        POLYGON 3460.930 950.940 3460.985 950.940 3460.930 950.885 ;
        RECT 3483.895 950.855 3518.220 951.000 ;
        RECT 3519.275 950.855 3558.090 951.000 ;
        RECT 3566.900 950.980 3568.975 951.000 ;
      LAYER met1 ;
        RECT 209.830 937.960 210.150 938.020 ;
        RECT 212.590 937.960 212.910 938.020 ;
        RECT 209.830 937.820 212.910 937.960 ;
        RECT 209.830 937.760 210.150 937.820 ;
        RECT 212.590 937.760 212.910 937.820 ;
        RECT 208.910 922.320 209.230 922.380 ;
        RECT 213.050 922.320 213.370 922.380 ;
        RECT 208.910 922.180 213.370 922.320 ;
        RECT 208.910 922.120 209.230 922.180 ;
        RECT 211.300 921.020 211.440 922.180 ;
        RECT 213.050 922.120 213.370 922.180 ;
        RECT 211.210 920.760 211.530 921.020 ;
      LAYER met1 ;
        RECT 29.910 907.885 68.725 908.000 ;
        RECT 69.780 907.885 104.105 908.000 ;
        RECT 108.520 907.855 110.250 908.000 ;
        RECT 119.365 907.885 142.810 908.000 ;
        RECT 3445.190 806.000 3468.635 806.115 ;
        RECT 3477.750 806.000 3479.480 806.145 ;
        RECT 3483.895 806.000 3518.220 806.115 ;
        RECT 3519.275 806.000 3558.090 806.115 ;
      LAYER met1 ;
        RECT 3367.270 791.760 3367.590 791.820 ;
        RECT 3370.030 791.760 3370.350 791.820 ;
        RECT 3376.930 791.760 3377.250 791.820 ;
        RECT 3367.270 791.620 3377.250 791.760 ;
        RECT 3367.270 791.560 3367.590 791.620 ;
        RECT 3370.030 791.560 3370.350 791.620 ;
        RECT 3376.930 791.560 3377.250 791.620 ;
        RECT 3367.730 776.120 3368.050 776.180 ;
        RECT 3376.930 776.120 3377.250 776.180 ;
        RECT 3367.730 775.980 3377.250 776.120 ;
        RECT 3367.730 775.920 3368.050 775.980 ;
        RECT 3376.930 775.920 3377.250 775.980 ;
        RECT 3368.650 734.640 3368.970 734.700 ;
        RECT 3369.570 734.640 3369.890 734.700 ;
        RECT 3376.930 734.640 3377.250 734.700 ;
        RECT 3368.650 734.500 3377.250 734.640 ;
        RECT 3368.650 734.440 3368.970 734.500 ;
        RECT 3369.570 734.440 3369.890 734.500 ;
        RECT 3376.930 734.440 3377.250 734.500 ;
      LAYER met1 ;
        RECT 3381.155 726.000 3588.000 806.000 ;
        RECT 3407.485 725.885 3413.015 726.000 ;
        RECT 3418.120 725.885 3423.725 726.000 ;
        RECT 3439.220 725.940 3482.580 726.000 ;
        RECT 3439.220 725.885 3460.930 725.940 ;
        POLYGON 3460.930 725.940 3460.985 725.940 3460.930 725.885 ;
        RECT 3483.895 725.855 3518.220 726.000 ;
        RECT 3519.275 725.855 3558.090 726.000 ;
        RECT 3566.900 725.980 3568.975 726.000 ;
        RECT 0.275 621.680 197.965 623.915 ;
        RECT 0.275 620.540 199.030 621.680 ;
        RECT 0.275 564.350 197.965 620.540 ;
        POLYGON 197.965 620.540 198.080 620.540 198.080 620.425 ;
        POLYGON 198.080 564.465 198.080 564.350 197.965 564.350 ;
        RECT 198.080 564.350 199.030 620.540 ;
      LAYER met1 ;
        RECT 212.590 607.480 212.910 607.540 ;
        RECT 220.870 607.480 221.190 607.540 ;
        RECT 212.590 607.340 221.190 607.480 ;
        RECT 212.590 607.280 212.910 607.340 ;
        RECT 220.870 607.280 221.190 607.340 ;
      LAYER met1 ;
        RECT 3445.190 580.000 3468.635 580.115 ;
        RECT 3477.750 580.000 3479.480 580.145 ;
        RECT 3483.895 580.000 3518.220 580.115 ;
        RECT 3519.275 580.000 3558.090 580.115 ;
      LAYER met1 ;
        RECT 3367.270 566.000 3367.590 566.060 ;
        RECT 3376.930 566.000 3377.250 566.060 ;
        RECT 3367.270 565.860 3377.250 566.000 ;
        RECT 3367.270 565.800 3367.590 565.860 ;
        RECT 3376.930 565.800 3377.250 565.860 ;
      LAYER met1 ;
        RECT 0.275 563.035 199.030 564.350 ;
        RECT 0.275 559.855 197.965 563.035 ;
        RECT 0.275 554.625 198.870 559.855 ;
        RECT 0.275 551.185 197.965 554.625 ;
      LAYER met1 ;
        RECT 3367.730 547.640 3368.050 547.700 ;
        RECT 3376.930 547.640 3377.250 547.700 ;
        RECT 3367.730 547.500 3377.250 547.640 ;
        RECT 3367.730 547.440 3368.050 547.500 ;
        RECT 3376.930 547.440 3377.250 547.500 ;
        RECT 3368.650 508.540 3368.970 508.600 ;
        RECT 3376.930 508.540 3377.250 508.600 ;
        RECT 3368.650 508.400 3377.250 508.540 ;
        RECT 3368.650 508.340 3368.970 508.400 ;
        RECT 3376.930 508.340 3377.250 508.400 ;
      LAYER met1 ;
        RECT 3381.155 500.000 3588.000 580.000 ;
        RECT 3407.485 499.885 3413.015 500.000 ;
        RECT 3418.120 499.885 3423.725 500.000 ;
        RECT 3439.220 499.940 3482.580 500.000 ;
        RECT 3439.220 499.885 3460.930 499.940 ;
        POLYGON 3460.930 499.940 3460.985 499.940 3460.930 499.885 ;
        RECT 3483.895 499.855 3518.220 500.000 ;
        RECT 3519.275 499.855 3558.090 500.000 ;
        RECT 3566.900 499.980 3568.975 500.000 ;
        RECT 159.640 425.935 163.510 426.195 ;
        RECT 159.640 421.935 204.500 425.935 ;
        POLYGON 204.500 425.935 208.500 421.935 204.500 421.935 ;
        RECT 159.640 416.200 208.500 421.935 ;
        RECT 159.640 415.245 163.510 416.200 ;
        RECT 0.160 396.565 197.965 415.000 ;
        RECT 198.780 396.565 208.500 416.200 ;
      LAYER met1 ;
        RECT 212.130 414.360 212.450 414.420 ;
        RECT 220.870 414.360 221.190 414.420 ;
        RECT 212.130 414.220 221.190 414.360 ;
        RECT 212.130 414.160 212.450 414.220 ;
        RECT 220.870 414.160 221.190 414.220 ;
      LAYER met1 ;
        RECT 0.160 360.495 208.500 396.565 ;
        RECT 0.160 356.655 198.000 360.495 ;
        RECT 198.980 358.655 208.500 360.495 ;
        POLYGON 198.980 358.655 200.980 358.655 200.980 356.655 ;
        RECT 200.980 356.655 206.500 358.655 ;
        POLYGON 206.500 358.655 208.500 358.655 206.500 356.655 ;
        RECT 0.160 340.120 197.965 356.655 ;
      LAYER met1 ;
        RECT 224.090 234.840 224.410 234.900 ;
        RECT 224.090 234.700 938.470 234.840 ;
        RECT 224.090 234.640 224.410 234.700 ;
        RECT 745.360 234.560 745.500 234.700 ;
        RECT 745.270 234.300 745.590 234.560 ;
        RECT 938.330 234.500 938.470 234.700 ;
        RECT 1004.340 234.700 1488.860 234.840 ;
        RECT 1004.340 234.560 1004.480 234.700 ;
        RECT 942.610 234.500 942.930 234.560 ;
        RECT 938.330 234.360 942.930 234.500 ;
        RECT 942.610 234.300 942.930 234.360 ;
        RECT 1004.250 234.300 1004.570 234.560 ;
        RECT 1204.440 234.500 1204.580 234.700 ;
        RECT 1488.720 234.560 1488.860 234.700 ;
        RECT 1547.140 234.700 1763.020 234.840 ;
        RECT 1547.140 234.560 1547.280 234.700 ;
        RECT 1762.880 234.560 1763.020 234.700 ;
        RECT 1821.300 234.700 2037.180 234.840 ;
        RECT 1821.300 234.560 1821.440 234.700 ;
        RECT 2037.040 234.560 2037.180 234.700 ;
        RECT 2095.460 234.700 2310.880 234.840 ;
        RECT 2095.460 234.560 2095.600 234.700 ;
        RECT 2310.740 234.560 2310.880 234.700 ;
        RECT 2369.160 234.700 2585.040 234.840 ;
        RECT 2369.160 234.560 2369.300 234.700 ;
        RECT 2584.900 234.560 2585.040 234.700 ;
        RECT 1281.170 234.500 1281.490 234.560 ;
        RECT 1204.440 234.360 1281.490 234.500 ;
        RECT 1281.170 234.300 1281.490 234.360 ;
        RECT 1488.630 234.300 1488.950 234.560 ;
        RECT 1547.050 234.300 1547.370 234.560 ;
        RECT 1762.790 234.300 1763.110 234.560 ;
        RECT 1821.210 234.300 1821.530 234.560 ;
        RECT 2036.950 234.300 2037.270 234.560 ;
        RECT 2095.370 234.300 2095.690 234.560 ;
        RECT 2310.650 234.300 2310.970 234.560 ;
        RECT 2369.070 234.300 2369.390 234.560 ;
        RECT 2584.810 234.300 2585.130 234.560 ;
        RECT 211.210 228.040 211.530 228.100 ;
        RECT 704.790 228.040 705.110 228.100 ;
        RECT 211.210 227.900 705.110 228.040 ;
        RECT 211.210 227.840 211.530 227.900 ;
        RECT 704.790 227.840 705.110 227.900 ;
        RECT 2618.850 228.040 2619.170 228.100 ;
        RECT 3367.730 228.040 3368.050 228.100 ;
        RECT 2618.850 227.900 3368.050 228.040 ;
        RECT 2618.850 227.840 2619.170 227.900 ;
        RECT 3367.730 227.840 3368.050 227.900 ;
        RECT 224.550 227.700 224.870 227.760 ;
        RECT 979.870 227.700 980.190 227.760 ;
        RECT 224.550 227.560 980.190 227.700 ;
        RECT 224.550 227.500 224.870 227.560 ;
        RECT 979.870 227.500 980.190 227.560 ;
        RECT 2593.550 227.700 2593.870 227.760 ;
        RECT 3368.650 227.700 3368.970 227.760 ;
        RECT 2593.550 227.560 3368.970 227.700 ;
        RECT 2593.550 227.500 2593.870 227.560 ;
        RECT 3368.650 227.500 3368.970 227.560 ;
        RECT 979.870 222.260 980.190 222.320 ;
        RECT 1522.670 222.260 1522.990 222.320 ;
        RECT 1531.410 222.260 1531.730 222.320 ;
        RECT 979.870 222.120 1531.730 222.260 ;
        RECT 979.870 222.060 980.190 222.120 ;
        RECT 1522.670 222.060 1522.990 222.120 ;
        RECT 1531.410 222.060 1531.730 222.120 ;
        RECT 2033.730 222.260 2034.050 222.320 ;
        RECT 2307.430 222.260 2307.750 222.320 ;
        RECT 2033.730 222.120 2307.750 222.260 ;
        RECT 2033.730 222.060 2034.050 222.120 ;
        RECT 2307.430 222.060 2307.750 222.120 ;
        RECT 2344.690 222.260 2345.010 222.320 ;
        RECT 2618.850 222.260 2619.170 222.320 ;
        RECT 2344.690 222.120 2619.170 222.260 ;
        RECT 2344.690 222.060 2345.010 222.120 ;
        RECT 2618.850 222.060 2619.170 222.120 ;
        RECT 1759.570 221.920 1759.890 221.980 ;
        RECT 1771.990 221.920 1772.310 221.980 ;
        RECT 1802.810 221.920 1803.130 221.980 ;
        RECT 1614.530 221.780 1904.470 221.920 ;
        RECT 942.610 221.580 942.930 221.640 ;
        RECT 964.230 221.580 964.550 221.640 ;
        RECT 1007.470 221.580 1007.790 221.640 ;
        RECT 1485.410 221.580 1485.730 221.640 ;
        RECT 1497.830 221.580 1498.150 221.640 ;
        RECT 1528.650 221.580 1528.970 221.640 ;
        RECT 1614.530 221.580 1614.670 221.780 ;
        RECT 1759.570 221.720 1759.890 221.780 ;
        RECT 1771.990 221.720 1772.310 221.780 ;
        RECT 1802.810 221.720 1803.130 221.780 ;
        RECT 942.610 221.440 1614.670 221.580 ;
        RECT 1904.330 221.580 1904.470 221.780 ;
        RECT 2033.730 221.580 2034.050 221.640 ;
        RECT 2344.690 221.580 2345.010 221.640 ;
        RECT 1904.330 221.440 2034.050 221.580 ;
        RECT 942.610 221.380 942.930 221.440 ;
        RECT 964.230 221.380 964.550 221.440 ;
        RECT 1007.470 221.380 1007.790 221.440 ;
        RECT 1485.410 221.380 1485.730 221.440 ;
        RECT 1497.830 221.380 1498.150 221.440 ;
        RECT 1528.650 221.380 1528.970 221.440 ;
        RECT 2033.730 221.380 2034.050 221.440 ;
        RECT 2097.530 221.440 2345.010 221.580 ;
        RECT 933.410 221.240 933.730 221.300 ;
        RECT 973.430 221.240 973.750 221.300 ;
        RECT 1796.830 221.240 1797.150 221.300 ;
        RECT 933.410 221.100 973.750 221.240 ;
        RECT 933.410 221.040 933.730 221.100 ;
        RECT 973.430 221.040 973.750 221.100 ;
        RECT 1750.000 221.100 1807.870 221.240 ;
        RECT 1476.210 220.900 1476.530 220.960 ;
        RECT 1516.230 220.900 1516.550 220.960 ;
        RECT 1476.210 220.760 1516.550 220.900 ;
        RECT 1476.210 220.700 1476.530 220.760 ;
        RECT 1516.230 220.700 1516.550 220.760 ;
        RECT 1531.410 220.900 1531.730 220.960 ;
        RECT 1750.000 220.900 1750.140 221.100 ;
        RECT 1796.830 221.040 1797.150 221.100 ;
        RECT 1531.410 220.760 1750.140 220.900 ;
        RECT 1750.370 220.900 1750.690 220.960 ;
        RECT 1790.390 220.900 1790.710 220.960 ;
        RECT 1750.370 220.760 1790.710 220.900 ;
        RECT 1807.730 220.900 1807.870 221.100 ;
        RECT 2070.990 220.900 2071.310 220.960 ;
        RECT 2097.530 220.900 2097.670 221.440 ;
        RECT 2344.690 221.380 2345.010 221.440 ;
        RECT 2307.430 221.240 2307.750 221.300 ;
        RECT 2581.590 221.240 2581.910 221.300 ;
        RECT 2593.550 221.240 2593.870 221.300 ;
        RECT 2307.430 221.100 2593.870 221.240 ;
        RECT 2307.430 221.040 2307.750 221.100 ;
        RECT 2581.590 221.040 2581.910 221.100 ;
        RECT 2593.550 221.040 2593.870 221.100 ;
        RECT 1807.730 220.760 2097.670 220.900 ;
        RECT 1531.410 220.700 1531.730 220.760 ;
        RECT 1750.370 220.700 1750.690 220.760 ;
        RECT 1790.390 220.700 1790.710 220.760 ;
        RECT 2070.990 220.700 2071.310 220.760 ;
        RECT 2899.450 213.760 2899.770 213.820 ;
        RECT 3367.270 213.760 3367.590 213.820 ;
        RECT 2899.450 213.620 3367.590 213.760 ;
        RECT 2899.450 213.560 2899.770 213.620 ;
        RECT 3367.270 213.560 3367.590 213.620 ;
        RECT 946.290 209.680 946.610 209.740 ;
        RECT 955.490 209.680 955.810 209.740 ;
        RECT 961.470 209.680 961.790 209.740 ;
        RECT 967.910 209.680 968.230 209.740 ;
        RECT 982.170 209.680 982.490 209.740 ;
        RECT 946.290 209.540 982.490 209.680 ;
        RECT 946.290 209.480 946.610 209.540 ;
        RECT 955.490 209.480 955.810 209.540 ;
        RECT 961.470 209.480 961.790 209.540 ;
        RECT 967.910 209.480 968.230 209.540 ;
        RECT 982.170 209.480 982.490 209.540 ;
        RECT 992.290 209.680 992.610 209.740 ;
        RECT 1000.570 209.680 1000.890 209.740 ;
        RECT 992.290 209.540 1000.890 209.680 ;
        RECT 992.290 209.480 992.610 209.540 ;
        RECT 1000.570 209.480 1000.890 209.540 ;
        RECT 1489.550 209.680 1489.870 209.740 ;
        RECT 1503.350 209.680 1503.670 209.740 ;
        RECT 1489.550 209.540 1503.670 209.680 ;
        RECT 1489.550 209.480 1489.870 209.540 ;
        RECT 1503.350 209.480 1503.670 209.540 ;
        RECT 1511.170 209.680 1511.490 209.740 ;
        RECT 1526.350 209.680 1526.670 209.740 ;
        RECT 1532.790 209.680 1533.110 209.740 ;
        RECT 1543.370 209.680 1543.690 209.740 ;
        RECT 1511.170 209.540 1543.690 209.680 ;
        RECT 1511.170 209.480 1511.490 209.540 ;
        RECT 1526.350 209.480 1526.670 209.540 ;
        RECT 1532.790 209.480 1533.110 209.540 ;
        RECT 1543.370 209.480 1543.690 209.540 ;
        RECT 1763.250 209.680 1763.570 209.740 ;
        RECT 1777.510 209.680 1777.830 209.740 ;
        RECT 1763.250 209.540 1777.830 209.680 ;
        RECT 1763.250 209.480 1763.570 209.540 ;
        RECT 1777.510 209.480 1777.830 209.540 ;
        RECT 1784.870 209.680 1785.190 209.740 ;
        RECT 1799.130 209.680 1799.450 209.740 ;
        RECT 1805.570 209.680 1805.890 209.740 ;
        RECT 1817.530 209.680 1817.850 209.740 ;
        RECT 1784.870 209.540 1817.850 209.680 ;
        RECT 1784.870 209.480 1785.190 209.540 ;
        RECT 1799.130 209.480 1799.450 209.540 ;
        RECT 1805.570 209.480 1805.890 209.540 ;
        RECT 1817.530 209.480 1817.850 209.540 ;
        RECT 2037.410 209.680 2037.730 209.740 ;
        RECT 2051.210 209.680 2051.530 209.740 ;
        RECT 2057.650 209.680 2057.970 209.740 ;
        RECT 2072.830 209.680 2073.150 209.740 ;
        RECT 2079.270 209.680 2079.590 209.740 ;
        RECT 2091.230 209.680 2091.550 209.740 ;
        RECT 2037.410 209.540 2091.550 209.680 ;
        RECT 2037.410 209.480 2037.730 209.540 ;
        RECT 2051.210 209.480 2051.530 209.540 ;
        RECT 2057.650 209.480 2057.970 209.540 ;
        RECT 2072.830 209.480 2073.150 209.540 ;
        RECT 2079.270 209.480 2079.590 209.540 ;
        RECT 2091.230 209.480 2091.550 209.540 ;
        RECT 2311.570 209.680 2311.890 209.740 ;
        RECT 2325.370 209.680 2325.690 209.740 ;
        RECT 2331.810 209.680 2332.130 209.740 ;
        RECT 2346.990 209.680 2347.310 209.740 ;
        RECT 2353.430 209.680 2353.750 209.740 ;
        RECT 2365.390 209.680 2365.710 209.740 ;
        RECT 2311.570 209.540 2365.710 209.680 ;
        RECT 2311.570 209.480 2311.890 209.540 ;
        RECT 2325.370 209.480 2325.690 209.540 ;
        RECT 2331.810 209.480 2332.130 209.540 ;
        RECT 2346.990 209.480 2347.310 209.540 ;
        RECT 2353.430 209.480 2353.750 209.540 ;
        RECT 2365.390 209.480 2365.710 209.540 ;
        RECT 2585.270 209.680 2585.590 209.740 ;
        RECT 2599.530 209.680 2599.850 209.740 ;
        RECT 2605.970 209.680 2606.290 209.740 ;
        RECT 2621.150 209.680 2621.470 209.740 ;
        RECT 2627.590 209.680 2627.910 209.740 ;
        RECT 2639.550 209.680 2639.870 209.740 ;
        RECT 2585.270 209.540 2639.870 209.680 ;
        RECT 2585.270 209.480 2585.590 209.540 ;
        RECT 2599.530 209.480 2599.850 209.540 ;
        RECT 2605.970 209.480 2606.290 209.540 ;
        RECT 2621.150 209.480 2621.470 209.540 ;
        RECT 2627.590 209.480 2627.910 209.540 ;
        RECT 2639.550 209.480 2639.870 209.540 ;
        RECT 735.610 209.340 735.930 209.400 ;
        RECT 2844.250 209.340 2844.570 209.400 ;
        RECT 2899.450 209.340 2899.770 209.400 ;
        RECT 735.610 209.200 2899.770 209.340 ;
        RECT 735.610 209.140 735.930 209.200 ;
        RECT 2844.250 209.140 2844.570 209.200 ;
        RECT 2899.450 209.140 2899.770 209.200 ;
        RECT 994.590 209.000 994.910 209.060 ;
        RECT 1538.770 209.000 1539.090 209.060 ;
        RECT 1812.470 209.000 1812.790 209.060 ;
        RECT 2086.630 209.000 2086.950 209.060 ;
        RECT 2360.790 209.000 2361.110 209.060 ;
        RECT 2633.570 209.000 2633.890 209.060 ;
        RECT 841.730 208.860 1904.470 209.000 ;
        RECT 468.810 207.640 469.130 207.700 ;
        RECT 841.730 207.640 841.870 208.860 ;
        RECT 994.590 208.800 994.910 208.860 ;
        RECT 1538.770 208.800 1539.090 208.860 ;
        RECT 1812.470 208.800 1812.790 208.860 ;
        RECT 468.810 207.500 841.870 207.640 ;
      LAYER met1 ;
        POLYGON 1199.065 208.500 1199.065 207.500 1198.065 207.500 ;
        RECT 1199.065 207.500 1262.345 208.500 ;
      LAYER met1 ;
        RECT 468.810 207.440 469.130 207.500 ;
      LAYER met1 ;
        POLYGON 1198.065 207.500 1198.065 207.440 1198.005 207.440 ;
        RECT 1198.065 207.440 1262.345 207.500 ;
        POLYGON 1198.005 207.440 1198.005 206.845 1197.410 206.845 ;
        RECT 1198.005 206.845 1262.345 207.440 ;
      LAYER met1 ;
        RECT 675.810 201.180 676.130 201.240 ;
        RECT 717.670 201.180 717.990 201.240 ;
        RECT 675.810 201.040 717.990 201.180 ;
        RECT 675.810 200.980 676.130 201.040 ;
        RECT 717.670 200.980 717.990 201.040 ;
        RECT 704.950 200.500 705.270 200.560 ;
        RECT 715.330 200.500 715.650 200.560 ;
        RECT 722.730 200.500 723.050 200.560 ;
        RECT 735.610 200.500 735.930 200.560 ;
        RECT 704.950 200.360 735.930 200.500 ;
        RECT 704.950 200.300 705.270 200.360 ;
        RECT 712.930 200.000 713.070 200.360 ;
        RECT 715.330 200.300 715.650 200.360 ;
        RECT 722.730 200.300 723.050 200.360 ;
        RECT 735.610 200.300 735.930 200.360 ;
      LAYER met1 ;
        RECT 663.000 199.390 704.700 199.815 ;
      LAYER met1 ;
        RECT 704.980 199.670 705.240 200.000 ;
      LAYER met1 ;
        RECT 705.520 199.390 706.565 199.815 ;
      LAYER met1 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met1 ;
        RECT 707.775 199.390 709.490 199.815 ;
      LAYER met1 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met1 ;
        RECT 710.700 199.390 712.585 199.815 ;
        RECT 398.320 198.080 456.965 199.030 ;
        RECT 398.320 197.965 399.460 198.080 ;
        POLYGON 399.460 198.080 399.575 198.080 399.460 197.965 ;
        POLYGON 455.535 198.080 455.650 198.080 455.650 197.965 ;
        RECT 455.650 197.965 456.965 198.080 ;
        RECT 395.380 0.275 468.815 197.965 ;
        RECT 663.000 189.745 712.585 199.390 ;
      LAYER met1 ;
        RECT 712.865 190.025 713.095 200.000 ;
      LAYER met1 ;
        RECT 713.375 199.390 715.060 199.815 ;
      LAYER met1 ;
        RECT 715.340 199.670 715.640 200.000 ;
      LAYER met1 ;
        RECT 715.920 199.390 722.585 199.815 ;
      LAYER met1 ;
        RECT 722.865 199.670 723.445 200.000 ;
      LAYER met1 ;
        RECT 723.725 199.390 725.175 199.815 ;
      LAYER met1 ;
        RECT 725.455 199.670 725.715 200.000 ;
      LAYER met1 ;
        RECT 725.995 199.390 738.000 199.815 ;
        RECT 713.375 189.745 738.000 199.390 ;
        RECT 663.000 104.105 738.000 189.745 ;
        RECT 932.000 180.515 1012.000 206.845 ;
        RECT 931.885 174.985 1012.000 180.515 ;
        RECT 932.000 169.880 1012.000 174.985 ;
        RECT 931.885 164.275 1012.000 169.880 ;
        RECT 932.000 148.780 1012.000 164.275 ;
        POLYGON 1197.410 206.845 1197.410 204.500 1195.065 204.500 ;
        RECT 1197.410 206.500 1262.345 206.845 ;
        POLYGON 1262.345 208.500 1264.345 206.500 1262.345 206.500 ;
      LAYER met1 ;
        RECT 1904.330 207.640 1904.470 208.860 ;
        RECT 2086.260 208.860 2086.950 209.000 ;
        RECT 2086.260 207.640 2086.400 208.860 ;
        RECT 2086.630 208.800 2086.950 208.860 ;
        RECT 2360.420 208.860 2361.110 209.000 ;
        RECT 2360.420 207.640 2360.560 208.860 ;
        RECT 2360.790 208.800 2361.110 208.860 ;
        RECT 2580.530 208.860 2633.890 209.000 ;
        RECT 2580.530 207.640 2580.670 208.860 ;
        RECT 2633.570 208.800 2633.890 208.860 ;
        RECT 1904.330 207.500 2580.670 207.640 ;
      LAYER met1 ;
        RECT 1197.410 204.500 1264.345 206.500 ;
        RECT 1195.065 200.980 1264.345 204.500 ;
        RECT 1195.065 198.980 1262.345 200.980 ;
        POLYGON 1262.345 200.980 1264.345 200.980 1262.345 198.980 ;
        RECT 1195.065 198.780 1260.505 198.980 ;
        RECT 1195.065 163.510 1204.800 198.780 ;
        RECT 1224.435 198.000 1260.505 198.780 ;
        RECT 1224.435 197.965 1264.345 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 931.885 142.810 1012.000 148.780 ;
        RECT 931.885 127.070 1012.115 142.810 ;
        POLYGON 931.885 127.070 931.940 127.070 931.940 127.015 ;
        RECT 931.940 119.365 1012.115 127.070 ;
        RECT 931.940 110.250 1012.000 119.365 ;
        RECT 931.940 108.520 1012.145 110.250 ;
        RECT 931.940 105.420 1012.000 108.520 ;
        RECT 932.000 104.105 1012.000 105.420 ;
        RECT 662.855 69.780 738.145 104.105 ;
        RECT 931.855 69.780 1012.115 104.105 ;
        RECT 663.000 68.725 738.000 69.780 ;
        RECT 932.000 68.725 1012.000 69.780 ;
        RECT 662.855 29.910 738.145 68.725 ;
        RECT 931.855 29.910 1012.115 68.725 ;
        RECT 663.000 0.790 738.000 29.910 ;
        RECT 932.000 21.100 1012.000 29.910 ;
        RECT 931.980 19.025 1012.000 21.100 ;
        RECT 932.000 0.000 1012.000 19.025 ;
        RECT 1206.000 0.160 1280.880 197.965 ;
        RECT 1475.000 180.515 1555.000 206.845 ;
        RECT 1749.000 180.515 1829.000 206.845 ;
        RECT 2023.000 180.515 2103.000 206.845 ;
        RECT 2297.000 180.515 2377.000 206.845 ;
        RECT 2571.000 180.515 2651.000 206.845 ;
        RECT 2849.320 198.080 2907.965 199.030 ;
        RECT 2849.320 197.965 2850.460 198.080 ;
        POLYGON 2850.460 198.080 2850.575 198.080 2850.460 197.965 ;
        POLYGON 2906.535 198.080 2906.650 198.080 2906.650 197.965 ;
        RECT 2906.650 197.965 2907.965 198.080 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.460 198.080 ;
        POLYGON 3119.460 198.080 3119.575 198.080 3119.460 197.965 ;
        POLYGON 3175.535 198.080 3175.650 198.080 3175.650 197.965 ;
        RECT 3175.650 197.965 3176.965 198.080 ;
        RECT 3180.145 197.965 3185.375 198.870 ;
        RECT 1474.885 174.985 1555.000 180.515 ;
        RECT 1748.885 174.985 1829.000 180.515 ;
        RECT 2022.885 174.985 2103.000 180.515 ;
        RECT 2296.885 174.985 2377.000 180.515 ;
        RECT 2570.885 174.985 2651.000 180.515 ;
        RECT 1475.000 169.880 1555.000 174.985 ;
        RECT 1749.000 169.880 1829.000 174.985 ;
        RECT 2023.000 169.880 2103.000 174.985 ;
        RECT 2297.000 169.880 2377.000 174.985 ;
        RECT 2571.000 169.880 2651.000 174.985 ;
        RECT 1474.885 164.275 1555.000 169.880 ;
        RECT 1748.885 164.275 1829.000 169.880 ;
        RECT 2022.885 164.275 2103.000 169.880 ;
        RECT 2296.885 164.275 2377.000 169.880 ;
        RECT 2570.885 164.275 2651.000 169.880 ;
        RECT 1475.000 148.780 1555.000 164.275 ;
        RECT 1749.000 148.780 1829.000 164.275 ;
        RECT 2023.000 148.780 2103.000 164.275 ;
        RECT 2297.000 148.780 2377.000 164.275 ;
        RECT 2571.000 148.780 2651.000 164.275 ;
        RECT 1474.885 142.810 1555.000 148.780 ;
        RECT 1748.885 142.810 1829.000 148.780 ;
        RECT 2022.885 142.810 2103.000 148.780 ;
        RECT 2296.885 142.810 2377.000 148.780 ;
        RECT 2570.885 142.810 2651.000 148.780 ;
        RECT 1474.885 127.070 1555.115 142.810 ;
        POLYGON 1474.885 127.070 1474.940 127.070 1474.940 127.015 ;
        RECT 1474.940 119.365 1555.115 127.070 ;
        RECT 1748.885 127.070 1829.115 142.810 ;
        POLYGON 1748.885 127.070 1748.940 127.070 1748.940 127.015 ;
        RECT 1748.940 119.365 1829.115 127.070 ;
        RECT 2022.885 127.070 2103.115 142.810 ;
        POLYGON 2022.885 127.070 2022.940 127.070 2022.940 127.015 ;
        RECT 2022.940 119.365 2103.115 127.070 ;
        RECT 2296.885 127.070 2377.115 142.810 ;
        POLYGON 2296.885 127.070 2296.940 127.070 2296.940 127.015 ;
        RECT 2296.940 119.365 2377.115 127.070 ;
        RECT 2570.885 127.070 2651.115 142.810 ;
        POLYGON 2570.885 127.070 2570.940 127.070 2570.940 127.015 ;
        RECT 2570.940 119.365 2651.115 127.070 ;
        RECT 1474.940 110.250 1555.000 119.365 ;
        RECT 1748.940 110.250 1829.000 119.365 ;
        RECT 2022.940 110.250 2103.000 119.365 ;
        RECT 2296.940 110.250 2377.000 119.365 ;
        RECT 2570.940 110.250 2651.000 119.365 ;
        RECT 1474.940 108.520 1555.145 110.250 ;
        RECT 1748.940 108.520 1829.145 110.250 ;
        RECT 2022.940 108.520 2103.145 110.250 ;
        RECT 2296.940 108.520 2377.145 110.250 ;
        RECT 2570.940 108.520 2651.145 110.250 ;
        RECT 1474.940 105.420 1555.000 108.520 ;
        RECT 1748.940 105.420 1829.000 108.520 ;
        RECT 2022.940 105.420 2103.000 108.520 ;
        RECT 2296.940 105.420 2377.000 108.520 ;
        RECT 2570.940 105.420 2651.000 108.520 ;
        RECT 1475.000 104.105 1555.000 105.420 ;
        RECT 1749.000 104.105 1829.000 105.420 ;
        RECT 2023.000 104.105 2103.000 105.420 ;
        RECT 2297.000 104.105 2377.000 105.420 ;
        RECT 2571.000 104.105 2651.000 105.420 ;
        RECT 1474.855 69.780 1555.115 104.105 ;
        RECT 1748.855 69.780 1829.115 104.105 ;
        RECT 2022.855 69.780 2103.115 104.105 ;
        RECT 2296.855 69.780 2377.115 104.105 ;
        RECT 2570.855 69.780 2651.115 104.105 ;
        RECT 1475.000 68.725 1555.000 69.780 ;
        RECT 1749.000 68.725 1829.000 69.780 ;
        RECT 2023.000 68.725 2103.000 69.780 ;
        RECT 2297.000 68.725 2377.000 69.780 ;
        RECT 2571.000 68.725 2651.000 69.780 ;
        RECT 1474.855 29.910 1555.115 68.725 ;
        RECT 1748.855 29.910 1829.115 68.725 ;
        RECT 2022.855 29.910 2103.115 68.725 ;
        RECT 2296.855 29.910 2377.115 68.725 ;
        RECT 2570.855 29.910 2651.115 68.725 ;
        RECT 1475.000 21.100 1555.000 29.910 ;
        RECT 1749.000 21.100 1829.000 29.910 ;
        RECT 2023.000 21.100 2103.000 29.910 ;
        RECT 2297.000 21.100 2377.000 29.910 ;
        RECT 2571.000 21.100 2651.000 29.910 ;
        RECT 1474.980 19.025 1555.000 21.100 ;
        RECT 1748.980 19.025 1829.000 21.100 ;
        RECT 2022.980 19.025 2103.000 21.100 ;
        RECT 2296.980 19.025 2377.000 21.100 ;
        RECT 2570.980 19.025 2651.000 21.100 ;
        RECT 1475.000 0.000 1555.000 19.025 ;
        RECT 1749.000 0.000 1829.000 19.025 ;
        RECT 2023.000 0.000 2103.000 19.025 ;
        RECT 2297.000 0.000 2377.000 19.025 ;
        RECT 2571.000 0.000 2651.000 19.025 ;
        RECT 2846.380 0.275 2919.815 197.965 ;
        RECT 3116.085 0.275 3188.815 197.965 ;
      LAYER via ;
        RECT 2925.240 4981.720 2925.500 4981.980 ;
        RECT 3373.740 4981.720 3374.000 4981.980 ;
        RECT 1780.300 4954.180 1780.560 4954.440 ;
        RECT 3367.760 4954.180 3368.020 4954.440 ;
        RECT 211.240 4950.780 211.500 4951.040 ;
        RECT 224.580 4950.440 224.840 4950.700 ;
        RECT 1718.200 4950.440 1718.460 4950.700 ;
        RECT 1780.300 4950.440 1780.560 4950.700 ;
        RECT 3367.300 4950.100 3367.560 4950.360 ;
        RECT 3367.760 4372.440 3368.020 4372.700 ;
        RECT 3376.960 4372.440 3377.220 4372.700 ;
        RECT 3367.300 4361.900 3367.560 4362.160 ;
        RECT 3368.220 4361.900 3368.480 4362.160 ;
        RECT 3376.960 4361.900 3377.220 4362.160 ;
        RECT 3369.140 4350.680 3369.400 4350.940 ;
        RECT 3376.960 4350.680 3377.220 4350.940 ;
        RECT 3367.300 4321.100 3367.560 4321.360 ;
        RECT 3376.960 4321.100 3377.220 4321.360 ;
        RECT 3369.140 4316.000 3369.400 4316.260 ;
        RECT 3376.960 4316.000 3377.220 4316.260 ;
        RECT 3376.500 4091.600 3376.760 4091.860 ;
        RECT 3388.000 4091.600 3388.260 4091.860 ;
        RECT 208.940 3988.580 209.200 3988.840 ;
        RECT 213.080 3988.580 213.340 3988.840 ;
        RECT 208.940 3956.620 209.200 3956.880 ;
        RECT 212.160 3956.620 212.420 3956.880 ;
        RECT 208.940 3941.320 209.200 3941.580 ;
        RECT 211.700 3941.320 211.960 3941.580 ;
        RECT 208.940 3936.220 209.200 3936.480 ;
        RECT 211.240 3935.200 211.500 3935.460 ;
        RECT 211.700 3934.860 211.960 3935.120 ;
        RECT 212.620 3934.860 212.880 3935.120 ;
        RECT 3367.760 3928.400 3368.020 3928.660 ;
        RECT 3376.960 3928.400 3377.220 3928.660 ;
        RECT 3368.220 3911.400 3368.480 3911.660 ;
        RECT 3376.960 3911.400 3377.220 3911.660 ;
        RECT 3376.040 3904.940 3376.300 3905.200 ;
        RECT 3376.960 3904.940 3377.220 3905.200 ;
        RECT 3367.300 3879.100 3367.560 3879.360 ;
        RECT 3376.960 3879.100 3377.220 3879.360 ;
        RECT 211.240 3787.980 211.500 3788.240 ;
        RECT 214.000 3787.980 214.260 3788.240 ;
        RECT 211.700 3787.640 211.960 3787.900 ;
        RECT 213.540 3787.640 213.800 3787.900 ;
        RECT 208.940 3777.100 209.200 3777.360 ;
        RECT 213.080 3777.100 213.340 3777.360 ;
        RECT 208.940 3738.340 209.200 3738.600 ;
        RECT 213.540 3738.340 213.800 3738.600 ;
        RECT 208.940 3719.980 209.200 3720.240 ;
        RECT 214.000 3719.980 214.260 3720.240 ;
        RECT 3367.760 3701.620 3368.020 3701.880 ;
        RECT 3369.140 3701.620 3369.400 3701.880 ;
        RECT 3376.960 3701.620 3377.220 3701.880 ;
        RECT 3368.220 3690.400 3368.480 3690.660 ;
        RECT 3376.960 3690.400 3377.220 3690.660 ;
        RECT 3367.300 3654.360 3367.560 3654.620 ;
        RECT 3370.060 3654.360 3370.320 3654.620 ;
        RECT 3376.960 3654.360 3377.220 3654.620 ;
        RECT 208.940 3561.200 209.200 3561.460 ;
        RECT 213.080 3561.200 213.340 3561.460 ;
        RECT 208.940 3519.720 209.200 3519.980 ;
        RECT 212.160 3519.720 212.420 3519.980 ;
        RECT 213.540 3519.720 213.800 3519.980 ;
        RECT 208.940 3504.080 209.200 3504.340 ;
        RECT 213.080 3504.080 213.340 3504.340 ;
        RECT 3367.300 3476.540 3367.560 3476.800 ;
        RECT 3369.140 3476.540 3369.400 3476.800 ;
        RECT 3376.960 3476.540 3377.220 3476.800 ;
        RECT 3369.600 3461.240 3369.860 3461.500 ;
        RECT 3376.960 3461.240 3377.220 3461.500 ;
        RECT 3367.760 3425.880 3368.020 3426.140 ;
        RECT 3370.060 3425.880 3370.320 3426.140 ;
        RECT 3376.960 3425.880 3377.220 3426.140 ;
        RECT 208.940 3340.540 209.200 3340.800 ;
        RECT 212.620 3340.540 212.880 3340.800 ;
        RECT 208.940 3305.180 209.200 3305.440 ;
        RECT 212.160 3305.180 212.420 3305.440 ;
        RECT 208.940 3293.280 209.200 3293.540 ;
        RECT 213.080 3293.280 213.340 3293.540 ;
        RECT 3367.300 3252.480 3367.560 3252.740 ;
        RECT 3376.960 3252.480 3377.220 3252.740 ;
        RECT 3367.300 3235.820 3367.560 3236.080 ;
        RECT 3368.220 3235.820 3368.480 3236.080 ;
        RECT 3367.300 3235.140 3367.560 3235.400 ;
        RECT 3369.600 3235.140 3369.860 3235.400 ;
        RECT 3376.960 3235.140 3377.220 3235.400 ;
        RECT 3376.040 3228.680 3376.300 3228.940 ;
        RECT 3376.960 3228.680 3377.220 3228.940 ;
        RECT 3367.760 3203.180 3368.020 3203.440 ;
        RECT 3376.960 3203.180 3377.220 3203.440 ;
        RECT 208.940 3124.640 209.200 3124.900 ;
        RECT 212.620 3124.640 212.880 3124.900 ;
        RECT 208.940 3092.340 209.200 3092.600 ;
        RECT 212.160 3092.340 212.420 3092.600 ;
        RECT 208.940 3077.380 209.200 3077.640 ;
        RECT 213.080 3077.380 213.340 3077.640 ;
        RECT 3368.220 3025.360 3368.480 3025.620 ;
        RECT 3376.960 3025.360 3377.220 3025.620 ;
        RECT 212.620 3015.840 212.880 3016.100 ;
        RECT 212.620 3014.820 212.880 3015.080 ;
        RECT 3367.300 3014.480 3367.560 3014.740 ;
        RECT 3376.960 3014.480 3377.220 3014.740 ;
        RECT 3367.760 2975.040 3368.020 2975.300 ;
        RECT 3376.960 2975.040 3377.220 2975.300 ;
        RECT 208.940 2908.400 209.200 2908.660 ;
        RECT 212.160 2908.400 212.420 2908.660 ;
        RECT 208.940 2876.100 209.200 2876.360 ;
        RECT 213.540 2876.100 213.800 2876.360 ;
        RECT 208.940 2861.140 209.200 2861.400 ;
        RECT 212.620 2861.140 212.880 2861.400 ;
        RECT 214.000 2861.140 214.260 2861.400 ;
        RECT 211.240 2855.700 211.500 2855.960 ;
        RECT 212.160 2855.700 212.420 2855.960 ;
        RECT 3368.220 2804.700 3368.480 2804.960 ;
        RECT 3376.960 2804.700 3377.220 2804.960 ;
        RECT 3367.300 2789.060 3367.560 2789.320 ;
        RECT 3376.960 2789.060 3377.220 2789.320 ;
        RECT 3376.040 2777.840 3376.300 2778.100 ;
        RECT 3376.960 2777.840 3377.220 2778.100 ;
        RECT 3367.760 2752.340 3368.020 2752.600 ;
        RECT 3376.960 2752.340 3377.220 2752.600 ;
        RECT 211.240 2715.280 211.500 2715.540 ;
        RECT 212.160 2715.280 212.420 2715.540 ;
        RECT 208.940 2697.260 209.200 2697.520 ;
        RECT 212.160 2697.260 212.420 2697.520 ;
        RECT 214.000 2697.260 214.260 2697.520 ;
        RECT 208.940 2655.780 209.200 2656.040 ;
        RECT 212.160 2655.780 212.420 2656.040 ;
        RECT 208.940 2640.140 209.200 2640.400 ;
        RECT 211.700 2640.140 211.960 2640.400 ;
        RECT 213.540 2640.140 213.800 2640.400 ;
        RECT 3376.500 2568.740 3376.760 2569.000 ;
        RECT 3388.460 2568.740 3388.720 2569.000 ;
        RECT 3373.740 2138.980 3374.000 2139.240 ;
        RECT 3387.540 2138.980 3387.800 2139.240 ;
        RECT 208.940 2054.660 209.200 2054.920 ;
        RECT 212.620 2054.660 212.880 2054.920 ;
        RECT 214.000 2054.660 214.260 2054.920 ;
        RECT 208.940 2022.360 209.200 2022.620 ;
        RECT 212.160 2022.360 212.420 2022.620 ;
        RECT 213.080 2022.360 213.340 2022.620 ;
        RECT 208.940 2004.000 209.200 2004.260 ;
        RECT 213.540 2004.000 213.800 2004.260 ;
        RECT 3367.760 1913.560 3368.020 1913.820 ;
        RECT 3376.960 1913.560 3377.220 1913.820 ;
        RECT 3368.680 1898.260 3368.940 1898.520 ;
        RECT 3376.960 1898.260 3377.220 1898.520 ;
        RECT 3367.300 1861.540 3367.560 1861.800 ;
        RECT 3369.600 1861.540 3369.860 1861.800 ;
        RECT 3376.960 1861.540 3377.220 1861.800 ;
        RECT 208.940 1847.600 209.200 1847.860 ;
        RECT 211.700 1847.600 211.960 1847.860 ;
        RECT 208.940 1843.180 209.200 1843.440 ;
        RECT 212.620 1843.180 212.880 1843.440 ;
        RECT 208.940 1812.920 209.200 1813.180 ;
        RECT 211.700 1812.920 211.960 1813.180 ;
        RECT 208.940 1803.400 209.200 1803.660 ;
        RECT 213.080 1803.400 213.340 1803.660 ;
        RECT 208.940 1786.060 209.200 1786.320 ;
        RECT 212.620 1786.060 212.880 1786.320 ;
        RECT 213.540 1786.060 213.800 1786.320 ;
        RECT 3367.760 1687.460 3368.020 1687.720 ;
        RECT 3376.960 1687.460 3377.220 1687.720 ;
        RECT 3368.680 1672.160 3368.940 1672.420 ;
        RECT 3370.060 1672.160 3370.320 1672.420 ;
        RECT 3376.960 1672.160 3377.220 1672.420 ;
        RECT 3369.600 1640.200 3369.860 1640.460 ;
        RECT 3376.960 1640.200 3377.220 1640.460 ;
        RECT 208.940 1627.280 209.200 1627.540 ;
        RECT 212.160 1627.280 212.420 1627.540 ;
        RECT 214.000 1627.280 214.260 1627.540 ;
        RECT 208.940 1585.800 209.200 1586.060 ;
        RECT 213.080 1585.800 213.340 1586.060 ;
        RECT 208.940 1570.160 209.200 1570.420 ;
        RECT 212.620 1570.160 212.880 1570.420 ;
        RECT 213.540 1570.160 213.800 1570.420 ;
        RECT 3367.300 1465.780 3367.560 1466.040 ;
        RECT 3376.960 1465.780 3377.220 1466.040 ;
        RECT 3367.760 1447.420 3368.020 1447.680 ;
        RECT 3370.060 1447.420 3370.320 1447.680 ;
        RECT 3376.960 1447.420 3377.220 1447.680 ;
        RECT 3369.600 1415.120 3369.860 1415.380 ;
        RECT 3376.960 1415.120 3377.220 1415.380 ;
        RECT 208.940 1406.620 209.200 1406.880 ;
        RECT 212.160 1406.620 212.420 1406.880 ;
        RECT 214.000 1406.620 214.260 1406.880 ;
        RECT 208.940 1372.620 209.200 1372.880 ;
        RECT 213.080 1372.620 213.340 1372.880 ;
        RECT 208.940 1359.360 209.200 1359.620 ;
        RECT 213.540 1359.360 213.800 1359.620 ;
        RECT 3367.300 1242.740 3367.560 1243.000 ;
        RECT 3370.060 1242.740 3370.320 1243.000 ;
        RECT 3376.960 1242.740 3377.220 1243.000 ;
        RECT 3367.760 1224.380 3368.020 1224.640 ;
        RECT 3376.960 1224.380 3377.220 1224.640 ;
        RECT 208.940 1190.380 209.200 1190.640 ;
        RECT 212.160 1190.380 212.420 1190.640 ;
        RECT 3369.600 1188.340 3369.860 1188.600 ;
        RECT 3376.960 1188.340 3377.220 1188.600 ;
        RECT 208.940 1158.420 209.200 1158.680 ;
        RECT 212.620 1158.420 212.880 1158.680 ;
        RECT 208.940 1143.120 209.200 1143.380 ;
        RECT 213.080 1143.120 213.340 1143.380 ;
        RECT 211.240 1137.340 211.500 1137.600 ;
        RECT 212.620 1137.340 212.880 1137.600 ;
        RECT 3370.060 1011.540 3370.320 1011.800 ;
        RECT 3376.960 1011.540 3377.220 1011.800 ;
        RECT 3367.760 996.240 3368.020 996.500 ;
        RECT 3376.960 996.240 3377.220 996.500 ;
        RECT 208.940 979.240 209.200 979.500 ;
        RECT 212.620 979.240 212.880 979.500 ;
        RECT 3369.600 959.520 3369.860 959.780 ;
        RECT 3376.960 959.520 3377.220 959.780 ;
        RECT 209.860 937.760 210.120 938.020 ;
        RECT 212.620 937.760 212.880 938.020 ;
        RECT 208.940 922.120 209.200 922.380 ;
        RECT 213.080 922.120 213.340 922.380 ;
        RECT 211.240 920.760 211.500 921.020 ;
        RECT 3367.300 791.560 3367.560 791.820 ;
        RECT 3370.060 791.560 3370.320 791.820 ;
        RECT 3376.960 791.560 3377.220 791.820 ;
        RECT 3367.760 775.920 3368.020 776.180 ;
        RECT 3376.960 775.920 3377.220 776.180 ;
        RECT 3368.680 734.440 3368.940 734.700 ;
        RECT 3369.600 734.440 3369.860 734.700 ;
        RECT 3376.960 734.440 3377.220 734.700 ;
        RECT 212.620 607.280 212.880 607.540 ;
        RECT 220.900 607.280 221.160 607.540 ;
        RECT 3367.300 565.800 3367.560 566.060 ;
        RECT 3376.960 565.800 3377.220 566.060 ;
        RECT 3367.760 547.440 3368.020 547.700 ;
        RECT 3376.960 547.440 3377.220 547.700 ;
        RECT 3368.680 508.340 3368.940 508.600 ;
        RECT 3376.960 508.340 3377.220 508.600 ;
        RECT 212.160 414.160 212.420 414.420 ;
        RECT 220.900 414.160 221.160 414.420 ;
        RECT 224.120 234.640 224.380 234.900 ;
        RECT 745.300 234.300 745.560 234.560 ;
        RECT 942.640 234.300 942.900 234.560 ;
        RECT 1004.280 234.300 1004.540 234.560 ;
        RECT 1281.200 234.300 1281.460 234.560 ;
        RECT 1488.660 234.300 1488.920 234.560 ;
        RECT 1547.080 234.300 1547.340 234.560 ;
        RECT 1762.820 234.300 1763.080 234.560 ;
        RECT 1821.240 234.300 1821.500 234.560 ;
        RECT 2036.980 234.300 2037.240 234.560 ;
        RECT 2095.400 234.300 2095.660 234.560 ;
        RECT 2310.680 234.300 2310.940 234.560 ;
        RECT 2369.100 234.300 2369.360 234.560 ;
        RECT 2584.840 234.300 2585.100 234.560 ;
        RECT 211.240 227.840 211.500 228.100 ;
        RECT 704.820 227.840 705.080 228.100 ;
        RECT 2618.880 227.840 2619.140 228.100 ;
        RECT 3367.760 227.840 3368.020 228.100 ;
        RECT 224.580 227.500 224.840 227.760 ;
        RECT 979.900 227.500 980.160 227.760 ;
        RECT 2593.580 227.500 2593.840 227.760 ;
        RECT 3368.680 227.500 3368.940 227.760 ;
        RECT 979.900 222.060 980.160 222.320 ;
        RECT 1522.700 222.060 1522.960 222.320 ;
        RECT 1531.440 222.060 1531.700 222.320 ;
        RECT 2033.760 222.060 2034.020 222.320 ;
        RECT 2307.460 222.060 2307.720 222.320 ;
        RECT 2344.720 222.060 2344.980 222.320 ;
        RECT 2618.880 222.060 2619.140 222.320 ;
        RECT 942.640 221.380 942.900 221.640 ;
        RECT 964.260 221.380 964.520 221.640 ;
        RECT 1007.500 221.380 1007.760 221.640 ;
        RECT 1485.440 221.380 1485.700 221.640 ;
        RECT 1497.860 221.380 1498.120 221.640 ;
        RECT 1528.680 221.380 1528.940 221.640 ;
        RECT 1759.600 221.720 1759.860 221.980 ;
        RECT 1772.020 221.720 1772.280 221.980 ;
        RECT 1802.840 221.720 1803.100 221.980 ;
        RECT 2033.760 221.380 2034.020 221.640 ;
        RECT 933.440 221.040 933.700 221.300 ;
        RECT 973.460 221.040 973.720 221.300 ;
        RECT 1476.240 220.700 1476.500 220.960 ;
        RECT 1516.260 220.700 1516.520 220.960 ;
        RECT 1531.440 220.700 1531.700 220.960 ;
        RECT 1796.860 221.040 1797.120 221.300 ;
        RECT 1750.400 220.700 1750.660 220.960 ;
        RECT 1790.420 220.700 1790.680 220.960 ;
        RECT 2071.020 220.700 2071.280 220.960 ;
        RECT 2344.720 221.380 2344.980 221.640 ;
        RECT 2307.460 221.040 2307.720 221.300 ;
        RECT 2581.620 221.040 2581.880 221.300 ;
        RECT 2593.580 221.040 2593.840 221.300 ;
        RECT 2899.480 213.560 2899.740 213.820 ;
        RECT 3367.300 213.560 3367.560 213.820 ;
        RECT 946.320 209.480 946.580 209.740 ;
        RECT 955.520 209.480 955.780 209.740 ;
        RECT 961.500 209.480 961.760 209.740 ;
        RECT 967.940 209.480 968.200 209.740 ;
        RECT 982.200 209.480 982.460 209.740 ;
        RECT 992.320 209.480 992.580 209.740 ;
        RECT 1000.600 209.480 1000.860 209.740 ;
        RECT 1489.580 209.480 1489.840 209.740 ;
        RECT 1503.380 209.480 1503.640 209.740 ;
        RECT 1511.200 209.480 1511.460 209.740 ;
        RECT 1526.380 209.480 1526.640 209.740 ;
        RECT 1532.820 209.480 1533.080 209.740 ;
        RECT 1543.400 209.480 1543.660 209.740 ;
        RECT 1763.280 209.480 1763.540 209.740 ;
        RECT 1777.540 209.480 1777.800 209.740 ;
        RECT 1784.900 209.480 1785.160 209.740 ;
        RECT 1799.160 209.480 1799.420 209.740 ;
        RECT 1805.600 209.480 1805.860 209.740 ;
        RECT 1817.560 209.480 1817.820 209.740 ;
        RECT 2037.440 209.480 2037.700 209.740 ;
        RECT 2051.240 209.480 2051.500 209.740 ;
        RECT 2057.680 209.480 2057.940 209.740 ;
        RECT 2072.860 209.480 2073.120 209.740 ;
        RECT 2079.300 209.480 2079.560 209.740 ;
        RECT 2091.260 209.480 2091.520 209.740 ;
        RECT 2311.600 209.480 2311.860 209.740 ;
        RECT 2325.400 209.480 2325.660 209.740 ;
        RECT 2331.840 209.480 2332.100 209.740 ;
        RECT 2347.020 209.480 2347.280 209.740 ;
        RECT 2353.460 209.480 2353.720 209.740 ;
        RECT 2365.420 209.480 2365.680 209.740 ;
        RECT 2585.300 209.480 2585.560 209.740 ;
        RECT 2599.560 209.480 2599.820 209.740 ;
        RECT 2606.000 209.480 2606.260 209.740 ;
        RECT 2621.180 209.480 2621.440 209.740 ;
        RECT 2627.620 209.480 2627.880 209.740 ;
        RECT 2639.580 209.480 2639.840 209.740 ;
        RECT 735.640 209.140 735.900 209.400 ;
        RECT 2844.280 209.140 2844.540 209.400 ;
        RECT 2899.480 209.140 2899.740 209.400 ;
        RECT 468.840 207.440 469.100 207.700 ;
        RECT 994.620 208.800 994.880 209.060 ;
        RECT 1538.800 208.800 1539.060 209.060 ;
        RECT 1812.500 208.800 1812.760 209.060 ;
        RECT 675.840 200.980 676.100 201.240 ;
        RECT 717.700 200.980 717.960 201.240 ;
        RECT 704.980 200.300 705.240 200.560 ;
        RECT 715.360 200.300 715.620 200.560 ;
        RECT 722.760 200.300 723.020 200.560 ;
        RECT 735.640 200.300 735.900 200.560 ;
        RECT 2086.660 208.800 2086.920 209.060 ;
        RECT 2360.820 208.800 2361.080 209.060 ;
        RECT 2633.600 208.800 2633.860 209.060 ;
      LAYER met2 ;
        RECT 385.250 5034.255 451.440 5036.855 ;
        RECT 642.250 5034.255 708.440 5036.855 ;
        RECT 899.250 5034.255 965.440 5036.855 ;
        RECT 1152.265 5013.940 1226.290 5183.075 ;
        RECT 1410.265 5013.940 1484.290 5183.075 ;
        RECT 1152.265 4990.335 1202.110 5013.940 ;
        RECT 1410.265 4990.335 1460.110 5013.940 ;
        RECT 1176.675 4990.035 1202.110 4990.335 ;
        RECT 1434.675 4990.035 1460.110 4990.335 ;
        RECT 1667.265 4990.035 1741.290 5183.075 ;
        RECT 1923.250 5034.255 1989.440 5036.855 ;
        RECT 2368.250 5034.255 2434.440 5036.855 ;
        RECT 2625.250 5034.255 2691.440 5036.855 ;
        RECT 2878.265 4990.035 2952.290 5183.075 ;
        RECT 3134.250 5034.255 3200.440 5036.855 ;
        RECT 1177.895 4988.000 1179.895 4989.920 ;
        RECT 1435.895 4988.000 1437.895 4989.920 ;
        RECT 1667.495 4988.000 1691.395 4990.035 ;
        RECT 1692.895 4988.000 1694.895 4989.920 ;
        RECT 1717.390 4988.000 1741.290 4990.035 ;
        RECT 2878.495 4988.000 2902.395 4990.035 ;
        RECT 2903.895 4988.000 2905.895 4989.920 ;
        RECT 2928.390 4988.000 2952.290 4990.035 ;
      LAYER met2 ;
        RECT 2925.230 4987.275 2925.510 4987.645 ;
        RECT 1718.190 4985.235 1718.470 4985.605 ;
        RECT 211.240 4950.750 211.500 4951.070 ;
      LAYER met2 ;
        RECT 151.145 4775.250 153.745 4841.440 ;
        RECT 0.035 4636.200 151.405 4645.935 ;
        RECT 153.765 4635.000 158.415 4646.140 ;
        RECT 160.165 4636.200 174.575 4645.935 ;
        RECT 0.035 4634.700 197.965 4635.000 ;
        RECT 0.035 4614.095 198.000 4634.700 ;
        RECT 0.035 4613.535 197.965 4614.095 ;
        RECT 0.035 4580.925 198.000 4613.535 ;
        RECT 0.035 4580.495 197.965 4580.925 ;
        RECT 0.035 4560.500 198.000 4580.495 ;
        RECT 0.035 4560.000 197.965 4560.500 ;
        RECT 153.800 4549.025 158.450 4560.000 ;
        RECT 4.925 4399.390 200.000 4423.290 ;
        RECT 4.925 4373.395 197.965 4399.390 ;
        RECT 198.080 4374.895 200.000 4376.895 ;
        RECT 4.925 4349.495 200.000 4373.395 ;
        RECT 4.925 4349.265 197.965 4349.495 ;
        RECT 4.925 4188.390 200.000 4212.290 ;
        RECT 4.925 4162.395 197.965 4188.390 ;
        RECT 198.080 4163.895 200.000 4165.895 ;
        RECT 4.925 4138.495 200.000 4162.395 ;
        RECT 4.925 4138.265 197.965 4138.495 ;
        RECT 0.000 4000.865 208.565 4001.915 ;
        RECT 0.000 4000.025 208.285 4000.865 ;
      LAYER met2 ;
        RECT 211.300 4000.850 211.440 4950.750 ;
        RECT 1718.260 4950.730 1718.400 4985.235 ;
        RECT 2925.300 4982.010 2925.440 4987.275 ;
        RECT 2925.240 4981.690 2925.500 4982.010 ;
        RECT 3373.740 4981.690 3374.000 4982.010 ;
        RECT 1780.300 4954.150 1780.560 4954.470 ;
        RECT 3367.760 4954.150 3368.020 4954.470 ;
        RECT 1780.360 4950.730 1780.500 4954.150 ;
        RECT 224.580 4950.410 224.840 4950.730 ;
        RECT 1718.200 4950.410 1718.460 4950.730 ;
        RECT 1780.300 4950.410 1780.560 4950.730 ;
        RECT 224.640 4443.670 224.780 4950.410 ;
        RECT 3367.300 4950.070 3367.560 4950.390 ;
        RECT 224.180 4443.530 224.780 4443.670 ;
        RECT 224.180 4350.485 224.320 4443.530 ;
        RECT 3367.360 4362.190 3367.500 4950.070 ;
        RECT 3367.820 4372.730 3367.960 4954.150 ;
        RECT 3367.760 4372.410 3368.020 4372.730 ;
        RECT 3367.300 4361.870 3367.560 4362.190 ;
        RECT 211.690 4350.115 211.970 4350.485 ;
        RECT 224.110 4350.115 224.390 4350.485 ;
        RECT 211.760 4029.670 211.900 4350.115 ;
        RECT 3367.300 4321.070 3367.560 4321.390 ;
        RECT 211.760 4029.530 212.360 4029.670 ;
        RECT 211.300 4000.710 211.900 4000.850 ;
        RECT 208.565 4000.515 210.965 4000.585 ;
        RECT 208.565 4000.375 211.440 4000.515 ;
        RECT 208.565 4000.305 210.965 4000.375 ;
      LAYER met2 ;
        RECT 0.000 3997.645 208.565 4000.025 ;
        RECT 0.000 3996.805 208.285 3997.645 ;
        RECT 0.000 3994.425 208.565 3996.805 ;
        RECT 0.000 3993.585 208.285 3994.425 ;
      LAYER met2 ;
        RECT 208.565 3993.865 210.965 3994.145 ;
      LAYER met2 ;
        RECT 0.000 3991.665 208.565 3993.585 ;
        RECT 0.000 3990.825 208.285 3991.665 ;
      LAYER met2 ;
        RECT 208.565 3991.105 210.965 3991.385 ;
      LAYER met2 ;
        RECT 0.000 3988.445 208.565 3990.825 ;
      LAYER met2 ;
        RECT 209.000 3988.870 209.140 3991.105 ;
        RECT 208.940 3988.550 209.200 3988.870 ;
      LAYER met2 ;
        RECT 0.000 3987.605 208.285 3988.445 ;
        RECT 0.000 3985.225 208.565 3987.605 ;
        RECT 0.000 3984.385 208.285 3985.225 ;
        RECT 0.000 3982.465 208.565 3984.385 ;
        RECT 0.000 3981.625 208.285 3982.465 ;
      LAYER met2 ;
        RECT 208.565 3981.905 210.965 3982.185 ;
      LAYER met2 ;
        RECT 0.000 3979.245 208.565 3981.625 ;
        RECT 0.000 3978.405 208.285 3979.245 ;
        RECT 0.000 3976.025 208.565 3978.405 ;
        RECT 0.000 3975.185 208.285 3976.025 ;
        RECT 0.000 3973.265 208.565 3975.185 ;
        RECT 0.000 3972.425 208.285 3973.265 ;
        RECT 0.000 3970.045 208.565 3972.425 ;
        RECT 0.000 3969.205 208.285 3970.045 ;
        RECT 0.000 3966.825 208.565 3969.205 ;
        RECT 0.000 3965.985 208.285 3966.825 ;
        RECT 0.000 3964.065 208.565 3965.985 ;
        RECT 0.000 3963.225 208.285 3964.065 ;
        RECT 0.000 3960.845 208.565 3963.225 ;
      LAYER met2 ;
        RECT 211.300 3961.410 211.440 4000.375 ;
        RECT 209.460 3961.270 211.440 3961.410 ;
      LAYER met2 ;
        RECT 0.000 3960.005 208.285 3960.845 ;
      LAYER met2 ;
        RECT 209.460 3960.565 209.600 3961.270 ;
        RECT 208.565 3960.285 210.965 3960.565 ;
      LAYER met2 ;
        RECT 0.000 3957.625 208.565 3960.005 ;
        RECT 0.000 3956.785 208.285 3957.625 ;
        RECT 0.000 3954.405 208.565 3956.785 ;
      LAYER met2 ;
        RECT 208.940 3956.590 209.200 3956.910 ;
      LAYER met2 ;
        RECT 0.000 3953.565 208.285 3954.405 ;
      LAYER met2 ;
        RECT 209.000 3954.125 209.140 3956.590 ;
        RECT 208.565 3953.845 210.965 3954.125 ;
        RECT 208.610 3953.790 209.140 3953.845 ;
      LAYER met2 ;
        RECT 0.000 3951.645 208.565 3953.565 ;
        RECT 0.000 3950.805 208.285 3951.645 ;
        RECT 0.000 3948.425 208.565 3950.805 ;
        RECT 0.000 3947.585 208.285 3948.425 ;
        RECT 0.000 3945.205 208.565 3947.585 ;
        RECT 0.000 3944.365 208.285 3945.205 ;
        RECT 0.000 3942.445 208.565 3944.365 ;
        RECT 0.000 3941.605 208.285 3942.445 ;
      LAYER met2 ;
        RECT 211.760 3941.610 211.900 4000.710 ;
        RECT 212.220 3956.910 212.360 4029.530 ;
        RECT 213.080 3988.550 213.340 3988.870 ;
        RECT 212.160 3956.590 212.420 3956.910 ;
      LAYER met2 ;
        RECT 0.000 3939.225 208.565 3941.605 ;
      LAYER met2 ;
        RECT 208.940 3941.290 209.200 3941.610 ;
        RECT 211.700 3941.290 211.960 3941.610 ;
      LAYER met2 ;
        RECT 0.000 3938.385 208.285 3939.225 ;
      LAYER met2 ;
        RECT 209.000 3938.970 209.140 3941.290 ;
        RECT 208.610 3938.945 209.140 3938.970 ;
        RECT 208.565 3938.665 210.965 3938.945 ;
      LAYER met2 ;
        RECT 0.000 3936.005 208.565 3938.385 ;
      LAYER met2 ;
        RECT 209.000 3936.510 209.140 3938.665 ;
        RECT 212.220 3936.930 212.360 3956.590 ;
        RECT 212.220 3936.790 212.820 3936.930 ;
        RECT 208.940 3936.190 209.200 3936.510 ;
      LAYER met2 ;
        RECT 0.000 3935.165 208.285 3936.005 ;
      LAYER met2 ;
        RECT 211.240 3935.170 211.500 3935.490 ;
      LAYER met2 ;
        RECT 0.000 3933.245 208.565 3935.165 ;
        RECT 0.000 3932.405 208.285 3933.245 ;
        RECT 0.000 3930.025 208.565 3932.405 ;
        RECT 0.000 3929.185 208.285 3930.025 ;
        RECT 0.000 3926.805 208.565 3929.185 ;
        RECT 0.000 3925.965 208.285 3926.805 ;
        RECT 0.000 3924.045 208.565 3925.965 ;
        RECT 0.000 3923.205 208.285 3924.045 ;
        RECT 0.000 3922.210 208.565 3923.205 ;
      LAYER met2 ;
        RECT 211.300 3788.270 211.440 3935.170 ;
        RECT 212.680 3935.150 212.820 3936.790 ;
        RECT 211.700 3934.830 211.960 3935.150 ;
        RECT 212.620 3934.830 212.880 3935.150 ;
        RECT 211.240 3787.950 211.500 3788.270 ;
        RECT 211.760 3787.930 211.900 3934.830 ;
        RECT 211.700 3787.610 211.960 3787.930 ;
      LAYER met2 ;
        RECT 0.000 3784.865 208.565 3785.915 ;
        RECT 0.000 3784.025 208.285 3784.865 ;
      LAYER met2 ;
        RECT 208.610 3784.585 211.440 3784.610 ;
        RECT 208.565 3784.470 211.440 3784.585 ;
        RECT 208.565 3784.305 210.965 3784.470 ;
      LAYER met2 ;
        RECT 0.000 3781.645 208.565 3784.025 ;
        RECT 0.000 3780.805 208.285 3781.645 ;
        RECT 0.000 3778.425 208.565 3780.805 ;
        RECT 0.000 3777.585 208.285 3778.425 ;
      LAYER met2 ;
        RECT 208.565 3777.865 210.965 3778.145 ;
      LAYER met2 ;
        RECT 0.000 3775.665 208.565 3777.585 ;
      LAYER met2 ;
        RECT 208.940 3777.070 209.200 3777.390 ;
      LAYER met2 ;
        RECT 0.000 3774.825 208.285 3775.665 ;
      LAYER met2 ;
        RECT 209.000 3775.385 209.140 3777.070 ;
        RECT 208.565 3775.105 210.965 3775.385 ;
      LAYER met2 ;
        RECT 0.000 3772.445 208.565 3774.825 ;
        RECT 0.000 3771.605 208.285 3772.445 ;
        RECT 0.000 3769.225 208.565 3771.605 ;
        RECT 0.000 3768.385 208.285 3769.225 ;
        RECT 0.000 3766.465 208.565 3768.385 ;
        RECT 0.000 3765.625 208.285 3766.465 ;
      LAYER met2 ;
        RECT 208.565 3765.905 210.965 3766.185 ;
      LAYER met2 ;
        RECT 0.000 3763.245 208.565 3765.625 ;
        RECT 0.000 3762.405 208.285 3763.245 ;
        RECT 0.000 3760.025 208.565 3762.405 ;
        RECT 0.000 3759.185 208.285 3760.025 ;
        RECT 0.000 3757.265 208.565 3759.185 ;
        RECT 0.000 3756.425 208.285 3757.265 ;
        RECT 0.000 3754.045 208.565 3756.425 ;
        RECT 0.000 3753.205 208.285 3754.045 ;
        RECT 0.000 3750.825 208.565 3753.205 ;
        RECT 0.000 3749.985 208.285 3750.825 ;
        RECT 0.000 3748.065 208.565 3749.985 ;
        RECT 0.000 3747.225 208.285 3748.065 ;
        RECT 0.000 3744.845 208.565 3747.225 ;
      LAYER met2 ;
        RECT 211.300 3745.170 211.440 3784.470 ;
        RECT 213.140 3777.390 213.280 3988.550 ;
        RECT 3367.360 3879.390 3367.500 4321.070 ;
        RECT 3367.820 3928.690 3367.960 4372.410 ;
        RECT 3368.220 4361.870 3368.480 4362.190 ;
        RECT 3367.760 3928.370 3368.020 3928.690 ;
        RECT 3367.300 3879.070 3367.560 3879.390 ;
        RECT 214.000 3787.950 214.260 3788.270 ;
        RECT 213.540 3787.610 213.800 3787.930 ;
        RECT 213.080 3777.070 213.340 3777.390 ;
        RECT 209.000 3745.030 211.440 3745.170 ;
      LAYER met2 ;
        RECT 0.000 3744.005 208.285 3744.845 ;
      LAYER met2 ;
        RECT 209.000 3744.565 209.140 3745.030 ;
        RECT 208.565 3744.285 210.965 3744.565 ;
      LAYER met2 ;
        RECT 0.000 3741.625 208.565 3744.005 ;
        RECT 0.000 3740.785 208.285 3741.625 ;
        RECT 0.000 3738.405 208.565 3740.785 ;
        RECT 0.000 3737.565 208.285 3738.405 ;
      LAYER met2 ;
        RECT 208.940 3738.310 209.200 3738.630 ;
        RECT 209.000 3738.125 209.140 3738.310 ;
        RECT 208.565 3737.845 210.965 3738.125 ;
      LAYER met2 ;
        RECT 0.000 3735.645 208.565 3737.565 ;
        RECT 0.000 3734.805 208.285 3735.645 ;
        RECT 0.000 3732.425 208.565 3734.805 ;
        RECT 0.000 3731.585 208.285 3732.425 ;
        RECT 0.000 3729.205 208.565 3731.585 ;
        RECT 0.000 3728.365 208.285 3729.205 ;
        RECT 0.000 3726.445 208.565 3728.365 ;
        RECT 0.000 3725.605 208.285 3726.445 ;
        RECT 0.000 3723.225 208.565 3725.605 ;
        RECT 0.000 3722.385 208.285 3723.225 ;
      LAYER met2 ;
        RECT 208.565 3722.665 210.965 3722.945 ;
      LAYER met2 ;
        RECT 0.000 3720.005 208.565 3722.385 ;
      LAYER met2 ;
        RECT 209.000 3720.270 209.140 3722.665 ;
      LAYER met2 ;
        RECT 0.000 3719.165 208.285 3720.005 ;
      LAYER met2 ;
        RECT 208.940 3719.950 209.200 3720.270 ;
      LAYER met2 ;
        RECT 0.000 3717.245 208.565 3719.165 ;
        RECT 0.000 3716.405 208.285 3717.245 ;
        RECT 0.000 3714.025 208.565 3716.405 ;
        RECT 0.000 3713.185 208.285 3714.025 ;
        RECT 0.000 3710.805 208.565 3713.185 ;
        RECT 0.000 3709.965 208.285 3710.805 ;
        RECT 0.000 3708.045 208.565 3709.965 ;
        RECT 0.000 3707.205 208.285 3708.045 ;
        RECT 0.000 3706.210 208.565 3707.205 ;
        RECT 0.000 3568.865 208.565 3569.915 ;
        RECT 0.000 3568.025 208.285 3568.865 ;
      LAYER met2 ;
        RECT 208.565 3568.515 210.965 3568.585 ;
        RECT 208.565 3568.375 211.440 3568.515 ;
        RECT 208.565 3568.305 210.965 3568.375 ;
      LAYER met2 ;
        RECT 0.000 3565.645 208.565 3568.025 ;
        RECT 0.000 3564.805 208.285 3565.645 ;
        RECT 0.000 3562.425 208.565 3564.805 ;
        RECT 0.000 3561.585 208.285 3562.425 ;
      LAYER met2 ;
        RECT 208.565 3561.865 210.965 3562.145 ;
      LAYER met2 ;
        RECT 0.000 3559.665 208.565 3561.585 ;
      LAYER met2 ;
        RECT 208.940 3561.170 209.200 3561.490 ;
      LAYER met2 ;
        RECT 0.000 3558.825 208.285 3559.665 ;
      LAYER met2 ;
        RECT 209.000 3559.385 209.140 3561.170 ;
        RECT 208.565 3559.105 210.965 3559.385 ;
      LAYER met2 ;
        RECT 0.000 3556.445 208.565 3558.825 ;
        RECT 0.000 3555.605 208.285 3556.445 ;
        RECT 0.000 3553.225 208.565 3555.605 ;
        RECT 0.000 3552.385 208.285 3553.225 ;
        RECT 0.000 3550.465 208.565 3552.385 ;
        RECT 0.000 3549.625 208.285 3550.465 ;
      LAYER met2 ;
        RECT 208.565 3549.905 210.965 3550.185 ;
      LAYER met2 ;
        RECT 0.000 3547.245 208.565 3549.625 ;
        RECT 0.000 3546.405 208.285 3547.245 ;
        RECT 0.000 3544.025 208.565 3546.405 ;
        RECT 0.000 3543.185 208.285 3544.025 ;
        RECT 0.000 3541.265 208.565 3543.185 ;
        RECT 0.000 3540.425 208.285 3541.265 ;
        RECT 0.000 3538.045 208.565 3540.425 ;
        RECT 0.000 3537.205 208.285 3538.045 ;
        RECT 0.000 3534.825 208.565 3537.205 ;
        RECT 0.000 3533.985 208.285 3534.825 ;
        RECT 0.000 3532.065 208.565 3533.985 ;
        RECT 0.000 3531.225 208.285 3532.065 ;
        RECT 0.000 3528.845 208.565 3531.225 ;
      LAYER met2 ;
        RECT 211.300 3530.970 211.440 3568.375 ;
        RECT 213.140 3561.490 213.280 3777.070 ;
        RECT 213.600 3738.630 213.740 3787.610 ;
        RECT 213.540 3738.310 213.800 3738.630 ;
        RECT 213.080 3561.170 213.340 3561.490 ;
        RECT 213.140 3546.670 213.280 3561.170 ;
        RECT 209.460 3530.830 211.440 3530.970 ;
        RECT 212.680 3546.530 213.280 3546.670 ;
      LAYER met2 ;
        RECT 0.000 3528.005 208.285 3528.845 ;
      LAYER met2 ;
        RECT 209.460 3528.565 209.600 3530.830 ;
        RECT 208.565 3528.285 210.965 3528.565 ;
      LAYER met2 ;
        RECT 0.000 3525.625 208.565 3528.005 ;
        RECT 0.000 3524.785 208.285 3525.625 ;
        RECT 0.000 3522.405 208.565 3524.785 ;
        RECT 0.000 3521.565 208.285 3522.405 ;
      LAYER met2 ;
        RECT 208.610 3522.125 209.140 3522.130 ;
        RECT 208.565 3521.845 210.965 3522.125 ;
      LAYER met2 ;
        RECT 0.000 3519.645 208.565 3521.565 ;
      LAYER met2 ;
        RECT 209.000 3520.010 209.140 3521.845 ;
        RECT 208.940 3519.690 209.200 3520.010 ;
        RECT 212.160 3519.690 212.420 3520.010 ;
      LAYER met2 ;
        RECT 0.000 3518.805 208.285 3519.645 ;
        RECT 0.000 3516.425 208.565 3518.805 ;
        RECT 0.000 3515.585 208.285 3516.425 ;
        RECT 0.000 3513.205 208.565 3515.585 ;
        RECT 0.000 3512.365 208.285 3513.205 ;
        RECT 0.000 3510.445 208.565 3512.365 ;
        RECT 0.000 3509.605 208.285 3510.445 ;
        RECT 0.000 3507.225 208.565 3509.605 ;
        RECT 0.000 3506.385 208.285 3507.225 ;
      LAYER met2 ;
        RECT 208.565 3506.665 210.965 3506.945 ;
      LAYER met2 ;
        RECT 0.000 3504.005 208.565 3506.385 ;
      LAYER met2 ;
        RECT 209.000 3504.370 209.140 3506.665 ;
        RECT 208.940 3504.050 209.200 3504.370 ;
      LAYER met2 ;
        RECT 0.000 3503.165 208.285 3504.005 ;
        RECT 0.000 3501.245 208.565 3503.165 ;
        RECT 0.000 3500.405 208.285 3501.245 ;
        RECT 0.000 3498.025 208.565 3500.405 ;
        RECT 0.000 3497.185 208.285 3498.025 ;
        RECT 0.000 3494.805 208.565 3497.185 ;
        RECT 0.000 3493.965 208.285 3494.805 ;
        RECT 0.000 3492.045 208.565 3493.965 ;
        RECT 0.000 3491.205 208.285 3492.045 ;
        RECT 0.000 3490.210 208.565 3491.205 ;
        RECT 0.000 3352.865 208.565 3353.915 ;
        RECT 0.000 3352.025 208.285 3352.865 ;
      LAYER met2 ;
        RECT 208.565 3352.515 210.965 3352.585 ;
        RECT 208.565 3352.375 211.440 3352.515 ;
        RECT 208.565 3352.305 210.965 3352.375 ;
      LAYER met2 ;
        RECT 0.000 3349.645 208.565 3352.025 ;
        RECT 0.000 3348.805 208.285 3349.645 ;
        RECT 0.000 3346.425 208.565 3348.805 ;
        RECT 0.000 3345.585 208.285 3346.425 ;
      LAYER met2 ;
        RECT 208.565 3345.865 210.965 3346.145 ;
      LAYER met2 ;
        RECT 0.000 3343.665 208.565 3345.585 ;
        RECT 0.000 3342.825 208.285 3343.665 ;
      LAYER met2 ;
        RECT 208.565 3343.105 210.965 3343.385 ;
      LAYER met2 ;
        RECT 0.000 3340.445 208.565 3342.825 ;
      LAYER met2 ;
        RECT 209.000 3340.830 209.140 3343.105 ;
        RECT 208.940 3340.510 209.200 3340.830 ;
      LAYER met2 ;
        RECT 0.000 3339.605 208.285 3340.445 ;
        RECT 0.000 3337.225 208.565 3339.605 ;
        RECT 0.000 3336.385 208.285 3337.225 ;
        RECT 0.000 3334.465 208.565 3336.385 ;
        RECT 0.000 3333.625 208.285 3334.465 ;
      LAYER met2 ;
        RECT 208.565 3333.905 210.965 3334.185 ;
      LAYER met2 ;
        RECT 0.000 3331.245 208.565 3333.625 ;
        RECT 0.000 3330.405 208.285 3331.245 ;
        RECT 0.000 3328.025 208.565 3330.405 ;
        RECT 0.000 3327.185 208.285 3328.025 ;
        RECT 0.000 3325.265 208.565 3327.185 ;
        RECT 0.000 3324.425 208.285 3325.265 ;
        RECT 0.000 3322.045 208.565 3324.425 ;
        RECT 0.000 3321.205 208.285 3322.045 ;
        RECT 0.000 3318.825 208.565 3321.205 ;
        RECT 0.000 3317.985 208.285 3318.825 ;
        RECT 0.000 3316.065 208.565 3317.985 ;
        RECT 0.000 3315.225 208.285 3316.065 ;
        RECT 0.000 3312.845 208.565 3315.225 ;
        RECT 0.000 3312.005 208.285 3312.845 ;
      LAYER met2 ;
        RECT 211.300 3312.690 211.440 3352.375 ;
        RECT 208.540 3312.550 211.440 3312.690 ;
        RECT 208.540 3312.425 210.965 3312.550 ;
        RECT 208.565 3312.285 210.965 3312.425 ;
      LAYER met2 ;
        RECT 0.000 3309.625 208.565 3312.005 ;
        RECT 0.000 3308.785 208.285 3309.625 ;
        RECT 0.000 3306.405 208.565 3308.785 ;
        RECT 0.000 3305.565 208.285 3306.405 ;
      LAYER met2 ;
        RECT 208.565 3305.845 210.965 3306.125 ;
      LAYER met2 ;
        RECT 0.000 3303.645 208.565 3305.565 ;
      LAYER met2 ;
        RECT 209.000 3305.470 209.140 3305.845 ;
        RECT 212.220 3305.470 212.360 3519.690 ;
        RECT 212.680 3340.830 212.820 3546.530 ;
        RECT 213.600 3520.010 213.740 3738.310 ;
        RECT 214.060 3720.270 214.200 3787.950 ;
        RECT 214.000 3719.950 214.260 3720.270 ;
        RECT 213.540 3519.690 213.800 3520.010 ;
        RECT 214.060 3504.450 214.200 3719.950 ;
        RECT 3367.360 3654.650 3367.500 3879.070 ;
        RECT 3367.820 3701.910 3367.960 3928.370 ;
        RECT 3368.280 3911.690 3368.420 4361.870 ;
        RECT 3369.140 4350.650 3369.400 4350.970 ;
        RECT 3369.200 4316.290 3369.340 4350.650 ;
        RECT 3369.140 4315.970 3369.400 4316.290 ;
        RECT 3368.220 3911.370 3368.480 3911.690 ;
        RECT 3367.760 3701.590 3368.020 3701.910 ;
        RECT 3368.280 3690.690 3368.420 3911.370 ;
        RECT 3369.140 3701.590 3369.400 3701.910 ;
        RECT 3368.220 3690.370 3368.480 3690.690 ;
        RECT 3367.300 3654.330 3367.560 3654.650 ;
        RECT 213.140 3504.370 214.200 3504.450 ;
        RECT 213.080 3504.310 214.200 3504.370 ;
        RECT 213.080 3504.050 213.340 3504.310 ;
        RECT 212.620 3340.510 212.880 3340.830 ;
        RECT 208.940 3305.150 209.200 3305.470 ;
        RECT 212.160 3305.150 212.420 3305.470 ;
      LAYER met2 ;
        RECT 0.000 3302.805 208.285 3303.645 ;
        RECT 0.000 3300.425 208.565 3302.805 ;
        RECT 0.000 3299.585 208.285 3300.425 ;
        RECT 0.000 3297.205 208.565 3299.585 ;
        RECT 0.000 3296.365 208.285 3297.205 ;
        RECT 0.000 3294.445 208.565 3296.365 ;
        RECT 0.000 3293.605 208.285 3294.445 ;
        RECT 0.000 3291.225 208.565 3293.605 ;
      LAYER met2 ;
        RECT 208.940 3293.250 209.200 3293.570 ;
      LAYER met2 ;
        RECT 0.000 3290.385 208.285 3291.225 ;
      LAYER met2 ;
        RECT 209.000 3290.945 209.140 3293.250 ;
        RECT 208.565 3290.665 210.965 3290.945 ;
      LAYER met2 ;
        RECT 0.000 3288.005 208.565 3290.385 ;
        RECT 0.000 3287.165 208.285 3288.005 ;
        RECT 0.000 3285.245 208.565 3287.165 ;
        RECT 0.000 3284.405 208.285 3285.245 ;
        RECT 0.000 3282.025 208.565 3284.405 ;
        RECT 0.000 3281.185 208.285 3282.025 ;
        RECT 0.000 3278.805 208.565 3281.185 ;
        RECT 0.000 3277.965 208.285 3278.805 ;
        RECT 0.000 3276.045 208.565 3277.965 ;
        RECT 0.000 3275.205 208.285 3276.045 ;
        RECT 0.000 3274.210 208.565 3275.205 ;
        RECT 0.000 3136.865 208.565 3137.915 ;
        RECT 0.000 3136.025 208.285 3136.865 ;
      LAYER met2 ;
        RECT 208.565 3136.570 210.965 3136.585 ;
        RECT 208.565 3136.430 211.440 3136.570 ;
        RECT 208.565 3136.305 210.965 3136.430 ;
      LAYER met2 ;
        RECT 0.000 3133.645 208.565 3136.025 ;
        RECT 0.000 3132.805 208.285 3133.645 ;
        RECT 0.000 3130.425 208.565 3132.805 ;
        RECT 0.000 3129.585 208.285 3130.425 ;
      LAYER met2 ;
        RECT 208.565 3129.865 210.965 3130.145 ;
      LAYER met2 ;
        RECT 0.000 3127.665 208.565 3129.585 ;
        RECT 0.000 3126.825 208.285 3127.665 ;
      LAYER met2 ;
        RECT 208.565 3127.105 210.965 3127.385 ;
      LAYER met2 ;
        RECT 0.000 3124.445 208.565 3126.825 ;
      LAYER met2 ;
        RECT 209.000 3124.930 209.140 3127.105 ;
        RECT 208.940 3124.610 209.200 3124.930 ;
      LAYER met2 ;
        RECT 0.000 3123.605 208.285 3124.445 ;
        RECT 0.000 3121.225 208.565 3123.605 ;
        RECT 0.000 3120.385 208.285 3121.225 ;
        RECT 0.000 3118.465 208.565 3120.385 ;
        RECT 0.000 3117.625 208.285 3118.465 ;
      LAYER met2 ;
        RECT 208.565 3117.905 210.965 3118.185 ;
      LAYER met2 ;
        RECT 0.000 3115.245 208.565 3117.625 ;
        RECT 0.000 3114.405 208.285 3115.245 ;
        RECT 0.000 3112.025 208.565 3114.405 ;
        RECT 0.000 3111.185 208.285 3112.025 ;
        RECT 0.000 3109.265 208.565 3111.185 ;
        RECT 0.000 3108.425 208.285 3109.265 ;
        RECT 0.000 3106.045 208.565 3108.425 ;
        RECT 0.000 3105.205 208.285 3106.045 ;
        RECT 0.000 3102.825 208.565 3105.205 ;
        RECT 0.000 3101.985 208.285 3102.825 ;
        RECT 0.000 3100.065 208.565 3101.985 ;
        RECT 0.000 3099.225 208.285 3100.065 ;
        RECT 0.000 3096.845 208.565 3099.225 ;
      LAYER met2 ;
        RECT 211.300 3097.130 211.440 3136.430 ;
        RECT 209.000 3096.990 211.440 3097.130 ;
      LAYER met2 ;
        RECT 0.000 3096.005 208.285 3096.845 ;
      LAYER met2 ;
        RECT 209.000 3096.565 209.140 3096.990 ;
        RECT 208.565 3096.285 210.965 3096.565 ;
      LAYER met2 ;
        RECT 0.000 3093.625 208.565 3096.005 ;
        RECT 0.000 3092.785 208.285 3093.625 ;
        RECT 0.000 3090.405 208.565 3092.785 ;
      LAYER met2 ;
        RECT 212.220 3092.630 212.360 3305.150 ;
        RECT 212.680 3124.930 212.820 3340.510 ;
        RECT 213.140 3293.570 213.280 3504.050 ;
        RECT 3367.300 3476.510 3367.560 3476.830 ;
        RECT 213.080 3293.250 213.340 3293.570 ;
        RECT 212.620 3124.610 212.880 3124.930 ;
        RECT 208.940 3092.310 209.200 3092.630 ;
        RECT 212.160 3092.310 212.420 3092.630 ;
      LAYER met2 ;
        RECT 0.000 3089.565 208.285 3090.405 ;
      LAYER met2 ;
        RECT 209.000 3090.125 209.140 3092.310 ;
        RECT 208.565 3089.845 210.965 3090.125 ;
      LAYER met2 ;
        RECT 0.000 3087.645 208.565 3089.565 ;
        RECT 0.000 3086.805 208.285 3087.645 ;
        RECT 0.000 3084.425 208.565 3086.805 ;
        RECT 0.000 3083.585 208.285 3084.425 ;
        RECT 0.000 3081.205 208.565 3083.585 ;
        RECT 0.000 3080.365 208.285 3081.205 ;
        RECT 0.000 3078.445 208.565 3080.365 ;
        RECT 0.000 3077.605 208.285 3078.445 ;
        RECT 0.000 3075.225 208.565 3077.605 ;
      LAYER met2 ;
        RECT 208.940 3077.350 209.200 3077.670 ;
      LAYER met2 ;
        RECT 0.000 3074.385 208.285 3075.225 ;
      LAYER met2 ;
        RECT 209.000 3074.945 209.140 3077.350 ;
        RECT 208.565 3074.665 210.965 3074.945 ;
      LAYER met2 ;
        RECT 0.000 3072.005 208.565 3074.385 ;
        RECT 0.000 3071.165 208.285 3072.005 ;
        RECT 0.000 3069.245 208.565 3071.165 ;
        RECT 0.000 3068.405 208.285 3069.245 ;
        RECT 0.000 3066.025 208.565 3068.405 ;
        RECT 0.000 3065.185 208.285 3066.025 ;
        RECT 0.000 3062.805 208.565 3065.185 ;
        RECT 0.000 3061.965 208.285 3062.805 ;
        RECT 0.000 3060.045 208.565 3061.965 ;
        RECT 0.000 3059.205 208.285 3060.045 ;
        RECT 0.000 3058.210 208.565 3059.205 ;
      LAYER met2 ;
        RECT 212.220 3015.530 212.360 3092.310 ;
        RECT 212.680 3016.130 212.820 3124.610 ;
        RECT 213.140 3077.670 213.280 3293.250 ;
        RECT 3367.360 3252.770 3367.500 3476.510 ;
        RECT 3368.280 3461.610 3368.420 3690.370 ;
        RECT 3369.200 3476.830 3369.340 3701.590 ;
        RECT 3370.060 3654.330 3370.320 3654.650 ;
        RECT 3369.140 3476.510 3369.400 3476.830 ;
        RECT 3368.280 3461.530 3369.800 3461.610 ;
        RECT 3368.280 3461.470 3369.860 3461.530 ;
        RECT 3369.600 3461.210 3369.860 3461.470 ;
        RECT 3367.760 3425.850 3368.020 3426.170 ;
        RECT 3367.300 3252.450 3367.560 3252.770 ;
        RECT 3367.360 3236.110 3367.500 3252.450 ;
        RECT 3367.300 3235.790 3367.560 3236.110 ;
        RECT 3367.300 3235.110 3367.560 3235.430 ;
        RECT 213.080 3077.350 213.340 3077.670 ;
        RECT 213.140 3063.670 213.280 3077.350 ;
        RECT 213.140 3063.530 214.200 3063.670 ;
        RECT 212.620 3015.810 212.880 3016.130 ;
        RECT 212.220 3015.390 213.280 3015.530 ;
        RECT 212.620 3014.790 212.880 3015.110 ;
        RECT 212.680 2925.670 212.820 3014.790 ;
        RECT 213.140 2967.070 213.280 3015.390 ;
        RECT 213.140 2966.930 213.740 2967.070 ;
        RECT 212.220 2925.530 212.820 2925.670 ;
      LAYER met2 ;
        RECT 0.000 2920.865 208.565 2921.915 ;
        RECT 0.000 2920.025 208.285 2920.865 ;
      LAYER met2 ;
        RECT 208.565 2920.515 210.965 2920.585 ;
        RECT 208.565 2920.375 211.440 2920.515 ;
        RECT 208.565 2920.305 210.965 2920.375 ;
      LAYER met2 ;
        RECT 0.000 2917.645 208.565 2920.025 ;
        RECT 0.000 2916.805 208.285 2917.645 ;
        RECT 0.000 2914.425 208.565 2916.805 ;
        RECT 0.000 2913.585 208.285 2914.425 ;
      LAYER met2 ;
        RECT 208.565 2913.865 210.965 2914.145 ;
      LAYER met2 ;
        RECT 0.000 2911.665 208.565 2913.585 ;
        RECT 0.000 2910.825 208.285 2911.665 ;
      LAYER met2 ;
        RECT 208.565 2911.105 210.965 2911.385 ;
      LAYER met2 ;
        RECT 0.000 2908.445 208.565 2910.825 ;
      LAYER met2 ;
        RECT 209.000 2908.690 209.140 2911.105 ;
      LAYER met2 ;
        RECT 0.000 2907.605 208.285 2908.445 ;
      LAYER met2 ;
        RECT 208.940 2908.370 209.200 2908.690 ;
      LAYER met2 ;
        RECT 0.000 2905.225 208.565 2907.605 ;
        RECT 0.000 2904.385 208.285 2905.225 ;
        RECT 0.000 2902.465 208.565 2904.385 ;
        RECT 0.000 2901.625 208.285 2902.465 ;
      LAYER met2 ;
        RECT 208.565 2901.905 210.965 2902.185 ;
      LAYER met2 ;
        RECT 0.000 2899.245 208.565 2901.625 ;
        RECT 0.000 2898.405 208.285 2899.245 ;
        RECT 0.000 2896.025 208.565 2898.405 ;
        RECT 0.000 2895.185 208.285 2896.025 ;
        RECT 0.000 2893.265 208.565 2895.185 ;
        RECT 0.000 2892.425 208.285 2893.265 ;
        RECT 0.000 2890.045 208.565 2892.425 ;
        RECT 0.000 2889.205 208.285 2890.045 ;
        RECT 0.000 2886.825 208.565 2889.205 ;
        RECT 0.000 2885.985 208.285 2886.825 ;
        RECT 0.000 2884.065 208.565 2885.985 ;
        RECT 0.000 2883.225 208.285 2884.065 ;
        RECT 0.000 2880.845 208.565 2883.225 ;
      LAYER met2 ;
        RECT 211.300 2880.890 211.440 2920.375 ;
        RECT 212.220 2908.690 212.360 2925.530 ;
        RECT 212.160 2908.370 212.420 2908.690 ;
      LAYER met2 ;
        RECT 0.000 2880.005 208.285 2880.845 ;
      LAYER met2 ;
        RECT 209.000 2880.750 211.440 2880.890 ;
        RECT 209.000 2880.565 209.140 2880.750 ;
        RECT 208.565 2880.285 210.965 2880.565 ;
      LAYER met2 ;
        RECT 0.000 2877.625 208.565 2880.005 ;
        RECT 0.000 2876.785 208.285 2877.625 ;
        RECT 0.000 2874.405 208.565 2876.785 ;
      LAYER met2 ;
        RECT 208.940 2876.070 209.200 2876.390 ;
      LAYER met2 ;
        RECT 0.000 2873.565 208.285 2874.405 ;
      LAYER met2 ;
        RECT 209.000 2874.125 209.140 2876.070 ;
        RECT 208.565 2873.845 210.965 2874.125 ;
      LAYER met2 ;
        RECT 0.000 2871.645 208.565 2873.565 ;
        RECT 0.000 2870.805 208.285 2871.645 ;
        RECT 0.000 2868.425 208.565 2870.805 ;
        RECT 0.000 2867.585 208.285 2868.425 ;
        RECT 0.000 2865.205 208.565 2867.585 ;
        RECT 0.000 2864.365 208.285 2865.205 ;
        RECT 0.000 2862.445 208.565 2864.365 ;
        RECT 0.000 2861.605 208.285 2862.445 ;
        RECT 0.000 2859.225 208.565 2861.605 ;
      LAYER met2 ;
        RECT 208.940 2861.110 209.200 2861.430 ;
      LAYER met2 ;
        RECT 0.000 2858.385 208.285 2859.225 ;
      LAYER met2 ;
        RECT 209.000 2858.945 209.140 2861.110 ;
        RECT 208.565 2858.665 210.965 2858.945 ;
      LAYER met2 ;
        RECT 0.000 2856.005 208.565 2858.385 ;
        RECT 0.000 2855.165 208.285 2856.005 ;
      LAYER met2 ;
        RECT 212.220 2855.990 212.360 2908.370 ;
        RECT 213.600 2876.390 213.740 2966.930 ;
        RECT 213.540 2876.070 213.800 2876.390 ;
        RECT 212.620 2861.110 212.880 2861.430 ;
        RECT 211.240 2855.670 211.500 2855.990 ;
        RECT 212.160 2855.670 212.420 2855.990 ;
      LAYER met2 ;
        RECT 0.000 2853.245 208.565 2855.165 ;
        RECT 0.000 2852.405 208.285 2853.245 ;
        RECT 0.000 2850.025 208.565 2852.405 ;
        RECT 0.000 2849.185 208.285 2850.025 ;
        RECT 0.000 2846.805 208.565 2849.185 ;
        RECT 0.000 2845.965 208.285 2846.805 ;
        RECT 0.000 2844.045 208.565 2845.965 ;
        RECT 0.000 2843.205 208.285 2844.045 ;
        RECT 0.000 2842.210 208.565 2843.205 ;
      LAYER met2 ;
        RECT 211.300 2715.570 211.440 2855.670 ;
        RECT 211.240 2715.250 211.500 2715.570 ;
        RECT 212.160 2715.250 212.420 2715.570 ;
      LAYER met2 ;
        RECT 0.000 2704.865 208.565 2705.915 ;
        RECT 0.000 2704.025 208.285 2704.865 ;
      LAYER met2 ;
        RECT 208.565 2704.515 210.965 2704.585 ;
        RECT 208.565 2704.375 211.440 2704.515 ;
        RECT 208.565 2704.305 210.965 2704.375 ;
      LAYER met2 ;
        RECT 0.000 2701.645 208.565 2704.025 ;
        RECT 0.000 2700.805 208.285 2701.645 ;
        RECT 0.000 2698.425 208.565 2700.805 ;
        RECT 0.000 2697.585 208.285 2698.425 ;
      LAYER met2 ;
        RECT 208.565 2697.865 210.965 2698.145 ;
      LAYER met2 ;
        RECT 0.000 2695.665 208.565 2697.585 ;
      LAYER met2 ;
        RECT 208.940 2697.230 209.200 2697.550 ;
      LAYER met2 ;
        RECT 0.000 2694.825 208.285 2695.665 ;
      LAYER met2 ;
        RECT 209.000 2695.385 209.140 2697.230 ;
        RECT 208.565 2695.105 210.965 2695.385 ;
      LAYER met2 ;
        RECT 0.000 2692.445 208.565 2694.825 ;
        RECT 0.000 2691.605 208.285 2692.445 ;
        RECT 0.000 2689.225 208.565 2691.605 ;
        RECT 0.000 2688.385 208.285 2689.225 ;
        RECT 0.000 2686.465 208.565 2688.385 ;
        RECT 0.000 2685.625 208.285 2686.465 ;
      LAYER met2 ;
        RECT 208.565 2685.905 210.965 2686.185 ;
      LAYER met2 ;
        RECT 0.000 2683.245 208.565 2685.625 ;
        RECT 0.000 2682.405 208.285 2683.245 ;
        RECT 0.000 2680.025 208.565 2682.405 ;
        RECT 0.000 2679.185 208.285 2680.025 ;
        RECT 0.000 2677.265 208.565 2679.185 ;
        RECT 0.000 2676.425 208.285 2677.265 ;
        RECT 0.000 2674.045 208.565 2676.425 ;
        RECT 0.000 2673.205 208.285 2674.045 ;
        RECT 0.000 2670.825 208.565 2673.205 ;
        RECT 0.000 2669.985 208.285 2670.825 ;
        RECT 0.000 2668.065 208.565 2669.985 ;
        RECT 0.000 2667.225 208.285 2668.065 ;
        RECT 0.000 2664.845 208.565 2667.225 ;
      LAYER met2 ;
        RECT 211.300 2665.330 211.440 2704.375 ;
        RECT 212.220 2697.550 212.360 2715.250 ;
        RECT 212.160 2697.230 212.420 2697.550 ;
        RECT 209.000 2665.190 211.440 2665.330 ;
      LAYER met2 ;
        RECT 0.000 2664.005 208.285 2664.845 ;
      LAYER met2 ;
        RECT 209.000 2664.565 209.140 2665.190 ;
        RECT 208.565 2664.285 210.965 2664.565 ;
      LAYER met2 ;
        RECT 0.000 2661.625 208.565 2664.005 ;
        RECT 0.000 2660.785 208.285 2661.625 ;
        RECT 0.000 2658.405 208.565 2660.785 ;
        RECT 0.000 2657.565 208.285 2658.405 ;
      LAYER met2 ;
        RECT 208.565 2657.845 210.965 2658.125 ;
      LAYER met2 ;
        RECT 0.000 2655.645 208.565 2657.565 ;
      LAYER met2 ;
        RECT 209.000 2656.070 209.140 2657.845 ;
        RECT 212.680 2657.170 212.820 2861.110 ;
        RECT 213.600 2773.870 213.740 2876.070 ;
        RECT 214.060 2861.430 214.200 3063.530 ;
        RECT 3367.360 3014.770 3367.500 3235.110 ;
        RECT 3367.820 3203.470 3367.960 3425.850 ;
        RECT 3368.220 3235.790 3368.480 3236.110 ;
        RECT 3367.760 3203.150 3368.020 3203.470 ;
        RECT 3367.300 3014.450 3367.560 3014.770 ;
        RECT 214.000 2861.110 214.260 2861.430 ;
        RECT 3367.360 2789.350 3367.500 3014.450 ;
        RECT 3367.820 2975.330 3367.960 3203.150 ;
        RECT 3368.280 3025.650 3368.420 3235.790 ;
        RECT 3369.660 3235.430 3369.800 3461.210 ;
        RECT 3370.120 3426.170 3370.260 3654.330 ;
        RECT 3370.060 3425.850 3370.320 3426.170 ;
        RECT 3369.600 3235.110 3369.860 3235.430 ;
        RECT 3368.220 3025.330 3368.480 3025.650 ;
        RECT 3367.760 2975.010 3368.020 2975.330 ;
        RECT 3367.300 2789.030 3367.560 2789.350 ;
        RECT 211.760 2657.030 212.820 2657.170 ;
        RECT 213.140 2773.730 213.740 2773.870 ;
        RECT 208.940 2655.750 209.200 2656.070 ;
      LAYER met2 ;
        RECT 0.000 2654.805 208.285 2655.645 ;
        RECT 0.000 2652.425 208.565 2654.805 ;
        RECT 0.000 2651.585 208.285 2652.425 ;
        RECT 0.000 2649.205 208.565 2651.585 ;
        RECT 0.000 2648.365 208.285 2649.205 ;
        RECT 0.000 2646.445 208.565 2648.365 ;
        RECT 0.000 2645.605 208.285 2646.445 ;
        RECT 0.000 2643.225 208.565 2645.605 ;
        RECT 0.000 2642.385 208.285 2643.225 ;
      LAYER met2 ;
        RECT 208.565 2642.665 210.965 2642.945 ;
      LAYER met2 ;
        RECT 0.000 2640.005 208.565 2642.385 ;
      LAYER met2 ;
        RECT 209.000 2640.430 209.140 2642.665 ;
        RECT 211.760 2640.430 211.900 2657.030 ;
        RECT 213.140 2656.490 213.280 2773.730 ;
        RECT 3367.820 2752.630 3367.960 2975.010 ;
        RECT 3368.280 2804.990 3368.420 3025.330 ;
        RECT 3368.220 2804.670 3368.480 2804.990 ;
        RECT 3367.760 2752.310 3368.020 2752.630 ;
        RECT 3367.820 2732.470 3367.960 2752.310 ;
        RECT 3367.360 2732.330 3367.960 2732.470 ;
        RECT 214.000 2697.230 214.260 2697.550 ;
        RECT 212.220 2656.350 213.280 2656.490 ;
        RECT 212.220 2656.070 212.360 2656.350 ;
        RECT 212.160 2655.750 212.420 2656.070 ;
        RECT 208.940 2640.110 209.200 2640.430 ;
        RECT 211.700 2640.110 211.960 2640.430 ;
      LAYER met2 ;
        RECT 0.000 2639.165 208.285 2640.005 ;
        RECT 0.000 2637.245 208.565 2639.165 ;
        RECT 0.000 2636.405 208.285 2637.245 ;
        RECT 0.000 2634.025 208.565 2636.405 ;
        RECT 0.000 2633.185 208.285 2634.025 ;
        RECT 0.000 2630.805 208.565 2633.185 ;
        RECT 0.000 2629.965 208.285 2630.805 ;
        RECT 0.000 2628.045 208.565 2629.965 ;
        RECT 0.000 2627.205 208.285 2628.045 ;
        RECT 0.000 2626.210 208.565 2627.205 ;
        RECT 4.925 2465.390 200.000 2489.290 ;
        RECT 4.925 2439.395 197.965 2465.390 ;
        RECT 198.080 2440.895 200.000 2442.895 ;
        RECT 4.925 2415.495 200.000 2439.395 ;
        RECT 4.925 2415.265 197.965 2415.495 ;
        RECT 0.035 2280.200 151.405 2289.935 ;
        RECT 153.765 2279.000 158.415 2290.140 ;
        RECT 160.165 2280.200 174.575 2289.935 ;
        RECT 0.035 2278.700 197.965 2279.000 ;
        RECT 0.035 2258.095 198.000 2278.700 ;
        RECT 0.035 2257.535 197.965 2258.095 ;
        RECT 0.035 2224.925 198.000 2257.535 ;
        RECT 0.035 2224.495 197.965 2224.925 ;
        RECT 0.035 2204.500 198.000 2224.495 ;
        RECT 0.035 2204.000 197.965 2204.500 ;
        RECT 153.800 2193.025 158.450 2204.000 ;
        RECT 0.000 2066.865 208.565 2067.915 ;
        RECT 0.000 2066.025 208.285 2066.865 ;
      LAYER met2 ;
        RECT 208.565 2066.515 210.965 2066.585 ;
        RECT 208.565 2066.375 211.440 2066.515 ;
        RECT 208.565 2066.305 210.965 2066.375 ;
      LAYER met2 ;
        RECT 0.000 2063.645 208.565 2066.025 ;
        RECT 0.000 2062.805 208.285 2063.645 ;
        RECT 0.000 2060.425 208.565 2062.805 ;
        RECT 0.000 2059.585 208.285 2060.425 ;
      LAYER met2 ;
        RECT 208.565 2059.865 210.965 2060.145 ;
      LAYER met2 ;
        RECT 0.000 2057.665 208.565 2059.585 ;
        RECT 0.000 2056.825 208.285 2057.665 ;
      LAYER met2 ;
        RECT 208.610 2057.385 209.140 2057.410 ;
        RECT 208.565 2057.105 210.965 2057.385 ;
      LAYER met2 ;
        RECT 0.000 2054.445 208.565 2056.825 ;
      LAYER met2 ;
        RECT 209.000 2054.950 209.140 2057.105 ;
        RECT 208.940 2054.630 209.200 2054.950 ;
      LAYER met2 ;
        RECT 0.000 2053.605 208.285 2054.445 ;
        RECT 0.000 2051.225 208.565 2053.605 ;
        RECT 0.000 2050.385 208.285 2051.225 ;
        RECT 0.000 2048.465 208.565 2050.385 ;
        RECT 0.000 2047.625 208.285 2048.465 ;
      LAYER met2 ;
        RECT 208.565 2047.905 210.965 2048.185 ;
      LAYER met2 ;
        RECT 0.000 2045.245 208.565 2047.625 ;
        RECT 0.000 2044.405 208.285 2045.245 ;
        RECT 0.000 2042.025 208.565 2044.405 ;
        RECT 0.000 2041.185 208.285 2042.025 ;
        RECT 0.000 2039.265 208.565 2041.185 ;
        RECT 0.000 2038.425 208.285 2039.265 ;
        RECT 0.000 2036.045 208.565 2038.425 ;
        RECT 0.000 2035.205 208.285 2036.045 ;
        RECT 0.000 2032.825 208.565 2035.205 ;
        RECT 0.000 2031.985 208.285 2032.825 ;
        RECT 0.000 2030.065 208.565 2031.985 ;
        RECT 0.000 2029.225 208.285 2030.065 ;
        RECT 0.000 2026.845 208.565 2029.225 ;
      LAYER met2 ;
        RECT 211.300 2027.490 211.440 2066.375 ;
        RECT 209.000 2027.350 211.440 2027.490 ;
      LAYER met2 ;
        RECT 0.000 2026.005 208.285 2026.845 ;
      LAYER met2 ;
        RECT 209.000 2026.565 209.140 2027.350 ;
        RECT 208.565 2026.285 210.965 2026.565 ;
      LAYER met2 ;
        RECT 0.000 2023.625 208.565 2026.005 ;
        RECT 0.000 2022.785 208.285 2023.625 ;
        RECT 0.000 2020.405 208.565 2022.785 ;
      LAYER met2 ;
        RECT 212.220 2022.650 212.360 2655.750 ;
        RECT 213.540 2640.110 213.800 2640.430 ;
        RECT 212.620 2054.630 212.880 2054.950 ;
        RECT 208.940 2022.330 209.200 2022.650 ;
        RECT 212.160 2022.330 212.420 2022.650 ;
      LAYER met2 ;
        RECT 0.000 2019.565 208.285 2020.405 ;
      LAYER met2 ;
        RECT 209.000 2020.125 209.140 2022.330 ;
        RECT 208.565 2019.845 210.965 2020.125 ;
      LAYER met2 ;
        RECT 0.000 2017.645 208.565 2019.565 ;
        RECT 0.000 2016.805 208.285 2017.645 ;
        RECT 0.000 2014.425 208.565 2016.805 ;
        RECT 0.000 2013.585 208.285 2014.425 ;
        RECT 0.000 2011.205 208.565 2013.585 ;
        RECT 0.000 2010.365 208.285 2011.205 ;
        RECT 0.000 2008.445 208.565 2010.365 ;
        RECT 0.000 2007.605 208.285 2008.445 ;
        RECT 0.000 2005.225 208.565 2007.605 ;
        RECT 0.000 2004.385 208.285 2005.225 ;
      LAYER met2 ;
        RECT 208.565 2004.665 210.965 2004.945 ;
      LAYER met2 ;
        RECT 0.000 2002.005 208.565 2004.385 ;
      LAYER met2 ;
        RECT 209.000 2004.290 209.140 2004.665 ;
        RECT 208.940 2003.970 209.200 2004.290 ;
      LAYER met2 ;
        RECT 0.000 2001.165 208.285 2002.005 ;
        RECT 0.000 1999.245 208.565 2001.165 ;
        RECT 0.000 1998.405 208.285 1999.245 ;
        RECT 0.000 1996.025 208.565 1998.405 ;
        RECT 0.000 1995.185 208.285 1996.025 ;
        RECT 0.000 1992.805 208.565 1995.185 ;
        RECT 0.000 1991.965 208.285 1992.805 ;
        RECT 0.000 1990.045 208.565 1991.965 ;
        RECT 0.000 1989.205 208.285 1990.045 ;
        RECT 0.000 1988.210 208.565 1989.205 ;
        RECT 0.000 1850.865 208.565 1851.915 ;
        RECT 0.000 1850.025 208.285 1850.865 ;
      LAYER met2 ;
        RECT 208.565 1850.305 210.965 1850.585 ;
      LAYER met2 ;
        RECT 0.000 1847.645 208.565 1850.025 ;
      LAYER met2 ;
        RECT 209.000 1847.890 209.140 1850.305 ;
      LAYER met2 ;
        RECT 0.000 1846.805 208.285 1847.645 ;
      LAYER met2 ;
        RECT 208.940 1847.570 209.200 1847.890 ;
        RECT 211.700 1847.570 211.960 1847.890 ;
      LAYER met2 ;
        RECT 0.000 1844.425 208.565 1846.805 ;
        RECT 0.000 1843.585 208.285 1844.425 ;
      LAYER met2 ;
        RECT 208.565 1843.865 210.965 1844.145 ;
      LAYER met2 ;
        RECT 0.000 1841.665 208.565 1843.585 ;
      LAYER met2 ;
        RECT 208.940 1843.150 209.200 1843.470 ;
      LAYER met2 ;
        RECT 0.000 1840.825 208.285 1841.665 ;
      LAYER met2 ;
        RECT 209.000 1841.385 209.140 1843.150 ;
        RECT 208.565 1841.105 210.965 1841.385 ;
      LAYER met2 ;
        RECT 0.000 1838.445 208.565 1840.825 ;
        RECT 0.000 1837.605 208.285 1838.445 ;
        RECT 0.000 1835.225 208.565 1837.605 ;
        RECT 0.000 1834.385 208.285 1835.225 ;
        RECT 0.000 1832.465 208.565 1834.385 ;
        RECT 0.000 1831.625 208.285 1832.465 ;
      LAYER met2 ;
        RECT 208.565 1831.905 210.965 1832.185 ;
      LAYER met2 ;
        RECT 0.000 1829.245 208.565 1831.625 ;
        RECT 0.000 1828.405 208.285 1829.245 ;
        RECT 0.000 1826.025 208.565 1828.405 ;
        RECT 0.000 1825.185 208.285 1826.025 ;
        RECT 0.000 1823.265 208.565 1825.185 ;
        RECT 0.000 1822.425 208.285 1823.265 ;
        RECT 0.000 1820.045 208.565 1822.425 ;
        RECT 0.000 1819.205 208.285 1820.045 ;
        RECT 0.000 1816.825 208.565 1819.205 ;
        RECT 0.000 1815.985 208.285 1816.825 ;
        RECT 0.000 1814.065 208.565 1815.985 ;
        RECT 0.000 1813.225 208.285 1814.065 ;
        RECT 0.000 1810.845 208.565 1813.225 ;
      LAYER met2 ;
        RECT 211.760 1813.210 211.900 1847.570 ;
        RECT 212.680 1843.470 212.820 2054.630 ;
        RECT 213.080 2022.330 213.340 2022.650 ;
        RECT 212.620 1843.150 212.880 1843.470 ;
        RECT 208.940 1812.890 209.200 1813.210 ;
        RECT 211.700 1812.890 211.960 1813.210 ;
      LAYER met2 ;
        RECT 0.000 1810.005 208.285 1810.845 ;
      LAYER met2 ;
        RECT 209.000 1810.570 209.140 1812.890 ;
        RECT 208.610 1810.565 209.140 1810.570 ;
        RECT 208.565 1810.285 210.965 1810.565 ;
      LAYER met2 ;
        RECT 0.000 1807.625 208.565 1810.005 ;
      LAYER met2 ;
        RECT 212.680 1807.870 212.820 1843.150 ;
        RECT 211.760 1807.730 212.820 1807.870 ;
      LAYER met2 ;
        RECT 0.000 1806.785 208.285 1807.625 ;
        RECT 0.000 1804.405 208.565 1806.785 ;
        RECT 0.000 1803.565 208.285 1804.405 ;
      LAYER met2 ;
        RECT 208.565 1803.845 210.965 1804.125 ;
        RECT 209.000 1803.690 209.140 1803.845 ;
      LAYER met2 ;
        RECT 0.000 1801.645 208.565 1803.565 ;
      LAYER met2 ;
        RECT 208.940 1803.370 209.200 1803.690 ;
      LAYER met2 ;
        RECT 0.000 1800.805 208.285 1801.645 ;
        RECT 0.000 1798.425 208.565 1800.805 ;
        RECT 0.000 1797.585 208.285 1798.425 ;
        RECT 0.000 1795.205 208.565 1797.585 ;
        RECT 0.000 1794.365 208.285 1795.205 ;
        RECT 0.000 1792.445 208.565 1794.365 ;
        RECT 0.000 1791.605 208.285 1792.445 ;
        RECT 0.000 1789.225 208.565 1791.605 ;
        RECT 0.000 1788.385 208.285 1789.225 ;
      LAYER met2 ;
        RECT 208.565 1788.665 210.965 1788.945 ;
      LAYER met2 ;
        RECT 0.000 1786.005 208.565 1788.385 ;
      LAYER met2 ;
        RECT 209.000 1786.350 209.140 1788.665 ;
        RECT 208.940 1786.030 209.200 1786.350 ;
      LAYER met2 ;
        RECT 0.000 1785.165 208.285 1786.005 ;
        RECT 0.000 1783.245 208.565 1785.165 ;
        RECT 0.000 1782.405 208.285 1783.245 ;
        RECT 0.000 1780.025 208.565 1782.405 ;
        RECT 0.000 1779.185 208.285 1780.025 ;
        RECT 0.000 1776.805 208.565 1779.185 ;
        RECT 0.000 1775.965 208.285 1776.805 ;
        RECT 0.000 1774.045 208.565 1775.965 ;
        RECT 0.000 1773.205 208.285 1774.045 ;
        RECT 0.000 1772.210 208.565 1773.205 ;
      LAYER met2 ;
        RECT 211.760 1711.270 211.900 1807.730 ;
        RECT 213.140 1803.690 213.280 2022.330 ;
        RECT 213.600 2004.290 213.740 2640.110 ;
        RECT 214.060 2054.950 214.200 2697.230 ;
        RECT 214.000 2054.630 214.260 2054.950 ;
        RECT 213.540 2003.970 213.800 2004.290 ;
        RECT 213.080 1803.370 213.340 1803.690 ;
        RECT 212.620 1786.030 212.880 1786.350 ;
        RECT 211.760 1711.130 212.360 1711.270 ;
      LAYER met2 ;
        RECT 0.000 1634.865 208.565 1635.915 ;
        RECT 0.000 1634.025 208.285 1634.865 ;
      LAYER met2 ;
        RECT 208.565 1634.305 210.965 1634.585 ;
      LAYER met2 ;
        RECT 0.000 1631.645 208.565 1634.025 ;
      LAYER met2 ;
        RECT 209.460 1633.770 209.600 1634.305 ;
        RECT 209.460 1633.630 211.440 1633.770 ;
      LAYER met2 ;
        RECT 0.000 1630.805 208.285 1631.645 ;
        RECT 0.000 1628.425 208.565 1630.805 ;
        RECT 0.000 1627.585 208.285 1628.425 ;
      LAYER met2 ;
        RECT 208.565 1627.865 210.965 1628.145 ;
      LAYER met2 ;
        RECT 0.000 1625.665 208.565 1627.585 ;
      LAYER met2 ;
        RECT 208.940 1627.250 209.200 1627.570 ;
      LAYER met2 ;
        RECT 0.000 1624.825 208.285 1625.665 ;
      LAYER met2 ;
        RECT 209.000 1625.385 209.140 1627.250 ;
        RECT 208.565 1625.105 210.965 1625.385 ;
      LAYER met2 ;
        RECT 0.000 1622.445 208.565 1624.825 ;
        RECT 0.000 1621.605 208.285 1622.445 ;
        RECT 0.000 1619.225 208.565 1621.605 ;
        RECT 0.000 1618.385 208.285 1619.225 ;
        RECT 0.000 1616.465 208.565 1618.385 ;
        RECT 0.000 1615.625 208.285 1616.465 ;
      LAYER met2 ;
        RECT 208.565 1615.905 210.965 1616.185 ;
      LAYER met2 ;
        RECT 0.000 1613.245 208.565 1615.625 ;
        RECT 0.000 1612.405 208.285 1613.245 ;
        RECT 0.000 1610.025 208.565 1612.405 ;
        RECT 0.000 1609.185 208.285 1610.025 ;
        RECT 0.000 1607.265 208.565 1609.185 ;
        RECT 0.000 1606.425 208.285 1607.265 ;
        RECT 0.000 1604.045 208.565 1606.425 ;
        RECT 0.000 1603.205 208.285 1604.045 ;
        RECT 0.000 1600.825 208.565 1603.205 ;
        RECT 0.000 1599.985 208.285 1600.825 ;
        RECT 0.000 1598.065 208.565 1599.985 ;
        RECT 0.000 1597.225 208.285 1598.065 ;
        RECT 0.000 1594.845 208.565 1597.225 ;
        RECT 0.000 1594.005 208.285 1594.845 ;
      LAYER met2 ;
        RECT 208.565 1594.495 210.965 1594.565 ;
        RECT 211.300 1594.495 211.440 1633.630 ;
        RECT 212.220 1627.570 212.360 1711.130 ;
        RECT 212.160 1627.250 212.420 1627.570 ;
        RECT 208.565 1594.355 211.440 1594.495 ;
        RECT 208.565 1594.285 210.965 1594.355 ;
      LAYER met2 ;
        RECT 0.000 1591.625 208.565 1594.005 ;
        RECT 0.000 1590.785 208.285 1591.625 ;
        RECT 0.000 1588.405 208.565 1590.785 ;
        RECT 0.000 1587.565 208.285 1588.405 ;
      LAYER met2 ;
        RECT 208.565 1587.845 210.965 1588.125 ;
      LAYER met2 ;
        RECT 0.000 1585.645 208.565 1587.565 ;
      LAYER met2 ;
        RECT 209.000 1586.090 209.140 1587.845 ;
        RECT 208.940 1585.770 209.200 1586.090 ;
      LAYER met2 ;
        RECT 0.000 1584.805 208.285 1585.645 ;
        RECT 0.000 1582.425 208.565 1584.805 ;
        RECT 0.000 1581.585 208.285 1582.425 ;
        RECT 0.000 1579.205 208.565 1581.585 ;
        RECT 0.000 1578.365 208.285 1579.205 ;
        RECT 0.000 1576.445 208.565 1578.365 ;
        RECT 0.000 1575.605 208.285 1576.445 ;
        RECT 0.000 1573.225 208.565 1575.605 ;
        RECT 0.000 1572.385 208.285 1573.225 ;
      LAYER met2 ;
        RECT 208.565 1572.665 210.965 1572.945 ;
      LAYER met2 ;
        RECT 0.000 1570.005 208.565 1572.385 ;
      LAYER met2 ;
        RECT 209.000 1570.450 209.140 1572.665 ;
        RECT 212.680 1570.450 212.820 1786.030 ;
        RECT 213.140 1586.090 213.280 1803.370 ;
        RECT 213.600 1786.350 213.740 2003.970 ;
        RECT 3367.360 1861.830 3367.500 2732.330 ;
        RECT 3373.800 2139.270 3373.940 4981.690 ;
      LAYER met2 ;
        RECT 3390.335 4813.325 3583.075 4837.735 ;
        RECT 3388.000 4810.105 3389.920 4812.105 ;
        RECT 3390.035 4787.890 3583.075 4813.325 ;
        RECT 3413.940 4763.710 3583.075 4787.890 ;
        RECT 3429.550 4613.000 3434.200 4623.975 ;
        RECT 3390.035 4612.500 3587.965 4613.000 ;
        RECT 3390.000 4592.505 3587.965 4612.500 ;
        RECT 3390.035 4592.075 3587.965 4592.505 ;
        RECT 3390.000 4559.465 3587.965 4592.075 ;
        RECT 3390.035 4558.905 3587.965 4559.465 ;
        RECT 3390.000 4538.300 3587.965 4558.905 ;
        RECT 3390.035 4538.000 3587.965 4538.300 ;
        RECT 3413.425 4527.065 3427.835 4536.800 ;
        RECT 3429.585 4526.860 3434.235 4538.000 ;
        RECT 3436.595 4527.065 3587.965 4536.800 ;
        RECT 3379.435 4390.795 3588.000 4391.790 ;
        RECT 3379.715 4389.955 3588.000 4390.795 ;
        RECT 3379.435 4388.035 3588.000 4389.955 ;
        RECT 3379.715 4387.195 3588.000 4388.035 ;
        RECT 3379.435 4384.815 3588.000 4387.195 ;
        RECT 3379.715 4383.975 3588.000 4384.815 ;
        RECT 3379.435 4381.595 3588.000 4383.975 ;
        RECT 3379.715 4380.755 3588.000 4381.595 ;
        RECT 3379.435 4378.835 3588.000 4380.755 ;
        RECT 3379.715 4377.995 3588.000 4378.835 ;
        RECT 3379.435 4375.615 3588.000 4377.995 ;
      LAYER met2 ;
        RECT 3377.035 4375.195 3379.435 4375.335 ;
        RECT 3377.020 4375.055 3379.435 4375.195 ;
        RECT 3377.020 4372.730 3377.160 4375.055 ;
      LAYER met2 ;
        RECT 3379.715 4374.775 3588.000 4375.615 ;
      LAYER met2 ;
        RECT 3376.960 4372.410 3377.220 4372.730 ;
      LAYER met2 ;
        RECT 3379.435 4372.395 3588.000 4374.775 ;
        RECT 3379.715 4371.555 3588.000 4372.395 ;
        RECT 3379.435 4369.635 3588.000 4371.555 ;
        RECT 3379.715 4368.795 3588.000 4369.635 ;
        RECT 3379.435 4366.415 3588.000 4368.795 ;
        RECT 3379.715 4365.575 3588.000 4366.415 ;
        RECT 3379.435 4363.195 3588.000 4365.575 ;
        RECT 3379.715 4362.355 3588.000 4363.195 ;
      LAYER met2 ;
        RECT 3376.960 4361.870 3377.220 4362.190 ;
        RECT 3377.020 4360.155 3377.160 4361.870 ;
      LAYER met2 ;
        RECT 3379.435 4360.435 3588.000 4362.355 ;
      LAYER met2 ;
        RECT 3377.020 4360.015 3379.435 4360.155 ;
        RECT 3377.035 4359.875 3379.435 4360.015 ;
      LAYER met2 ;
        RECT 3379.715 4359.595 3588.000 4360.435 ;
        RECT 3379.435 4357.215 3588.000 4359.595 ;
        RECT 3379.715 4356.375 3588.000 4357.215 ;
        RECT 3379.435 4353.995 3588.000 4356.375 ;
      LAYER met2 ;
        RECT 3377.035 4353.700 3379.435 4353.715 ;
        RECT 3377.020 4353.435 3379.435 4353.700 ;
        RECT 3377.020 4350.970 3377.160 4353.435 ;
      LAYER met2 ;
        RECT 3379.715 4353.155 3588.000 4353.995 ;
      LAYER met2 ;
        RECT 3376.960 4350.650 3377.220 4350.970 ;
      LAYER met2 ;
        RECT 3379.435 4350.775 3588.000 4353.155 ;
        RECT 3379.715 4349.935 3588.000 4350.775 ;
        RECT 3379.435 4348.015 3588.000 4349.935 ;
        RECT 3379.715 4347.175 3588.000 4348.015 ;
        RECT 3379.435 4344.795 3588.000 4347.175 ;
        RECT 3379.715 4343.955 3588.000 4344.795 ;
        RECT 3379.435 4341.575 3588.000 4343.955 ;
        RECT 3379.715 4340.735 3588.000 4341.575 ;
        RECT 3379.435 4338.815 3588.000 4340.735 ;
        RECT 3379.715 4337.975 3588.000 4338.815 ;
        RECT 3379.435 4335.595 3588.000 4337.975 ;
        RECT 3379.715 4334.755 3588.000 4335.595 ;
        RECT 3379.435 4332.375 3588.000 4334.755 ;
      LAYER met2 ;
        RECT 3377.035 4331.815 3379.435 4332.095 ;
      LAYER met2 ;
        RECT 3379.715 4331.535 3588.000 4332.375 ;
        RECT 3379.435 4329.615 3588.000 4331.535 ;
        RECT 3379.715 4328.775 3588.000 4329.615 ;
        RECT 3379.435 4326.395 3588.000 4328.775 ;
        RECT 3379.715 4325.555 3588.000 4326.395 ;
        RECT 3379.435 4323.175 3588.000 4325.555 ;
      LAYER met2 ;
        RECT 3377.035 4322.755 3379.435 4322.895 ;
        RECT 3377.020 4322.615 3379.435 4322.755 ;
        RECT 3377.020 4321.390 3377.160 4322.615 ;
      LAYER met2 ;
        RECT 3379.715 4322.335 3588.000 4323.175 ;
      LAYER met2 ;
        RECT 3376.960 4321.070 3377.220 4321.390 ;
      LAYER met2 ;
        RECT 3379.435 4320.415 3588.000 4322.335 ;
      LAYER met2 ;
        RECT 3377.035 4319.855 3379.435 4320.135 ;
      LAYER met2 ;
        RECT 3379.715 4319.575 3588.000 4320.415 ;
        RECT 3379.435 4317.195 3588.000 4319.575 ;
        RECT 3379.715 4316.355 3588.000 4317.195 ;
      LAYER met2 ;
        RECT 3376.960 4315.970 3377.220 4316.290 ;
        RECT 3377.020 4313.695 3377.160 4315.970 ;
      LAYER met2 ;
        RECT 3379.435 4313.975 3588.000 4316.355 ;
      LAYER met2 ;
        RECT 3377.020 4313.580 3379.435 4313.695 ;
        RECT 3377.035 4313.415 3379.435 4313.580 ;
      LAYER met2 ;
        RECT 3379.715 4313.135 3588.000 4313.975 ;
        RECT 3379.435 4312.085 3588.000 4313.135 ;
        RECT 3390.035 4166.505 3583.075 4166.735 ;
        RECT 3388.000 4142.605 3583.075 4166.505 ;
        RECT 3388.000 4139.105 3389.920 4141.105 ;
        RECT 3390.035 4116.610 3583.075 4142.605 ;
        RECT 3388.000 4092.710 3583.075 4116.610 ;
      LAYER met2 ;
        RECT 3376.500 4091.570 3376.760 4091.890 ;
        RECT 3387.990 4091.715 3388.270 4092.085 ;
        RECT 3388.000 4091.570 3388.260 4091.715 ;
        RECT 3376.560 3933.070 3376.700 4091.570 ;
      LAYER met2 ;
        RECT 3379.435 3944.795 3588.000 3945.790 ;
        RECT 3379.715 3943.955 3588.000 3944.795 ;
        RECT 3379.435 3942.035 3588.000 3943.955 ;
        RECT 3379.715 3941.195 3588.000 3942.035 ;
        RECT 3379.435 3938.815 3588.000 3941.195 ;
        RECT 3379.715 3937.975 3588.000 3938.815 ;
        RECT 3379.435 3935.595 3588.000 3937.975 ;
        RECT 3379.715 3934.755 3588.000 3935.595 ;
      LAYER met2 ;
        RECT 3375.640 3932.930 3376.700 3933.070 ;
        RECT 3375.640 3644.530 3375.780 3932.930 ;
      LAYER met2 ;
        RECT 3379.435 3932.835 3588.000 3934.755 ;
        RECT 3379.715 3931.995 3588.000 3932.835 ;
        RECT 3379.435 3929.615 3588.000 3931.995 ;
      LAYER met2 ;
        RECT 3377.035 3929.195 3379.435 3929.335 ;
        RECT 3377.020 3929.055 3379.435 3929.195 ;
        RECT 3377.020 3928.690 3377.160 3929.055 ;
      LAYER met2 ;
        RECT 3379.715 3928.775 3588.000 3929.615 ;
      LAYER met2 ;
        RECT 3376.960 3928.370 3377.220 3928.690 ;
      LAYER met2 ;
        RECT 3379.435 3926.395 3588.000 3928.775 ;
        RECT 3379.715 3925.555 3588.000 3926.395 ;
        RECT 3379.435 3923.635 3588.000 3925.555 ;
        RECT 3379.715 3922.795 3588.000 3923.635 ;
        RECT 3379.435 3920.415 3588.000 3922.795 ;
        RECT 3379.715 3919.575 3588.000 3920.415 ;
        RECT 3379.435 3917.195 3588.000 3919.575 ;
        RECT 3379.715 3916.355 3588.000 3917.195 ;
        RECT 3379.435 3914.435 3588.000 3916.355 ;
      LAYER met2 ;
        RECT 3377.035 3914.015 3379.435 3914.155 ;
        RECT 3377.020 3913.875 3379.435 3914.015 ;
        RECT 3377.020 3911.690 3377.160 3913.875 ;
      LAYER met2 ;
        RECT 3379.715 3913.595 3588.000 3914.435 ;
      LAYER met2 ;
        RECT 3376.960 3911.370 3377.220 3911.690 ;
      LAYER met2 ;
        RECT 3379.435 3911.215 3588.000 3913.595 ;
        RECT 3379.715 3910.375 3588.000 3911.215 ;
        RECT 3379.435 3907.995 3588.000 3910.375 ;
      LAYER met2 ;
        RECT 3377.035 3907.620 3379.435 3907.715 ;
        RECT 3377.020 3907.435 3379.435 3907.620 ;
        RECT 3377.020 3905.230 3377.160 3907.435 ;
      LAYER met2 ;
        RECT 3379.715 3907.155 3588.000 3907.995 ;
      LAYER met2 ;
        RECT 3376.040 3904.910 3376.300 3905.230 ;
        RECT 3376.960 3904.910 3377.220 3905.230 ;
        RECT 3376.100 3867.570 3376.240 3904.910 ;
      LAYER met2 ;
        RECT 3379.435 3904.775 3588.000 3907.155 ;
        RECT 3379.715 3903.935 3588.000 3904.775 ;
        RECT 3379.435 3902.015 3588.000 3903.935 ;
        RECT 3379.715 3901.175 3588.000 3902.015 ;
        RECT 3379.435 3898.795 3588.000 3901.175 ;
        RECT 3379.715 3897.955 3588.000 3898.795 ;
        RECT 3379.435 3895.575 3588.000 3897.955 ;
        RECT 3379.715 3894.735 3588.000 3895.575 ;
        RECT 3379.435 3892.815 3588.000 3894.735 ;
        RECT 3379.715 3891.975 3588.000 3892.815 ;
        RECT 3379.435 3889.595 3588.000 3891.975 ;
        RECT 3379.715 3888.755 3588.000 3889.595 ;
        RECT 3379.435 3886.375 3588.000 3888.755 ;
      LAYER met2 ;
        RECT 3377.035 3885.815 3379.435 3886.095 ;
      LAYER met2 ;
        RECT 3379.715 3885.535 3588.000 3886.375 ;
        RECT 3379.435 3883.615 3588.000 3885.535 ;
        RECT 3379.715 3882.775 3588.000 3883.615 ;
        RECT 3379.435 3880.395 3588.000 3882.775 ;
        RECT 3379.715 3879.555 3588.000 3880.395 ;
      LAYER met2 ;
        RECT 3376.960 3879.070 3377.220 3879.390 ;
        RECT 3377.020 3876.895 3377.160 3879.070 ;
      LAYER met2 ;
        RECT 3379.435 3877.175 3588.000 3879.555 ;
      LAYER met2 ;
        RECT 3377.020 3876.755 3379.435 3876.895 ;
        RECT 3377.035 3876.615 3379.435 3876.755 ;
      LAYER met2 ;
        RECT 3379.715 3876.335 3588.000 3877.175 ;
        RECT 3379.435 3874.415 3588.000 3876.335 ;
      LAYER met2 ;
        RECT 3377.035 3873.855 3379.435 3874.135 ;
      LAYER met2 ;
        RECT 3379.715 3873.575 3588.000 3874.415 ;
        RECT 3379.435 3871.195 3588.000 3873.575 ;
        RECT 3379.715 3870.355 3588.000 3871.195 ;
        RECT 3379.435 3867.975 3588.000 3870.355 ;
      LAYER met2 ;
        RECT 3377.035 3867.570 3379.435 3867.695 ;
        RECT 3376.100 3867.430 3379.435 3867.570 ;
        RECT 3377.035 3867.415 3379.435 3867.430 ;
      LAYER met2 ;
        RECT 3379.715 3867.135 3588.000 3867.975 ;
        RECT 3379.435 3866.085 3588.000 3867.135 ;
        RECT 3379.435 3719.795 3588.000 3720.790 ;
        RECT 3379.715 3718.955 3588.000 3719.795 ;
        RECT 3379.435 3717.035 3588.000 3718.955 ;
        RECT 3379.715 3716.195 3588.000 3717.035 ;
        RECT 3379.435 3713.815 3588.000 3716.195 ;
        RECT 3379.715 3712.975 3588.000 3713.815 ;
        RECT 3379.435 3710.595 3588.000 3712.975 ;
        RECT 3379.715 3709.755 3588.000 3710.595 ;
        RECT 3379.435 3707.835 3588.000 3709.755 ;
        RECT 3379.715 3706.995 3588.000 3707.835 ;
        RECT 3379.435 3704.615 3588.000 3706.995 ;
      LAYER met2 ;
        RECT 3377.035 3704.300 3379.435 3704.335 ;
        RECT 3377.020 3704.055 3379.435 3704.300 ;
        RECT 3377.020 3701.910 3377.160 3704.055 ;
      LAYER met2 ;
        RECT 3379.715 3703.775 3588.000 3704.615 ;
      LAYER met2 ;
        RECT 3376.960 3701.590 3377.220 3701.910 ;
      LAYER met2 ;
        RECT 3379.435 3701.395 3588.000 3703.775 ;
        RECT 3379.715 3700.555 3588.000 3701.395 ;
        RECT 3379.435 3698.635 3588.000 3700.555 ;
        RECT 3379.715 3697.795 3588.000 3698.635 ;
        RECT 3379.435 3695.415 3588.000 3697.795 ;
        RECT 3379.715 3694.575 3588.000 3695.415 ;
        RECT 3379.435 3692.195 3588.000 3694.575 ;
        RECT 3379.715 3691.355 3588.000 3692.195 ;
      LAYER met2 ;
        RECT 3376.960 3690.370 3377.220 3690.690 ;
        RECT 3377.020 3689.155 3377.160 3690.370 ;
      LAYER met2 ;
        RECT 3379.435 3689.435 3588.000 3691.355 ;
      LAYER met2 ;
        RECT 3377.020 3689.015 3379.435 3689.155 ;
        RECT 3377.035 3688.875 3379.435 3689.015 ;
      LAYER met2 ;
        RECT 3379.715 3688.595 3588.000 3689.435 ;
        RECT 3379.435 3686.215 3588.000 3688.595 ;
        RECT 3379.715 3685.375 3588.000 3686.215 ;
        RECT 3379.435 3682.995 3588.000 3685.375 ;
      LAYER met2 ;
        RECT 3377.035 3682.610 3379.435 3682.715 ;
        RECT 3376.560 3682.470 3379.435 3682.610 ;
        RECT 3376.560 3645.210 3376.700 3682.470 ;
        RECT 3377.035 3682.435 3379.435 3682.470 ;
      LAYER met2 ;
        RECT 3379.715 3682.155 3588.000 3682.995 ;
        RECT 3379.435 3679.775 3588.000 3682.155 ;
        RECT 3379.715 3678.935 3588.000 3679.775 ;
        RECT 3379.435 3677.015 3588.000 3678.935 ;
        RECT 3379.715 3676.175 3588.000 3677.015 ;
        RECT 3379.435 3673.795 3588.000 3676.175 ;
        RECT 3379.715 3672.955 3588.000 3673.795 ;
        RECT 3379.435 3670.575 3588.000 3672.955 ;
        RECT 3379.715 3669.735 3588.000 3670.575 ;
        RECT 3379.435 3667.815 3588.000 3669.735 ;
        RECT 3379.715 3666.975 3588.000 3667.815 ;
        RECT 3379.435 3664.595 3588.000 3666.975 ;
        RECT 3379.715 3663.755 3588.000 3664.595 ;
        RECT 3379.435 3661.375 3588.000 3663.755 ;
      LAYER met2 ;
        RECT 3377.035 3660.815 3379.435 3661.095 ;
      LAYER met2 ;
        RECT 3379.715 3660.535 3588.000 3661.375 ;
        RECT 3379.435 3658.615 3588.000 3660.535 ;
        RECT 3379.715 3657.775 3588.000 3658.615 ;
        RECT 3379.435 3655.395 3588.000 3657.775 ;
      LAYER met2 ;
        RECT 3376.960 3654.330 3377.220 3654.650 ;
      LAYER met2 ;
        RECT 3379.715 3654.555 3588.000 3655.395 ;
      LAYER met2 ;
        RECT 3377.020 3651.895 3377.160 3654.330 ;
      LAYER met2 ;
        RECT 3379.435 3652.175 3588.000 3654.555 ;
      LAYER met2 ;
        RECT 3377.020 3651.755 3379.435 3651.895 ;
        RECT 3377.035 3651.615 3379.435 3651.755 ;
      LAYER met2 ;
        RECT 3379.715 3651.335 3588.000 3652.175 ;
        RECT 3379.435 3649.415 3588.000 3651.335 ;
      LAYER met2 ;
        RECT 3377.035 3648.855 3379.435 3649.135 ;
      LAYER met2 ;
        RECT 3379.715 3648.575 3588.000 3649.415 ;
        RECT 3379.435 3646.195 3588.000 3648.575 ;
        RECT 3379.715 3645.355 3588.000 3646.195 ;
      LAYER met2 ;
        RECT 3376.560 3645.070 3377.160 3645.210 ;
        RECT 3375.640 3644.390 3376.700 3644.530 ;
        RECT 3376.560 3505.270 3376.700 3644.390 ;
        RECT 3377.020 3642.695 3377.160 3645.070 ;
      LAYER met2 ;
        RECT 3379.435 3642.975 3588.000 3645.355 ;
      LAYER met2 ;
        RECT 3377.020 3642.420 3379.435 3642.695 ;
        RECT 3377.035 3642.415 3379.435 3642.420 ;
      LAYER met2 ;
        RECT 3379.715 3642.135 3588.000 3642.975 ;
        RECT 3379.435 3641.085 3588.000 3642.135 ;
      LAYER met2 ;
        RECT 3375.640 3505.130 3376.700 3505.270 ;
        RECT 3375.640 3408.670 3375.780 3505.130 ;
      LAYER met2 ;
        RECT 3379.435 3494.795 3588.000 3495.790 ;
        RECT 3379.715 3493.955 3588.000 3494.795 ;
        RECT 3379.435 3492.035 3588.000 3493.955 ;
        RECT 3379.715 3491.195 3588.000 3492.035 ;
        RECT 3379.435 3488.815 3588.000 3491.195 ;
        RECT 3379.715 3487.975 3588.000 3488.815 ;
        RECT 3379.435 3485.595 3588.000 3487.975 ;
        RECT 3379.715 3484.755 3588.000 3485.595 ;
        RECT 3379.435 3482.835 3588.000 3484.755 ;
        RECT 3379.715 3481.995 3588.000 3482.835 ;
        RECT 3379.435 3479.615 3588.000 3481.995 ;
      LAYER met2 ;
        RECT 3377.035 3479.220 3379.435 3479.335 ;
        RECT 3377.020 3479.055 3379.435 3479.220 ;
        RECT 3377.020 3476.830 3377.160 3479.055 ;
      LAYER met2 ;
        RECT 3379.715 3478.775 3588.000 3479.615 ;
      LAYER met2 ;
        RECT 3376.960 3476.510 3377.220 3476.830 ;
      LAYER met2 ;
        RECT 3379.435 3476.395 3588.000 3478.775 ;
        RECT 3379.715 3475.555 3588.000 3476.395 ;
        RECT 3379.435 3473.635 3588.000 3475.555 ;
        RECT 3379.715 3472.795 3588.000 3473.635 ;
        RECT 3379.435 3470.415 3588.000 3472.795 ;
        RECT 3379.715 3469.575 3588.000 3470.415 ;
        RECT 3379.435 3467.195 3588.000 3469.575 ;
        RECT 3379.715 3466.355 3588.000 3467.195 ;
        RECT 3379.435 3464.435 3588.000 3466.355 ;
      LAYER met2 ;
        RECT 3377.035 3464.015 3379.435 3464.155 ;
        RECT 3377.020 3463.875 3379.435 3464.015 ;
        RECT 3377.020 3461.530 3377.160 3463.875 ;
      LAYER met2 ;
        RECT 3379.715 3463.595 3588.000 3464.435 ;
      LAYER met2 ;
        RECT 3376.960 3461.210 3377.220 3461.530 ;
      LAYER met2 ;
        RECT 3379.435 3461.215 3588.000 3463.595 ;
        RECT 3379.715 3460.375 3588.000 3461.215 ;
      LAYER met2 ;
        RECT 3376.560 3458.070 3377.160 3458.210 ;
        RECT 3376.560 3417.625 3376.700 3458.070 ;
        RECT 3377.020 3457.715 3377.160 3458.070 ;
      LAYER met2 ;
        RECT 3379.435 3457.995 3588.000 3460.375 ;
      LAYER met2 ;
        RECT 3377.020 3457.460 3379.435 3457.715 ;
        RECT 3377.035 3457.435 3379.435 3457.460 ;
      LAYER met2 ;
        RECT 3379.715 3457.155 3588.000 3457.995 ;
        RECT 3379.435 3454.775 3588.000 3457.155 ;
        RECT 3379.715 3453.935 3588.000 3454.775 ;
        RECT 3379.435 3452.015 3588.000 3453.935 ;
        RECT 3379.715 3451.175 3588.000 3452.015 ;
        RECT 3379.435 3448.795 3588.000 3451.175 ;
        RECT 3379.715 3447.955 3588.000 3448.795 ;
        RECT 3379.435 3445.575 3588.000 3447.955 ;
        RECT 3379.715 3444.735 3588.000 3445.575 ;
        RECT 3379.435 3442.815 3588.000 3444.735 ;
        RECT 3379.715 3441.975 3588.000 3442.815 ;
        RECT 3379.435 3439.595 3588.000 3441.975 ;
        RECT 3379.715 3438.755 3588.000 3439.595 ;
        RECT 3379.435 3436.375 3588.000 3438.755 ;
      LAYER met2 ;
        RECT 3377.035 3435.815 3379.435 3436.095 ;
      LAYER met2 ;
        RECT 3379.715 3435.535 3588.000 3436.375 ;
        RECT 3379.435 3433.615 3588.000 3435.535 ;
        RECT 3379.715 3432.775 3588.000 3433.615 ;
        RECT 3379.435 3430.395 3588.000 3432.775 ;
        RECT 3379.715 3429.555 3588.000 3430.395 ;
        RECT 3379.435 3427.175 3588.000 3429.555 ;
      LAYER met2 ;
        RECT 3377.035 3426.860 3379.435 3426.895 ;
        RECT 3377.020 3426.615 3379.435 3426.860 ;
        RECT 3377.020 3426.170 3377.160 3426.615 ;
      LAYER met2 ;
        RECT 3379.715 3426.335 3588.000 3427.175 ;
      LAYER met2 ;
        RECT 3376.960 3425.850 3377.220 3426.170 ;
      LAYER met2 ;
        RECT 3379.435 3424.415 3588.000 3426.335 ;
      LAYER met2 ;
        RECT 3377.035 3423.855 3379.435 3424.135 ;
      LAYER met2 ;
        RECT 3379.715 3423.575 3588.000 3424.415 ;
        RECT 3379.435 3421.195 3588.000 3423.575 ;
        RECT 3379.715 3420.355 3588.000 3421.195 ;
        RECT 3379.435 3417.975 3588.000 3420.355 ;
      LAYER met2 ;
        RECT 3377.035 3417.625 3379.435 3417.695 ;
        RECT 3376.560 3417.485 3379.435 3417.625 ;
        RECT 3377.035 3417.415 3379.435 3417.485 ;
      LAYER met2 ;
        RECT 3379.715 3417.135 3588.000 3417.975 ;
        RECT 3379.435 3416.085 3588.000 3417.135 ;
      LAYER met2 ;
        RECT 3375.640 3408.530 3376.700 3408.670 ;
        RECT 3376.560 3256.870 3376.700 3408.530 ;
      LAYER met2 ;
        RECT 3379.435 3268.795 3588.000 3269.790 ;
        RECT 3379.715 3267.955 3588.000 3268.795 ;
        RECT 3379.435 3266.035 3588.000 3267.955 ;
        RECT 3379.715 3265.195 3588.000 3266.035 ;
        RECT 3379.435 3262.815 3588.000 3265.195 ;
        RECT 3379.715 3261.975 3588.000 3262.815 ;
        RECT 3379.435 3259.595 3588.000 3261.975 ;
        RECT 3379.715 3258.755 3588.000 3259.595 ;
      LAYER met2 ;
        RECT 3375.640 3256.730 3376.700 3256.870 ;
      LAYER met2 ;
        RECT 3379.435 3256.835 3588.000 3258.755 ;
      LAYER met2 ;
        RECT 3375.640 3160.270 3375.780 3256.730 ;
      LAYER met2 ;
        RECT 3379.715 3255.995 3588.000 3256.835 ;
        RECT 3379.435 3253.615 3588.000 3255.995 ;
      LAYER met2 ;
        RECT 3377.035 3253.195 3379.435 3253.335 ;
        RECT 3377.020 3253.055 3379.435 3253.195 ;
        RECT 3377.020 3252.770 3377.160 3253.055 ;
      LAYER met2 ;
        RECT 3379.715 3252.775 3588.000 3253.615 ;
      LAYER met2 ;
        RECT 3376.960 3252.450 3377.220 3252.770 ;
      LAYER met2 ;
        RECT 3379.435 3250.395 3588.000 3252.775 ;
        RECT 3379.715 3249.555 3588.000 3250.395 ;
        RECT 3379.435 3247.635 3588.000 3249.555 ;
        RECT 3379.715 3246.795 3588.000 3247.635 ;
        RECT 3379.435 3244.415 3588.000 3246.795 ;
        RECT 3379.715 3243.575 3588.000 3244.415 ;
        RECT 3379.435 3241.195 3588.000 3243.575 ;
        RECT 3379.715 3240.355 3588.000 3241.195 ;
        RECT 3379.435 3238.435 3588.000 3240.355 ;
      LAYER met2 ;
        RECT 3377.035 3238.015 3379.435 3238.155 ;
        RECT 3377.020 3237.875 3379.435 3238.015 ;
        RECT 3377.020 3235.430 3377.160 3237.875 ;
      LAYER met2 ;
        RECT 3379.715 3237.595 3588.000 3238.435 ;
      LAYER met2 ;
        RECT 3376.960 3235.110 3377.220 3235.430 ;
      LAYER met2 ;
        RECT 3379.435 3235.215 3588.000 3237.595 ;
        RECT 3379.715 3234.375 3588.000 3235.215 ;
        RECT 3379.435 3231.995 3588.000 3234.375 ;
      LAYER met2 ;
        RECT 3377.035 3231.700 3379.435 3231.715 ;
        RECT 3377.020 3231.435 3379.435 3231.700 ;
        RECT 3377.020 3228.970 3377.160 3231.435 ;
      LAYER met2 ;
        RECT 3379.715 3231.155 3588.000 3231.995 ;
      LAYER met2 ;
        RECT 3376.040 3228.650 3376.300 3228.970 ;
        RECT 3376.960 3228.650 3377.220 3228.970 ;
      LAYER met2 ;
        RECT 3379.435 3228.775 3588.000 3231.155 ;
      LAYER met2 ;
        RECT 3376.100 3191.650 3376.240 3228.650 ;
      LAYER met2 ;
        RECT 3379.715 3227.935 3588.000 3228.775 ;
        RECT 3379.435 3226.015 3588.000 3227.935 ;
        RECT 3379.715 3225.175 3588.000 3226.015 ;
        RECT 3379.435 3222.795 3588.000 3225.175 ;
        RECT 3379.715 3221.955 3588.000 3222.795 ;
        RECT 3379.435 3219.575 3588.000 3221.955 ;
        RECT 3379.715 3218.735 3588.000 3219.575 ;
        RECT 3379.435 3216.815 3588.000 3218.735 ;
        RECT 3379.715 3215.975 3588.000 3216.815 ;
        RECT 3379.435 3213.595 3588.000 3215.975 ;
        RECT 3379.715 3212.755 3588.000 3213.595 ;
        RECT 3379.435 3210.375 3588.000 3212.755 ;
      LAYER met2 ;
        RECT 3377.035 3209.815 3379.435 3210.095 ;
      LAYER met2 ;
        RECT 3379.715 3209.535 3588.000 3210.375 ;
        RECT 3379.435 3207.615 3588.000 3209.535 ;
        RECT 3379.715 3206.775 3588.000 3207.615 ;
        RECT 3379.435 3204.395 3588.000 3206.775 ;
        RECT 3379.715 3203.555 3588.000 3204.395 ;
      LAYER met2 ;
        RECT 3376.960 3203.150 3377.220 3203.470 ;
        RECT 3377.020 3200.895 3377.160 3203.150 ;
      LAYER met2 ;
        RECT 3379.435 3201.175 3588.000 3203.555 ;
      LAYER met2 ;
        RECT 3377.020 3200.755 3379.435 3200.895 ;
        RECT 3377.035 3200.615 3379.435 3200.755 ;
      LAYER met2 ;
        RECT 3379.715 3200.335 3588.000 3201.175 ;
        RECT 3379.435 3198.415 3588.000 3200.335 ;
      LAYER met2 ;
        RECT 3377.035 3197.855 3379.435 3198.135 ;
      LAYER met2 ;
        RECT 3379.715 3197.575 3588.000 3198.415 ;
        RECT 3379.435 3195.195 3588.000 3197.575 ;
        RECT 3379.715 3194.355 3588.000 3195.195 ;
        RECT 3379.435 3191.975 3588.000 3194.355 ;
      LAYER met2 ;
        RECT 3377.035 3191.650 3379.435 3191.695 ;
        RECT 3376.100 3191.510 3379.435 3191.650 ;
        RECT 3377.035 3191.415 3379.435 3191.510 ;
      LAYER met2 ;
        RECT 3379.715 3191.135 3588.000 3191.975 ;
        RECT 3379.435 3190.085 3588.000 3191.135 ;
      LAYER met2 ;
        RECT 3375.640 3160.130 3376.700 3160.270 ;
        RECT 3376.560 3063.670 3376.700 3160.130 ;
        RECT 3375.640 3063.530 3376.700 3063.670 ;
        RECT 3375.640 2968.610 3375.780 3063.530 ;
      LAYER met2 ;
        RECT 3379.435 3043.795 3588.000 3044.790 ;
        RECT 3379.715 3042.955 3588.000 3043.795 ;
        RECT 3379.435 3041.035 3588.000 3042.955 ;
        RECT 3379.715 3040.195 3588.000 3041.035 ;
        RECT 3379.435 3037.815 3588.000 3040.195 ;
        RECT 3379.715 3036.975 3588.000 3037.815 ;
        RECT 3379.435 3034.595 3588.000 3036.975 ;
        RECT 3379.715 3033.755 3588.000 3034.595 ;
        RECT 3379.435 3031.835 3588.000 3033.755 ;
        RECT 3379.715 3030.995 3588.000 3031.835 ;
        RECT 3379.435 3028.615 3588.000 3030.995 ;
      LAYER met2 ;
        RECT 3377.035 3028.195 3379.435 3028.335 ;
        RECT 3377.020 3028.055 3379.435 3028.195 ;
        RECT 3377.020 3025.650 3377.160 3028.055 ;
      LAYER met2 ;
        RECT 3379.715 3027.775 3588.000 3028.615 ;
      LAYER met2 ;
        RECT 3376.960 3025.330 3377.220 3025.650 ;
      LAYER met2 ;
        RECT 3379.435 3025.395 3588.000 3027.775 ;
        RECT 3379.715 3024.555 3588.000 3025.395 ;
        RECT 3379.435 3022.635 3588.000 3024.555 ;
        RECT 3379.715 3021.795 3588.000 3022.635 ;
        RECT 3379.435 3019.415 3588.000 3021.795 ;
        RECT 3379.715 3018.575 3588.000 3019.415 ;
        RECT 3379.435 3016.195 3588.000 3018.575 ;
        RECT 3379.715 3015.355 3588.000 3016.195 ;
      LAYER met2 ;
        RECT 3376.960 3014.450 3377.220 3014.770 ;
        RECT 3377.020 3013.155 3377.160 3014.450 ;
      LAYER met2 ;
        RECT 3379.435 3013.435 3588.000 3015.355 ;
      LAYER met2 ;
        RECT 3377.020 3013.015 3379.435 3013.155 ;
        RECT 3377.035 3012.875 3379.435 3013.015 ;
      LAYER met2 ;
        RECT 3379.715 3012.595 3588.000 3013.435 ;
        RECT 3379.435 3010.215 3588.000 3012.595 ;
        RECT 3379.715 3009.375 3588.000 3010.215 ;
        RECT 3379.435 3006.995 3588.000 3009.375 ;
      LAYER met2 ;
        RECT 3377.035 3006.690 3379.435 3006.715 ;
        RECT 3376.560 3006.550 3379.435 3006.690 ;
        RECT 3376.560 2969.290 3376.700 3006.550 ;
        RECT 3377.035 3006.435 3379.435 3006.550 ;
      LAYER met2 ;
        RECT 3379.715 3006.155 3588.000 3006.995 ;
        RECT 3379.435 3003.775 3588.000 3006.155 ;
        RECT 3379.715 3002.935 3588.000 3003.775 ;
        RECT 3379.435 3001.015 3588.000 3002.935 ;
        RECT 3379.715 3000.175 3588.000 3001.015 ;
        RECT 3379.435 2997.795 3588.000 3000.175 ;
        RECT 3379.715 2996.955 3588.000 2997.795 ;
        RECT 3379.435 2994.575 3588.000 2996.955 ;
        RECT 3379.715 2993.735 3588.000 2994.575 ;
        RECT 3379.435 2991.815 3588.000 2993.735 ;
        RECT 3379.715 2990.975 3588.000 2991.815 ;
        RECT 3379.435 2988.595 3588.000 2990.975 ;
        RECT 3379.715 2987.755 3588.000 2988.595 ;
        RECT 3379.435 2985.375 3588.000 2987.755 ;
      LAYER met2 ;
        RECT 3377.035 2984.815 3379.435 2985.095 ;
      LAYER met2 ;
        RECT 3379.715 2984.535 3588.000 2985.375 ;
        RECT 3379.435 2982.615 3588.000 2984.535 ;
        RECT 3379.715 2981.775 3588.000 2982.615 ;
        RECT 3379.435 2979.395 3588.000 2981.775 ;
        RECT 3379.715 2978.555 3588.000 2979.395 ;
        RECT 3379.435 2976.175 3588.000 2978.555 ;
      LAYER met2 ;
        RECT 3377.035 2975.755 3379.435 2975.895 ;
        RECT 3377.020 2975.615 3379.435 2975.755 ;
        RECT 3377.020 2975.330 3377.160 2975.615 ;
      LAYER met2 ;
        RECT 3379.715 2975.335 3588.000 2976.175 ;
      LAYER met2 ;
        RECT 3376.960 2975.010 3377.220 2975.330 ;
      LAYER met2 ;
        RECT 3379.435 2973.415 3588.000 2975.335 ;
      LAYER met2 ;
        RECT 3377.035 2972.855 3379.435 2973.135 ;
      LAYER met2 ;
        RECT 3379.715 2972.575 3588.000 2973.415 ;
        RECT 3379.435 2970.195 3588.000 2972.575 ;
        RECT 3379.715 2969.355 3588.000 2970.195 ;
      LAYER met2 ;
        RECT 3376.560 2969.150 3377.160 2969.290 ;
        RECT 3375.640 2968.470 3376.700 2968.610 ;
        RECT 3376.560 2870.470 3376.700 2968.470 ;
        RECT 3377.020 2966.695 3377.160 2969.150 ;
      LAYER met2 ;
        RECT 3379.435 2966.975 3588.000 2969.355 ;
      LAYER met2 ;
        RECT 3377.020 2966.500 3379.435 2966.695 ;
        RECT 3377.035 2966.415 3379.435 2966.500 ;
      LAYER met2 ;
        RECT 3379.715 2966.135 3588.000 2966.975 ;
        RECT 3379.435 2965.085 3588.000 2966.135 ;
      LAYER met2 ;
        RECT 3375.640 2870.330 3376.700 2870.470 ;
        RECT 3375.640 2732.470 3375.780 2870.330 ;
      LAYER met2 ;
        RECT 3379.435 2817.795 3588.000 2818.790 ;
        RECT 3379.715 2816.955 3588.000 2817.795 ;
        RECT 3379.435 2815.035 3588.000 2816.955 ;
        RECT 3379.715 2814.195 3588.000 2815.035 ;
        RECT 3379.435 2811.815 3588.000 2814.195 ;
        RECT 3379.715 2810.975 3588.000 2811.815 ;
        RECT 3379.435 2808.595 3588.000 2810.975 ;
        RECT 3379.715 2807.755 3588.000 2808.595 ;
        RECT 3379.435 2805.835 3588.000 2807.755 ;
        RECT 3379.715 2804.995 3588.000 2805.835 ;
      LAYER met2 ;
        RECT 3376.960 2804.670 3377.220 2804.990 ;
        RECT 3377.020 2802.335 3377.160 2804.670 ;
      LAYER met2 ;
        RECT 3379.435 2802.615 3588.000 2804.995 ;
      LAYER met2 ;
        RECT 3377.020 2802.195 3379.435 2802.335 ;
        RECT 3377.035 2802.055 3379.435 2802.195 ;
      LAYER met2 ;
        RECT 3379.715 2801.775 3588.000 2802.615 ;
        RECT 3379.435 2799.395 3588.000 2801.775 ;
        RECT 3379.715 2798.555 3588.000 2799.395 ;
        RECT 3379.435 2796.635 3588.000 2798.555 ;
        RECT 3379.715 2795.795 3588.000 2796.635 ;
        RECT 3379.435 2793.415 3588.000 2795.795 ;
        RECT 3379.715 2792.575 3588.000 2793.415 ;
        RECT 3379.435 2790.195 3588.000 2792.575 ;
        RECT 3379.715 2789.355 3588.000 2790.195 ;
      LAYER met2 ;
        RECT 3376.960 2789.030 3377.220 2789.350 ;
        RECT 3377.020 2787.155 3377.160 2789.030 ;
      LAYER met2 ;
        RECT 3379.435 2787.435 3588.000 2789.355 ;
      LAYER met2 ;
        RECT 3377.020 2786.980 3379.435 2787.155 ;
        RECT 3377.035 2786.875 3379.435 2786.980 ;
      LAYER met2 ;
        RECT 3379.715 2786.595 3588.000 2787.435 ;
        RECT 3379.435 2784.215 3588.000 2786.595 ;
        RECT 3379.715 2783.375 3588.000 2784.215 ;
        RECT 3379.435 2780.995 3588.000 2783.375 ;
      LAYER met2 ;
        RECT 3377.035 2780.575 3379.435 2780.715 ;
        RECT 3377.020 2780.435 3379.435 2780.575 ;
        RECT 3377.020 2778.130 3377.160 2780.435 ;
      LAYER met2 ;
        RECT 3379.715 2780.155 3588.000 2780.995 ;
      LAYER met2 ;
        RECT 3376.040 2777.810 3376.300 2778.130 ;
        RECT 3376.960 2777.810 3377.220 2778.130 ;
        RECT 3376.100 2740.625 3376.240 2777.810 ;
      LAYER met2 ;
        RECT 3379.435 2777.775 3588.000 2780.155 ;
        RECT 3379.715 2776.935 3588.000 2777.775 ;
        RECT 3379.435 2775.015 3588.000 2776.935 ;
        RECT 3379.715 2774.175 3588.000 2775.015 ;
        RECT 3379.435 2771.795 3588.000 2774.175 ;
        RECT 3379.715 2770.955 3588.000 2771.795 ;
        RECT 3379.435 2768.575 3588.000 2770.955 ;
        RECT 3379.715 2767.735 3588.000 2768.575 ;
        RECT 3379.435 2765.815 3588.000 2767.735 ;
        RECT 3379.715 2764.975 3588.000 2765.815 ;
        RECT 3379.435 2762.595 3588.000 2764.975 ;
        RECT 3379.715 2761.755 3588.000 2762.595 ;
        RECT 3379.435 2759.375 3588.000 2761.755 ;
      LAYER met2 ;
        RECT 3377.035 2758.815 3379.435 2759.095 ;
      LAYER met2 ;
        RECT 3379.715 2758.535 3588.000 2759.375 ;
        RECT 3379.435 2756.615 3588.000 2758.535 ;
        RECT 3379.715 2755.775 3588.000 2756.615 ;
        RECT 3379.435 2753.395 3588.000 2755.775 ;
      LAYER met2 ;
        RECT 3376.960 2752.310 3377.220 2752.630 ;
      LAYER met2 ;
        RECT 3379.715 2752.555 3588.000 2753.395 ;
      LAYER met2 ;
        RECT 3377.020 2749.895 3377.160 2752.310 ;
      LAYER met2 ;
        RECT 3379.435 2750.175 3588.000 2752.555 ;
      LAYER met2 ;
        RECT 3377.020 2749.755 3379.435 2749.895 ;
        RECT 3377.035 2749.615 3379.435 2749.755 ;
      LAYER met2 ;
        RECT 3379.715 2749.335 3588.000 2750.175 ;
        RECT 3379.435 2747.415 3588.000 2749.335 ;
      LAYER met2 ;
        RECT 3377.035 2746.855 3379.435 2747.135 ;
      LAYER met2 ;
        RECT 3379.715 2746.575 3588.000 2747.415 ;
        RECT 3379.435 2744.195 3588.000 2746.575 ;
        RECT 3379.715 2743.355 3588.000 2744.195 ;
        RECT 3379.435 2740.975 3588.000 2743.355 ;
      LAYER met2 ;
        RECT 3377.035 2740.625 3379.435 2740.695 ;
        RECT 3376.100 2740.485 3379.435 2740.625 ;
        RECT 3377.035 2740.415 3379.435 2740.485 ;
      LAYER met2 ;
        RECT 3379.715 2740.135 3588.000 2740.975 ;
        RECT 3379.435 2739.085 3588.000 2740.135 ;
      LAYER met2 ;
        RECT 3375.640 2732.330 3376.700 2732.470 ;
        RECT 3376.560 2569.030 3376.700 2732.330 ;
      LAYER met2 ;
        RECT 3390.035 2593.505 3583.075 2593.735 ;
        RECT 3388.000 2569.605 3583.075 2593.505 ;
      LAYER met2 ;
        RECT 3376.500 2568.710 3376.760 2569.030 ;
        RECT 3388.460 2568.885 3388.720 2569.030 ;
        RECT 3388.450 2568.515 3388.730 2568.885 ;
      LAYER met2 ;
        RECT 3388.000 2566.105 3389.920 2568.105 ;
        RECT 3390.035 2543.610 3583.075 2569.605 ;
        RECT 3388.000 2519.710 3583.075 2543.610 ;
        RECT 3429.550 2374.000 3434.200 2384.975 ;
        RECT 3390.035 2373.500 3587.965 2374.000 ;
        RECT 3390.000 2353.505 3587.965 2373.500 ;
        RECT 3390.035 2353.075 3587.965 2353.505 ;
        RECT 3390.000 2320.465 3587.965 2353.075 ;
        RECT 3390.035 2319.905 3587.965 2320.465 ;
        RECT 3390.000 2299.300 3587.965 2319.905 ;
        RECT 3390.035 2299.000 3587.965 2299.300 ;
        RECT 3413.425 2288.065 3427.835 2297.800 ;
        RECT 3429.585 2287.860 3434.235 2299.000 ;
        RECT 3436.595 2288.065 3587.965 2297.800 ;
        RECT 3390.035 2152.505 3583.075 2152.735 ;
      LAYER met2 ;
        RECT 3373.740 2138.950 3374.000 2139.270 ;
        RECT 3387.540 2138.950 3387.800 2139.270 ;
        RECT 3387.600 2128.245 3387.740 2138.950 ;
      LAYER met2 ;
        RECT 3388.000 2128.605 3583.075 2152.505 ;
      LAYER met2 ;
        RECT 3387.530 2127.875 3387.810 2128.245 ;
      LAYER met2 ;
        RECT 3388.000 2125.105 3389.920 2127.105 ;
        RECT 3390.035 2102.610 3583.075 2128.605 ;
        RECT 3388.000 2078.710 3583.075 2102.610 ;
        RECT 3379.435 1931.795 3588.000 1932.790 ;
        RECT 3379.715 1930.955 3588.000 1931.795 ;
        RECT 3379.435 1929.035 3588.000 1930.955 ;
        RECT 3379.715 1928.195 3588.000 1929.035 ;
        RECT 3379.435 1925.815 3588.000 1928.195 ;
        RECT 3379.715 1924.975 3588.000 1925.815 ;
        RECT 3379.435 1922.595 3588.000 1924.975 ;
        RECT 3379.715 1921.755 3588.000 1922.595 ;
        RECT 3379.435 1919.835 3588.000 1921.755 ;
        RECT 3379.715 1918.995 3588.000 1919.835 ;
        RECT 3379.435 1916.615 3588.000 1918.995 ;
      LAYER met2 ;
        RECT 3377.035 1916.195 3379.435 1916.335 ;
        RECT 3377.020 1916.055 3379.435 1916.195 ;
        RECT 3377.020 1913.850 3377.160 1916.055 ;
      LAYER met2 ;
        RECT 3379.715 1915.775 3588.000 1916.615 ;
      LAYER met2 ;
        RECT 3367.760 1913.530 3368.020 1913.850 ;
        RECT 3376.960 1913.530 3377.220 1913.850 ;
        RECT 3367.300 1861.510 3367.560 1861.830 ;
        RECT 213.540 1786.030 213.800 1786.350 ;
        RECT 3367.820 1687.750 3367.960 1913.530 ;
      LAYER met2 ;
        RECT 3379.435 1913.395 3588.000 1915.775 ;
        RECT 3379.715 1912.555 3588.000 1913.395 ;
        RECT 3379.435 1910.635 3588.000 1912.555 ;
        RECT 3379.715 1909.795 3588.000 1910.635 ;
        RECT 3379.435 1907.415 3588.000 1909.795 ;
        RECT 3379.715 1906.575 3588.000 1907.415 ;
        RECT 3379.435 1904.195 3588.000 1906.575 ;
        RECT 3379.715 1903.355 3588.000 1904.195 ;
        RECT 3379.435 1901.435 3588.000 1903.355 ;
      LAYER met2 ;
        RECT 3377.035 1900.940 3379.435 1901.155 ;
        RECT 3377.020 1900.875 3379.435 1900.940 ;
        RECT 3377.020 1898.550 3377.160 1900.875 ;
      LAYER met2 ;
        RECT 3379.715 1900.595 3588.000 1901.435 ;
      LAYER met2 ;
        RECT 3368.680 1898.230 3368.940 1898.550 ;
        RECT 3376.960 1898.230 3377.220 1898.550 ;
        RECT 3367.760 1687.430 3368.020 1687.750 ;
        RECT 214.000 1627.250 214.260 1627.570 ;
        RECT 213.080 1585.770 213.340 1586.090 ;
        RECT 208.940 1570.130 209.200 1570.450 ;
        RECT 212.620 1570.130 212.880 1570.450 ;
      LAYER met2 ;
        RECT 0.000 1569.165 208.285 1570.005 ;
        RECT 0.000 1567.245 208.565 1569.165 ;
        RECT 0.000 1566.405 208.285 1567.245 ;
        RECT 0.000 1564.025 208.565 1566.405 ;
        RECT 0.000 1563.185 208.285 1564.025 ;
        RECT 0.000 1560.805 208.565 1563.185 ;
        RECT 0.000 1559.965 208.285 1560.805 ;
        RECT 0.000 1558.045 208.565 1559.965 ;
        RECT 0.000 1557.205 208.285 1558.045 ;
        RECT 0.000 1556.210 208.565 1557.205 ;
        RECT 0.000 1418.865 208.565 1419.915 ;
        RECT 0.000 1418.025 208.285 1418.865 ;
      LAYER met2 ;
        RECT 208.565 1418.515 210.965 1418.585 ;
        RECT 208.565 1418.375 211.440 1418.515 ;
        RECT 208.565 1418.305 210.965 1418.375 ;
      LAYER met2 ;
        RECT 0.000 1415.645 208.565 1418.025 ;
        RECT 0.000 1414.805 208.285 1415.645 ;
        RECT 0.000 1412.425 208.565 1414.805 ;
        RECT 0.000 1411.585 208.285 1412.425 ;
      LAYER met2 ;
        RECT 208.565 1411.865 210.965 1412.145 ;
      LAYER met2 ;
        RECT 0.000 1409.665 208.565 1411.585 ;
        RECT 0.000 1408.825 208.285 1409.665 ;
      LAYER met2 ;
        RECT 208.565 1409.105 210.965 1409.385 ;
      LAYER met2 ;
        RECT 0.000 1406.445 208.565 1408.825 ;
      LAYER met2 ;
        RECT 209.000 1406.910 209.140 1409.105 ;
        RECT 208.940 1406.590 209.200 1406.910 ;
      LAYER met2 ;
        RECT 0.000 1405.605 208.285 1406.445 ;
        RECT 0.000 1403.225 208.565 1405.605 ;
        RECT 0.000 1402.385 208.285 1403.225 ;
        RECT 0.000 1400.465 208.565 1402.385 ;
        RECT 0.000 1399.625 208.285 1400.465 ;
      LAYER met2 ;
        RECT 208.565 1399.905 210.965 1400.185 ;
      LAYER met2 ;
        RECT 0.000 1397.245 208.565 1399.625 ;
        RECT 0.000 1396.405 208.285 1397.245 ;
        RECT 0.000 1394.025 208.565 1396.405 ;
        RECT 0.000 1393.185 208.285 1394.025 ;
        RECT 0.000 1391.265 208.565 1393.185 ;
        RECT 0.000 1390.425 208.285 1391.265 ;
        RECT 0.000 1388.045 208.565 1390.425 ;
        RECT 0.000 1387.205 208.285 1388.045 ;
        RECT 0.000 1384.825 208.565 1387.205 ;
        RECT 0.000 1383.985 208.285 1384.825 ;
        RECT 0.000 1382.065 208.565 1383.985 ;
        RECT 0.000 1381.225 208.285 1382.065 ;
        RECT 0.000 1378.845 208.565 1381.225 ;
        RECT 0.000 1378.005 208.285 1378.845 ;
      LAYER met2 ;
        RECT 208.565 1378.495 210.965 1378.565 ;
        RECT 211.300 1378.495 211.440 1418.375 ;
        RECT 212.160 1406.590 212.420 1406.910 ;
        RECT 208.565 1378.355 211.440 1378.495 ;
        RECT 208.565 1378.285 210.965 1378.355 ;
      LAYER met2 ;
        RECT 0.000 1375.625 208.565 1378.005 ;
        RECT 0.000 1374.785 208.285 1375.625 ;
        RECT 0.000 1372.405 208.565 1374.785 ;
      LAYER met2 ;
        RECT 208.940 1372.590 209.200 1372.910 ;
      LAYER met2 ;
        RECT 0.000 1371.565 208.285 1372.405 ;
      LAYER met2 ;
        RECT 209.000 1372.125 209.140 1372.590 ;
        RECT 208.565 1371.845 210.965 1372.125 ;
        RECT 208.610 1371.830 209.140 1371.845 ;
      LAYER met2 ;
        RECT 0.000 1369.645 208.565 1371.565 ;
        RECT 0.000 1368.805 208.285 1369.645 ;
        RECT 0.000 1366.425 208.565 1368.805 ;
        RECT 0.000 1365.585 208.285 1366.425 ;
        RECT 0.000 1363.205 208.565 1365.585 ;
        RECT 0.000 1362.365 208.285 1363.205 ;
        RECT 0.000 1360.445 208.565 1362.365 ;
        RECT 0.000 1359.605 208.285 1360.445 ;
        RECT 0.000 1357.225 208.565 1359.605 ;
      LAYER met2 ;
        RECT 208.940 1359.330 209.200 1359.650 ;
      LAYER met2 ;
        RECT 0.000 1356.385 208.285 1357.225 ;
      LAYER met2 ;
        RECT 209.000 1357.010 209.140 1359.330 ;
        RECT 208.610 1356.945 209.140 1357.010 ;
        RECT 208.565 1356.665 210.965 1356.945 ;
      LAYER met2 ;
        RECT 0.000 1354.005 208.565 1356.385 ;
        RECT 0.000 1353.165 208.285 1354.005 ;
        RECT 0.000 1351.245 208.565 1353.165 ;
        RECT 0.000 1350.405 208.285 1351.245 ;
        RECT 0.000 1348.025 208.565 1350.405 ;
        RECT 0.000 1347.185 208.285 1348.025 ;
        RECT 0.000 1344.805 208.565 1347.185 ;
        RECT 0.000 1343.965 208.285 1344.805 ;
        RECT 0.000 1342.045 208.565 1343.965 ;
        RECT 0.000 1341.205 208.285 1342.045 ;
        RECT 0.000 1340.210 208.565 1341.205 ;
        RECT 0.000 1202.865 208.565 1203.915 ;
        RECT 0.000 1202.025 208.285 1202.865 ;
      LAYER met2 ;
        RECT 208.610 1202.585 211.440 1202.650 ;
        RECT 208.565 1202.510 211.440 1202.585 ;
        RECT 208.565 1202.305 210.965 1202.510 ;
      LAYER met2 ;
        RECT 0.000 1199.645 208.565 1202.025 ;
        RECT 0.000 1198.805 208.285 1199.645 ;
        RECT 0.000 1196.425 208.565 1198.805 ;
        RECT 0.000 1195.585 208.285 1196.425 ;
      LAYER met2 ;
        RECT 208.565 1195.865 210.965 1196.145 ;
      LAYER met2 ;
        RECT 0.000 1193.665 208.565 1195.585 ;
        RECT 0.000 1192.825 208.285 1193.665 ;
      LAYER met2 ;
        RECT 208.565 1193.105 210.965 1193.385 ;
      LAYER met2 ;
        RECT 0.000 1190.445 208.565 1192.825 ;
      LAYER met2 ;
        RECT 209.000 1190.670 209.140 1193.105 ;
      LAYER met2 ;
        RECT 0.000 1189.605 208.285 1190.445 ;
      LAYER met2 ;
        RECT 208.940 1190.350 209.200 1190.670 ;
      LAYER met2 ;
        RECT 0.000 1187.225 208.565 1189.605 ;
        RECT 0.000 1186.385 208.285 1187.225 ;
      LAYER met2 ;
        RECT 208.565 1186.665 210.965 1186.945 ;
      LAYER met2 ;
        RECT 0.000 1184.465 208.565 1186.385 ;
        RECT 0.000 1183.625 208.285 1184.465 ;
      LAYER met2 ;
        RECT 208.565 1183.905 210.965 1184.185 ;
      LAYER met2 ;
        RECT 0.000 1181.245 208.565 1183.625 ;
        RECT 0.000 1180.405 208.285 1181.245 ;
        RECT 0.000 1178.025 208.565 1180.405 ;
        RECT 0.000 1177.185 208.285 1178.025 ;
      LAYER met2 ;
        RECT 208.565 1177.465 210.965 1177.745 ;
      LAYER met2 ;
        RECT 0.000 1175.265 208.565 1177.185 ;
        RECT 0.000 1174.425 208.285 1175.265 ;
        RECT 0.000 1172.045 208.565 1174.425 ;
        RECT 0.000 1171.205 208.285 1172.045 ;
        RECT 0.000 1168.825 208.565 1171.205 ;
        RECT 0.000 1167.985 208.285 1168.825 ;
        RECT 0.000 1166.065 208.565 1167.985 ;
        RECT 0.000 1165.225 208.285 1166.065 ;
        RECT 0.000 1162.845 208.565 1165.225 ;
      LAYER met2 ;
        RECT 211.300 1163.210 211.440 1202.510 ;
        RECT 212.220 1190.670 212.360 1406.590 ;
        RECT 213.140 1372.910 213.280 1585.770 ;
        RECT 213.540 1570.130 213.800 1570.450 ;
        RECT 213.080 1372.650 213.340 1372.910 ;
        RECT 212.680 1372.590 213.340 1372.650 ;
        RECT 212.680 1372.510 213.280 1372.590 ;
        RECT 212.160 1190.350 212.420 1190.670 ;
        RECT 209.000 1163.070 211.440 1163.210 ;
      LAYER met2 ;
        RECT 0.000 1162.005 208.285 1162.845 ;
      LAYER met2 ;
        RECT 209.000 1162.565 209.140 1163.070 ;
        RECT 208.565 1162.285 210.965 1162.565 ;
      LAYER met2 ;
        RECT 0.000 1159.625 208.565 1162.005 ;
        RECT 0.000 1158.785 208.285 1159.625 ;
        RECT 0.000 1156.405 208.565 1158.785 ;
      LAYER met2 ;
        RECT 208.940 1158.390 209.200 1158.710 ;
      LAYER met2 ;
        RECT 0.000 1155.565 208.285 1156.405 ;
      LAYER met2 ;
        RECT 209.000 1156.125 209.140 1158.390 ;
        RECT 208.565 1155.845 210.965 1156.125 ;
      LAYER met2 ;
        RECT 0.000 1153.645 208.565 1155.565 ;
        RECT 0.000 1152.805 208.285 1153.645 ;
        RECT 0.000 1150.425 208.565 1152.805 ;
        RECT 0.000 1149.585 208.285 1150.425 ;
        RECT 0.000 1147.205 208.565 1149.585 ;
        RECT 0.000 1146.365 208.285 1147.205 ;
        RECT 0.000 1144.445 208.565 1146.365 ;
        RECT 0.000 1143.605 208.285 1144.445 ;
        RECT 0.000 1141.225 208.565 1143.605 ;
      LAYER met2 ;
        RECT 208.940 1143.090 209.200 1143.410 ;
      LAYER met2 ;
        RECT 0.000 1140.385 208.285 1141.225 ;
      LAYER met2 ;
        RECT 209.000 1140.945 209.140 1143.090 ;
        RECT 208.565 1140.665 210.965 1140.945 ;
        RECT 208.610 1140.630 209.140 1140.665 ;
      LAYER met2 ;
        RECT 0.000 1138.005 208.565 1140.385 ;
        RECT 0.000 1137.165 208.285 1138.005 ;
      LAYER met2 ;
        RECT 211.240 1137.310 211.500 1137.630 ;
      LAYER met2 ;
        RECT 0.000 1135.245 208.565 1137.165 ;
        RECT 0.000 1134.405 208.285 1135.245 ;
        RECT 0.000 1132.025 208.565 1134.405 ;
        RECT 0.000 1131.185 208.285 1132.025 ;
        RECT 0.000 1128.805 208.565 1131.185 ;
        RECT 0.000 1127.965 208.285 1128.805 ;
        RECT 0.000 1126.045 208.565 1127.965 ;
        RECT 0.000 1125.205 208.285 1126.045 ;
        RECT 0.000 1124.210 208.565 1125.205 ;
        RECT 0.000 986.865 208.565 987.915 ;
      LAYER met2 ;
        RECT 211.300 987.090 211.440 1137.310 ;
        RECT 212.220 1131.670 212.360 1190.350 ;
        RECT 212.680 1158.710 212.820 1372.510 ;
        RECT 213.600 1359.650 213.740 1570.130 ;
        RECT 214.060 1406.910 214.200 1627.250 ;
        RECT 3367.820 1476.670 3367.960 1687.430 ;
        RECT 3368.740 1672.450 3368.880 1898.230 ;
      LAYER met2 ;
        RECT 3379.435 1898.215 3588.000 1900.595 ;
        RECT 3379.715 1897.375 3588.000 1898.215 ;
        RECT 3379.435 1894.995 3588.000 1897.375 ;
      LAYER met2 ;
        RECT 3377.035 1894.645 3379.435 1894.715 ;
        RECT 3376.560 1894.505 3379.435 1894.645 ;
        RECT 3369.600 1861.510 3369.860 1861.830 ;
        RECT 3368.680 1672.130 3368.940 1672.450 ;
        RECT 3369.660 1640.490 3369.800 1861.510 ;
        RECT 3376.560 1854.625 3376.700 1894.505 ;
        RECT 3377.035 1894.435 3379.435 1894.505 ;
      LAYER met2 ;
        RECT 3379.715 1894.155 3588.000 1894.995 ;
        RECT 3379.435 1891.775 3588.000 1894.155 ;
        RECT 3379.715 1890.935 3588.000 1891.775 ;
        RECT 3379.435 1889.015 3588.000 1890.935 ;
        RECT 3379.715 1888.175 3588.000 1889.015 ;
        RECT 3379.435 1885.795 3588.000 1888.175 ;
        RECT 3379.715 1884.955 3588.000 1885.795 ;
        RECT 3379.435 1882.575 3588.000 1884.955 ;
        RECT 3379.715 1881.735 3588.000 1882.575 ;
        RECT 3379.435 1879.815 3588.000 1881.735 ;
      LAYER met2 ;
        RECT 3377.035 1879.255 3379.435 1879.535 ;
      LAYER met2 ;
        RECT 3379.715 1878.975 3588.000 1879.815 ;
        RECT 3379.435 1876.595 3588.000 1878.975 ;
        RECT 3379.715 1875.755 3588.000 1876.595 ;
        RECT 3379.435 1873.375 3588.000 1875.755 ;
      LAYER met2 ;
        RECT 3377.035 1872.815 3379.435 1873.095 ;
      LAYER met2 ;
        RECT 3379.715 1872.535 3588.000 1873.375 ;
        RECT 3379.435 1870.615 3588.000 1872.535 ;
      LAYER met2 ;
        RECT 3377.035 1870.055 3379.435 1870.335 ;
      LAYER met2 ;
        RECT 3379.715 1869.775 3588.000 1870.615 ;
        RECT 3379.435 1867.395 3588.000 1869.775 ;
        RECT 3379.715 1866.555 3588.000 1867.395 ;
        RECT 3379.435 1864.175 3588.000 1866.555 ;
      LAYER met2 ;
        RECT 3377.035 1863.755 3379.435 1863.895 ;
        RECT 3377.020 1863.615 3379.435 1863.755 ;
        RECT 3377.020 1861.830 3377.160 1863.615 ;
      LAYER met2 ;
        RECT 3379.715 1863.335 3588.000 1864.175 ;
      LAYER met2 ;
        RECT 3376.960 1861.510 3377.220 1861.830 ;
      LAYER met2 ;
        RECT 3379.435 1861.415 3588.000 1863.335 ;
      LAYER met2 ;
        RECT 3377.035 1860.855 3379.435 1861.135 ;
      LAYER met2 ;
        RECT 3379.715 1860.575 3588.000 1861.415 ;
        RECT 3379.435 1858.195 3588.000 1860.575 ;
        RECT 3379.715 1857.355 3588.000 1858.195 ;
        RECT 3379.435 1854.975 3588.000 1857.355 ;
      LAYER met2 ;
        RECT 3377.035 1854.625 3379.435 1854.695 ;
        RECT 3376.560 1854.485 3379.435 1854.625 ;
        RECT 3377.035 1854.415 3379.435 1854.485 ;
      LAYER met2 ;
        RECT 3379.715 1854.135 3588.000 1854.975 ;
        RECT 3379.435 1853.085 3588.000 1854.135 ;
        RECT 3379.435 1705.795 3588.000 1706.790 ;
        RECT 3379.715 1704.955 3588.000 1705.795 ;
        RECT 3379.435 1703.035 3588.000 1704.955 ;
        RECT 3379.715 1702.195 3588.000 1703.035 ;
        RECT 3379.435 1699.815 3588.000 1702.195 ;
        RECT 3379.715 1698.975 3588.000 1699.815 ;
        RECT 3379.435 1696.595 3588.000 1698.975 ;
        RECT 3379.715 1695.755 3588.000 1696.595 ;
        RECT 3379.435 1693.835 3588.000 1695.755 ;
        RECT 3379.715 1692.995 3588.000 1693.835 ;
        RECT 3379.435 1690.615 3588.000 1692.995 ;
      LAYER met2 ;
        RECT 3377.035 1690.140 3379.435 1690.335 ;
        RECT 3377.020 1690.055 3379.435 1690.140 ;
        RECT 3377.020 1687.750 3377.160 1690.055 ;
      LAYER met2 ;
        RECT 3379.715 1689.775 3588.000 1690.615 ;
      LAYER met2 ;
        RECT 3376.960 1687.430 3377.220 1687.750 ;
      LAYER met2 ;
        RECT 3379.435 1687.395 3588.000 1689.775 ;
        RECT 3379.715 1686.555 3588.000 1687.395 ;
        RECT 3379.435 1684.635 3588.000 1686.555 ;
        RECT 3379.715 1683.795 3588.000 1684.635 ;
        RECT 3379.435 1681.415 3588.000 1683.795 ;
        RECT 3379.715 1680.575 3588.000 1681.415 ;
        RECT 3379.435 1678.195 3588.000 1680.575 ;
        RECT 3379.715 1677.355 3588.000 1678.195 ;
        RECT 3379.435 1675.435 3588.000 1677.355 ;
      LAYER met2 ;
        RECT 3377.035 1675.015 3379.435 1675.155 ;
        RECT 3377.020 1674.875 3379.435 1675.015 ;
        RECT 3377.020 1672.450 3377.160 1674.875 ;
      LAYER met2 ;
        RECT 3379.715 1674.595 3588.000 1675.435 ;
      LAYER met2 ;
        RECT 3370.060 1672.130 3370.320 1672.450 ;
        RECT 3376.960 1672.130 3377.220 1672.450 ;
      LAYER met2 ;
        RECT 3379.435 1672.215 3588.000 1674.595 ;
      LAYER met2 ;
        RECT 3369.600 1640.170 3369.860 1640.490 ;
        RECT 3367.360 1476.530 3367.960 1476.670 ;
        RECT 3367.360 1466.070 3367.500 1476.530 ;
        RECT 3367.300 1465.750 3367.560 1466.070 ;
        RECT 214.000 1406.590 214.260 1406.910 ;
        RECT 213.540 1359.330 213.800 1359.650 ;
        RECT 213.600 1228.270 213.740 1359.330 ;
        RECT 3367.360 1243.030 3367.500 1465.750 ;
        RECT 3367.760 1447.390 3368.020 1447.710 ;
        RECT 3367.300 1242.710 3367.560 1243.030 ;
        RECT 213.140 1228.130 213.740 1228.270 ;
        RECT 212.620 1158.390 212.880 1158.710 ;
        RECT 212.680 1137.630 212.820 1158.390 ;
        RECT 213.140 1143.410 213.280 1228.130 ;
        RECT 3367.820 1224.670 3367.960 1447.390 ;
        RECT 3369.660 1415.410 3369.800 1640.170 ;
        RECT 3370.120 1447.710 3370.260 1672.130 ;
      LAYER met2 ;
        RECT 3379.715 1671.375 3588.000 1672.215 ;
        RECT 3379.435 1668.995 3588.000 1671.375 ;
      LAYER met2 ;
        RECT 3377.035 1668.645 3379.435 1668.715 ;
        RECT 3376.560 1668.505 3379.435 1668.645 ;
        RECT 3376.560 1628.625 3376.700 1668.505 ;
        RECT 3377.035 1668.435 3379.435 1668.505 ;
      LAYER met2 ;
        RECT 3379.715 1668.155 3588.000 1668.995 ;
        RECT 3379.435 1665.775 3588.000 1668.155 ;
        RECT 3379.715 1664.935 3588.000 1665.775 ;
        RECT 3379.435 1663.015 3588.000 1664.935 ;
        RECT 3379.715 1662.175 3588.000 1663.015 ;
        RECT 3379.435 1659.795 3588.000 1662.175 ;
        RECT 3379.715 1658.955 3588.000 1659.795 ;
        RECT 3379.435 1656.575 3588.000 1658.955 ;
        RECT 3379.715 1655.735 3588.000 1656.575 ;
        RECT 3379.435 1653.815 3588.000 1655.735 ;
      LAYER met2 ;
        RECT 3377.035 1653.255 3379.435 1653.535 ;
      LAYER met2 ;
        RECT 3379.715 1652.975 3588.000 1653.815 ;
        RECT 3379.435 1650.595 3588.000 1652.975 ;
        RECT 3379.715 1649.755 3588.000 1650.595 ;
        RECT 3379.435 1647.375 3588.000 1649.755 ;
      LAYER met2 ;
        RECT 3377.035 1646.815 3379.435 1647.095 ;
      LAYER met2 ;
        RECT 3379.715 1646.535 3588.000 1647.375 ;
        RECT 3379.435 1644.615 3588.000 1646.535 ;
      LAYER met2 ;
        RECT 3377.035 1644.055 3379.435 1644.335 ;
      LAYER met2 ;
        RECT 3379.715 1643.775 3588.000 1644.615 ;
        RECT 3379.435 1641.395 3588.000 1643.775 ;
        RECT 3379.715 1640.555 3588.000 1641.395 ;
      LAYER met2 ;
        RECT 3376.960 1640.170 3377.220 1640.490 ;
        RECT 3377.020 1637.895 3377.160 1640.170 ;
      LAYER met2 ;
        RECT 3379.435 1638.175 3588.000 1640.555 ;
      LAYER met2 ;
        RECT 3377.020 1637.780 3379.435 1637.895 ;
        RECT 3377.035 1637.615 3379.435 1637.780 ;
      LAYER met2 ;
        RECT 3379.715 1637.335 3588.000 1638.175 ;
        RECT 3379.435 1635.415 3588.000 1637.335 ;
      LAYER met2 ;
        RECT 3377.035 1634.855 3379.435 1635.135 ;
      LAYER met2 ;
        RECT 3379.715 1634.575 3588.000 1635.415 ;
        RECT 3379.435 1632.195 3588.000 1634.575 ;
        RECT 3379.715 1631.355 3588.000 1632.195 ;
        RECT 3379.435 1628.975 3588.000 1631.355 ;
      LAYER met2 ;
        RECT 3377.035 1628.625 3379.435 1628.695 ;
        RECT 3376.560 1628.485 3379.435 1628.625 ;
        RECT 3377.035 1628.415 3379.435 1628.485 ;
      LAYER met2 ;
        RECT 3379.715 1628.135 3588.000 1628.975 ;
        RECT 3379.435 1627.085 3588.000 1628.135 ;
        RECT 3379.435 1480.795 3588.000 1481.790 ;
        RECT 3379.715 1479.955 3588.000 1480.795 ;
        RECT 3379.435 1478.035 3588.000 1479.955 ;
        RECT 3379.715 1477.195 3588.000 1478.035 ;
        RECT 3379.435 1474.815 3588.000 1477.195 ;
        RECT 3379.715 1473.975 3588.000 1474.815 ;
        RECT 3379.435 1471.595 3588.000 1473.975 ;
        RECT 3379.715 1470.755 3588.000 1471.595 ;
        RECT 3379.435 1468.835 3588.000 1470.755 ;
        RECT 3379.715 1467.995 3588.000 1468.835 ;
      LAYER met2 ;
        RECT 3376.960 1465.750 3377.220 1466.070 ;
        RECT 3377.020 1465.335 3377.160 1465.750 ;
      LAYER met2 ;
        RECT 3379.435 1465.615 3588.000 1467.995 ;
      LAYER met2 ;
        RECT 3377.020 1465.060 3379.435 1465.335 ;
        RECT 3377.035 1465.055 3379.435 1465.060 ;
      LAYER met2 ;
        RECT 3379.715 1464.775 3588.000 1465.615 ;
        RECT 3379.435 1462.395 3588.000 1464.775 ;
        RECT 3379.715 1461.555 3588.000 1462.395 ;
        RECT 3379.435 1459.635 3588.000 1461.555 ;
        RECT 3379.715 1458.795 3588.000 1459.635 ;
        RECT 3379.435 1456.415 3588.000 1458.795 ;
        RECT 3379.715 1455.575 3588.000 1456.415 ;
        RECT 3379.435 1453.195 3588.000 1455.575 ;
        RECT 3379.715 1452.355 3588.000 1453.195 ;
        RECT 3379.435 1450.435 3588.000 1452.355 ;
      LAYER met2 ;
        RECT 3377.035 1450.100 3379.435 1450.155 ;
        RECT 3377.020 1449.875 3379.435 1450.100 ;
        RECT 3377.020 1447.710 3377.160 1449.875 ;
      LAYER met2 ;
        RECT 3379.715 1449.595 3588.000 1450.435 ;
      LAYER met2 ;
        RECT 3370.060 1447.390 3370.320 1447.710 ;
        RECT 3376.960 1447.390 3377.220 1447.710 ;
      LAYER met2 ;
        RECT 3379.435 1447.215 3588.000 1449.595 ;
        RECT 3379.715 1446.375 3588.000 1447.215 ;
        RECT 3379.435 1443.995 3588.000 1446.375 ;
      LAYER met2 ;
        RECT 3377.035 1443.645 3379.435 1443.715 ;
        RECT 3376.560 1443.505 3379.435 1443.645 ;
        RECT 3369.600 1415.090 3369.860 1415.410 ;
        RECT 3369.660 1380.070 3369.800 1415.090 ;
        RECT 3376.560 1403.625 3376.700 1443.505 ;
        RECT 3377.035 1443.435 3379.435 1443.505 ;
      LAYER met2 ;
        RECT 3379.715 1443.155 3588.000 1443.995 ;
        RECT 3379.435 1440.775 3588.000 1443.155 ;
        RECT 3379.715 1439.935 3588.000 1440.775 ;
        RECT 3379.435 1438.015 3588.000 1439.935 ;
        RECT 3379.715 1437.175 3588.000 1438.015 ;
        RECT 3379.435 1434.795 3588.000 1437.175 ;
        RECT 3379.715 1433.955 3588.000 1434.795 ;
        RECT 3379.435 1431.575 3588.000 1433.955 ;
        RECT 3379.715 1430.735 3588.000 1431.575 ;
        RECT 3379.435 1428.815 3588.000 1430.735 ;
      LAYER met2 ;
        RECT 3377.035 1428.255 3379.435 1428.535 ;
      LAYER met2 ;
        RECT 3379.715 1427.975 3588.000 1428.815 ;
        RECT 3379.435 1425.595 3588.000 1427.975 ;
        RECT 3379.715 1424.755 3588.000 1425.595 ;
        RECT 3379.435 1422.375 3588.000 1424.755 ;
      LAYER met2 ;
        RECT 3377.035 1421.815 3379.435 1422.095 ;
      LAYER met2 ;
        RECT 3379.715 1421.535 3588.000 1422.375 ;
        RECT 3379.435 1419.615 3588.000 1421.535 ;
      LAYER met2 ;
        RECT 3377.035 1419.055 3379.435 1419.335 ;
      LAYER met2 ;
        RECT 3379.715 1418.775 3588.000 1419.615 ;
        RECT 3379.435 1416.395 3588.000 1418.775 ;
        RECT 3379.715 1415.555 3588.000 1416.395 ;
      LAYER met2 ;
        RECT 3376.960 1415.090 3377.220 1415.410 ;
        RECT 3377.020 1412.895 3377.160 1415.090 ;
      LAYER met2 ;
        RECT 3379.435 1413.175 3588.000 1415.555 ;
      LAYER met2 ;
        RECT 3377.020 1412.700 3379.435 1412.895 ;
        RECT 3377.035 1412.615 3379.435 1412.700 ;
      LAYER met2 ;
        RECT 3379.715 1412.335 3588.000 1413.175 ;
        RECT 3379.435 1410.415 3588.000 1412.335 ;
      LAYER met2 ;
        RECT 3377.035 1409.855 3379.435 1410.135 ;
      LAYER met2 ;
        RECT 3379.715 1409.575 3588.000 1410.415 ;
        RECT 3379.435 1407.195 3588.000 1409.575 ;
        RECT 3379.715 1406.355 3588.000 1407.195 ;
        RECT 3379.435 1403.975 3588.000 1406.355 ;
      LAYER met2 ;
        RECT 3377.035 1403.625 3379.435 1403.695 ;
        RECT 3376.560 1403.485 3379.435 1403.625 ;
        RECT 3377.035 1403.415 3379.435 1403.485 ;
      LAYER met2 ;
        RECT 3379.715 1403.135 3588.000 1403.975 ;
        RECT 3379.435 1402.085 3588.000 1403.135 ;
      LAYER met2 ;
        RECT 3368.740 1379.930 3369.800 1380.070 ;
        RECT 3368.740 1324.870 3368.880 1379.930 ;
        RECT 3368.740 1324.730 3369.800 1324.870 ;
        RECT 3367.760 1224.350 3368.020 1224.670 ;
        RECT 213.080 1143.090 213.340 1143.410 ;
        RECT 212.620 1137.310 212.880 1137.630 ;
        RECT 212.220 1131.530 212.820 1131.670 ;
        RECT 211.300 986.950 211.900 987.090 ;
      LAYER met2 ;
        RECT 0.000 986.025 208.285 986.865 ;
      LAYER met2 ;
        RECT 208.565 986.410 210.965 986.585 ;
        RECT 208.565 986.305 211.440 986.410 ;
        RECT 208.610 986.270 211.440 986.305 ;
      LAYER met2 ;
        RECT 0.000 983.645 208.565 986.025 ;
        RECT 0.000 982.805 208.285 983.645 ;
        RECT 0.000 980.425 208.565 982.805 ;
        RECT 0.000 979.585 208.285 980.425 ;
      LAYER met2 ;
        RECT 208.565 979.865 210.965 980.145 ;
      LAYER met2 ;
        RECT 0.000 977.665 208.565 979.585 ;
      LAYER met2 ;
        RECT 208.940 979.210 209.200 979.530 ;
      LAYER met2 ;
        RECT 0.000 976.825 208.285 977.665 ;
      LAYER met2 ;
        RECT 209.000 977.385 209.140 979.210 ;
        RECT 208.565 977.105 210.965 977.385 ;
      LAYER met2 ;
        RECT 0.000 974.445 208.565 976.825 ;
        RECT 0.000 973.605 208.285 974.445 ;
        RECT 0.000 971.225 208.565 973.605 ;
        RECT 0.000 970.385 208.285 971.225 ;
      LAYER met2 ;
        RECT 208.565 970.665 210.965 970.945 ;
      LAYER met2 ;
        RECT 0.000 968.465 208.565 970.385 ;
        RECT 0.000 967.625 208.285 968.465 ;
      LAYER met2 ;
        RECT 208.565 967.905 210.965 968.185 ;
      LAYER met2 ;
        RECT 0.000 965.245 208.565 967.625 ;
        RECT 0.000 964.405 208.285 965.245 ;
        RECT 0.000 962.025 208.565 964.405 ;
        RECT 0.000 961.185 208.285 962.025 ;
      LAYER met2 ;
        RECT 208.565 961.465 210.965 961.745 ;
      LAYER met2 ;
        RECT 0.000 959.265 208.565 961.185 ;
        RECT 0.000 958.425 208.285 959.265 ;
        RECT 0.000 956.045 208.565 958.425 ;
        RECT 0.000 955.205 208.285 956.045 ;
        RECT 0.000 952.825 208.565 955.205 ;
        RECT 0.000 951.985 208.285 952.825 ;
        RECT 0.000 950.065 208.565 951.985 ;
        RECT 0.000 949.225 208.285 950.065 ;
        RECT 0.000 946.845 208.565 949.225 ;
      LAYER met2 ;
        RECT 211.300 946.970 211.440 986.270 ;
      LAYER met2 ;
        RECT 0.000 946.005 208.285 946.845 ;
      LAYER met2 ;
        RECT 209.460 946.830 211.440 946.970 ;
        RECT 209.460 946.565 209.600 946.830 ;
        RECT 208.565 946.285 210.965 946.565 ;
      LAYER met2 ;
        RECT 0.000 943.625 208.565 946.005 ;
        RECT 0.000 942.785 208.285 943.625 ;
        RECT 0.000 940.405 208.565 942.785 ;
      LAYER met2 ;
        RECT 211.760 940.850 211.900 986.950 ;
        RECT 212.680 979.530 212.820 1131.530 ;
        RECT 212.620 979.210 212.880 979.530 ;
        RECT 209.460 940.710 211.900 940.850 ;
      LAYER met2 ;
        RECT 0.000 939.565 208.285 940.405 ;
      LAYER met2 ;
        RECT 209.460 940.170 209.600 940.710 ;
        RECT 208.610 940.125 209.600 940.170 ;
        RECT 209.920 940.125 210.060 940.710 ;
        RECT 208.565 939.845 210.965 940.125 ;
      LAYER met2 ;
        RECT 0.000 937.645 208.565 939.565 ;
      LAYER met2 ;
        RECT 209.920 938.050 210.060 939.845 ;
        RECT 212.680 938.470 212.820 979.210 ;
        RECT 212.220 938.330 212.820 938.470 ;
        RECT 209.860 937.730 210.120 938.050 ;
      LAYER met2 ;
        RECT 0.000 936.805 208.285 937.645 ;
        RECT 0.000 934.425 208.565 936.805 ;
        RECT 0.000 933.585 208.285 934.425 ;
        RECT 0.000 931.205 208.565 933.585 ;
        RECT 0.000 930.365 208.285 931.205 ;
        RECT 0.000 928.445 208.565 930.365 ;
        RECT 0.000 927.605 208.285 928.445 ;
        RECT 0.000 925.225 208.565 927.605 ;
        RECT 0.000 924.385 208.285 925.225 ;
      LAYER met2 ;
        RECT 208.565 924.665 210.965 924.945 ;
      LAYER met2 ;
        RECT 0.000 922.005 208.565 924.385 ;
      LAYER met2 ;
        RECT 209.000 922.410 209.140 924.665 ;
        RECT 208.940 922.090 209.200 922.410 ;
      LAYER met2 ;
        RECT 0.000 921.165 208.285 922.005 ;
        RECT 0.000 919.245 208.565 921.165 ;
      LAYER met2 ;
        RECT 211.240 920.730 211.500 921.050 ;
      LAYER met2 ;
        RECT 0.000 918.405 208.285 919.245 ;
        RECT 0.000 916.025 208.565 918.405 ;
        RECT 0.000 915.185 208.285 916.025 ;
        RECT 0.000 912.805 208.565 915.185 ;
        RECT 0.000 911.965 208.285 912.805 ;
        RECT 0.000 910.045 208.565 911.965 ;
        RECT 0.000 909.205 208.285 910.045 ;
        RECT 0.000 908.210 208.565 909.205 ;
        RECT 4.925 601.390 200.000 625.290 ;
        RECT 4.925 575.395 197.965 601.390 ;
        RECT 198.080 576.895 200.000 578.895 ;
        RECT 4.925 551.495 200.000 575.395 ;
        RECT 4.925 551.265 197.965 551.495 ;
        RECT 153.765 415.000 158.415 426.140 ;
        RECT 159.640 415.245 163.510 426.195 ;
        RECT 3.570 414.700 197.965 415.000 ;
        RECT 3.570 394.095 198.000 414.700 ;
        RECT 3.570 393.535 197.965 394.095 ;
        RECT 3.570 360.925 198.000 393.535 ;
        RECT 3.570 360.495 197.965 360.925 ;
        RECT 3.570 340.500 198.000 360.495 ;
        RECT 3.570 340.490 197.965 340.500 ;
      LAYER met2 ;
        RECT 211.300 228.130 211.440 920.730 ;
        RECT 212.220 414.450 212.360 938.330 ;
        RECT 212.620 937.730 212.880 938.050 ;
        RECT 212.680 607.570 212.820 937.730 ;
        RECT 213.140 922.410 213.280 1143.090 ;
        RECT 3367.820 996.530 3367.960 1224.350 ;
        RECT 3369.660 1188.630 3369.800 1324.730 ;
      LAYER met2 ;
        RECT 3379.435 1255.795 3588.000 1256.790 ;
        RECT 3379.715 1254.955 3588.000 1255.795 ;
        RECT 3379.435 1253.035 3588.000 1254.955 ;
        RECT 3379.715 1252.195 3588.000 1253.035 ;
        RECT 3379.435 1249.815 3588.000 1252.195 ;
        RECT 3379.715 1248.975 3588.000 1249.815 ;
        RECT 3379.435 1246.595 3588.000 1248.975 ;
        RECT 3379.715 1245.755 3588.000 1246.595 ;
        RECT 3379.435 1243.835 3588.000 1245.755 ;
      LAYER met2 ;
        RECT 3370.060 1242.710 3370.320 1243.030 ;
        RECT 3376.960 1242.710 3377.220 1243.030 ;
      LAYER met2 ;
        RECT 3379.715 1242.995 3588.000 1243.835 ;
      LAYER met2 ;
        RECT 3369.600 1188.310 3369.860 1188.630 ;
        RECT 3367.760 996.210 3368.020 996.530 ;
        RECT 213.080 922.090 213.340 922.410 ;
        RECT 3367.300 791.530 3367.560 791.850 ;
        RECT 212.620 607.250 212.880 607.570 ;
        RECT 220.900 607.250 221.160 607.570 ;
        RECT 220.960 552.685 221.100 607.250 ;
        RECT 3367.360 566.090 3367.500 791.530 ;
        RECT 3367.820 776.210 3367.960 996.210 ;
        RECT 3369.660 959.810 3369.800 1188.310 ;
        RECT 3370.120 1011.830 3370.260 1242.710 ;
        RECT 3377.020 1240.335 3377.160 1242.710 ;
      LAYER met2 ;
        RECT 3379.435 1240.615 3588.000 1242.995 ;
      LAYER met2 ;
        RECT 3377.020 1240.195 3379.435 1240.335 ;
        RECT 3377.035 1240.055 3379.435 1240.195 ;
      LAYER met2 ;
        RECT 3379.715 1239.775 3588.000 1240.615 ;
        RECT 3379.435 1237.395 3588.000 1239.775 ;
        RECT 3379.715 1236.555 3588.000 1237.395 ;
        RECT 3379.435 1234.635 3588.000 1236.555 ;
        RECT 3379.715 1233.795 3588.000 1234.635 ;
        RECT 3379.435 1231.415 3588.000 1233.795 ;
        RECT 3379.715 1230.575 3588.000 1231.415 ;
        RECT 3379.435 1228.195 3588.000 1230.575 ;
        RECT 3379.715 1227.355 3588.000 1228.195 ;
        RECT 3379.435 1225.435 3588.000 1227.355 ;
      LAYER met2 ;
        RECT 3377.035 1225.020 3379.435 1225.155 ;
        RECT 3377.020 1224.875 3379.435 1225.020 ;
        RECT 3377.020 1224.670 3377.160 1224.875 ;
        RECT 3376.960 1224.350 3377.220 1224.670 ;
      LAYER met2 ;
        RECT 3379.715 1224.595 3588.000 1225.435 ;
        RECT 3379.435 1222.215 3588.000 1224.595 ;
        RECT 3379.715 1221.375 3588.000 1222.215 ;
        RECT 3379.435 1218.995 3588.000 1221.375 ;
      LAYER met2 ;
        RECT 3377.035 1218.645 3379.435 1218.715 ;
        RECT 3376.560 1218.505 3379.435 1218.645 ;
        RECT 3376.560 1178.625 3376.700 1218.505 ;
        RECT 3377.035 1218.435 3379.435 1218.505 ;
      LAYER met2 ;
        RECT 3379.715 1218.155 3588.000 1218.995 ;
        RECT 3379.435 1215.775 3588.000 1218.155 ;
        RECT 3379.715 1214.935 3588.000 1215.775 ;
        RECT 3379.435 1213.015 3588.000 1214.935 ;
        RECT 3379.715 1212.175 3588.000 1213.015 ;
        RECT 3379.435 1209.795 3588.000 1212.175 ;
        RECT 3379.715 1208.955 3588.000 1209.795 ;
        RECT 3379.435 1206.575 3588.000 1208.955 ;
        RECT 3379.715 1205.735 3588.000 1206.575 ;
        RECT 3379.435 1203.815 3588.000 1205.735 ;
      LAYER met2 ;
        RECT 3377.035 1203.255 3379.435 1203.535 ;
      LAYER met2 ;
        RECT 3379.715 1202.975 3588.000 1203.815 ;
        RECT 3379.435 1200.595 3588.000 1202.975 ;
        RECT 3379.715 1199.755 3588.000 1200.595 ;
        RECT 3379.435 1197.375 3588.000 1199.755 ;
      LAYER met2 ;
        RECT 3377.035 1196.815 3379.435 1197.095 ;
      LAYER met2 ;
        RECT 3379.715 1196.535 3588.000 1197.375 ;
        RECT 3379.435 1194.615 3588.000 1196.535 ;
      LAYER met2 ;
        RECT 3377.035 1194.055 3379.435 1194.335 ;
      LAYER met2 ;
        RECT 3379.715 1193.775 3588.000 1194.615 ;
        RECT 3379.435 1191.395 3588.000 1193.775 ;
        RECT 3379.715 1190.555 3588.000 1191.395 ;
      LAYER met2 ;
        RECT 3376.960 1188.310 3377.220 1188.630 ;
        RECT 3377.020 1187.895 3377.160 1188.310 ;
      LAYER met2 ;
        RECT 3379.435 1188.175 3588.000 1190.555 ;
      LAYER met2 ;
        RECT 3377.020 1187.620 3379.435 1187.895 ;
        RECT 3377.035 1187.615 3379.435 1187.620 ;
      LAYER met2 ;
        RECT 3379.715 1187.335 3588.000 1188.175 ;
        RECT 3379.435 1185.415 3588.000 1187.335 ;
      LAYER met2 ;
        RECT 3377.035 1184.855 3379.435 1185.135 ;
      LAYER met2 ;
        RECT 3379.715 1184.575 3588.000 1185.415 ;
        RECT 3379.435 1182.195 3588.000 1184.575 ;
        RECT 3379.715 1181.355 3588.000 1182.195 ;
        RECT 3379.435 1178.975 3588.000 1181.355 ;
      LAYER met2 ;
        RECT 3377.035 1178.625 3379.435 1178.695 ;
        RECT 3376.560 1178.485 3379.435 1178.625 ;
        RECT 3377.035 1178.415 3379.435 1178.485 ;
      LAYER met2 ;
        RECT 3379.715 1178.135 3588.000 1178.975 ;
        RECT 3379.435 1177.085 3588.000 1178.135 ;
        RECT 3379.435 1029.795 3588.000 1030.790 ;
        RECT 3379.715 1028.955 3588.000 1029.795 ;
        RECT 3379.435 1027.035 3588.000 1028.955 ;
        RECT 3379.715 1026.195 3588.000 1027.035 ;
        RECT 3379.435 1023.815 3588.000 1026.195 ;
        RECT 3379.715 1022.975 3588.000 1023.815 ;
        RECT 3379.435 1020.595 3588.000 1022.975 ;
        RECT 3379.715 1019.755 3588.000 1020.595 ;
        RECT 3379.435 1017.835 3588.000 1019.755 ;
        RECT 3379.715 1016.995 3588.000 1017.835 ;
        RECT 3379.435 1014.615 3588.000 1016.995 ;
      LAYER met2 ;
        RECT 3377.035 1014.220 3379.435 1014.335 ;
        RECT 3377.020 1014.055 3379.435 1014.220 ;
        RECT 3377.020 1011.830 3377.160 1014.055 ;
      LAYER met2 ;
        RECT 3379.715 1013.775 3588.000 1014.615 ;
      LAYER met2 ;
        RECT 3370.060 1011.510 3370.320 1011.830 ;
        RECT 3376.960 1011.510 3377.220 1011.830 ;
        RECT 3369.600 959.490 3369.860 959.810 ;
        RECT 3367.760 775.890 3368.020 776.210 ;
        RECT 3367.300 565.770 3367.560 566.090 ;
        RECT 220.890 552.315 221.170 552.685 ;
        RECT 224.110 552.315 224.390 552.685 ;
        RECT 224.180 552.070 224.320 552.315 ;
        RECT 224.180 551.930 224.780 552.070 ;
        RECT 212.160 414.130 212.420 414.450 ;
        RECT 220.900 414.130 221.160 414.450 ;
        RECT 220.960 359.565 221.100 414.130 ;
        RECT 220.890 359.195 221.170 359.565 ;
        RECT 224.110 359.195 224.390 359.565 ;
        RECT 224.180 234.930 224.320 359.195 ;
        RECT 224.120 234.610 224.380 234.930 ;
        RECT 211.240 227.810 211.500 228.130 ;
        RECT 224.640 227.790 224.780 551.930 ;
        RECT 745.300 234.270 745.560 234.590 ;
        RECT 942.640 234.270 942.900 234.590 ;
        RECT 1004.280 234.270 1004.540 234.590 ;
        RECT 1281.200 234.270 1281.460 234.590 ;
        RECT 1488.660 234.270 1488.920 234.590 ;
        RECT 1547.080 234.270 1547.340 234.590 ;
        RECT 1762.820 234.270 1763.080 234.590 ;
        RECT 1821.240 234.270 1821.500 234.590 ;
        RECT 2036.980 234.270 2037.240 234.590 ;
        RECT 2095.400 234.270 2095.660 234.590 ;
        RECT 2310.680 234.270 2310.940 234.590 ;
        RECT 2369.100 234.270 2369.360 234.590 ;
        RECT 2584.840 234.270 2585.100 234.590 ;
        RECT 704.820 227.810 705.080 228.130 ;
        RECT 224.580 227.470 224.840 227.790 ;
        RECT 468.840 207.410 469.100 207.730 ;
        RECT 468.900 201.125 469.040 207.410 ;
        RECT 675.840 201.125 676.100 201.270 ;
        RECT 468.830 200.755 469.110 201.125 ;
        RECT 675.830 200.755 676.110 201.125 ;
        RECT 704.880 201.010 705.020 227.810 ;
        RECT 735.640 209.110 735.900 209.430 ;
        RECT 717.700 201.125 717.960 201.270 ;
        RECT 704.880 200.870 705.180 201.010 ;
        RECT 705.040 200.590 705.180 200.870 ;
        RECT 715.390 200.755 715.670 201.125 ;
        RECT 717.690 200.755 717.970 201.125 ;
        RECT 715.420 200.590 715.560 200.755 ;
        RECT 735.700 200.590 735.840 209.110 ;
        RECT 745.360 201.805 745.500 234.270 ;
        RECT 942.700 221.670 942.840 234.270 ;
        RECT 979.900 227.470 980.160 227.790 ;
        RECT 979.960 222.350 980.100 227.470 ;
        RECT 979.900 222.030 980.160 222.350 ;
        RECT 942.640 221.350 942.900 221.670 ;
        RECT 964.260 221.350 964.520 221.670 ;
        RECT 933.440 221.010 933.700 221.330 ;
        RECT 933.500 210.965 933.640 221.010 ;
        RECT 942.700 210.965 942.840 221.350 ;
        RECT 964.320 210.965 964.460 221.350 ;
        RECT 973.460 221.010 973.720 221.330 ;
        RECT 973.520 210.965 973.660 221.010 ;
        RECT 979.960 210.965 980.100 222.030 ;
        RECT 1004.340 210.965 1004.480 234.270 ;
        RECT 1007.500 221.350 1007.760 221.670 ;
        RECT 1007.560 210.965 1007.700 221.350 ;
        RECT 933.415 208.565 933.695 210.965 ;
        RECT 939.855 208.565 940.135 210.965 ;
        RECT 942.615 208.565 942.895 210.965 ;
        RECT 945.835 209.170 946.115 210.965 ;
        RECT 946.320 209.450 946.580 209.770 ;
        RECT 946.380 209.170 946.520 209.450 ;
        RECT 945.835 209.030 946.520 209.170 ;
        RECT 945.835 208.565 946.115 209.030 ;
        RECT 949.055 208.565 949.335 210.965 ;
        RECT 951.815 208.565 952.095 210.965 ;
        RECT 955.035 209.170 955.315 210.965 ;
        RECT 955.520 209.450 955.780 209.770 ;
        RECT 955.580 209.170 955.720 209.450 ;
        RECT 955.035 209.030 955.720 209.170 ;
        RECT 955.035 208.565 955.315 209.030 ;
        RECT 958.255 208.565 958.535 210.965 ;
        RECT 961.015 209.170 961.295 210.965 ;
        RECT 961.500 209.450 961.760 209.770 ;
        RECT 961.560 209.170 961.700 209.450 ;
        RECT 961.015 209.030 961.700 209.170 ;
        RECT 961.015 208.565 961.295 209.030 ;
        RECT 964.235 208.565 964.515 210.965 ;
        RECT 967.455 209.170 967.735 210.965 ;
        RECT 967.940 209.450 968.200 209.770 ;
        RECT 968.000 209.170 968.140 209.450 ;
        RECT 967.455 209.030 968.140 209.170 ;
        RECT 967.455 208.565 967.735 209.030 ;
        RECT 973.435 208.565 973.715 210.965 ;
        RECT 979.875 208.565 980.155 210.965 ;
        RECT 982.200 209.450 982.460 209.770 ;
        RECT 982.260 209.170 982.400 209.450 ;
        RECT 982.635 209.170 982.915 210.965 ;
        RECT 985.855 209.170 986.135 210.965 ;
        RECT 989.075 209.170 989.355 210.965 ;
        RECT 991.835 209.170 992.115 210.965 ;
        RECT 992.320 209.450 992.580 209.770 ;
        RECT 992.380 209.170 992.520 209.450 ;
        RECT 995.055 209.170 995.335 210.965 ;
        RECT 1000.600 209.450 1000.860 209.770 ;
        RECT 982.260 209.030 992.520 209.170 ;
        RECT 994.680 209.090 995.335 209.170 ;
        RECT 994.620 209.030 995.335 209.090 ;
        RECT 1000.660 209.170 1000.800 209.450 ;
        RECT 1001.035 209.170 1001.315 210.965 ;
        RECT 1004.255 209.170 1004.535 210.965 ;
        RECT 1000.660 209.030 1004.535 209.170 ;
        RECT 982.635 208.565 982.915 209.030 ;
        RECT 985.855 208.565 986.135 209.030 ;
        RECT 989.075 208.565 989.355 209.030 ;
        RECT 991.835 208.565 992.115 209.030 ;
        RECT 994.620 208.770 994.880 209.030 ;
        RECT 995.055 208.565 995.335 209.030 ;
        RECT 1001.035 208.565 1001.315 209.030 ;
        RECT 1004.255 208.565 1004.535 209.030 ;
        RECT 1007.475 208.565 1007.755 210.965 ;
        RECT 1010.235 208.565 1010.515 210.965 ;
      LAYER met2 ;
        RECT 932.085 208.285 933.135 208.565 ;
        RECT 933.975 208.285 936.355 208.565 ;
        RECT 937.195 208.285 939.575 208.565 ;
        RECT 940.415 208.285 942.335 208.565 ;
        RECT 943.175 208.285 945.555 208.565 ;
        RECT 946.395 208.285 948.775 208.565 ;
        RECT 949.615 208.285 951.535 208.565 ;
        RECT 952.375 208.285 954.755 208.565 ;
        RECT 955.595 208.285 957.975 208.565 ;
        RECT 958.815 208.285 960.735 208.565 ;
        RECT 961.575 208.285 963.955 208.565 ;
        RECT 964.795 208.285 967.175 208.565 ;
        RECT 968.015 208.285 969.935 208.565 ;
        RECT 970.775 208.285 973.155 208.565 ;
        RECT 973.995 208.285 976.375 208.565 ;
        RECT 977.215 208.285 979.595 208.565 ;
        RECT 980.435 208.285 982.355 208.565 ;
        RECT 983.195 208.285 985.575 208.565 ;
        RECT 986.415 208.285 988.795 208.565 ;
        RECT 989.635 208.285 991.555 208.565 ;
        RECT 992.395 208.285 994.775 208.565 ;
        RECT 995.615 208.285 997.995 208.565 ;
        RECT 998.835 208.285 1000.755 208.565 ;
        RECT 1001.595 208.285 1003.975 208.565 ;
        RECT 1004.815 208.285 1007.195 208.565 ;
        RECT 1008.035 208.285 1009.955 208.565 ;
        RECT 1010.795 208.285 1011.790 208.565 ;
      LAYER met2 ;
        RECT 745.290 201.435 745.570 201.805 ;
        RECT 704.980 200.270 705.240 200.590 ;
        RECT 715.360 200.270 715.620 200.590 ;
        RECT 722.760 200.270 723.020 200.590 ;
        RECT 735.640 200.270 735.900 200.590 ;
        RECT 705.040 200.000 705.180 200.270 ;
        RECT 715.420 200.000 715.560 200.270 ;
        RECT 722.820 200.000 722.960 200.270 ;
      LAYER met2 ;
        RECT 394.710 197.965 418.610 200.000 ;
        RECT 441.105 198.080 443.105 200.000 ;
        RECT 444.605 197.965 468.505 200.000 ;
        RECT 663.085 199.390 664.485 200.000 ;
      LAYER met2 ;
        RECT 664.765 199.670 665.785 200.000 ;
      LAYER met2 ;
        RECT 666.065 199.390 704.700 200.000 ;
        RECT 663.085 199.080 704.700 199.390 ;
      LAYER met2 ;
        RECT 704.980 199.360 705.240 200.000 ;
      LAYER met2 ;
        RECT 705.520 199.390 706.565 200.000 ;
      LAYER met2 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met2 ;
        RECT 707.775 199.390 708.055 200.000 ;
      LAYER met2 ;
        RECT 708.335 199.670 709.065 200.000 ;
      LAYER met2 ;
        RECT 709.345 199.390 709.490 200.000 ;
      LAYER met2 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met2 ;
        RECT 710.700 199.390 715.060 200.000 ;
        RECT 705.520 199.080 715.060 199.390 ;
        RECT 394.710 4.925 468.735 197.965 ;
        RECT 663.085 196.020 715.060 199.080 ;
        RECT 663.085 195.735 714.775 196.020 ;
      LAYER met2 ;
        RECT 715.340 195.755 715.640 200.000 ;
      LAYER met2 ;
        RECT 715.920 198.310 716.495 200.000 ;
      LAYER met2 ;
        RECT 716.775 198.590 717.925 200.000 ;
      LAYER met2 ;
        RECT 718.205 199.155 718.810 200.000 ;
      LAYER met2 ;
        RECT 719.090 199.435 720.755 200.000 ;
      LAYER met2 ;
        RECT 721.035 199.155 722.585 200.000 ;
      LAYER met2 ;
        RECT 722.820 199.580 723.445 200.000 ;
      LAYER met2 ;
        RECT 718.205 198.735 722.585 199.155 ;
      LAYER met2 ;
        RECT 722.865 199.015 723.445 199.580 ;
      LAYER met2 ;
        RECT 723.725 198.735 725.175 200.000 ;
        RECT 718.205 198.310 725.175 198.735 ;
        RECT 715.920 198.250 725.175 198.310 ;
        RECT 725.995 199.390 728.825 200.000 ;
      LAYER met2 ;
        RECT 729.105 199.670 729.575 200.000 ;
      LAYER met2 ;
        RECT 729.855 199.390 737.660 200.000 ;
        RECT 725.995 198.250 737.660 199.390 ;
        RECT 715.920 196.845 737.660 198.250 ;
        RECT 715.920 196.485 722.475 196.845 ;
        RECT 727.600 196.705 737.660 196.845 ;
        RECT 715.920 196.215 722.205 196.485 ;
      LAYER met2 ;
        RECT 722.755 196.425 727.320 196.565 ;
        RECT 722.755 196.355 727.650 196.425 ;
      LAYER met2 ;
        RECT 727.930 196.375 737.660 196.705 ;
      LAYER met2 ;
        RECT 722.755 196.305 727.180 196.355 ;
      LAYER met2 ;
        RECT 715.920 196.035 721.835 196.215 ;
      LAYER met2 ;
        RECT 722.755 196.205 723.115 196.305 ;
        RECT 723.125 196.205 723.225 196.305 ;
        RECT 727.070 196.235 727.305 196.305 ;
        RECT 727.320 196.235 727.650 196.355 ;
      LAYER met2 ;
        RECT 716.220 195.845 721.835 196.035 ;
      LAYER met2 ;
        RECT 722.485 196.165 722.755 196.205 ;
        RECT 722.855 196.165 723.125 196.205 ;
        RECT 722.485 196.025 723.125 196.165 ;
        RECT 727.070 196.095 727.650 196.235 ;
        RECT 727.070 196.070 727.305 196.095 ;
        RECT 722.485 195.935 722.755 196.025 ;
        RECT 722.855 195.935 723.125 196.025 ;
        RECT 715.340 195.740 715.940 195.755 ;
      LAYER met2 ;
        RECT 663.085 195.380 708.600 195.735 ;
      LAYER met2 ;
        RECT 715.055 195.455 715.940 195.740 ;
      LAYER met2 ;
        RECT 716.220 195.735 721.725 195.845 ;
      LAYER met2 ;
        RECT 722.115 195.565 722.855 195.935 ;
      LAYER met2 ;
        RECT 723.505 195.925 726.790 196.025 ;
        RECT 723.405 195.790 726.790 195.925 ;
      LAYER met2 ;
        RECT 727.305 195.955 727.625 196.070 ;
        RECT 727.650 195.955 727.995 196.095 ;
      LAYER met2 ;
        RECT 728.275 196.030 737.660 196.375 ;
      LAYER met2 ;
        RECT 727.305 195.815 727.995 195.955 ;
      LAYER met2 ;
        RECT 723.405 195.655 727.025 195.790 ;
      LAYER met2 ;
        RECT 727.305 195.750 727.625 195.815 ;
        RECT 727.650 195.750 727.995 195.815 ;
        RECT 722.005 195.455 722.485 195.565 ;
      LAYER met2 ;
        RECT 663.085 195.050 708.270 195.380 ;
      LAYER met2 ;
        RECT 708.880 195.315 722.485 195.455 ;
        RECT 708.880 195.245 709.235 195.315 ;
        RECT 715.340 195.245 715.640 195.315 ;
        RECT 722.115 195.245 722.485 195.315 ;
      LAYER met2 ;
        RECT 723.135 195.470 727.025 195.655 ;
      LAYER met2 ;
        RECT 727.625 195.675 727.955 195.750 ;
        RECT 727.995 195.675 728.265 195.750 ;
      LAYER met2 ;
        RECT 723.135 195.285 727.345 195.470 ;
      LAYER met2 ;
        RECT 727.625 195.425 728.265 195.675 ;
        RECT 727.625 195.420 727.955 195.425 ;
        RECT 708.880 195.195 722.485 195.245 ;
        RECT 708.880 195.100 709.235 195.195 ;
        RECT 709.250 195.100 709.345 195.195 ;
      LAYER met2 ;
        RECT 722.765 195.140 727.345 195.285 ;
      LAYER met2 ;
        RECT 708.550 195.055 708.880 195.100 ;
        RECT 708.920 195.055 709.250 195.100 ;
      LAYER met2 ;
        RECT 663.085 189.305 708.140 195.050 ;
      LAYER met2 ;
        RECT 708.550 194.845 709.250 195.055 ;
      LAYER met2 ;
        RECT 722.765 194.915 727.725 195.140 ;
      LAYER met2 ;
        RECT 708.550 194.770 708.880 194.845 ;
        RECT 708.920 194.770 709.250 194.845 ;
      LAYER met2 ;
        RECT 709.625 194.820 727.725 194.915 ;
      LAYER met2 ;
        RECT 708.420 194.640 708.550 194.770 ;
        RECT 708.680 194.640 708.920 194.770 ;
        RECT 708.420 194.530 708.920 194.640 ;
      LAYER met2 ;
        RECT 663.085 189.115 707.950 189.305 ;
        RECT 663.085 184.635 707.690 189.115 ;
      LAYER met2 ;
        RECT 708.420 189.025 708.680 194.530 ;
      LAYER met2 ;
        RECT 709.530 194.490 727.725 194.820 ;
        RECT 709.200 194.250 727.725 194.490 ;
      LAYER met2 ;
        RECT 708.230 188.915 708.680 189.025 ;
        RECT 708.230 188.835 708.420 188.915 ;
        RECT 708.600 188.835 708.680 188.915 ;
      LAYER met2 ;
        RECT 708.960 191.420 727.725 194.250 ;
        RECT 708.960 191.080 727.385 191.420 ;
      LAYER met2 ;
        RECT 728.005 191.140 728.265 195.425 ;
      LAYER met2 ;
        RECT 708.960 190.880 727.185 191.080 ;
      LAYER met2 ;
        RECT 727.665 190.890 728.265 191.140 ;
      LAYER met2 ;
        RECT 708.960 190.550 726.855 190.880 ;
      LAYER met2 ;
        RECT 727.665 190.800 728.005 190.890 ;
        RECT 728.035 190.800 728.265 190.890 ;
        RECT 727.465 190.750 727.665 190.800 ;
        RECT 727.835 190.750 728.035 190.800 ;
        RECT 727.465 190.680 728.035 190.750 ;
        RECT 727.465 190.600 727.665 190.680 ;
        RECT 727.835 190.600 728.035 190.680 ;
        RECT 707.970 188.465 708.600 188.835 ;
      LAYER met2 ;
        RECT 708.960 188.555 726.595 190.550 ;
      LAYER met2 ;
        RECT 727.135 190.540 727.465 190.600 ;
        RECT 727.505 190.540 727.835 190.600 ;
        RECT 727.135 190.400 727.835 190.540 ;
      LAYER met2 ;
        RECT 728.545 190.520 737.660 196.030 ;
      LAYER met2 ;
        RECT 727.135 190.270 727.465 190.400 ;
        RECT 727.505 190.270 727.835 190.400 ;
      LAYER met2 ;
        RECT 728.315 190.320 737.660 190.520 ;
        RECT 663.085 184.300 707.355 184.635 ;
      LAYER met2 ;
        RECT 707.970 184.355 708.230 188.465 ;
      LAYER met2 ;
        RECT 708.880 188.185 726.595 188.555 ;
        RECT 663.085 179.225 707.095 184.300 ;
      LAYER met2 ;
        RECT 707.635 184.105 708.230 184.355 ;
        RECT 707.635 184.020 707.970 184.105 ;
        RECT 708.005 184.020 708.230 184.105 ;
        RECT 707.375 183.650 708.005 184.020 ;
      LAYER met2 ;
        RECT 708.510 183.740 726.595 188.185 ;
      LAYER met2 ;
        RECT 707.375 179.505 707.635 183.650 ;
      LAYER met2 ;
        RECT 708.285 183.370 726.595 183.740 ;
        RECT 707.915 179.225 726.595 183.370 ;
        RECT 663.085 172.420 726.595 179.225 ;
      LAYER met2 ;
        RECT 726.875 189.900 727.505 190.270 ;
      LAYER met2 ;
        RECT 728.115 189.990 737.660 190.320 ;
      LAYER met2 ;
        RECT 726.875 173.390 727.135 189.900 ;
      LAYER met2 ;
        RECT 727.785 189.620 737.660 189.990 ;
        RECT 727.415 173.670 737.660 189.620 ;
      LAYER met2 ;
        RECT 726.875 172.700 727.350 173.390 ;
      LAYER met2 ;
        RECT 663.085 172.345 726.810 172.420 ;
        RECT 663.085 169.195 726.595 172.345 ;
      LAYER met2 ;
        RECT 727.090 172.065 727.350 172.700 ;
        RECT 726.875 171.855 727.350 172.065 ;
        RECT 726.875 171.850 727.090 171.855 ;
        RECT 726.875 171.375 727.350 171.850 ;
      LAYER met2 ;
        RECT 663.085 169.050 726.450 169.195 ;
        RECT 663.085 168.825 726.225 169.050 ;
      LAYER met2 ;
        RECT 726.875 168.915 727.135 171.375 ;
      LAYER met2 ;
        RECT 727.630 171.095 737.660 173.670 ;
        RECT 663.085 164.260 726.200 168.825 ;
      LAYER met2 ;
        RECT 726.730 168.770 727.135 168.915 ;
        RECT 726.505 168.735 726.730 168.770 ;
        RECT 726.875 168.735 727.135 168.770 ;
        RECT 726.505 168.665 727.135 168.735 ;
        RECT 726.505 168.545 726.730 168.665 ;
        RECT 726.875 168.545 727.135 168.665 ;
        RECT 726.480 168.520 726.505 168.545 ;
        RECT 726.740 168.520 726.875 168.545 ;
        RECT 726.480 168.410 726.875 168.520 ;
      LAYER met2 ;
        RECT 663.085 163.440 725.570 164.260 ;
      LAYER met2 ;
        RECT 726.480 163.980 726.740 168.410 ;
      LAYER met2 ;
        RECT 727.415 168.265 737.660 171.095 ;
        RECT 727.155 168.130 737.660 168.265 ;
      LAYER met2 ;
        RECT 725.850 163.720 726.740 163.980 ;
      LAYER met2 ;
        RECT 727.020 163.440 737.660 168.130 ;
        RECT 663.085 0.790 737.660 163.440 ;
        RECT 932.085 0.000 1011.790 208.285 ;
        RECT 1206.300 197.965 1226.905 198.000 ;
        RECT 1227.465 197.965 1260.075 198.000 ;
        RECT 1260.505 197.965 1280.500 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 1206.000 158.415 1280.500 197.965 ;
      LAYER met2 ;
        RECT 1281.260 197.725 1281.400 234.270 ;
        RECT 1485.440 221.350 1485.700 221.670 ;
        RECT 1476.240 220.670 1476.500 220.990 ;
        RECT 1476.300 210.965 1476.440 220.670 ;
        RECT 1485.500 210.965 1485.640 221.350 ;
        RECT 1488.720 210.965 1488.860 234.270 ;
        RECT 1522.700 222.030 1522.960 222.350 ;
        RECT 1531.440 222.030 1531.700 222.350 ;
        RECT 1497.860 221.350 1498.120 221.670 ;
        RECT 1497.920 210.965 1498.060 221.350 ;
        RECT 1516.260 220.670 1516.520 220.990 ;
        RECT 1516.320 210.965 1516.460 220.670 ;
        RECT 1522.760 210.965 1522.900 222.030 ;
        RECT 1528.680 221.350 1528.940 221.670 ;
        RECT 1528.740 210.965 1528.880 221.350 ;
        RECT 1531.500 220.990 1531.640 222.030 ;
        RECT 1531.440 220.670 1531.700 220.990 ;
        RECT 1547.140 210.965 1547.280 234.270 ;
        RECT 1759.600 221.690 1759.860 222.010 ;
        RECT 1750.400 220.670 1750.660 220.990 ;
        RECT 1750.460 210.965 1750.600 220.670 ;
        RECT 1759.660 210.965 1759.800 221.690 ;
        RECT 1762.880 210.965 1763.020 234.270 ;
        RECT 1772.020 221.690 1772.280 222.010 ;
        RECT 1802.840 221.690 1803.100 222.010 ;
        RECT 1772.080 210.965 1772.220 221.690 ;
        RECT 1796.860 221.010 1797.120 221.330 ;
        RECT 1790.420 220.670 1790.680 220.990 ;
        RECT 1790.480 210.965 1790.620 220.670 ;
        RECT 1796.920 210.965 1797.060 221.010 ;
        RECT 1802.900 210.965 1803.040 221.690 ;
        RECT 1821.300 210.965 1821.440 234.270 ;
        RECT 2033.760 222.030 2034.020 222.350 ;
        RECT 2033.820 221.670 2033.960 222.030 ;
        RECT 2024.550 221.155 2024.830 221.525 ;
        RECT 2033.760 221.350 2034.020 221.670 ;
        RECT 2024.620 210.965 2024.760 221.155 ;
        RECT 2033.820 210.965 2033.960 221.350 ;
        RECT 2037.040 210.965 2037.180 234.270 ;
        RECT 2064.570 221.155 2064.850 221.525 ;
        RECT 2064.640 210.965 2064.780 221.155 ;
        RECT 2071.020 220.670 2071.280 220.990 ;
        RECT 2071.080 210.965 2071.220 220.670 ;
        RECT 2095.460 210.965 2095.600 234.270 ;
        RECT 2307.460 222.030 2307.720 222.350 ;
        RECT 2298.250 221.155 2298.530 221.525 ;
        RECT 2307.520 221.330 2307.660 222.030 ;
        RECT 2298.320 210.965 2298.460 221.155 ;
        RECT 2307.460 221.010 2307.720 221.330 ;
        RECT 2307.520 210.965 2307.660 221.010 ;
        RECT 2310.740 210.965 2310.880 234.270 ;
        RECT 2344.720 222.030 2344.980 222.350 ;
        RECT 2344.780 221.670 2344.920 222.030 ;
        RECT 2338.270 221.155 2338.550 221.525 ;
        RECT 2344.720 221.350 2344.980 221.670 ;
        RECT 2338.340 210.965 2338.480 221.155 ;
        RECT 2344.780 210.965 2344.920 221.350 ;
        RECT 2369.160 210.965 2369.300 234.270 ;
        RECT 2572.410 221.155 2572.690 221.525 ;
        RECT 2572.480 210.965 2572.620 221.155 ;
        RECT 2581.620 221.010 2581.880 221.330 ;
        RECT 2581.680 210.965 2581.820 221.010 ;
        RECT 2584.900 210.965 2585.040 234.270 ;
        RECT 2618.880 227.810 2619.140 228.130 ;
        RECT 2593.580 227.470 2593.840 227.790 ;
        RECT 2593.640 221.330 2593.780 227.470 ;
        RECT 2618.940 222.350 2619.080 227.810 ;
        RECT 2612.430 221.835 2612.710 222.205 ;
        RECT 2618.880 222.030 2619.140 222.350 ;
        RECT 2593.580 221.010 2593.840 221.330 ;
        RECT 2612.500 210.965 2612.640 221.835 ;
        RECT 2618.940 210.965 2619.080 222.030 ;
        RECT 3367.360 213.850 3367.500 565.770 ;
        RECT 3367.820 547.730 3367.960 775.890 ;
        RECT 3369.660 734.730 3369.800 959.490 ;
        RECT 3370.120 791.850 3370.260 1011.510 ;
      LAYER met2 ;
        RECT 3379.435 1011.395 3588.000 1013.775 ;
        RECT 3379.715 1010.555 3588.000 1011.395 ;
        RECT 3379.435 1008.635 3588.000 1010.555 ;
        RECT 3379.715 1007.795 3588.000 1008.635 ;
        RECT 3379.435 1005.415 3588.000 1007.795 ;
        RECT 3379.715 1004.575 3588.000 1005.415 ;
        RECT 3379.435 1002.195 3588.000 1004.575 ;
        RECT 3379.715 1001.355 3588.000 1002.195 ;
        RECT 3379.435 999.435 3588.000 1001.355 ;
      LAYER met2 ;
        RECT 3377.035 999.015 3379.435 999.155 ;
        RECT 3377.020 998.875 3379.435 999.015 ;
        RECT 3377.020 996.530 3377.160 998.875 ;
      LAYER met2 ;
        RECT 3379.715 998.595 3588.000 999.435 ;
      LAYER met2 ;
        RECT 3376.960 996.210 3377.220 996.530 ;
      LAYER met2 ;
        RECT 3379.435 996.215 3588.000 998.595 ;
        RECT 3379.715 995.375 3588.000 996.215 ;
      LAYER met2 ;
        RECT 3376.560 993.070 3377.160 993.210 ;
        RECT 3376.560 952.625 3376.700 993.070 ;
        RECT 3377.020 992.715 3377.160 993.070 ;
      LAYER met2 ;
        RECT 3379.435 992.995 3588.000 995.375 ;
      LAYER met2 ;
        RECT 3377.020 992.460 3379.435 992.715 ;
        RECT 3377.035 992.435 3379.435 992.460 ;
      LAYER met2 ;
        RECT 3379.715 992.155 3588.000 992.995 ;
        RECT 3379.435 989.775 3588.000 992.155 ;
        RECT 3379.715 988.935 3588.000 989.775 ;
        RECT 3379.435 987.015 3588.000 988.935 ;
        RECT 3379.715 986.175 3588.000 987.015 ;
        RECT 3379.435 983.795 3588.000 986.175 ;
        RECT 3379.715 982.955 3588.000 983.795 ;
        RECT 3379.435 980.575 3588.000 982.955 ;
        RECT 3379.715 979.735 3588.000 980.575 ;
        RECT 3379.435 977.815 3588.000 979.735 ;
      LAYER met2 ;
        RECT 3377.035 977.255 3379.435 977.535 ;
      LAYER met2 ;
        RECT 3379.715 976.975 3588.000 977.815 ;
        RECT 3379.435 974.595 3588.000 976.975 ;
        RECT 3379.715 973.755 3588.000 974.595 ;
        RECT 3379.435 971.375 3588.000 973.755 ;
      LAYER met2 ;
        RECT 3377.035 970.815 3379.435 971.095 ;
      LAYER met2 ;
        RECT 3379.715 970.535 3588.000 971.375 ;
        RECT 3379.435 968.615 3588.000 970.535 ;
      LAYER met2 ;
        RECT 3377.035 968.055 3379.435 968.335 ;
      LAYER met2 ;
        RECT 3379.715 967.775 3588.000 968.615 ;
        RECT 3379.435 965.395 3588.000 967.775 ;
        RECT 3379.715 964.555 3588.000 965.395 ;
        RECT 3379.435 962.175 3588.000 964.555 ;
      LAYER met2 ;
        RECT 3377.035 961.860 3379.435 961.895 ;
        RECT 3377.020 961.615 3379.435 961.860 ;
        RECT 3377.020 959.810 3377.160 961.615 ;
      LAYER met2 ;
        RECT 3379.715 961.335 3588.000 962.175 ;
      LAYER met2 ;
        RECT 3376.960 959.490 3377.220 959.810 ;
      LAYER met2 ;
        RECT 3379.435 959.415 3588.000 961.335 ;
      LAYER met2 ;
        RECT 3377.035 958.855 3379.435 959.135 ;
      LAYER met2 ;
        RECT 3379.715 958.575 3588.000 959.415 ;
        RECT 3379.435 956.195 3588.000 958.575 ;
        RECT 3379.715 955.355 3588.000 956.195 ;
        RECT 3379.435 952.975 3588.000 955.355 ;
      LAYER met2 ;
        RECT 3377.035 952.625 3379.435 952.695 ;
        RECT 3376.560 952.485 3379.435 952.625 ;
        RECT 3377.035 952.415 3379.435 952.485 ;
      LAYER met2 ;
        RECT 3379.715 952.135 3588.000 952.975 ;
        RECT 3379.435 951.085 3588.000 952.135 ;
        RECT 3379.435 804.795 3588.000 805.790 ;
        RECT 3379.715 803.955 3588.000 804.795 ;
        RECT 3379.435 802.035 3588.000 803.955 ;
        RECT 3379.715 801.195 3588.000 802.035 ;
        RECT 3379.435 798.815 3588.000 801.195 ;
        RECT 3379.715 797.975 3588.000 798.815 ;
        RECT 3379.435 795.595 3588.000 797.975 ;
        RECT 3379.715 794.755 3588.000 795.595 ;
        RECT 3379.435 792.835 3588.000 794.755 ;
        RECT 3379.715 791.995 3588.000 792.835 ;
      LAYER met2 ;
        RECT 3370.060 791.530 3370.320 791.850 ;
        RECT 3376.960 791.530 3377.220 791.850 ;
        RECT 3377.020 789.335 3377.160 791.530 ;
      LAYER met2 ;
        RECT 3379.435 789.615 3588.000 791.995 ;
      LAYER met2 ;
        RECT 3377.020 789.140 3379.435 789.335 ;
        RECT 3377.035 789.055 3379.435 789.140 ;
      LAYER met2 ;
        RECT 3379.715 788.775 3588.000 789.615 ;
        RECT 3379.435 786.395 3588.000 788.775 ;
        RECT 3379.715 785.555 3588.000 786.395 ;
        RECT 3379.435 783.635 3588.000 785.555 ;
        RECT 3379.715 782.795 3588.000 783.635 ;
        RECT 3379.435 780.415 3588.000 782.795 ;
        RECT 3379.715 779.575 3588.000 780.415 ;
        RECT 3379.435 777.195 3588.000 779.575 ;
        RECT 3379.715 776.355 3588.000 777.195 ;
      LAYER met2 ;
        RECT 3376.960 775.890 3377.220 776.210 ;
        RECT 3377.020 774.155 3377.160 775.890 ;
      LAYER met2 ;
        RECT 3379.435 774.435 3588.000 776.355 ;
      LAYER met2 ;
        RECT 3377.020 774.015 3379.435 774.155 ;
        RECT 3377.035 773.875 3379.435 774.015 ;
      LAYER met2 ;
        RECT 3379.715 773.595 3588.000 774.435 ;
        RECT 3379.435 771.215 3588.000 773.595 ;
        RECT 3379.715 770.375 3588.000 771.215 ;
        RECT 3379.435 767.995 3588.000 770.375 ;
      LAYER met2 ;
        RECT 3377.035 767.645 3379.435 767.715 ;
        RECT 3376.560 767.505 3379.435 767.645 ;
        RECT 3368.680 734.410 3368.940 734.730 ;
        RECT 3369.600 734.410 3369.860 734.730 ;
        RECT 3367.760 547.410 3368.020 547.730 ;
        RECT 3367.820 228.130 3367.960 547.410 ;
        RECT 3368.740 508.630 3368.880 734.410 ;
        RECT 3376.560 727.625 3376.700 767.505 ;
        RECT 3377.035 767.435 3379.435 767.505 ;
      LAYER met2 ;
        RECT 3379.715 767.155 3588.000 767.995 ;
        RECT 3379.435 764.775 3588.000 767.155 ;
        RECT 3379.715 763.935 3588.000 764.775 ;
        RECT 3379.435 762.015 3588.000 763.935 ;
        RECT 3379.715 761.175 3588.000 762.015 ;
        RECT 3379.435 758.795 3588.000 761.175 ;
        RECT 3379.715 757.955 3588.000 758.795 ;
        RECT 3379.435 755.575 3588.000 757.955 ;
        RECT 3379.715 754.735 3588.000 755.575 ;
        RECT 3379.435 752.815 3588.000 754.735 ;
      LAYER met2 ;
        RECT 3377.035 752.255 3379.435 752.535 ;
      LAYER met2 ;
        RECT 3379.715 751.975 3588.000 752.815 ;
        RECT 3379.435 749.595 3588.000 751.975 ;
        RECT 3379.715 748.755 3588.000 749.595 ;
        RECT 3379.435 746.375 3588.000 748.755 ;
      LAYER met2 ;
        RECT 3377.035 745.815 3379.435 746.095 ;
      LAYER met2 ;
        RECT 3379.715 745.535 3588.000 746.375 ;
        RECT 3379.435 743.615 3588.000 745.535 ;
      LAYER met2 ;
        RECT 3377.035 743.055 3379.435 743.335 ;
      LAYER met2 ;
        RECT 3379.715 742.775 3588.000 743.615 ;
        RECT 3379.435 740.395 3588.000 742.775 ;
        RECT 3379.715 739.555 3588.000 740.395 ;
        RECT 3379.435 737.175 3588.000 739.555 ;
      LAYER met2 ;
        RECT 3377.035 736.780 3379.435 736.895 ;
        RECT 3377.020 736.615 3379.435 736.780 ;
        RECT 3377.020 734.730 3377.160 736.615 ;
      LAYER met2 ;
        RECT 3379.715 736.335 3588.000 737.175 ;
      LAYER met2 ;
        RECT 3376.960 734.410 3377.220 734.730 ;
      LAYER met2 ;
        RECT 3379.435 734.415 3588.000 736.335 ;
      LAYER met2 ;
        RECT 3377.035 733.855 3379.435 734.135 ;
      LAYER met2 ;
        RECT 3379.715 733.575 3588.000 734.415 ;
        RECT 3379.435 731.195 3588.000 733.575 ;
        RECT 3379.715 730.355 3588.000 731.195 ;
        RECT 3379.435 727.975 3588.000 730.355 ;
      LAYER met2 ;
        RECT 3377.035 727.625 3379.435 727.695 ;
        RECT 3376.560 727.485 3379.435 727.625 ;
        RECT 3377.035 727.415 3379.435 727.485 ;
      LAYER met2 ;
        RECT 3379.715 727.135 3588.000 727.975 ;
        RECT 3379.435 726.085 3588.000 727.135 ;
        RECT 3379.435 578.795 3588.000 579.790 ;
        RECT 3379.715 577.955 3588.000 578.795 ;
        RECT 3379.435 576.035 3588.000 577.955 ;
        RECT 3379.715 575.195 3588.000 576.035 ;
        RECT 3379.435 572.815 3588.000 575.195 ;
        RECT 3379.715 571.975 3588.000 572.815 ;
        RECT 3379.435 569.595 3588.000 571.975 ;
        RECT 3379.715 568.755 3588.000 569.595 ;
        RECT 3379.435 566.835 3588.000 568.755 ;
      LAYER met2 ;
        RECT 3376.960 565.770 3377.220 566.090 ;
      LAYER met2 ;
        RECT 3379.715 565.995 3588.000 566.835 ;
      LAYER met2 ;
        RECT 3377.020 563.335 3377.160 565.770 ;
      LAYER met2 ;
        RECT 3379.435 563.615 3588.000 565.995 ;
      LAYER met2 ;
        RECT 3377.020 563.195 3379.435 563.335 ;
        RECT 3377.035 563.055 3379.435 563.195 ;
      LAYER met2 ;
        RECT 3379.715 562.775 3588.000 563.615 ;
        RECT 3379.435 560.395 3588.000 562.775 ;
        RECT 3379.715 559.555 3588.000 560.395 ;
        RECT 3379.435 557.635 3588.000 559.555 ;
        RECT 3379.715 556.795 3588.000 557.635 ;
        RECT 3379.435 554.415 3588.000 556.795 ;
        RECT 3379.715 553.575 3588.000 554.415 ;
        RECT 3379.435 551.195 3588.000 553.575 ;
        RECT 3379.715 550.355 3588.000 551.195 ;
        RECT 3379.435 548.435 3588.000 550.355 ;
      LAYER met2 ;
        RECT 3377.035 548.015 3379.435 548.155 ;
        RECT 3377.020 547.875 3379.435 548.015 ;
        RECT 3377.020 547.730 3377.160 547.875 ;
        RECT 3376.960 547.410 3377.220 547.730 ;
      LAYER met2 ;
        RECT 3379.715 547.595 3588.000 548.435 ;
        RECT 3379.435 545.215 3588.000 547.595 ;
        RECT 3379.715 544.375 3588.000 545.215 ;
        RECT 3379.435 541.995 3588.000 544.375 ;
      LAYER met2 ;
        RECT 3377.035 541.690 3379.435 541.715 ;
        RECT 3376.560 541.550 3379.435 541.690 ;
        RECT 3368.680 508.310 3368.940 508.630 ;
        RECT 3367.760 227.810 3368.020 228.130 ;
        RECT 3368.740 227.790 3368.880 508.310 ;
        RECT 3376.560 501.570 3376.700 541.550 ;
        RECT 3377.035 541.435 3379.435 541.550 ;
      LAYER met2 ;
        RECT 3379.715 541.155 3588.000 541.995 ;
        RECT 3379.435 538.775 3588.000 541.155 ;
        RECT 3379.715 537.935 3588.000 538.775 ;
        RECT 3379.435 536.015 3588.000 537.935 ;
        RECT 3379.715 535.175 3588.000 536.015 ;
        RECT 3379.435 532.795 3588.000 535.175 ;
        RECT 3379.715 531.955 3588.000 532.795 ;
        RECT 3379.435 529.575 3588.000 531.955 ;
        RECT 3379.715 528.735 3588.000 529.575 ;
        RECT 3379.435 526.815 3588.000 528.735 ;
      LAYER met2 ;
        RECT 3377.035 526.255 3379.435 526.535 ;
      LAYER met2 ;
        RECT 3379.715 525.975 3588.000 526.815 ;
        RECT 3379.435 523.595 3588.000 525.975 ;
        RECT 3379.715 522.755 3588.000 523.595 ;
        RECT 3379.435 520.375 3588.000 522.755 ;
      LAYER met2 ;
        RECT 3377.035 519.815 3379.435 520.095 ;
      LAYER met2 ;
        RECT 3379.715 519.535 3588.000 520.375 ;
        RECT 3379.435 517.615 3588.000 519.535 ;
      LAYER met2 ;
        RECT 3377.035 517.055 3379.435 517.335 ;
      LAYER met2 ;
        RECT 3379.715 516.775 3588.000 517.615 ;
        RECT 3379.435 514.395 3588.000 516.775 ;
        RECT 3379.715 513.555 3588.000 514.395 ;
        RECT 3379.435 511.175 3588.000 513.555 ;
      LAYER met2 ;
        RECT 3377.035 510.755 3379.435 510.895 ;
        RECT 3377.020 510.615 3379.435 510.755 ;
        RECT 3377.020 508.630 3377.160 510.615 ;
      LAYER met2 ;
        RECT 3379.715 510.335 3588.000 511.175 ;
      LAYER met2 ;
        RECT 3376.960 508.310 3377.220 508.630 ;
      LAYER met2 ;
        RECT 3379.435 508.415 3588.000 510.335 ;
      LAYER met2 ;
        RECT 3377.035 507.855 3379.435 508.135 ;
      LAYER met2 ;
        RECT 3379.715 507.575 3588.000 508.415 ;
        RECT 3379.435 505.195 3588.000 507.575 ;
        RECT 3379.715 504.355 3588.000 505.195 ;
        RECT 3379.435 501.975 3588.000 504.355 ;
      LAYER met2 ;
        RECT 3377.035 501.570 3379.435 501.695 ;
        RECT 3376.560 501.430 3379.435 501.570 ;
        RECT 3377.035 501.415 3379.435 501.430 ;
      LAYER met2 ;
        RECT 3379.715 501.135 3588.000 501.975 ;
        RECT 3379.435 500.085 3588.000 501.135 ;
      LAYER met2 ;
        RECT 3368.680 227.470 3368.940 227.790 ;
        RECT 2899.480 213.530 2899.740 213.850 ;
        RECT 3367.300 213.530 3367.560 213.850 ;
        RECT 1476.300 209.030 1476.695 210.965 ;
        RECT 1476.415 208.565 1476.695 209.030 ;
        RECT 1479.635 208.565 1479.915 210.965 ;
        RECT 1482.855 208.565 1483.135 210.965 ;
        RECT 1485.500 209.030 1485.895 210.965 ;
        RECT 1488.720 209.170 1489.115 210.965 ;
        RECT 1489.580 209.450 1489.840 209.770 ;
        RECT 1489.640 209.170 1489.780 209.450 ;
        RECT 1488.720 209.030 1489.780 209.170 ;
        RECT 1485.615 208.565 1485.895 209.030 ;
        RECT 1488.835 208.565 1489.115 209.030 ;
        RECT 1492.055 208.565 1492.335 210.965 ;
        RECT 1494.815 208.565 1495.095 210.965 ;
        RECT 1497.920 209.030 1498.315 210.965 ;
        RECT 1498.035 208.565 1498.315 209.030 ;
        RECT 1501.255 208.565 1501.535 210.965 ;
        RECT 1503.380 209.450 1503.640 209.770 ;
        RECT 1503.440 209.170 1503.580 209.450 ;
        RECT 1504.015 209.170 1504.295 210.965 ;
        RECT 1507.235 209.170 1507.515 210.965 ;
        RECT 1510.455 209.170 1510.735 210.965 ;
        RECT 1511.200 209.450 1511.460 209.770 ;
        RECT 1511.260 209.170 1511.400 209.450 ;
        RECT 1503.440 209.030 1511.400 209.170 ;
        RECT 1516.320 209.030 1516.715 210.965 ;
        RECT 1522.760 209.030 1523.155 210.965 ;
        RECT 1504.015 208.565 1504.295 209.030 ;
        RECT 1507.235 208.565 1507.515 209.030 ;
        RECT 1510.455 208.565 1510.735 209.030 ;
        RECT 1516.435 208.565 1516.715 209.030 ;
        RECT 1522.875 208.565 1523.155 209.030 ;
        RECT 1525.635 209.170 1525.915 210.965 ;
        RECT 1526.380 209.450 1526.640 209.770 ;
        RECT 1526.440 209.170 1526.580 209.450 ;
        RECT 1525.635 209.030 1526.580 209.170 ;
        RECT 1528.740 209.030 1529.135 210.965 ;
        RECT 1525.635 208.565 1525.915 209.030 ;
        RECT 1528.855 208.565 1529.135 209.030 ;
        RECT 1532.075 209.170 1532.355 210.965 ;
        RECT 1532.820 209.450 1533.080 209.770 ;
        RECT 1532.880 209.170 1533.020 209.450 ;
        RECT 1532.075 209.030 1533.020 209.170 ;
        RECT 1538.055 209.170 1538.335 210.965 ;
        RECT 1543.400 209.450 1543.660 209.770 ;
        RECT 1543.460 209.170 1543.600 209.450 ;
        RECT 1544.035 209.170 1544.315 210.965 ;
        RECT 1547.140 209.170 1547.535 210.965 ;
        RECT 1538.055 209.090 1539.000 209.170 ;
        RECT 1538.055 209.030 1539.060 209.090 ;
        RECT 1543.460 209.030 1547.535 209.170 ;
        RECT 1532.075 208.565 1532.355 209.030 ;
        RECT 1538.055 208.565 1538.335 209.030 ;
        RECT 1538.800 208.770 1539.060 209.030 ;
        RECT 1544.035 208.565 1544.315 209.030 ;
        RECT 1547.255 208.565 1547.535 209.030 ;
        RECT 1553.235 208.565 1553.515 210.965 ;
        RECT 1750.415 208.565 1750.695 210.965 ;
        RECT 1753.635 208.565 1753.915 210.965 ;
        RECT 1756.855 208.565 1757.135 210.965 ;
        RECT 1759.615 208.565 1759.895 210.965 ;
        RECT 1762.835 209.850 1763.115 210.965 ;
        RECT 1762.835 209.770 1763.480 209.850 ;
        RECT 1762.835 209.710 1763.540 209.770 ;
        RECT 1762.835 208.565 1763.115 209.710 ;
        RECT 1763.280 209.450 1763.540 209.710 ;
        RECT 1766.055 208.565 1766.335 210.965 ;
        RECT 1768.815 208.565 1769.095 210.965 ;
        RECT 1772.035 208.565 1772.315 210.965 ;
        RECT 1775.255 208.565 1775.535 210.965 ;
        RECT 1777.540 209.450 1777.800 209.770 ;
        RECT 1777.600 209.170 1777.740 209.450 ;
        RECT 1778.015 209.170 1778.295 210.965 ;
        RECT 1781.235 209.170 1781.515 210.965 ;
        RECT 1784.455 209.170 1784.735 210.965 ;
        RECT 1784.900 209.450 1785.160 209.770 ;
        RECT 1784.960 209.170 1785.100 209.450 ;
        RECT 1777.600 209.030 1785.100 209.170 ;
        RECT 1778.015 208.565 1778.295 209.030 ;
        RECT 1781.235 208.565 1781.515 209.030 ;
        RECT 1784.455 208.565 1784.735 209.030 ;
        RECT 1790.435 208.565 1790.715 210.965 ;
        RECT 1796.875 208.565 1797.155 210.965 ;
        RECT 1799.160 209.450 1799.420 209.770 ;
        RECT 1799.220 209.170 1799.360 209.450 ;
        RECT 1799.635 209.170 1799.915 210.965 ;
        RECT 1799.220 209.030 1799.915 209.170 ;
        RECT 1799.635 208.565 1799.915 209.030 ;
        RECT 1802.855 208.565 1803.135 210.965 ;
        RECT 1805.600 209.450 1805.860 209.770 ;
        RECT 1805.660 209.170 1805.800 209.450 ;
        RECT 1806.075 209.170 1806.355 210.965 ;
        RECT 1805.660 209.030 1806.355 209.170 ;
        RECT 1806.075 208.565 1806.355 209.030 ;
        RECT 1812.055 209.170 1812.335 210.965 ;
        RECT 1817.560 209.450 1817.820 209.770 ;
        RECT 1817.620 209.170 1817.760 209.450 ;
        RECT 1818.035 209.170 1818.315 210.965 ;
        RECT 1821.255 209.170 1821.535 210.965 ;
        RECT 1812.055 209.090 1812.700 209.170 ;
        RECT 1812.055 209.030 1812.760 209.090 ;
        RECT 1817.620 209.030 1821.535 209.170 ;
        RECT 1812.055 208.565 1812.335 209.030 ;
        RECT 1812.500 208.770 1812.760 209.030 ;
        RECT 1818.035 208.565 1818.315 209.030 ;
        RECT 1821.255 208.565 1821.535 209.030 ;
        RECT 1827.235 208.565 1827.515 210.965 ;
        RECT 2024.415 209.100 2024.760 210.965 ;
        RECT 2024.415 208.565 2024.695 209.100 ;
        RECT 2030.855 208.565 2031.135 210.965 ;
        RECT 2033.615 209.100 2033.960 210.965 ;
        RECT 2036.835 209.850 2037.180 210.965 ;
        RECT 2036.835 209.770 2037.640 209.850 ;
        RECT 2036.835 209.710 2037.700 209.770 ;
        RECT 2036.835 209.100 2037.180 209.710 ;
        RECT 2037.440 209.450 2037.700 209.710 ;
        RECT 2033.615 208.565 2033.895 209.100 ;
        RECT 2036.835 208.565 2037.115 209.100 ;
        RECT 2040.055 208.565 2040.335 210.965 ;
        RECT 2042.815 208.565 2043.095 210.965 ;
        RECT 2049.255 208.565 2049.535 210.965 ;
        RECT 2051.240 209.450 2051.500 209.770 ;
        RECT 2051.300 209.170 2051.440 209.450 ;
        RECT 2052.015 209.170 2052.295 210.965 ;
        RECT 2057.680 209.450 2057.940 209.770 ;
        RECT 2051.300 209.030 2052.295 209.170 ;
        RECT 2057.740 209.170 2057.880 209.450 ;
        RECT 2058.455 209.170 2058.735 210.965 ;
        RECT 2057.740 209.030 2058.735 209.170 ;
        RECT 2052.015 208.565 2052.295 209.030 ;
        RECT 2058.455 208.565 2058.735 209.030 ;
        RECT 2064.435 209.100 2064.780 210.965 ;
        RECT 2070.875 209.100 2071.220 210.965 ;
        RECT 2072.860 209.450 2073.120 209.770 ;
        RECT 2072.920 209.170 2073.060 209.450 ;
        RECT 2073.635 209.170 2073.915 210.965 ;
        RECT 2079.300 209.450 2079.560 209.770 ;
        RECT 2064.435 208.565 2064.715 209.100 ;
        RECT 2070.875 208.565 2071.155 209.100 ;
        RECT 2072.920 209.030 2073.915 209.170 ;
        RECT 2079.360 209.170 2079.500 209.450 ;
        RECT 2080.075 209.170 2080.355 210.965 ;
        RECT 2079.360 209.030 2080.355 209.170 ;
        RECT 2073.635 208.565 2073.915 209.030 ;
        RECT 2080.075 208.565 2080.355 209.030 ;
        RECT 2086.055 209.170 2086.335 210.965 ;
        RECT 2091.260 209.450 2091.520 209.770 ;
        RECT 2091.320 209.170 2091.460 209.450 ;
        RECT 2092.035 209.170 2092.315 210.965 ;
        RECT 2095.255 209.170 2095.600 210.965 ;
        RECT 2086.055 209.090 2086.860 209.170 ;
        RECT 2091.320 209.100 2095.600 209.170 ;
        RECT 2086.055 209.030 2086.920 209.090 ;
        RECT 2091.320 209.030 2095.535 209.100 ;
        RECT 2086.055 208.565 2086.335 209.030 ;
        RECT 2086.660 208.770 2086.920 209.030 ;
        RECT 2092.035 208.565 2092.315 209.030 ;
        RECT 2095.255 208.565 2095.535 209.030 ;
        RECT 2101.235 208.565 2101.515 210.965 ;
        RECT 2298.320 209.030 2298.695 210.965 ;
        RECT 2298.415 208.565 2298.695 209.030 ;
        RECT 2304.855 208.565 2305.135 210.965 ;
        RECT 2307.520 209.030 2307.895 210.965 ;
        RECT 2310.740 209.170 2311.115 210.965 ;
        RECT 2311.600 209.450 2311.860 209.770 ;
        RECT 2311.660 209.170 2311.800 209.450 ;
        RECT 2310.740 209.030 2311.800 209.170 ;
        RECT 2307.615 208.565 2307.895 209.030 ;
        RECT 2310.835 208.565 2311.115 209.030 ;
        RECT 2314.055 208.565 2314.335 210.965 ;
        RECT 2316.815 208.565 2317.095 210.965 ;
        RECT 2323.255 208.565 2323.535 210.965 ;
        RECT 2325.400 209.450 2325.660 209.770 ;
        RECT 2325.460 209.170 2325.600 209.450 ;
        RECT 2326.015 209.170 2326.295 210.965 ;
        RECT 2331.840 209.450 2332.100 209.770 ;
        RECT 2325.460 209.030 2326.295 209.170 ;
        RECT 2331.900 209.170 2332.040 209.450 ;
        RECT 2332.455 209.170 2332.735 210.965 ;
        RECT 2331.900 209.030 2332.735 209.170 ;
        RECT 2338.340 209.030 2338.715 210.965 ;
        RECT 2344.780 209.030 2345.155 210.965 ;
        RECT 2347.020 209.450 2347.280 209.770 ;
        RECT 2347.080 209.170 2347.220 209.450 ;
        RECT 2347.635 209.170 2347.915 210.965 ;
        RECT 2353.460 209.450 2353.720 209.770 ;
        RECT 2347.080 209.030 2347.915 209.170 ;
        RECT 2353.520 209.170 2353.660 209.450 ;
        RECT 2354.075 209.170 2354.355 210.965 ;
        RECT 2353.520 209.030 2354.355 209.170 ;
        RECT 2326.015 208.565 2326.295 209.030 ;
        RECT 2332.455 208.565 2332.735 209.030 ;
        RECT 2338.435 208.565 2338.715 209.030 ;
        RECT 2344.875 208.565 2345.155 209.030 ;
        RECT 2347.635 208.565 2347.915 209.030 ;
        RECT 2354.075 208.565 2354.355 209.030 ;
        RECT 2360.055 209.170 2360.335 210.965 ;
        RECT 2365.420 209.450 2365.680 209.770 ;
        RECT 2365.480 209.170 2365.620 209.450 ;
        RECT 2366.035 209.170 2366.315 210.965 ;
        RECT 2369.160 209.170 2369.535 210.965 ;
        RECT 2360.055 209.090 2361.020 209.170 ;
        RECT 2360.055 209.030 2361.080 209.090 ;
        RECT 2365.480 209.030 2369.535 209.170 ;
        RECT 2360.055 208.565 2360.335 209.030 ;
        RECT 2360.820 208.770 2361.080 209.030 ;
        RECT 2366.035 208.565 2366.315 209.030 ;
        RECT 2369.255 208.565 2369.535 209.030 ;
        RECT 2375.235 208.565 2375.515 210.965 ;
        RECT 2572.415 208.565 2572.695 210.965 ;
        RECT 2578.855 208.565 2579.135 210.965 ;
        RECT 2581.615 208.565 2581.895 210.965 ;
        RECT 2584.835 209.850 2585.115 210.965 ;
        RECT 2584.835 209.770 2585.500 209.850 ;
        RECT 2584.835 209.710 2585.560 209.770 ;
        RECT 2584.835 208.565 2585.115 209.710 ;
        RECT 2585.300 209.450 2585.560 209.710 ;
        RECT 2588.055 208.565 2588.335 210.965 ;
        RECT 2590.815 208.565 2591.095 210.965 ;
        RECT 2597.255 208.565 2597.535 210.965 ;
        RECT 2599.560 209.450 2599.820 209.770 ;
        RECT 2599.620 209.170 2599.760 209.450 ;
        RECT 2600.015 209.170 2600.295 210.965 ;
        RECT 2606.000 209.450 2606.260 209.770 ;
        RECT 2599.620 209.030 2600.295 209.170 ;
        RECT 2606.060 209.170 2606.200 209.450 ;
        RECT 2606.455 209.170 2606.735 210.965 ;
        RECT 2606.060 209.030 2606.735 209.170 ;
        RECT 2600.015 208.565 2600.295 209.030 ;
        RECT 2606.455 208.565 2606.735 209.030 ;
        RECT 2612.435 208.565 2612.715 210.965 ;
        RECT 2618.875 208.565 2619.155 210.965 ;
        RECT 2621.180 209.450 2621.440 209.770 ;
        RECT 2621.240 209.170 2621.380 209.450 ;
        RECT 2621.635 209.170 2621.915 210.965 ;
        RECT 2627.620 209.450 2627.880 209.770 ;
        RECT 2621.240 209.030 2621.915 209.170 ;
        RECT 2627.680 209.170 2627.820 209.450 ;
        RECT 2628.075 209.170 2628.355 210.965 ;
        RECT 2634.055 209.170 2634.335 210.965 ;
        RECT 2639.580 209.450 2639.840 209.770 ;
        RECT 2627.680 209.030 2628.355 209.170 ;
        RECT 2633.660 209.090 2634.335 209.170 ;
        RECT 2621.635 208.565 2621.915 209.030 ;
        RECT 2628.075 208.565 2628.355 209.030 ;
        RECT 2633.600 209.030 2634.335 209.090 ;
        RECT 2639.640 209.170 2639.780 209.450 ;
        RECT 2640.035 209.170 2640.315 210.965 ;
        RECT 2643.255 209.170 2643.535 210.965 ;
        RECT 2639.640 209.030 2643.535 209.170 ;
        RECT 2633.600 208.770 2633.860 209.030 ;
        RECT 2634.055 208.565 2634.335 209.030 ;
        RECT 2640.035 208.565 2640.315 209.030 ;
        RECT 2643.255 208.565 2643.535 209.030 ;
        RECT 2649.235 208.565 2649.515 210.965 ;
        RECT 2899.540 209.430 2899.680 213.530 ;
        RECT 2844.280 209.110 2844.540 209.430 ;
        RECT 2899.480 209.110 2899.740 209.430 ;
      LAYER met2 ;
        RECT 1475.085 208.285 1476.135 208.565 ;
        RECT 1476.975 208.285 1479.355 208.565 ;
        RECT 1480.195 208.285 1482.575 208.565 ;
        RECT 1483.415 208.285 1485.335 208.565 ;
        RECT 1486.175 208.285 1488.555 208.565 ;
        RECT 1489.395 208.285 1491.775 208.565 ;
        RECT 1492.615 208.285 1494.535 208.565 ;
        RECT 1495.375 208.285 1497.755 208.565 ;
        RECT 1498.595 208.285 1500.975 208.565 ;
        RECT 1501.815 208.285 1503.735 208.565 ;
        RECT 1504.575 208.285 1506.955 208.565 ;
        RECT 1507.795 208.285 1510.175 208.565 ;
        RECT 1511.015 208.285 1512.935 208.565 ;
        RECT 1513.775 208.285 1516.155 208.565 ;
        RECT 1516.995 208.285 1519.375 208.565 ;
        RECT 1520.215 208.285 1522.595 208.565 ;
        RECT 1523.435 208.285 1525.355 208.565 ;
        RECT 1526.195 208.285 1528.575 208.565 ;
        RECT 1529.415 208.285 1531.795 208.565 ;
        RECT 1532.635 208.285 1534.555 208.565 ;
        RECT 1535.395 208.285 1537.775 208.565 ;
        RECT 1538.615 208.285 1540.995 208.565 ;
        RECT 1541.835 208.285 1543.755 208.565 ;
        RECT 1544.595 208.285 1546.975 208.565 ;
        RECT 1547.815 208.285 1550.195 208.565 ;
        RECT 1551.035 208.285 1552.955 208.565 ;
        RECT 1553.795 208.285 1554.790 208.565 ;
      LAYER met2 ;
        RECT 1281.190 197.355 1281.470 197.725 ;
      LAYER met2 ;
        RECT 1194.860 153.765 1280.500 158.415 ;
        RECT 1206.000 3.570 1280.500 153.765 ;
        RECT 1475.085 0.000 1554.790 208.285 ;
        RECT 1749.085 208.285 1750.135 208.565 ;
        RECT 1750.975 208.285 1753.355 208.565 ;
        RECT 1754.195 208.285 1756.575 208.565 ;
        RECT 1757.415 208.285 1759.335 208.565 ;
        RECT 1760.175 208.285 1762.555 208.565 ;
        RECT 1763.395 208.285 1765.775 208.565 ;
        RECT 1766.615 208.285 1768.535 208.565 ;
        RECT 1769.375 208.285 1771.755 208.565 ;
        RECT 1772.595 208.285 1774.975 208.565 ;
        RECT 1775.815 208.285 1777.735 208.565 ;
        RECT 1778.575 208.285 1780.955 208.565 ;
        RECT 1781.795 208.285 1784.175 208.565 ;
        RECT 1785.015 208.285 1786.935 208.565 ;
        RECT 1787.775 208.285 1790.155 208.565 ;
        RECT 1790.995 208.285 1793.375 208.565 ;
        RECT 1794.215 208.285 1796.595 208.565 ;
        RECT 1797.435 208.285 1799.355 208.565 ;
        RECT 1800.195 208.285 1802.575 208.565 ;
        RECT 1803.415 208.285 1805.795 208.565 ;
        RECT 1806.635 208.285 1808.555 208.565 ;
        RECT 1809.395 208.285 1811.775 208.565 ;
        RECT 1812.615 208.285 1814.995 208.565 ;
        RECT 1815.835 208.285 1817.755 208.565 ;
        RECT 1818.595 208.285 1820.975 208.565 ;
        RECT 1821.815 208.285 1824.195 208.565 ;
        RECT 1825.035 208.285 1826.955 208.565 ;
        RECT 1827.795 208.285 1828.790 208.565 ;
        RECT 1749.085 0.000 1828.790 208.285 ;
        RECT 2023.085 208.285 2024.135 208.565 ;
        RECT 2024.975 208.285 2027.355 208.565 ;
        RECT 2028.195 208.285 2030.575 208.565 ;
        RECT 2031.415 208.285 2033.335 208.565 ;
        RECT 2034.175 208.285 2036.555 208.565 ;
        RECT 2037.395 208.285 2039.775 208.565 ;
        RECT 2040.615 208.285 2042.535 208.565 ;
        RECT 2043.375 208.285 2045.755 208.565 ;
        RECT 2046.595 208.285 2048.975 208.565 ;
        RECT 2049.815 208.285 2051.735 208.565 ;
        RECT 2052.575 208.285 2054.955 208.565 ;
        RECT 2055.795 208.285 2058.175 208.565 ;
        RECT 2059.015 208.285 2060.935 208.565 ;
        RECT 2061.775 208.285 2064.155 208.565 ;
        RECT 2064.995 208.285 2067.375 208.565 ;
        RECT 2068.215 208.285 2070.595 208.565 ;
        RECT 2071.435 208.285 2073.355 208.565 ;
        RECT 2074.195 208.285 2076.575 208.565 ;
        RECT 2077.415 208.285 2079.795 208.565 ;
        RECT 2080.635 208.285 2082.555 208.565 ;
        RECT 2083.395 208.285 2085.775 208.565 ;
        RECT 2086.615 208.285 2088.995 208.565 ;
        RECT 2089.835 208.285 2091.755 208.565 ;
        RECT 2092.595 208.285 2094.975 208.565 ;
        RECT 2095.815 208.285 2098.195 208.565 ;
        RECT 2099.035 208.285 2100.955 208.565 ;
        RECT 2101.795 208.285 2102.790 208.565 ;
        RECT 2023.085 0.000 2102.790 208.285 ;
        RECT 2297.085 208.285 2298.135 208.565 ;
        RECT 2298.975 208.285 2301.355 208.565 ;
        RECT 2302.195 208.285 2304.575 208.565 ;
        RECT 2305.415 208.285 2307.335 208.565 ;
        RECT 2308.175 208.285 2310.555 208.565 ;
        RECT 2311.395 208.285 2313.775 208.565 ;
        RECT 2314.615 208.285 2316.535 208.565 ;
        RECT 2317.375 208.285 2319.755 208.565 ;
        RECT 2320.595 208.285 2322.975 208.565 ;
        RECT 2323.815 208.285 2325.735 208.565 ;
        RECT 2326.575 208.285 2328.955 208.565 ;
        RECT 2329.795 208.285 2332.175 208.565 ;
        RECT 2333.015 208.285 2334.935 208.565 ;
        RECT 2335.775 208.285 2338.155 208.565 ;
        RECT 2338.995 208.285 2341.375 208.565 ;
        RECT 2342.215 208.285 2344.595 208.565 ;
        RECT 2345.435 208.285 2347.355 208.565 ;
        RECT 2348.195 208.285 2350.575 208.565 ;
        RECT 2351.415 208.285 2353.795 208.565 ;
        RECT 2354.635 208.285 2356.555 208.565 ;
        RECT 2357.395 208.285 2359.775 208.565 ;
        RECT 2360.615 208.285 2362.995 208.565 ;
        RECT 2363.835 208.285 2365.755 208.565 ;
        RECT 2366.595 208.285 2368.975 208.565 ;
        RECT 2369.815 208.285 2372.195 208.565 ;
        RECT 2373.035 208.285 2374.955 208.565 ;
        RECT 2375.795 208.285 2376.790 208.565 ;
        RECT 2297.085 0.000 2376.790 208.285 ;
        RECT 2571.085 208.285 2572.135 208.565 ;
        RECT 2572.975 208.285 2575.355 208.565 ;
        RECT 2576.195 208.285 2578.575 208.565 ;
        RECT 2579.415 208.285 2581.335 208.565 ;
        RECT 2582.175 208.285 2584.555 208.565 ;
        RECT 2585.395 208.285 2587.775 208.565 ;
        RECT 2588.615 208.285 2590.535 208.565 ;
        RECT 2591.375 208.285 2593.755 208.565 ;
        RECT 2594.595 208.285 2596.975 208.565 ;
        RECT 2597.815 208.285 2599.735 208.565 ;
        RECT 2600.575 208.285 2602.955 208.565 ;
        RECT 2603.795 208.285 2606.175 208.565 ;
        RECT 2607.015 208.285 2608.935 208.565 ;
        RECT 2609.775 208.285 2612.155 208.565 ;
        RECT 2612.995 208.285 2615.375 208.565 ;
        RECT 2616.215 208.285 2618.595 208.565 ;
        RECT 2619.435 208.285 2621.355 208.565 ;
        RECT 2622.195 208.285 2624.575 208.565 ;
        RECT 2625.415 208.285 2627.795 208.565 ;
        RECT 2628.635 208.285 2630.555 208.565 ;
        RECT 2631.395 208.285 2633.775 208.565 ;
        RECT 2634.615 208.285 2636.995 208.565 ;
        RECT 2637.835 208.285 2639.755 208.565 ;
        RECT 2640.595 208.285 2642.975 208.565 ;
        RECT 2643.815 208.285 2646.195 208.565 ;
        RECT 2647.035 208.285 2648.955 208.565 ;
        RECT 2649.795 208.285 2650.790 208.565 ;
        RECT 2571.085 0.000 2650.790 208.285 ;
      LAYER met2 ;
        RECT 2844.340 198.405 2844.480 209.110 ;
        RECT 2844.270 198.035 2844.550 198.405 ;
      LAYER met2 ;
        RECT 2845.710 197.965 2869.610 200.000 ;
        RECT 2892.105 198.080 2894.105 200.000 ;
        RECT 2895.605 197.965 2919.505 200.000 ;
        RECT 3114.710 197.965 3138.610 200.000 ;
        RECT 3161.105 198.080 3163.105 200.000 ;
        RECT 3164.605 197.965 3188.505 200.000 ;
        RECT 2845.710 4.925 2919.735 197.965 ;
        RECT 3114.710 4.925 3188.735 197.965 ;
      LAYER via2 ;
        RECT 2925.230 4987.320 2925.510 4987.600 ;
        RECT 1718.190 4985.280 1718.470 4985.560 ;
        RECT 211.690 4350.160 211.970 4350.440 ;
        RECT 224.110 4350.160 224.390 4350.440 ;
        RECT 3387.990 4091.760 3388.270 4092.040 ;
        RECT 3388.450 2568.560 3388.730 2568.840 ;
        RECT 3387.530 2127.920 3387.810 2128.200 ;
        RECT 220.890 552.360 221.170 552.640 ;
        RECT 224.110 552.360 224.390 552.640 ;
        RECT 220.890 359.240 221.170 359.520 ;
        RECT 224.110 359.240 224.390 359.520 ;
        RECT 468.830 200.800 469.110 201.080 ;
        RECT 675.830 200.800 676.110 201.080 ;
        RECT 715.390 200.800 715.670 201.080 ;
        RECT 717.690 200.800 717.970 201.080 ;
        RECT 745.290 201.480 745.570 201.760 ;
        RECT 2024.550 221.200 2024.830 221.480 ;
        RECT 2064.570 221.200 2064.850 221.480 ;
        RECT 2298.250 221.200 2298.530 221.480 ;
        RECT 2338.270 221.200 2338.550 221.480 ;
        RECT 2572.410 221.200 2572.690 221.480 ;
        RECT 2612.430 221.880 2612.710 222.160 ;
        RECT 1281.190 197.400 1281.470 197.680 ;
        RECT 2844.270 198.080 2844.550 198.360 ;
      LAYER met3 ;
        RECT 381.455 5070.750 455.250 5161.315 ;
        RECT 381.455 5002.905 405.320 5070.750 ;
        RECT 431.120 5002.905 455.250 5070.750 ;
        RECT 638.455 5070.750 712.250 5161.315 ;
        RECT 638.455 5002.905 662.320 5070.750 ;
        RECT 688.120 5002.905 712.250 5070.750 ;
        RECT 895.455 5070.750 969.250 5161.315 ;
        RECT 895.455 5002.905 919.320 5070.750 ;
        RECT 945.120 5002.905 969.250 5070.750 ;
        RECT 1105.000 5004.085 1274.000 5188.000 ;
        RECT 1363.000 5004.085 1532.000 5188.000 ;
        RECT 1667.240 5014.250 1741.290 5188.000 ;
        RECT 1919.455 5070.750 1993.250 5161.315 ;
      LAYER met3 ;
        RECT 1105.000 4988.000 1176.395 5003.685 ;
      LAYER met3 ;
        RECT 1176.795 4999.730 1201.990 5004.085 ;
        RECT 1176.795 4991.125 1189.490 4999.730 ;
        RECT 1176.795 4990.725 1177.495 4991.125 ;
        RECT 1189.295 4990.725 1189.490 4991.125 ;
      LAYER met3 ;
        RECT 1177.895 4988.000 1188.895 4990.725 ;
        RECT 1189.890 4988.000 1200.890 4999.330 ;
      LAYER met3 ;
        RECT 1201.290 4990.725 1201.990 4999.730 ;
      LAYER met3 ;
        RECT 1363.000 4988.000 1434.395 5003.685 ;
      LAYER met3 ;
        RECT 1434.795 4999.730 1459.990 5004.085 ;
        RECT 1434.795 4991.125 1447.490 4999.730 ;
        RECT 1434.795 4990.725 1435.495 4991.125 ;
        RECT 1447.295 4990.725 1447.490 4991.125 ;
      LAYER met3 ;
        RECT 1435.895 4988.000 1446.895 4990.725 ;
        RECT 1447.890 4988.000 1458.890 4999.330 ;
      LAYER met3 ;
        RECT 1459.290 4990.725 1459.990 4999.730 ;
      LAYER met3 ;
        RECT 1667.495 4988.000 1691.395 5013.850 ;
      LAYER met3 ;
        RECT 1691.795 4990.035 1716.990 5014.250 ;
        RECT 1692.895 4988.000 1703.895 4990.035 ;
        RECT 1704.890 4988.000 1715.890 4990.035 ;
      LAYER met3 ;
        RECT 1717.390 4988.000 1741.290 5013.850 ;
      LAYER met3 ;
        RECT 1919.455 5002.905 1943.320 5070.750 ;
        RECT 1969.120 5002.905 1993.250 5070.750 ;
        RECT 2364.455 5070.750 2438.250 5161.315 ;
        RECT 2364.455 5002.905 2388.320 5070.750 ;
        RECT 2414.120 5002.905 2438.250 5070.750 ;
        RECT 2621.455 5070.750 2695.250 5161.315 ;
        RECT 2621.455 5002.905 2645.320 5070.750 ;
        RECT 2671.120 5002.905 2695.250 5070.750 ;
        RECT 2878.240 5025.160 2952.290 5183.100 ;
        RECT 3130.455 5070.750 3204.250 5161.315 ;
        RECT 2878.240 5020.915 2927.990 5025.160 ;
      LAYER met3 ;
        RECT 2878.495 4988.000 2902.395 5020.515 ;
      LAYER met3 ;
        RECT 2902.795 4990.035 2927.990 5020.915 ;
        RECT 2903.895 4988.000 2914.895 4990.035 ;
        RECT 2915.890 4988.000 2926.890 4990.035 ;
      LAYER met3 ;
        RECT 2928.390 4988.000 2952.290 5024.760 ;
      LAYER met3 ;
        RECT 3130.455 5002.905 3154.320 5070.750 ;
        RECT 3180.120 5002.905 3204.250 5070.750 ;
      LAYER met3 ;
        RECT 1717.950 4985.585 1718.250 4988.000 ;
        RECT 2925.205 4987.610 2925.535 4987.625 ;
        RECT 2928.670 4987.610 2928.970 4988.000 ;
        RECT 2925.205 4987.310 2928.970 4987.610 ;
        RECT 2925.205 4987.295 2925.535 4987.310 ;
        RECT 1717.950 4985.270 1718.495 4985.585 ;
        RECT 1718.165 4985.255 1718.495 4985.270 ;
      LAYER met3 ;
        RECT 26.685 4821.120 185.095 4845.250 ;
        RECT 26.685 4795.320 117.250 4821.120 ;
      LAYER met3 ;
        RECT 3388.000 4813.605 3403.685 4885.000 ;
      LAYER met3 ;
        RECT 3404.085 4813.205 3588.000 4885.000 ;
        RECT 3390.725 4812.505 3588.000 4813.205 ;
      LAYER met3 ;
        RECT 3388.000 4801.105 3390.725 4812.105 ;
      LAYER met3 ;
        RECT 3391.125 4800.705 3588.000 4812.505 ;
        RECT 3390.725 4800.510 3588.000 4800.705 ;
        RECT 26.685 4771.455 185.095 4795.320 ;
      LAYER met3 ;
        RECT 3388.000 4789.110 3399.330 4800.110 ;
      LAYER met3 ;
        RECT 3399.730 4788.710 3588.000 4800.510 ;
        RECT 3390.725 4788.010 3588.000 4788.710 ;
        RECT 3404.085 4716.000 3588.000 4788.010 ;
        RECT 0.035 4636.200 24.250 4645.935 ;
        RECT 153.765 4635.605 158.415 4646.140 ;
        RECT 169.550 4636.200 174.200 4645.935 ;
        RECT 0.035 4610.355 190.700 4635.000 ;
      LAYER met3 ;
        RECT 191.100 4610.755 198.000 4634.700 ;
      LAYER met3 ;
        RECT 3429.550 4613.895 3434.200 4623.975 ;
        RECT 3390.035 4612.900 3587.965 4613.000 ;
        RECT 0.035 4609.255 197.965 4610.355 ;
        RECT 0.035 4598.380 198.000 4609.255 ;
        RECT 0.035 4596.880 197.965 4598.380 ;
        RECT 0.035 4586.000 198.000 4596.880 ;
      LAYER met3 ;
        RECT 3390.000 4588.500 3396.900 4612.500 ;
      LAYER met3 ;
        RECT 3397.300 4588.100 3587.965 4612.900 ;
        RECT 3390.035 4587.000 3587.965 4588.100 ;
        RECT 0.035 4584.900 197.965 4586.000 ;
        RECT 0.035 4560.100 190.700 4584.900 ;
      LAYER met3 ;
        RECT 191.100 4560.500 198.000 4584.500 ;
      LAYER met3 ;
        RECT 3390.000 4576.120 3587.965 4587.000 ;
        RECT 3390.035 4574.620 3587.965 4576.120 ;
        RECT 3390.000 4563.745 3587.965 4574.620 ;
        RECT 3390.035 4562.645 3587.965 4563.745 ;
        RECT 0.035 4560.000 197.965 4560.100 ;
        RECT 153.800 4549.025 158.450 4559.105 ;
      LAYER met3 ;
        RECT 3390.000 4538.300 3396.900 4562.245 ;
      LAYER met3 ;
        RECT 3397.300 4538.000 3587.965 4562.645 ;
        RECT 3413.800 4527.065 3418.450 4536.800 ;
        RECT 3429.585 4526.860 3434.235 4537.395 ;
        RECT 3563.750 4527.065 3587.965 4536.800 ;
        RECT 0.000 4398.990 179.800 4423.290 ;
      LAYER met3 ;
        RECT 180.200 4399.390 200.000 4423.290 ;
      LAYER met3 ;
        RECT 0.000 4397.890 197.965 4398.990 ;
        RECT 0.000 4386.890 200.000 4397.890 ;
        RECT 0.000 4385.895 197.965 4386.890 ;
        RECT 0.000 4374.895 200.000 4385.895 ;
        RECT 0.000 4373.795 197.965 4374.895 ;
        RECT 0.000 4349.240 179.800 4373.795 ;
      LAYER met3 ;
        RECT 180.200 4350.450 200.000 4373.395 ;
        RECT 211.665 4350.450 211.995 4350.465 ;
        RECT 224.085 4350.450 224.415 4350.465 ;
        RECT 180.200 4350.150 224.415 4350.450 ;
        RECT 180.200 4349.495 200.000 4350.150 ;
        RECT 211.665 4350.135 211.995 4350.150 ;
        RECT 224.085 4350.135 224.415 4350.150 ;
      LAYER met3 ;
        RECT 3386.690 4312.430 3588.000 4391.690 ;
        RECT 4.900 4187.990 162.840 4212.290 ;
      LAYER met3 ;
        RECT 163.240 4188.390 200.000 4212.290 ;
      LAYER met3 ;
        RECT 4.900 4186.890 197.965 4187.990 ;
        RECT 4.900 4175.890 200.000 4186.890 ;
        RECT 4.900 4174.895 197.965 4175.890 ;
        RECT 4.900 4163.895 200.000 4174.895 ;
        RECT 4.900 4162.795 197.965 4163.895 ;
        RECT 4.900 4138.240 167.085 4162.795 ;
      LAYER met3 ;
        RECT 167.485 4138.495 200.000 4162.395 ;
        RECT 3388.000 4142.605 3402.960 4166.505 ;
      LAYER met3 ;
        RECT 3403.360 4142.205 3588.000 4166.760 ;
        RECT 3390.035 4141.105 3588.000 4142.205 ;
        RECT 3388.000 4130.105 3588.000 4141.105 ;
        RECT 3390.035 4129.110 3588.000 4130.105 ;
        RECT 3388.000 4118.110 3588.000 4129.110 ;
        RECT 3390.035 4117.010 3588.000 4118.110 ;
      LAYER met3 ;
        RECT 3388.000 4092.710 3402.960 4116.610 ;
      LAYER met3 ;
        RECT 3403.360 4092.710 3588.000 4117.010 ;
      LAYER met3 ;
        RECT 3387.965 4092.050 3388.295 4092.065 ;
        RECT 3388.670 4092.050 3388.970 4092.710 ;
        RECT 3387.965 4091.750 3388.970 4092.050 ;
        RECT 3387.965 4091.735 3388.295 4091.750 ;
      LAYER met3 ;
        RECT 0.000 3922.310 201.310 4001.570 ;
        RECT 3386.690 3866.430 3588.000 3945.690 ;
        RECT 0.000 3706.310 201.310 3785.570 ;
        RECT 3386.690 3641.430 3588.000 3720.690 ;
        RECT 0.000 3490.310 201.310 3569.570 ;
        RECT 3386.690 3416.430 3588.000 3495.690 ;
        RECT 0.000 3274.310 201.310 3353.570 ;
        RECT 3386.690 3190.430 3588.000 3269.690 ;
        RECT 0.000 3058.310 201.310 3137.570 ;
        RECT 3386.690 2965.430 3588.000 3044.690 ;
        RECT 0.000 2842.310 201.310 2921.570 ;
        RECT 3386.690 2739.430 3588.000 2818.690 ;
        RECT 0.000 2626.310 201.310 2705.570 ;
      LAYER met3 ;
        RECT 3388.000 2569.605 3402.960 2593.505 ;
        RECT 3388.670 2568.865 3388.970 2569.605 ;
      LAYER met3 ;
        RECT 3403.360 2569.205 3588.000 2593.760 ;
      LAYER met3 ;
        RECT 3388.425 2568.550 3388.970 2568.865 ;
        RECT 3388.425 2568.535 3388.755 2568.550 ;
      LAYER met3 ;
        RECT 3390.035 2568.105 3588.000 2569.205 ;
        RECT 3388.000 2557.105 3588.000 2568.105 ;
        RECT 3390.035 2556.110 3588.000 2557.105 ;
        RECT 3388.000 2545.110 3588.000 2556.110 ;
        RECT 3390.035 2544.010 3588.000 2545.110 ;
      LAYER met3 ;
        RECT 3388.000 2519.710 3402.960 2543.610 ;
      LAYER met3 ;
        RECT 3403.360 2519.710 3588.000 2544.010 ;
        RECT 0.000 2464.990 184.640 2489.290 ;
      LAYER met3 ;
        RECT 185.040 2465.390 200.000 2489.290 ;
      LAYER met3 ;
        RECT 0.000 2463.890 197.965 2464.990 ;
        RECT 0.000 2452.890 200.000 2463.890 ;
        RECT 0.000 2451.895 197.965 2452.890 ;
        RECT 0.000 2440.895 200.000 2451.895 ;
        RECT 0.000 2439.795 197.965 2440.895 ;
        RECT 0.000 2415.240 184.640 2439.795 ;
      LAYER met3 ;
        RECT 185.040 2415.495 200.000 2439.395 ;
      LAYER met3 ;
        RECT 3429.550 2374.895 3434.200 2384.975 ;
        RECT 3390.035 2373.900 3587.965 2374.000 ;
        RECT 3430.000 2349.100 3587.965 2373.900 ;
        RECT 3390.035 2348.000 3587.965 2349.100 ;
        RECT 3390.000 2337.120 3587.965 2348.000 ;
        RECT 3390.035 2335.620 3587.965 2337.120 ;
        RECT 3390.000 2324.745 3587.965 2335.620 ;
        RECT 3390.035 2323.645 3587.965 2324.745 ;
      LAYER met3 ;
        RECT 3390.000 2299.300 3429.600 2323.245 ;
      LAYER met3 ;
        RECT 3430.000 2299.000 3587.965 2323.645 ;
        RECT 0.035 2280.200 24.250 2289.935 ;
        RECT 153.765 2279.605 158.415 2290.140 ;
        RECT 169.550 2280.200 174.200 2289.935 ;
        RECT 3413.800 2288.065 3418.450 2297.800 ;
        RECT 3429.585 2287.860 3434.235 2298.395 ;
        RECT 3563.750 2288.065 3587.965 2297.800 ;
        RECT 0.035 2254.355 158.000 2279.000 ;
      LAYER met3 ;
        RECT 158.400 2254.755 198.000 2278.700 ;
      LAYER met3 ;
        RECT 0.035 2253.255 197.965 2254.355 ;
        RECT 0.035 2242.380 198.000 2253.255 ;
        RECT 0.035 2240.880 197.965 2242.380 ;
        RECT 0.035 2230.000 198.000 2240.880 ;
        RECT 0.035 2228.900 197.965 2230.000 ;
        RECT 0.035 2204.100 158.000 2228.900 ;
        RECT 0.035 2204.000 197.965 2204.100 ;
        RECT 153.800 2193.025 158.450 2203.105 ;
      LAYER met3 ;
        RECT 3388.000 2128.605 3420.515 2152.505 ;
        RECT 3387.505 2128.210 3387.835 2128.225 ;
        RECT 3388.670 2128.210 3388.970 2128.605 ;
        RECT 3387.505 2127.910 3388.970 2128.210 ;
      LAYER met3 ;
        RECT 3420.915 2128.205 3583.100 2152.760 ;
      LAYER met3 ;
        RECT 3387.505 2127.895 3387.835 2127.910 ;
      LAYER met3 ;
        RECT 3390.035 2127.105 3583.100 2128.205 ;
        RECT 3388.000 2116.105 3583.100 2127.105 ;
        RECT 3390.035 2115.110 3583.100 2116.105 ;
        RECT 3388.000 2104.110 3583.100 2115.110 ;
        RECT 3390.035 2103.010 3583.100 2104.110 ;
      LAYER met3 ;
        RECT 3388.000 2078.710 3424.760 2102.610 ;
      LAYER met3 ;
        RECT 3425.160 2078.710 3583.100 2103.010 ;
        RECT 0.000 1988.310 201.310 2067.570 ;
        RECT 3386.690 1853.430 3588.000 1932.690 ;
        RECT 0.000 1772.310 201.310 1851.570 ;
        RECT 0.000 1556.310 201.310 1635.570 ;
        RECT 3386.690 1627.430 3588.000 1706.690 ;
        RECT 0.000 1340.310 201.310 1419.570 ;
        RECT 3386.690 1402.430 3588.000 1481.690 ;
        RECT 0.000 1124.310 201.310 1203.570 ;
        RECT 3386.690 1177.430 3588.000 1256.690 ;
        RECT 0.000 908.310 201.310 987.570 ;
        RECT 3386.690 951.430 3588.000 1030.690 ;
        RECT 3386.690 726.430 3588.000 805.690 ;
        RECT 0.000 600.990 179.800 625.290 ;
      LAYER met3 ;
        RECT 180.200 601.390 200.000 625.290 ;
      LAYER met3 ;
        RECT 0.000 599.890 197.965 600.990 ;
        RECT 0.000 588.890 200.000 599.890 ;
        RECT 0.000 587.895 197.965 588.890 ;
        RECT 0.000 576.895 200.000 587.895 ;
        RECT 0.000 575.795 197.965 576.895 ;
        RECT 0.000 551.240 179.800 575.795 ;
      LAYER met3 ;
        RECT 180.200 552.650 200.000 575.395 ;
        RECT 220.865 552.650 221.195 552.665 ;
        RECT 224.085 552.650 224.415 552.665 ;
        RECT 180.200 552.350 224.415 552.650 ;
        RECT 180.200 551.495 200.000 552.350 ;
        RECT 220.865 552.335 221.195 552.350 ;
        RECT 224.085 552.335 224.415 552.350 ;
      LAYER met3 ;
        RECT 3386.690 500.430 3588.000 579.690 ;
        RECT 153.765 415.605 158.415 426.140 ;
        RECT 159.805 415.440 163.270 426.140 ;
        RECT 4.395 390.355 190.700 415.000 ;
      LAYER met3 ;
        RECT 191.100 390.755 198.000 414.700 ;
      LAYER met3 ;
        RECT 4.395 389.255 197.965 390.355 ;
        RECT 4.395 378.380 198.000 389.255 ;
        RECT 4.395 376.880 197.965 378.380 ;
        RECT 4.395 366.000 198.000 376.880 ;
        RECT 4.395 364.900 197.965 366.000 ;
        RECT 4.395 340.490 190.700 364.900 ;
      LAYER met3 ;
        RECT 191.100 359.530 198.000 364.500 ;
        RECT 220.865 359.530 221.195 359.545 ;
        RECT 224.085 359.530 224.415 359.545 ;
        RECT 191.100 359.230 224.415 359.530 ;
        RECT 191.100 340.500 198.000 359.230 ;
        RECT 220.865 359.215 221.195 359.230 ;
        RECT 224.085 359.215 224.415 359.230 ;
        RECT 2612.405 222.170 2612.735 222.185 ;
        RECT 2580.450 221.870 2612.735 222.170 ;
        RECT 2024.525 221.490 2024.855 221.505 ;
        RECT 2064.545 221.490 2064.875 221.505 ;
        RECT 2024.525 221.190 2064.875 221.490 ;
        RECT 2024.525 221.175 2024.855 221.190 ;
        RECT 2064.545 221.175 2064.875 221.190 ;
        RECT 2298.225 221.490 2298.555 221.505 ;
        RECT 2338.245 221.490 2338.575 221.505 ;
        RECT 2298.225 221.190 2338.575 221.490 ;
        RECT 2298.225 221.175 2298.555 221.190 ;
        RECT 2338.245 221.175 2338.575 221.190 ;
        RECT 2572.385 221.490 2572.715 221.505 ;
        RECT 2580.450 221.490 2580.750 221.870 ;
        RECT 2612.405 221.855 2612.735 221.870 ;
        RECT 2572.385 221.190 2580.750 221.490 ;
        RECT 2572.385 221.175 2572.715 221.190 ;
        RECT 745.265 201.770 745.595 201.785 ;
        RECT 729.190 201.470 745.595 201.770 ;
        RECT 468.805 201.090 469.135 201.105 ;
        RECT 675.805 201.090 676.135 201.105 ;
        RECT 455.710 200.790 469.135 201.090 ;
        RECT 455.710 200.000 456.010 200.790 ;
        RECT 468.805 200.775 469.135 200.790 ;
        RECT 665.470 200.790 676.135 201.090 ;
        RECT 665.470 200.000 665.770 200.790 ;
        RECT 675.805 200.775 676.135 200.790 ;
        RECT 715.365 201.090 715.695 201.105 ;
        RECT 717.665 201.090 717.995 201.105 ;
        RECT 715.365 200.790 717.290 201.090 ;
        RECT 715.365 200.775 715.695 200.790 ;
        RECT 716.990 200.000 717.290 200.790 ;
        RECT 717.665 200.790 720.050 201.090 ;
        RECT 717.665 200.775 717.995 200.790 ;
        RECT 719.750 200.000 720.050 200.790 ;
        RECT 729.190 200.070 729.490 201.470 ;
        RECT 745.265 201.455 745.595 201.470 ;
        RECT 729.100 200.000 729.490 200.070 ;
        RECT 238.000 164.765 256.010 180.085 ;
        RECT 258.000 164.765 276.010 180.085 ;
        RECT 278.000 164.765 296.010 180.085 ;
        RECT 298.000 164.765 316.010 180.085 ;
        RECT 318.000 164.765 336.010 180.085 ;
        RECT 338.000 164.765 356.010 180.085 ;
        RECT 394.710 163.240 418.610 200.000 ;
      LAYER met3 ;
        RECT 420.110 197.965 431.110 200.000 ;
        RECT 432.105 197.965 443.105 200.000 ;
        RECT 419.010 167.085 444.205 197.965 ;
      LAYER met3 ;
        RECT 444.605 167.485 468.505 200.000 ;
      LAYER met3 ;
        RECT 419.010 162.840 468.760 167.085 ;
      LAYER met3 ;
        RECT 507.000 164.765 525.010 180.085 ;
        RECT 527.000 164.765 545.010 180.085 ;
        RECT 547.000 164.765 565.010 180.085 ;
        RECT 567.000 164.765 585.010 180.085 ;
        RECT 587.000 164.765 605.010 180.085 ;
        RECT 607.000 164.765 625.010 180.085 ;
      LAYER met3 ;
        RECT 394.710 4.900 468.760 162.840 ;
        RECT 663.300 151.080 664.340 199.375 ;
        RECT 663.300 133.400 663.675 151.080 ;
      LAYER met3 ;
        RECT 664.740 150.680 665.810 200.000 ;
        RECT 664.075 135.400 665.810 150.680 ;
      LAYER met3 ;
        RECT 666.210 188.690 707.935 199.375 ;
        RECT 709.465 193.730 716.375 199.375 ;
        RECT 709.465 192.265 714.910 193.730 ;
      LAYER met3 ;
        RECT 716.775 193.330 717.925 200.000 ;
      LAYER met3 ;
        RECT 709.465 191.985 714.630 192.265 ;
        RECT 709.465 190.555 713.550 191.985 ;
      LAYER met3 ;
        RECT 715.310 191.950 717.925 193.330 ;
        RECT 715.310 191.865 716.875 191.950 ;
        RECT 716.940 191.865 717.925 191.950 ;
      LAYER met3 ;
        RECT 718.325 196.465 718.690 199.375 ;
      LAYER met3 ;
        RECT 719.090 196.865 720.755 200.000 ;
      LAYER met3 ;
        RECT 721.155 196.465 728.680 199.375 ;
      LAYER met3 ;
        RECT 715.030 191.800 715.310 191.865 ;
        RECT 715.395 191.800 716.940 191.865 ;
        RECT 715.030 191.650 716.940 191.800 ;
        RECT 715.030 191.585 716.575 191.650 ;
        RECT 716.660 191.585 716.940 191.650 ;
      LAYER met3 ;
        RECT 709.765 190.255 713.550 190.555 ;
        RECT 666.210 184.830 708.700 188.690 ;
        RECT 710.230 187.335 713.550 190.255 ;
      LAYER met3 ;
        RECT 713.950 191.500 715.030 191.585 ;
        RECT 715.095 191.500 716.660 191.585 ;
        RECT 713.950 190.020 716.660 191.500 ;
      LAYER met3 ;
        RECT 718.325 191.465 728.680 196.465 ;
        RECT 717.340 191.185 728.680 191.465 ;
      LAYER met3 ;
        RECT 713.950 187.735 715.095 190.020 ;
      LAYER met3 ;
        RECT 717.060 189.620 728.680 191.185 ;
        RECT 715.495 187.335 728.680 189.620 ;
        RECT 710.230 184.830 728.680 187.335 ;
        RECT 666.210 183.015 728.680 184.830 ;
      LAYER met3 ;
        RECT 729.080 184.215 729.600 200.000 ;
      LAYER met3 ;
        RECT 730.000 184.615 737.035 199.375 ;
        RECT 730.210 184.405 737.035 184.615 ;
      LAYER met3 ;
        RECT 729.080 184.005 729.810 184.215 ;
        RECT 729.080 183.555 730.260 184.005 ;
      LAYER met3 ;
        RECT 730.660 183.955 737.035 184.405 ;
      LAYER met3 ;
        RECT 729.080 183.415 729.670 183.555 ;
        RECT 729.680 183.415 730.710 183.555 ;
      LAYER met3 ;
        RECT 731.110 183.505 737.035 183.955 ;
      LAYER met3 ;
        RECT 729.670 183.105 730.710 183.415 ;
      LAYER met3 ;
        RECT 666.210 182.555 729.270 183.015 ;
      LAYER met3 ;
        RECT 729.670 182.955 731.225 183.105 ;
      LAYER met3 ;
        RECT 666.210 181.980 729.730 182.555 ;
      LAYER met3 ;
        RECT 730.130 182.380 731.225 182.955 ;
      LAYER met3 ;
        RECT 666.210 169.105 730.305 181.980 ;
        RECT 666.210 168.520 729.720 169.105 ;
      LAYER met3 ;
        RECT 730.705 168.705 731.225 182.380 ;
      LAYER met3 ;
        RECT 666.210 167.805 729.005 168.520 ;
      LAYER met3 ;
        RECT 730.120 168.195 731.225 168.705 ;
        RECT 730.120 168.120 730.775 168.195 ;
        RECT 730.850 168.120 731.225 168.195 ;
        RECT 729.405 168.045 730.120 168.120 ;
        RECT 730.135 168.045 730.850 168.120 ;
      LAYER met3 ;
        RECT 666.210 167.220 728.420 167.805 ;
      LAYER met3 ;
        RECT 729.405 167.445 730.850 168.045 ;
      LAYER met3 ;
        RECT 731.625 167.720 737.035 183.505 ;
      LAYER met3 ;
        RECT 729.405 167.405 730.120 167.445 ;
        RECT 730.135 167.405 730.850 167.445 ;
        RECT 728.820 167.295 729.405 167.405 ;
        RECT 729.445 167.295 730.135 167.405 ;
      LAYER met3 ;
        RECT 666.210 167.005 728.205 167.220 ;
        RECT 666.210 165.475 715.325 167.005 ;
      LAYER met3 ;
        RECT 728.820 166.845 730.135 167.295 ;
      LAYER met3 ;
        RECT 731.250 167.005 737.035 167.720 ;
      LAYER met3 ;
        RECT 728.820 166.820 729.425 166.845 ;
        RECT 729.550 166.820 730.135 166.845 ;
        RECT 728.605 166.695 728.820 166.820 ;
        RECT 728.845 166.695 729.550 166.820 ;
        RECT 728.605 166.605 729.550 166.695 ;
        RECT 715.725 166.305 729.550 166.605 ;
      LAYER met3 ;
        RECT 730.535 166.420 737.035 167.005 ;
      LAYER met3 ;
        RECT 715.725 166.300 728.885 166.305 ;
        RECT 729.030 166.300 729.550 166.305 ;
        RECT 715.725 165.875 729.030 166.300 ;
      LAYER met3 ;
        RECT 729.950 165.900 737.035 166.420 ;
        RECT 729.430 165.475 737.035 165.900 ;
        RECT 666.210 135.800 737.035 165.475 ;
      LAYER met3 ;
        RECT 776.000 164.765 794.010 180.085 ;
        RECT 796.000 164.765 814.010 180.085 ;
        RECT 816.000 164.765 834.010 180.085 ;
        RECT 836.000 164.765 854.010 180.085 ;
        RECT 856.000 164.765 874.010 180.085 ;
        RECT 876.000 164.765 894.010 180.085 ;
        RECT 664.075 133.800 667.410 135.400 ;
      LAYER met3 ;
        RECT 667.810 134.200 737.035 135.800 ;
        RECT 663.300 131.800 665.410 133.400 ;
      LAYER met3 ;
        RECT 665.810 132.400 668.810 133.800 ;
      LAYER met3 ;
        RECT 669.210 132.800 737.035 134.200 ;
      LAYER met3 ;
        RECT 665.810 132.250 669.745 132.400 ;
        RECT 665.810 132.200 667.410 132.250 ;
        RECT 667.510 132.200 669.745 132.250 ;
      LAYER met3 ;
        RECT 663.300 130.515 667.010 131.800 ;
      LAYER met3 ;
        RECT 667.410 131.465 669.745 132.200 ;
      LAYER met3 ;
        RECT 670.145 131.865 737.035 132.800 ;
      LAYER met3 ;
        RECT 667.410 131.350 669.710 131.465 ;
        RECT 669.745 131.350 670.610 131.465 ;
        RECT 667.410 131.050 670.610 131.350 ;
        RECT 667.410 130.915 668.695 131.050 ;
        RECT 668.710 130.915 670.610 131.050 ;
      LAYER met3 ;
        RECT 671.010 131.000 737.035 131.865 ;
      LAYER met3 ;
        RECT 668.695 130.600 670.610 130.915 ;
      LAYER met3 ;
        RECT 663.300 129.565 668.295 130.515 ;
      LAYER met3 ;
        RECT 668.695 130.000 671.960 130.600 ;
        RECT 668.695 129.965 669.645 130.000 ;
        RECT 669.760 129.965 671.960 130.000 ;
      LAYER met3 ;
        RECT 663.300 128.600 669.245 129.565 ;
      LAYER met3 ;
        RECT 669.645 129.250 671.960 129.965 ;
      LAYER met3 ;
        RECT 672.360 129.650 737.035 131.000 ;
      LAYER met3 ;
        RECT 669.645 129.100 673.140 129.250 ;
        RECT 669.645 129.000 670.610 129.100 ;
        RECT 670.660 129.000 673.140 129.100 ;
      LAYER met3 ;
        RECT 663.300 127.390 670.210 128.600 ;
      LAYER met3 ;
        RECT 670.610 127.920 673.140 129.000 ;
        RECT 670.610 127.790 671.820 127.920 ;
        RECT 671.840 127.790 673.140 127.920 ;
        RECT 671.820 127.600 673.140 127.790 ;
      LAYER met3 ;
        RECT 663.300 127.200 671.420 127.390 ;
        RECT 663.300 104.955 671.610 127.200 ;
      LAYER met3 ;
        RECT 672.010 105.355 673.140 127.600 ;
      LAYER met3 ;
        RECT 673.540 104.955 737.035 129.650 ;
        RECT 663.300 0.000 737.035 104.955 ;
        RECT 932.430 0.000 1011.690 201.310 ;
      LAYER met3 ;
        RECT 1050.000 164.765 1068.010 180.085 ;
        RECT 1070.000 164.765 1088.010 180.085 ;
        RECT 1090.000 164.765 1108.010 180.085 ;
        RECT 1110.000 164.765 1128.010 180.085 ;
        RECT 1130.000 164.765 1148.010 180.085 ;
        RECT 1150.000 164.765 1168.010 180.085 ;
      LAYER met3 ;
        RECT 1194.860 159.805 1205.560 163.270 ;
        RECT 1194.860 153.765 1205.395 158.415 ;
      LAYER met3 ;
        RECT 1206.300 158.400 1230.245 198.000 ;
      LAYER met3 ;
        RECT 1231.745 197.965 1242.620 198.000 ;
        RECT 1244.120 197.965 1255.000 198.000 ;
        RECT 1230.645 158.000 1256.100 197.965 ;
      LAYER met3 ;
        RECT 1256.500 197.690 1280.500 198.000 ;
        RECT 1281.165 197.690 1281.495 197.705 ;
        RECT 1256.500 197.390 1281.495 197.690 ;
        RECT 1256.500 158.400 1280.500 197.390 ;
        RECT 1281.165 197.375 1281.495 197.390 ;
        RECT 1319.000 164.765 1337.010 180.085 ;
        RECT 1339.000 164.765 1357.010 180.085 ;
        RECT 1359.000 164.765 1377.010 180.085 ;
        RECT 1379.000 164.765 1397.010 180.085 ;
        RECT 1399.000 164.765 1417.010 180.085 ;
        RECT 1419.000 164.765 1437.010 180.085 ;
      LAYER met3 ;
        RECT 1206.000 4.395 1280.500 158.000 ;
        RECT 1475.430 0.000 1554.690 201.310 ;
      LAYER met3 ;
        RECT 1593.000 164.765 1611.010 180.085 ;
        RECT 1613.000 164.765 1631.010 180.085 ;
        RECT 1633.000 164.765 1651.010 180.085 ;
        RECT 1653.000 164.765 1671.010 180.085 ;
        RECT 1673.000 164.765 1691.010 180.085 ;
        RECT 1693.000 164.765 1711.010 180.085 ;
      LAYER met3 ;
        RECT 1749.430 0.000 1828.690 201.310 ;
      LAYER met3 ;
        RECT 1867.000 164.765 1885.010 180.085 ;
        RECT 1887.000 164.765 1905.010 180.085 ;
        RECT 1907.000 164.765 1925.010 180.085 ;
        RECT 1927.000 164.765 1945.010 180.085 ;
        RECT 1947.000 164.765 1965.010 180.085 ;
        RECT 1967.000 164.765 1985.010 180.085 ;
      LAYER met3 ;
        RECT 2023.430 0.000 2102.690 201.310 ;
      LAYER met3 ;
        RECT 2141.000 164.765 2159.010 180.085 ;
        RECT 2161.000 164.765 2179.010 180.085 ;
        RECT 2181.000 164.765 2199.010 180.085 ;
        RECT 2201.000 164.765 2219.010 180.085 ;
        RECT 2221.000 164.765 2239.010 180.085 ;
        RECT 2241.000 164.765 2259.010 180.085 ;
      LAYER met3 ;
        RECT 2297.430 0.000 2376.690 201.310 ;
      LAYER met3 ;
        RECT 2415.000 164.765 2433.010 180.085 ;
        RECT 2435.000 164.765 2453.010 180.085 ;
        RECT 2455.000 164.765 2473.010 180.085 ;
        RECT 2475.000 164.765 2493.010 180.085 ;
        RECT 2495.000 164.765 2513.010 180.085 ;
        RECT 2515.000 164.765 2533.010 180.085 ;
      LAYER met3 ;
        RECT 2571.430 0.000 2650.690 201.310 ;
      LAYER met3 ;
        RECT 2844.245 198.370 2844.575 198.385 ;
        RECT 2845.710 198.370 2869.610 200.000 ;
        RECT 2844.245 198.070 2869.610 198.370 ;
        RECT 2844.245 198.055 2844.575 198.070 ;
        RECT 2689.000 164.765 2707.010 180.085 ;
        RECT 2709.000 164.765 2727.010 180.085 ;
        RECT 2729.000 164.765 2747.010 180.085 ;
        RECT 2749.000 164.765 2767.010 180.085 ;
        RECT 2769.000 164.765 2787.010 180.085 ;
        RECT 2789.000 164.765 2807.010 180.085 ;
        RECT 2845.710 174.150 2869.610 198.070 ;
      LAYER met3 ;
        RECT 2871.110 197.965 2882.110 200.000 ;
        RECT 2883.105 197.965 2894.105 200.000 ;
        RECT 2870.010 173.750 2895.205 197.965 ;
      LAYER met3 ;
        RECT 2895.605 174.150 2919.505 200.000 ;
        RECT 3114.710 185.040 3138.610 200.000 ;
      LAYER met3 ;
        RECT 3140.110 197.965 3151.110 200.000 ;
        RECT 3152.105 197.965 3163.105 200.000 ;
        RECT 3139.010 184.640 3164.205 197.965 ;
      LAYER met3 ;
        RECT 3164.605 185.040 3188.505 200.000 ;
      LAYER met3 ;
        RECT 2845.710 0.000 2919.760 173.750 ;
      LAYER met3 ;
        RECT 2958.000 164.765 2976.010 180.085 ;
        RECT 2978.000 164.765 2996.010 180.085 ;
        RECT 2998.000 164.765 3016.010 180.085 ;
        RECT 3018.000 164.765 3036.010 180.085 ;
        RECT 3038.000 164.765 3056.010 180.085 ;
        RECT 3058.000 164.765 3076.010 180.085 ;
      LAYER met3 ;
        RECT 3114.710 0.000 3188.760 184.640 ;
      LAYER met3 ;
        RECT 3227.000 164.765 3245.010 180.085 ;
        RECT 3247.000 164.765 3265.010 180.085 ;
        RECT 3267.000 164.765 3285.010 180.085 ;
        RECT 3287.000 164.765 3305.010 180.085 ;
        RECT 3307.000 164.765 3325.010 180.085 ;
        RECT 3327.000 164.765 3345.010 180.085 ;
      LAYER via3 ;
        RECT 238.230 175.875 255.720 179.885 ;
        RECT 238.260 164.935 255.910 167.885 ;
        RECT 258.230 175.875 275.720 179.885 ;
        RECT 258.260 164.935 275.910 167.885 ;
        RECT 278.230 175.875 295.720 179.885 ;
        RECT 278.260 164.935 295.910 167.885 ;
        RECT 298.230 175.875 315.720 179.885 ;
        RECT 298.260 164.935 315.910 167.885 ;
        RECT 318.230 175.875 335.720 179.885 ;
        RECT 318.260 164.935 335.910 167.885 ;
        RECT 338.230 175.875 355.720 179.885 ;
        RECT 338.260 164.935 355.910 167.885 ;
        RECT 507.230 175.875 524.720 179.885 ;
        RECT 507.260 164.935 524.910 167.885 ;
        RECT 527.230 175.875 544.720 179.885 ;
        RECT 527.260 164.935 544.910 167.885 ;
        RECT 547.230 175.875 564.720 179.885 ;
        RECT 547.260 164.935 564.910 167.885 ;
        RECT 567.230 175.875 584.720 179.885 ;
        RECT 567.260 164.935 584.910 167.885 ;
        RECT 587.230 175.875 604.720 179.885 ;
        RECT 587.260 164.935 604.910 167.885 ;
        RECT 607.230 175.875 624.720 179.885 ;
        RECT 607.260 164.935 624.910 167.885 ;
        RECT 776.230 175.875 793.720 179.885 ;
        RECT 776.260 164.935 793.910 167.885 ;
        RECT 796.230 175.875 813.720 179.885 ;
        RECT 796.260 164.935 813.910 167.885 ;
        RECT 816.230 175.875 833.720 179.885 ;
        RECT 816.260 164.935 833.910 167.885 ;
        RECT 836.230 175.875 853.720 179.885 ;
        RECT 836.260 164.935 853.910 167.885 ;
        RECT 856.230 175.875 873.720 179.885 ;
        RECT 856.260 164.935 873.910 167.885 ;
        RECT 876.230 175.875 893.720 179.885 ;
        RECT 876.260 164.935 893.910 167.885 ;
        RECT 1050.230 175.875 1067.720 179.885 ;
        RECT 1050.260 164.935 1067.910 167.885 ;
        RECT 1070.230 175.875 1087.720 179.885 ;
        RECT 1070.260 164.935 1087.910 167.885 ;
        RECT 1090.230 175.875 1107.720 179.885 ;
        RECT 1090.260 164.935 1107.910 167.885 ;
        RECT 1110.230 175.875 1127.720 179.885 ;
        RECT 1110.260 164.935 1127.910 167.885 ;
        RECT 1130.230 175.875 1147.720 179.885 ;
        RECT 1130.260 164.935 1147.910 167.885 ;
        RECT 1150.230 175.875 1167.720 179.885 ;
        RECT 1150.260 164.935 1167.910 167.885 ;
        RECT 1319.230 175.875 1336.720 179.885 ;
        RECT 1319.260 164.935 1336.910 167.885 ;
        RECT 1339.230 175.875 1356.720 179.885 ;
        RECT 1339.260 164.935 1356.910 167.885 ;
        RECT 1359.230 175.875 1376.720 179.885 ;
        RECT 1359.260 164.935 1376.910 167.885 ;
        RECT 1379.230 175.875 1396.720 179.885 ;
        RECT 1379.260 164.935 1396.910 167.885 ;
        RECT 1399.230 175.875 1416.720 179.885 ;
        RECT 1399.260 164.935 1416.910 167.885 ;
        RECT 1419.230 175.875 1436.720 179.885 ;
        RECT 1419.260 164.935 1436.910 167.885 ;
        RECT 1593.230 175.875 1610.720 179.885 ;
        RECT 1593.260 164.935 1610.910 167.885 ;
        RECT 1613.230 175.875 1630.720 179.885 ;
        RECT 1613.260 164.935 1630.910 167.885 ;
        RECT 1633.230 175.875 1650.720 179.885 ;
        RECT 1633.260 164.935 1650.910 167.885 ;
        RECT 1653.230 175.875 1670.720 179.885 ;
        RECT 1653.260 164.935 1670.910 167.885 ;
        RECT 1673.230 175.875 1690.720 179.885 ;
        RECT 1673.260 164.935 1690.910 167.885 ;
        RECT 1693.230 175.875 1710.720 179.885 ;
        RECT 1693.260 164.935 1710.910 167.885 ;
        RECT 1867.230 175.875 1884.720 179.885 ;
        RECT 1867.260 164.935 1884.910 167.885 ;
        RECT 1887.230 175.875 1904.720 179.885 ;
        RECT 1887.260 164.935 1904.910 167.885 ;
        RECT 1907.230 175.875 1924.720 179.885 ;
        RECT 1907.260 164.935 1924.910 167.885 ;
        RECT 1927.230 175.875 1944.720 179.885 ;
        RECT 1927.260 164.935 1944.910 167.885 ;
        RECT 1947.230 175.875 1964.720 179.885 ;
        RECT 1947.260 164.935 1964.910 167.885 ;
        RECT 1967.230 175.875 1984.720 179.885 ;
        RECT 1967.260 164.935 1984.910 167.885 ;
        RECT 2141.230 175.875 2158.720 179.885 ;
        RECT 2141.260 164.935 2158.910 167.885 ;
        RECT 2161.230 175.875 2178.720 179.885 ;
        RECT 2161.260 164.935 2178.910 167.885 ;
        RECT 2181.230 175.875 2198.720 179.885 ;
        RECT 2181.260 164.935 2198.910 167.885 ;
        RECT 2201.230 175.875 2218.720 179.885 ;
        RECT 2201.260 164.935 2218.910 167.885 ;
        RECT 2221.230 175.875 2238.720 179.885 ;
        RECT 2221.260 164.935 2238.910 167.885 ;
        RECT 2241.230 175.875 2258.720 179.885 ;
        RECT 2241.260 164.935 2258.910 167.885 ;
        RECT 2415.230 175.875 2432.720 179.885 ;
        RECT 2415.260 164.935 2432.910 167.885 ;
        RECT 2435.230 175.875 2452.720 179.885 ;
        RECT 2435.260 164.935 2452.910 167.885 ;
        RECT 2455.230 175.875 2472.720 179.885 ;
        RECT 2455.260 164.935 2472.910 167.885 ;
        RECT 2475.230 175.875 2492.720 179.885 ;
        RECT 2475.260 164.935 2492.910 167.885 ;
        RECT 2495.230 175.875 2512.720 179.885 ;
        RECT 2495.260 164.935 2512.910 167.885 ;
        RECT 2515.230 175.875 2532.720 179.885 ;
        RECT 2515.260 164.935 2532.910 167.885 ;
        RECT 2689.230 175.875 2706.720 179.885 ;
        RECT 2689.260 164.935 2706.910 167.885 ;
        RECT 2709.230 175.875 2726.720 179.885 ;
        RECT 2709.260 164.935 2726.910 167.885 ;
        RECT 2729.230 175.875 2746.720 179.885 ;
        RECT 2729.260 164.935 2746.910 167.885 ;
        RECT 2749.230 175.875 2766.720 179.885 ;
        RECT 2749.260 164.935 2766.910 167.885 ;
        RECT 2769.230 175.875 2786.720 179.885 ;
        RECT 2769.260 164.935 2786.910 167.885 ;
        RECT 2789.230 175.875 2806.720 179.885 ;
        RECT 2958.230 175.875 2975.720 179.885 ;
        RECT 2789.260 164.935 2806.910 167.885 ;
        RECT 2958.260 164.935 2975.910 167.885 ;
        RECT 2978.230 175.875 2995.720 179.885 ;
        RECT 2978.260 164.935 2995.910 167.885 ;
        RECT 2998.230 175.875 3015.720 179.885 ;
        RECT 2998.260 164.935 3015.910 167.885 ;
        RECT 3018.230 175.875 3035.720 179.885 ;
        RECT 3018.260 164.935 3035.910 167.885 ;
        RECT 3038.230 175.875 3055.720 179.885 ;
        RECT 3038.260 164.935 3055.910 167.885 ;
        RECT 3058.230 175.875 3075.720 179.885 ;
        RECT 3058.260 164.935 3075.910 167.885 ;
        RECT 3227.230 175.875 3244.720 179.885 ;
        RECT 3227.260 164.935 3244.910 167.885 ;
        RECT 3247.230 175.875 3264.720 179.885 ;
        RECT 3247.260 164.935 3264.910 167.885 ;
        RECT 3267.230 175.875 3284.720 179.885 ;
        RECT 3267.260 164.935 3284.910 167.885 ;
        RECT 3287.230 175.875 3304.720 179.885 ;
        RECT 3287.260 164.935 3304.910 167.885 ;
        RECT 3307.230 175.875 3324.720 179.885 ;
        RECT 3307.260 164.935 3324.910 167.885 ;
        RECT 3327.230 175.875 3344.720 179.885 ;
        RECT 3327.260 164.935 3344.910 167.885 ;
      LAYER met4 ;
        RECT 0.000 5163.385 202.330 5188.000 ;
      LAYER met4 ;
        RECT 202.730 5163.785 204.000 5188.000 ;
      LAYER met4 ;
        RECT 0.000 5083.400 202.745 5163.385 ;
        RECT 204.000 5083.400 381.000 5188.000 ;
      LAYER met4 ;
        RECT 381.000 5163.785 382.270 5188.000 ;
      LAYER met4 ;
        RECT 382.670 5163.385 454.330 5188.000 ;
      LAYER met4 ;
        RECT 454.730 5163.785 456.000 5188.000 ;
      LAYER met4 ;
        RECT 381.965 5083.400 455.035 5163.385 ;
        RECT 456.000 5083.400 638.000 5188.000 ;
      LAYER met4 ;
        RECT 638.000 5163.785 639.270 5188.000 ;
      LAYER met4 ;
        RECT 639.670 5163.385 711.330 5188.000 ;
      LAYER met4 ;
        RECT 711.730 5163.785 713.000 5188.000 ;
      LAYER met4 ;
        RECT 638.965 5083.400 712.035 5163.385 ;
        RECT 713.000 5083.400 895.000 5188.000 ;
      LAYER met4 ;
        RECT 895.000 5163.785 896.270 5188.000 ;
      LAYER met4 ;
        RECT 896.670 5163.385 968.330 5188.000 ;
      LAYER met4 ;
        RECT 968.730 5163.785 970.000 5188.000 ;
      LAYER met4 ;
        RECT 895.965 5083.400 969.035 5163.385 ;
        RECT 970.000 5083.400 1105.000 5188.000 ;
      LAYER met4 ;
        RECT 1105.000 5163.785 1153.205 5188.000 ;
      LAYER met4 ;
        RECT 1153.605 5163.385 1230.485 5188.000 ;
      LAYER met4 ;
        RECT 1230.885 5163.785 1274.000 5188.000 ;
      LAYER met4 ;
        RECT 1152.240 5083.400 1230.885 5163.385 ;
        RECT 1274.000 5083.400 1363.000 5188.000 ;
      LAYER met4 ;
        RECT 1363.000 5163.785 1411.205 5188.000 ;
      LAYER met4 ;
        RECT 1411.605 5163.385 1488.485 5188.000 ;
      LAYER met4 ;
        RECT 1488.885 5163.785 1532.000 5188.000 ;
      LAYER met4 ;
        RECT 1410.240 5083.400 1488.885 5163.385 ;
        RECT 1532.000 5083.400 1667.000 5188.000 ;
      LAYER met4 ;
        RECT 1667.000 5163.785 1668.270 5188.000 ;
      LAYER met4 ;
        RECT 1668.670 5163.385 1740.330 5188.000 ;
      LAYER met4 ;
        RECT 1740.730 5163.785 1742.000 5188.000 ;
      LAYER met4 ;
        RECT 1742.000 5163.785 1919.000 5188.000 ;
      LAYER met4 ;
        RECT 1919.000 5163.785 1920.270 5188.000 ;
      LAYER met4 ;
        RECT 1667.965 5083.400 1741.035 5163.385 ;
        RECT 1742.000 5083.400 1909.000 5163.785 ;
        RECT 1914.000 5083.400 1919.000 5163.785 ;
        RECT 1920.670 5163.385 1992.330 5188.000 ;
      LAYER met4 ;
        RECT 1992.730 5163.785 1994.000 5188.000 ;
      LAYER met4 ;
        RECT 1919.965 5083.400 1993.035 5163.385 ;
        RECT 1994.000 5083.400 2364.000 5188.000 ;
      LAYER met4 ;
        RECT 2364.000 5163.785 2365.270 5188.000 ;
      LAYER met4 ;
        RECT 2365.670 5163.385 2437.330 5188.000 ;
      LAYER met4 ;
        RECT 2437.730 5163.785 2439.000 5188.000 ;
      LAYER met4 ;
        RECT 2364.965 5083.400 2438.035 5163.385 ;
        RECT 2439.000 5083.400 2621.000 5188.000 ;
      LAYER met4 ;
        RECT 2621.000 5163.785 2622.270 5188.000 ;
      LAYER met4 ;
        RECT 2622.670 5163.385 2694.330 5188.000 ;
      LAYER met4 ;
        RECT 2694.730 5163.785 2696.000 5188.000 ;
      LAYER met4 ;
        RECT 2621.965 5083.400 2695.035 5163.385 ;
        RECT 2696.000 5083.400 2878.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.000 5163.785 2879.270 5188.000 ;
      LAYER met4 ;
        RECT 2879.670 5163.385 2951.330 5188.000 ;
      LAYER met4 ;
        RECT 2951.730 5163.785 2953.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.965 5083.400 2952.035 5163.385 ;
        RECT 2953.000 5083.400 3130.000 5188.000 ;
      LAYER met4 ;
        RECT 3130.000 5163.785 3131.270 5188.000 ;
      LAYER met4 ;
        RECT 3131.670 5163.385 3203.330 5188.000 ;
      LAYER met4 ;
        RECT 3203.730 5163.785 3205.000 5188.000 ;
      LAYER met4 ;
        RECT 3205.000 5163.385 3388.000 5188.000 ;
      LAYER met4 ;
        RECT 3388.000 5163.785 3389.435 5188.000 ;
      LAYER met4 ;
        RECT 3389.835 5163.385 3588.000 5188.000 ;
        RECT 3130.965 5083.400 3204.035 5163.385 ;
        RECT 3205.000 5083.400 3588.000 5163.385 ;
        RECT 0.000 5057.635 201.745 5083.400 ;
      LAYER met4 ;
        RECT 202.145 5058.035 382.270 5083.000 ;
      LAYER met4 ;
        RECT 382.670 5057.635 454.330 5083.400 ;
      LAYER met4 ;
        RECT 454.730 5058.035 639.270 5083.000 ;
      LAYER met4 ;
        RECT 639.670 5057.635 711.330 5083.400 ;
      LAYER met4 ;
        RECT 711.730 5058.035 896.270 5083.000 ;
      LAYER met4 ;
        RECT 896.670 5057.635 968.330 5083.400 ;
      LAYER met4 ;
        RECT 968.730 5058.035 1152.715 5083.000 ;
      LAYER met4 ;
        RECT 1153.115 5057.635 1230.485 5083.400 ;
      LAYER met4 ;
        RECT 1230.885 5058.035 1410.715 5083.000 ;
      LAYER met4 ;
        RECT 1411.115 5057.635 1488.485 5083.400 ;
      LAYER met4 ;
        RECT 1488.885 5058.035 1668.270 5083.000 ;
      LAYER met4 ;
        RECT 1668.670 5057.635 1740.330 5083.400 ;
      LAYER met4 ;
        RECT 1740.730 5058.035 1920.270 5083.000 ;
      LAYER met4 ;
        RECT 1920.670 5057.635 1992.330 5083.400 ;
      LAYER met4 ;
        RECT 1992.730 5058.035 2365.270 5083.000 ;
      LAYER met4 ;
        RECT 2365.670 5057.635 2437.330 5083.400 ;
      LAYER met4 ;
        RECT 2437.730 5058.035 2622.270 5083.000 ;
      LAYER met4 ;
        RECT 2622.670 5057.635 2694.330 5083.400 ;
      LAYER met4 ;
        RECT 2694.730 5058.035 2879.270 5083.000 ;
      LAYER met4 ;
        RECT 2879.670 5057.635 2951.330 5083.400 ;
      LAYER met4 ;
        RECT 2951.730 5058.035 3131.270 5083.000 ;
      LAYER met4 ;
        RECT 3131.670 5057.635 3203.330 5083.400 ;
      LAYER met4 ;
        RECT 3203.730 5058.035 3390.645 5083.000 ;
      LAYER met4 ;
        RECT 3391.045 5057.635 3588.000 5083.400 ;
        RECT 0.000 5056.935 202.745 5057.635 ;
        RECT 204.000 5056.935 381.000 5057.635 ;
        RECT 381.965 5056.935 455.035 5057.635 ;
        RECT 456.000 5056.935 638.000 5057.635 ;
        RECT 638.965 5056.935 712.035 5057.635 ;
        RECT 713.000 5056.935 895.000 5057.635 ;
        RECT 895.965 5056.935 969.035 5057.635 ;
        RECT 970.000 5056.935 1105.000 5057.635 ;
        RECT 1152.240 5056.935 1230.885 5057.635 ;
        RECT 1274.000 5056.935 1363.000 5057.635 ;
        RECT 1410.240 5056.935 1488.885 5057.635 ;
        RECT 1532.000 5056.935 1667.000 5057.635 ;
        RECT 1667.965 5056.935 1741.035 5057.635 ;
        RECT 1742.000 5056.935 1909.000 5057.635 ;
        RECT 1914.000 5056.935 1919.000 5057.635 ;
        RECT 1919.965 5056.935 1993.035 5057.635 ;
        RECT 1994.000 5056.935 2364.000 5057.635 ;
        RECT 2364.965 5056.935 2438.035 5057.635 ;
        RECT 2439.000 5056.935 2621.000 5057.635 ;
        RECT 2621.965 5056.935 2695.035 5057.635 ;
        RECT 2696.000 5056.935 2878.000 5057.635 ;
        RECT 2878.965 5056.935 2952.035 5057.635 ;
        RECT 2953.000 5056.935 3130.000 5057.635 ;
        RECT 3130.965 5056.935 3204.035 5057.635 ;
        RECT 3205.000 5056.935 3588.000 5057.635 ;
        RECT 0.000 5051.685 202.330 5056.935 ;
      LAYER met4 ;
        RECT 202.730 5052.085 382.270 5056.535 ;
      LAYER met4 ;
        RECT 382.670 5051.685 454.330 5056.935 ;
      LAYER met4 ;
        RECT 454.730 5052.085 639.270 5056.535 ;
      LAYER met4 ;
        RECT 639.670 5051.685 711.330 5056.935 ;
      LAYER met4 ;
        RECT 711.730 5052.085 896.270 5056.535 ;
      LAYER met4 ;
        RECT 896.670 5051.685 968.330 5056.935 ;
      LAYER met4 ;
        RECT 968.730 5052.085 1152.715 5056.535 ;
      LAYER met4 ;
        RECT 1153.115 5051.685 1230.485 5056.935 ;
      LAYER met4 ;
        RECT 1230.885 5052.085 1410.715 5056.535 ;
      LAYER met4 ;
        RECT 1411.115 5051.685 1488.485 5056.935 ;
      LAYER met4 ;
        RECT 1488.885 5052.085 1668.270 5056.535 ;
      LAYER met4 ;
        RECT 1668.670 5051.685 1740.330 5056.935 ;
      LAYER met4 ;
        RECT 1740.730 5052.085 1920.270 5056.535 ;
      LAYER met4 ;
        RECT 1920.670 5051.685 1992.330 5056.935 ;
      LAYER met4 ;
        RECT 1992.730 5052.085 2365.270 5056.535 ;
      LAYER met4 ;
        RECT 2365.670 5051.685 2437.330 5056.935 ;
      LAYER met4 ;
        RECT 2437.730 5052.085 2622.270 5056.535 ;
      LAYER met4 ;
        RECT 2622.670 5051.685 2694.330 5056.935 ;
      LAYER met4 ;
        RECT 2694.730 5052.085 2879.270 5056.535 ;
      LAYER met4 ;
        RECT 2879.670 5051.685 2951.330 5056.935 ;
      LAYER met4 ;
        RECT 2951.730 5052.085 3131.270 5056.535 ;
      LAYER met4 ;
        RECT 3131.670 5051.685 3203.330 5056.935 ;
      LAYER met4 ;
        RECT 3203.730 5052.085 3389.480 5056.535 ;
      LAYER met4 ;
        RECT 3389.880 5051.685 3588.000 5056.935 ;
        RECT 0.000 5051.085 202.745 5051.685 ;
        RECT 204.000 5051.085 381.000 5051.685 ;
        RECT 381.965 5051.085 455.035 5051.685 ;
        RECT 456.000 5051.085 638.000 5051.685 ;
        RECT 638.965 5051.085 712.035 5051.685 ;
        RECT 713.000 5051.085 895.000 5051.685 ;
        RECT 895.965 5051.085 969.035 5051.685 ;
        RECT 970.000 5051.085 1105.000 5051.685 ;
        RECT 1152.240 5051.085 1230.885 5051.685 ;
        RECT 1274.000 5051.085 1363.000 5051.685 ;
        RECT 1410.240 5051.085 1488.885 5051.685 ;
        RECT 1532.000 5051.085 1667.000 5051.685 ;
        RECT 1667.965 5051.085 1741.035 5051.685 ;
        RECT 1742.000 5051.085 1909.000 5051.685 ;
        RECT 1914.000 5051.085 1919.000 5051.685 ;
        RECT 1919.965 5051.085 1993.035 5051.685 ;
        RECT 1994.000 5051.085 2364.000 5051.685 ;
        RECT 2364.965 5051.085 2438.035 5051.685 ;
        RECT 2439.000 5051.085 2621.000 5051.685 ;
        RECT 2621.965 5051.085 2695.035 5051.685 ;
        RECT 2696.000 5051.085 2878.000 5051.685 ;
        RECT 2878.965 5051.085 2952.035 5051.685 ;
        RECT 2953.000 5051.085 3130.000 5051.685 ;
        RECT 3130.965 5051.085 3204.035 5051.685 ;
        RECT 3205.000 5051.085 3588.000 5051.685 ;
        RECT 0.000 5045.835 202.330 5051.085 ;
      LAYER met4 ;
        RECT 202.730 5046.235 382.270 5050.685 ;
      LAYER met4 ;
        RECT 382.670 5045.835 454.330 5051.085 ;
      LAYER met4 ;
        RECT 454.730 5046.235 639.270 5050.685 ;
      LAYER met4 ;
        RECT 639.670 5045.835 711.330 5051.085 ;
      LAYER met4 ;
        RECT 711.730 5046.235 896.270 5050.685 ;
      LAYER met4 ;
        RECT 896.670 5045.835 968.330 5051.085 ;
      LAYER met4 ;
        RECT 968.730 5046.235 1152.715 5050.685 ;
      LAYER met4 ;
        RECT 1153.115 5045.835 1230.485 5051.085 ;
      LAYER met4 ;
        RECT 1230.885 5046.235 1410.715 5050.685 ;
      LAYER met4 ;
        RECT 1411.115 5045.835 1488.485 5051.085 ;
      LAYER met4 ;
        RECT 1488.885 5046.235 1668.270 5050.685 ;
      LAYER met4 ;
        RECT 1668.670 5045.835 1740.330 5051.085 ;
      LAYER met4 ;
        RECT 1740.730 5046.235 1920.270 5050.685 ;
      LAYER met4 ;
        RECT 1920.670 5045.835 1992.330 5051.085 ;
      LAYER met4 ;
        RECT 1992.730 5046.235 2365.270 5050.685 ;
      LAYER met4 ;
        RECT 2365.670 5045.835 2437.330 5051.085 ;
      LAYER met4 ;
        RECT 2437.730 5046.235 2622.270 5050.685 ;
      LAYER met4 ;
        RECT 2622.670 5045.835 2694.330 5051.085 ;
      LAYER met4 ;
        RECT 2694.730 5046.235 2879.270 5050.685 ;
      LAYER met4 ;
        RECT 2879.670 5045.835 2951.330 5051.085 ;
      LAYER met4 ;
        RECT 2951.730 5046.235 3131.270 5050.685 ;
      LAYER met4 ;
        RECT 3131.670 5045.835 3203.330 5051.085 ;
      LAYER met4 ;
        RECT 3203.730 5046.235 3389.625 5050.685 ;
      LAYER met4 ;
        RECT 3390.025 5045.835 3588.000 5051.085 ;
        RECT 0.000 5045.135 202.745 5045.835 ;
        RECT 204.000 5045.135 381.000 5045.835 ;
        RECT 381.965 5045.135 455.035 5045.835 ;
        RECT 456.000 5045.135 638.000 5045.835 ;
        RECT 638.965 5045.135 712.035 5045.835 ;
        RECT 713.000 5045.135 895.000 5045.835 ;
        RECT 895.965 5045.135 969.035 5045.835 ;
        RECT 970.000 5045.135 1105.000 5045.835 ;
        RECT 1152.240 5045.135 1230.885 5045.835 ;
        RECT 1274.000 5045.135 1363.000 5045.835 ;
        RECT 1410.240 5045.135 1488.885 5045.835 ;
        RECT 1532.000 5045.135 1667.000 5045.835 ;
        RECT 1667.965 5045.135 1741.035 5045.835 ;
        RECT 1742.000 5045.135 1909.000 5045.835 ;
        RECT 1914.000 5045.135 1919.000 5045.835 ;
        RECT 1919.965 5045.135 1993.035 5045.835 ;
        RECT 1994.000 5045.135 2364.000 5045.835 ;
        RECT 2364.965 5045.135 2438.035 5045.835 ;
        RECT 2439.000 5045.135 2621.000 5045.835 ;
        RECT 2621.965 5045.135 2695.035 5045.835 ;
        RECT 2696.000 5045.135 2878.000 5045.835 ;
        RECT 2878.965 5045.135 2952.035 5045.835 ;
        RECT 2953.000 5045.135 3130.000 5045.835 ;
        RECT 3130.965 5045.135 3204.035 5045.835 ;
        RECT 3205.000 5045.135 3588.000 5045.835 ;
        RECT 0.000 5044.005 176.425 5045.135 ;
      LAYER met4 ;
        RECT 176.825 5044.405 1909.000 5044.735 ;
        RECT 1914.000 5044.405 2879.270 5044.735 ;
      LAYER met4 ;
        RECT 2879.670 5044.505 2951.330 5045.135 ;
      LAYER met4 ;
        RECT 2951.730 5044.405 3411.175 5044.735 ;
      LAYER met4 ;
        RECT 0.000 5040.725 176.690 5044.005 ;
      LAYER met4 ;
        RECT 177.090 5041.125 3410.910 5044.105 ;
      LAYER met4 ;
        RECT 3411.575 5044.005 3588.000 5045.135 ;
        RECT 0.000 5039.245 182.045 5040.725 ;
      LAYER met4 ;
        RECT 182.445 5039.645 204.000 5040.825 ;
      LAYER met4 ;
        RECT 204.000 5039.645 381.000 5040.825 ;
      LAYER met4 ;
        RECT 381.000 5039.645 382.270 5040.825 ;
      LAYER met4 ;
        RECT 382.670 5039.745 454.330 5040.725 ;
      LAYER met4 ;
        RECT 454.730 5039.645 456.000 5040.825 ;
      LAYER met4 ;
        RECT 456.000 5039.645 638.000 5040.825 ;
      LAYER met4 ;
        RECT 638.000 5039.645 639.270 5040.825 ;
      LAYER met4 ;
        RECT 639.670 5039.745 711.330 5040.725 ;
      LAYER met4 ;
        RECT 711.730 5039.645 713.000 5040.825 ;
      LAYER met4 ;
        RECT 713.000 5039.645 895.000 5040.825 ;
      LAYER met4 ;
        RECT 895.000 5039.645 896.270 5040.825 ;
      LAYER met4 ;
        RECT 896.670 5039.745 968.330 5040.725 ;
      LAYER met4 ;
        RECT 968.730 5039.645 970.000 5040.825 ;
      LAYER met4 ;
        RECT 970.000 5039.645 1105.000 5040.825 ;
      LAYER met4 ;
        RECT 1105.000 5039.645 1152.240 5040.825 ;
      LAYER met4 ;
        RECT 1152.640 5039.745 1230.485 5040.725 ;
      LAYER met4 ;
        RECT 1230.885 5039.645 1274.000 5040.825 ;
      LAYER met4 ;
        RECT 1274.000 5039.645 1363.000 5040.825 ;
      LAYER met4 ;
        RECT 1363.000 5039.645 1410.240 5040.825 ;
      LAYER met4 ;
        RECT 1410.640 5039.745 1488.485 5040.725 ;
      LAYER met4 ;
        RECT 1488.885 5039.645 1532.000 5040.825 ;
      LAYER met4 ;
        RECT 1532.000 5039.645 1667.000 5040.825 ;
      LAYER met4 ;
        RECT 1667.000 5039.645 1668.270 5040.825 ;
      LAYER met4 ;
        RECT 1668.670 5039.745 1740.330 5040.725 ;
      LAYER met4 ;
        RECT 1740.730 5039.645 1742.000 5040.825 ;
      LAYER met4 ;
        RECT 1742.000 5039.645 1909.000 5040.825 ;
        RECT 1914.000 5039.645 1919.000 5040.825 ;
      LAYER met4 ;
        RECT 1919.000 5039.645 1920.270 5040.825 ;
      LAYER met4 ;
        RECT 1920.670 5039.745 1992.330 5040.725 ;
      LAYER met4 ;
        RECT 1992.730 5039.645 1994.000 5040.825 ;
      LAYER met4 ;
        RECT 1994.000 5039.645 2364.000 5040.825 ;
      LAYER met4 ;
        RECT 2364.000 5039.645 2365.270 5040.825 ;
      LAYER met4 ;
        RECT 2365.670 5039.745 2437.330 5040.725 ;
      LAYER met4 ;
        RECT 2437.730 5039.645 2439.000 5040.825 ;
      LAYER met4 ;
        RECT 2439.000 5039.645 2621.000 5040.825 ;
      LAYER met4 ;
        RECT 2621.000 5039.645 2622.270 5040.825 ;
      LAYER met4 ;
        RECT 2622.670 5039.745 2694.330 5040.725 ;
      LAYER met4 ;
        RECT 2694.730 5039.645 2696.000 5040.825 ;
      LAYER met4 ;
        RECT 2696.000 5039.645 2878.000 5040.825 ;
      LAYER met4 ;
        RECT 2878.000 5039.645 2879.270 5040.825 ;
      LAYER met4 ;
        RECT 2879.670 5039.745 2951.330 5040.725 ;
      LAYER met4 ;
        RECT 2951.730 5039.645 2953.000 5040.825 ;
      LAYER met4 ;
        RECT 2953.000 5039.645 3130.000 5040.825 ;
      LAYER met4 ;
        RECT 3130.000 5039.645 3131.270 5040.825 ;
      LAYER met4 ;
        RECT 3131.670 5039.745 3203.330 5040.725 ;
      LAYER met4 ;
        RECT 3203.730 5039.645 3205.000 5040.825 ;
      LAYER met4 ;
        RECT 3205.000 5039.645 3388.000 5040.825 ;
      LAYER met4 ;
        RECT 3388.000 5039.645 3409.550 5040.825 ;
      LAYER met4 ;
        RECT 3411.310 5040.725 3588.000 5044.005 ;
        RECT 0.000 5036.465 182.725 5039.245 ;
        RECT 0.000 5035.335 180.025 5036.465 ;
      LAYER met4 ;
        RECT 183.125 5036.365 3408.935 5039.345 ;
      LAYER met4 ;
        RECT 3409.950 5039.245 3588.000 5040.725 ;
      LAYER met4 ;
        RECT 180.425 5035.735 1909.000 5036.065 ;
        RECT 1914.000 5035.735 2879.270 5036.065 ;
      LAYER met4 ;
        RECT 2879.670 5035.335 2951.330 5035.965 ;
      LAYER met4 ;
        RECT 2951.730 5035.735 3407.575 5036.065 ;
      LAYER met4 ;
        RECT 3409.335 5035.965 3588.000 5039.245 ;
        RECT 3407.975 5035.335 3588.000 5035.965 ;
        RECT 0.000 5034.635 202.745 5035.335 ;
        RECT 381.965 5034.635 455.035 5035.335 ;
        RECT 638.965 5034.635 712.035 5035.335 ;
        RECT 895.965 5034.635 969.035 5035.335 ;
        RECT 1152.240 5034.635 1230.885 5035.335 ;
        RECT 1410.240 5034.635 1488.885 5035.335 ;
        RECT 1667.965 5034.635 1741.035 5035.335 ;
        RECT 1919.965 5034.635 1993.035 5035.335 ;
        RECT 2364.965 5034.635 2438.035 5035.335 ;
        RECT 2621.965 5034.635 2695.035 5035.335 ;
        RECT 2878.965 5034.635 2952.035 5035.335 ;
        RECT 3130.965 5034.635 3204.035 5035.335 ;
        RECT 3388.000 5034.635 3588.000 5035.335 ;
        RECT 0.000 5029.185 202.330 5034.635 ;
      LAYER met4 ;
        RECT 202.730 5029.585 382.270 5034.235 ;
      LAYER met4 ;
        RECT 382.670 5029.185 454.330 5034.635 ;
      LAYER met4 ;
        RECT 454.730 5029.585 639.270 5034.235 ;
      LAYER met4 ;
        RECT 639.670 5029.185 711.330 5034.635 ;
      LAYER met4 ;
        RECT 711.730 5029.585 896.270 5034.235 ;
      LAYER met4 ;
        RECT 896.670 5029.185 968.330 5034.635 ;
      LAYER met4 ;
        RECT 968.730 5029.585 1152.250 5034.235 ;
      LAYER met4 ;
        RECT 1152.650 5029.185 1230.485 5034.635 ;
      LAYER met4 ;
        RECT 1230.885 5029.585 1410.250 5034.235 ;
      LAYER met4 ;
        RECT 1410.650 5029.185 1488.485 5034.635 ;
      LAYER met4 ;
        RECT 1488.885 5029.585 1668.270 5034.235 ;
      LAYER met4 ;
        RECT 1668.670 5029.185 1740.330 5034.635 ;
      LAYER met4 ;
        RECT 1740.730 5029.585 1914.000 5034.235 ;
        RECT 1919.000 5029.585 1920.270 5034.235 ;
      LAYER met4 ;
        RECT 1920.670 5029.185 1992.330 5034.635 ;
      LAYER met4 ;
        RECT 1992.730 5029.585 2365.270 5034.235 ;
      LAYER met4 ;
        RECT 2365.670 5029.185 2437.330 5034.635 ;
      LAYER met4 ;
        RECT 2437.730 5029.585 2622.270 5034.235 ;
      LAYER met4 ;
        RECT 2622.670 5029.185 2694.330 5034.635 ;
      LAYER met4 ;
        RECT 2694.730 5029.585 2879.270 5034.235 ;
      LAYER met4 ;
        RECT 2879.670 5029.185 2951.330 5034.635 ;
      LAYER met4 ;
        RECT 2951.730 5029.585 3131.270 5034.235 ;
      LAYER met4 ;
        RECT 3131.670 5029.185 3203.330 5034.635 ;
      LAYER met4 ;
        RECT 3203.730 5029.585 3389.475 5034.235 ;
      LAYER met4 ;
        RECT 3389.875 5029.185 3588.000 5034.635 ;
        RECT 0.000 5028.585 202.745 5029.185 ;
        RECT 381.965 5028.585 455.035 5029.185 ;
        RECT 638.965 5028.585 712.035 5029.185 ;
        RECT 895.965 5028.585 969.035 5029.185 ;
        RECT 1152.240 5028.585 1230.885 5029.185 ;
        RECT 1410.240 5028.585 1488.885 5029.185 ;
        RECT 1667.965 5028.585 1741.035 5029.185 ;
        RECT 1919.965 5028.585 1993.035 5029.185 ;
        RECT 2364.965 5028.585 2438.035 5029.185 ;
        RECT 2621.965 5028.585 2695.035 5029.185 ;
        RECT 2878.965 5028.585 2952.035 5029.185 ;
        RECT 3130.965 5028.585 3204.035 5029.185 ;
        RECT 3388.000 5028.585 3588.000 5029.185 ;
        RECT 0.000 5024.335 202.330 5028.585 ;
      LAYER met4 ;
        RECT 202.730 5024.735 382.270 5028.185 ;
      LAYER met4 ;
        RECT 382.670 5024.335 454.330 5028.585 ;
      LAYER met4 ;
        RECT 454.730 5024.735 639.270 5028.185 ;
      LAYER met4 ;
        RECT 639.670 5024.335 711.330 5028.585 ;
      LAYER met4 ;
        RECT 711.730 5024.735 896.270 5028.185 ;
      LAYER met4 ;
        RECT 896.670 5024.335 968.330 5028.585 ;
      LAYER met4 ;
        RECT 968.730 5024.735 1152.715 5028.185 ;
      LAYER met4 ;
        RECT 1153.115 5024.335 1230.485 5028.585 ;
      LAYER met4 ;
        RECT 1230.885 5024.735 1410.715 5028.185 ;
      LAYER met4 ;
        RECT 1411.115 5024.335 1488.485 5028.585 ;
      LAYER met4 ;
        RECT 1488.885 5024.735 1668.270 5028.185 ;
      LAYER met4 ;
        RECT 1668.670 5024.335 1740.330 5028.585 ;
      LAYER met4 ;
        RECT 1740.730 5024.735 1909.000 5028.185 ;
        RECT 1914.000 5024.735 1920.270 5028.185 ;
      LAYER met4 ;
        RECT 1920.670 5024.335 1992.330 5028.585 ;
      LAYER met4 ;
        RECT 1992.730 5024.735 2365.270 5028.185 ;
      LAYER met4 ;
        RECT 2365.670 5024.335 2437.330 5028.585 ;
      LAYER met4 ;
        RECT 2437.730 5024.735 2622.270 5028.185 ;
      LAYER met4 ;
        RECT 2622.670 5024.335 2694.330 5028.585 ;
      LAYER met4 ;
        RECT 2694.730 5024.735 2879.270 5028.185 ;
      LAYER met4 ;
        RECT 2879.670 5024.335 2951.330 5028.585 ;
      LAYER met4 ;
        RECT 2951.730 5024.735 3131.270 5028.185 ;
      LAYER met4 ;
        RECT 3131.670 5024.335 3203.330 5028.585 ;
      LAYER met4 ;
        RECT 3203.730 5024.735 3389.335 5028.185 ;
      LAYER met4 ;
        RECT 3389.735 5024.335 3588.000 5028.585 ;
        RECT 0.000 5023.735 202.745 5024.335 ;
        RECT 381.965 5023.735 455.035 5024.335 ;
        RECT 638.965 5023.735 712.035 5024.335 ;
        RECT 895.965 5023.735 969.035 5024.335 ;
        RECT 1152.240 5023.735 1230.885 5024.335 ;
        RECT 1410.240 5023.735 1488.885 5024.335 ;
        RECT 1667.965 5023.735 1741.035 5024.335 ;
        RECT 1919.965 5023.735 1993.035 5024.335 ;
        RECT 2364.965 5023.735 2438.035 5024.335 ;
        RECT 2621.965 5023.735 2695.035 5024.335 ;
        RECT 2878.965 5023.735 2952.035 5024.335 ;
        RECT 3130.965 5023.735 3204.035 5024.335 ;
        RECT 3388.000 5023.735 3588.000 5024.335 ;
        RECT 0.000 5019.485 202.330 5023.735 ;
      LAYER met4 ;
        RECT 202.730 5019.885 382.270 5023.335 ;
      LAYER met4 ;
        RECT 382.670 5019.485 454.330 5023.735 ;
      LAYER met4 ;
        RECT 454.730 5019.885 639.270 5023.335 ;
      LAYER met4 ;
        RECT 639.670 5019.485 711.330 5023.735 ;
      LAYER met4 ;
        RECT 711.730 5019.885 896.270 5023.335 ;
      LAYER met4 ;
        RECT 896.670 5019.485 968.330 5023.735 ;
      LAYER met4 ;
        RECT 968.730 5019.885 1152.715 5023.335 ;
      LAYER met4 ;
        RECT 1153.115 5019.485 1230.485 5023.735 ;
      LAYER met4 ;
        RECT 1230.885 5019.885 1410.715 5023.335 ;
      LAYER met4 ;
        RECT 1411.115 5019.485 1488.485 5023.735 ;
      LAYER met4 ;
        RECT 1488.885 5019.885 1668.270 5023.335 ;
      LAYER met4 ;
        RECT 1668.670 5019.485 1740.330 5023.735 ;
      LAYER met4 ;
        RECT 1740.730 5019.885 1920.270 5023.335 ;
      LAYER met4 ;
        RECT 1920.670 5019.485 1992.330 5023.735 ;
      LAYER met4 ;
        RECT 1992.730 5019.885 2365.270 5023.335 ;
      LAYER met4 ;
        RECT 2365.670 5019.485 2437.330 5023.735 ;
      LAYER met4 ;
        RECT 2437.730 5019.885 2622.270 5023.335 ;
      LAYER met4 ;
        RECT 2622.670 5019.485 2694.330 5023.735 ;
      LAYER met4 ;
        RECT 2694.730 5019.885 2879.270 5023.335 ;
      LAYER met4 ;
        RECT 2879.670 5019.485 2951.330 5023.735 ;
      LAYER met4 ;
        RECT 2951.730 5019.885 3131.270 5023.335 ;
      LAYER met4 ;
        RECT 3131.670 5019.485 3203.330 5023.735 ;
      LAYER met4 ;
        RECT 3203.730 5019.885 3389.385 5023.335 ;
      LAYER met4 ;
        RECT 3389.785 5019.485 3588.000 5023.735 ;
        RECT 0.000 5018.885 202.745 5019.485 ;
        RECT 381.965 5018.885 455.035 5019.485 ;
        RECT 638.965 5018.885 712.035 5019.485 ;
        RECT 895.965 5018.885 969.035 5019.485 ;
        RECT 1152.240 5018.885 1230.885 5019.485 ;
        RECT 1410.240 5018.885 1488.885 5019.485 ;
        RECT 1667.965 5018.885 1741.035 5019.485 ;
        RECT 1919.965 5018.885 1993.035 5019.485 ;
        RECT 2364.965 5018.885 2438.035 5019.485 ;
        RECT 2621.965 5018.885 2695.035 5019.485 ;
        RECT 2878.965 5018.885 2952.035 5019.485 ;
        RECT 3130.965 5018.885 3204.035 5019.485 ;
        RECT 3388.000 5018.885 3588.000 5019.485 ;
        RECT 0.000 5013.435 202.330 5018.885 ;
      LAYER met4 ;
        RECT 202.730 5013.835 382.270 5018.485 ;
      LAYER met4 ;
        RECT 382.670 5013.435 454.330 5018.885 ;
      LAYER met4 ;
        RECT 454.730 5013.835 639.270 5018.485 ;
      LAYER met4 ;
        RECT 639.670 5013.435 711.330 5018.885 ;
      LAYER met4 ;
        RECT 711.730 5013.835 896.270 5018.485 ;
      LAYER met4 ;
        RECT 896.670 5013.435 968.330 5018.885 ;
      LAYER met4 ;
        RECT 968.730 5013.835 1152.715 5018.485 ;
      LAYER met4 ;
        RECT 1153.115 5013.435 1230.485 5018.885 ;
      LAYER met4 ;
        RECT 1230.885 5013.835 1410.715 5018.485 ;
      LAYER met4 ;
        RECT 1411.115 5013.435 1488.485 5018.885 ;
      LAYER met4 ;
        RECT 1488.885 5013.835 1668.270 5018.485 ;
      LAYER met4 ;
        RECT 1668.670 5013.435 1740.330 5018.885 ;
      LAYER met4 ;
        RECT 1740.730 5013.835 1920.270 5018.485 ;
      LAYER met4 ;
        RECT 1920.670 5013.435 1992.330 5018.885 ;
      LAYER met4 ;
        RECT 1992.730 5013.835 2365.270 5018.485 ;
      LAYER met4 ;
        RECT 2365.670 5013.435 2437.330 5018.885 ;
      LAYER met4 ;
        RECT 2437.730 5013.835 2622.270 5018.485 ;
      LAYER met4 ;
        RECT 2622.670 5013.435 2694.330 5018.885 ;
      LAYER met4 ;
        RECT 2694.730 5013.835 2879.270 5018.485 ;
      LAYER met4 ;
        RECT 2879.670 5013.435 2951.330 5018.885 ;
      LAYER met4 ;
        RECT 2951.730 5013.835 3131.270 5018.485 ;
      LAYER met4 ;
        RECT 3131.670 5013.435 3203.330 5018.885 ;
      LAYER met4 ;
        RECT 3203.730 5013.835 3389.600 5018.485 ;
      LAYER met4 ;
        RECT 3390.000 5013.435 3588.000 5018.885 ;
        RECT 0.000 5012.835 202.745 5013.435 ;
        RECT 381.965 5012.835 455.035 5013.435 ;
        RECT 638.965 5012.835 712.035 5013.435 ;
        RECT 895.965 5012.835 969.035 5013.435 ;
        RECT 1152.240 5012.835 1230.885 5013.435 ;
        RECT 1410.240 5012.835 1488.885 5013.435 ;
        RECT 1667.965 5012.835 1741.035 5013.435 ;
        RECT 1919.965 5012.835 1993.035 5013.435 ;
        RECT 2364.965 5012.835 2438.035 5013.435 ;
        RECT 2621.965 5012.835 2695.035 5013.435 ;
        RECT 2878.965 5012.835 2952.035 5013.435 ;
        RECT 3130.965 5012.835 3204.035 5013.435 ;
        RECT 3388.000 5012.835 3588.000 5013.435 ;
        RECT 0.000 5011.575 202.330 5012.835 ;
        RECT 0.000 4991.045 142.865 5011.575 ;
        RECT 143.995 5011.310 202.330 5011.575 ;
        RECT 0.000 4989.835 104.600 4991.045 ;
      LAYER met4 ;
        RECT 0.000 4988.000 24.215 4989.435 ;
      LAYER met4 ;
        RECT 24.615 4988.000 104.600 4989.835 ;
        RECT 0.000 4846.000 104.600 4988.000 ;
      LAYER met4 ;
        RECT 0.000 4844.730 24.215 4846.000 ;
      LAYER met4 ;
        RECT 24.615 4844.330 104.600 4845.035 ;
      LAYER met4 ;
        RECT 105.000 4844.730 129.965 4990.645 ;
      LAYER met4 ;
        RECT 130.365 4990.025 142.865 4991.045 ;
        RECT 130.365 4989.880 136.915 4990.025 ;
        RECT 130.365 4846.000 131.065 4989.880 ;
        RECT 130.365 4844.330 131.065 4845.035 ;
      LAYER met4 ;
        RECT 131.465 4844.730 135.915 4989.480 ;
      LAYER met4 ;
        RECT 136.315 4846.000 136.915 4989.880 ;
        RECT 136.315 4844.330 136.915 4845.035 ;
      LAYER met4 ;
        RECT 137.315 4844.730 141.765 4989.625 ;
      LAYER met4 ;
        RECT 142.165 4846.000 142.865 4990.025 ;
        RECT 142.165 4844.330 142.865 4845.035 ;
        RECT 0.000 4772.670 142.865 4844.330 ;
      LAYER met4 ;
        RECT 0.000 4771.000 24.215 4772.270 ;
      LAYER met4 ;
        RECT 24.615 4771.965 104.600 4772.670 ;
        RECT 0.000 4635.000 104.600 4771.000 ;
      LAYER met4 ;
        RECT 0.000 4633.730 24.215 4635.000 ;
      LAYER met4 ;
        RECT 24.215 4634.785 24.250 4635.000 ;
        RECT 24.615 4633.330 104.600 4635.000 ;
      LAYER met4 ;
        RECT 105.000 4633.730 129.965 4772.270 ;
      LAYER met4 ;
        RECT 130.365 4771.965 131.065 4772.670 ;
        RECT 130.365 4633.330 131.065 4771.000 ;
      LAYER met4 ;
        RECT 131.465 4633.730 135.915 4772.270 ;
      LAYER met4 ;
        RECT 136.315 4771.965 136.915 4772.670 ;
        RECT 136.315 4633.330 136.915 4771.000 ;
      LAYER met4 ;
        RECT 137.315 4633.730 141.765 4772.270 ;
      LAYER met4 ;
        RECT 142.165 4771.965 142.865 4772.670 ;
        RECT 142.165 4633.330 142.865 4771.000 ;
        RECT 0.000 4561.670 142.865 4633.330 ;
      LAYER met4 ;
        RECT 0.000 4560.000 24.215 4561.270 ;
      LAYER met4 ;
        RECT 24.615 4560.000 104.600 4561.670 ;
        RECT 0.000 4424.000 104.600 4560.000 ;
      LAYER met4 ;
        RECT 0.000 4422.730 24.215 4424.000 ;
      LAYER met4 ;
        RECT 24.615 4422.330 104.600 4423.035 ;
      LAYER met4 ;
        RECT 105.000 4422.730 129.965 4561.270 ;
      LAYER met4 ;
        RECT 130.365 4424.000 131.065 4561.670 ;
        RECT 130.365 4422.330 131.065 4423.035 ;
      LAYER met4 ;
        RECT 131.465 4422.730 135.915 4561.270 ;
      LAYER met4 ;
        RECT 136.315 4424.000 136.915 4561.670 ;
        RECT 136.315 4422.330 136.915 4423.035 ;
      LAYER met4 ;
        RECT 137.315 4422.730 141.765 4561.270 ;
      LAYER met4 ;
        RECT 142.165 4424.000 142.865 4561.670 ;
        RECT 142.165 4422.330 142.865 4423.035 ;
        RECT 0.000 4350.670 142.865 4422.330 ;
      LAYER met4 ;
        RECT 0.000 4349.000 24.215 4350.270 ;
      LAYER met4 ;
        RECT 24.615 4349.965 104.600 4350.670 ;
        RECT 0.000 4213.000 104.600 4349.000 ;
      LAYER met4 ;
        RECT 0.000 4211.730 24.215 4213.000 ;
      LAYER met4 ;
        RECT 24.615 4211.330 104.600 4212.035 ;
      LAYER met4 ;
        RECT 105.000 4211.730 129.965 4350.270 ;
      LAYER met4 ;
        RECT 130.365 4349.965 131.065 4350.670 ;
        RECT 130.365 4213.000 131.065 4349.000 ;
        RECT 130.365 4211.330 131.065 4212.035 ;
      LAYER met4 ;
        RECT 131.465 4211.730 135.915 4350.270 ;
      LAYER met4 ;
        RECT 136.315 4349.965 136.915 4350.670 ;
        RECT 136.315 4213.000 136.915 4349.000 ;
        RECT 136.315 4211.330 136.915 4212.035 ;
      LAYER met4 ;
        RECT 137.315 4211.730 141.765 4350.270 ;
      LAYER met4 ;
        RECT 142.165 4349.965 142.865 4350.670 ;
        RECT 142.165 4213.000 142.865 4349.000 ;
        RECT 142.165 4211.330 142.865 4212.035 ;
      LAYER met4 ;
        RECT 143.265 4211.730 143.595 5011.175 ;
      LAYER met4 ;
        RECT 0.000 4139.670 143.495 4211.330 ;
      LAYER met4 ;
        RECT 0.000 4138.000 24.215 4139.270 ;
      LAYER met4 ;
        RECT 24.615 4138.965 104.600 4139.670 ;
        RECT 0.000 4002.000 104.600 4138.000 ;
      LAYER met4 ;
        RECT 0.000 4000.730 24.215 4002.000 ;
      LAYER met4 ;
        RECT 24.615 4000.330 104.600 4000.970 ;
      LAYER met4 ;
        RECT 105.000 4000.730 129.965 4139.270 ;
      LAYER met4 ;
        RECT 130.365 4138.965 131.065 4139.670 ;
        RECT 130.365 4002.000 131.065 4138.000 ;
        RECT 130.365 4000.330 131.065 4000.970 ;
      LAYER met4 ;
        RECT 131.465 4000.730 135.915 4139.270 ;
      LAYER met4 ;
        RECT 136.315 4138.965 136.915 4139.670 ;
        RECT 136.315 4002.000 136.915 4138.000 ;
        RECT 136.315 4000.330 136.915 4000.970 ;
      LAYER met4 ;
        RECT 137.315 4000.730 141.765 4139.270 ;
      LAYER met4 ;
        RECT 142.165 4138.965 142.865 4139.670 ;
        RECT 142.165 4002.000 142.865 4138.000 ;
        RECT 142.165 4000.330 142.865 4000.970 ;
        RECT 0.000 3968.690 142.865 4000.330 ;
      LAYER met4 ;
        RECT 143.265 3969.090 143.595 4139.270 ;
      LAYER met4 ;
        RECT 0.000 3960.360 143.495 3968.690 ;
      LAYER met4 ;
        RECT 143.895 3960.760 146.875 5010.910 ;
      LAYER met4 ;
        RECT 147.275 5009.950 202.330 5011.310 ;
      LAYER met4 ;
        RECT 147.175 4988.000 148.355 5009.550 ;
      LAYER met4 ;
        RECT 148.755 5009.335 202.330 5009.950 ;
        RECT 147.175 4846.000 148.355 4988.000 ;
      LAYER met4 ;
        RECT 147.175 4844.730 148.355 4846.000 ;
      LAYER met4 ;
        RECT 147.275 4772.670 148.255 4844.330 ;
      LAYER met4 ;
        RECT 147.175 4771.000 148.355 4772.270 ;
      LAYER met4 ;
        RECT 147.175 4635.000 148.355 4771.000 ;
      LAYER met4 ;
        RECT 147.175 4633.730 148.355 4635.000 ;
      LAYER met4 ;
        RECT 147.275 4561.670 148.255 4633.330 ;
      LAYER met4 ;
        RECT 147.175 4560.000 148.355 4561.270 ;
      LAYER met4 ;
        RECT 147.175 4424.000 148.355 4560.000 ;
      LAYER met4 ;
        RECT 147.175 4422.730 148.355 4424.000 ;
      LAYER met4 ;
        RECT 147.275 4350.670 148.255 4422.330 ;
      LAYER met4 ;
        RECT 147.175 4349.000 148.355 4350.270 ;
      LAYER met4 ;
        RECT 147.175 4213.000 148.355 4349.000 ;
      LAYER met4 ;
        RECT 147.175 4211.730 148.355 4213.000 ;
      LAYER met4 ;
        RECT 147.275 4139.670 148.255 4211.330 ;
      LAYER met4 ;
        RECT 147.175 4138.000 148.355 4139.270 ;
      LAYER met4 ;
        RECT 147.175 4002.000 148.355 4138.000 ;
      LAYER met4 ;
        RECT 147.175 4000.730 148.355 4002.000 ;
      LAYER met4 ;
        RECT 147.275 3976.065 148.255 4000.330 ;
      LAYER met4 ;
        RECT 148.655 3976.465 151.635 5008.935 ;
      LAYER met4 ;
        RECT 152.035 5007.975 202.330 5009.335 ;
      LAYER met4 ;
        RECT 151.935 4211.730 152.265 5007.575 ;
      LAYER met4 ;
        RECT 152.665 5007.385 202.330 5007.975 ;
      LAYER met4 ;
        RECT 202.730 5007.785 382.270 5012.435 ;
      LAYER met4 ;
        RECT 382.670 5007.385 454.330 5012.835 ;
      LAYER met4 ;
        RECT 454.730 5007.785 639.270 5012.435 ;
      LAYER met4 ;
        RECT 639.670 5007.385 711.330 5012.835 ;
      LAYER met4 ;
        RECT 711.730 5007.785 896.270 5012.435 ;
      LAYER met4 ;
        RECT 896.670 5007.385 968.330 5012.835 ;
      LAYER met4 ;
        RECT 968.730 5007.785 1152.715 5012.435 ;
      LAYER met4 ;
        RECT 1153.115 5007.385 1225.805 5012.835 ;
      LAYER met4 ;
        RECT 1226.205 5007.785 1410.715 5012.435 ;
      LAYER met4 ;
        RECT 1411.115 5007.385 1483.805 5012.835 ;
      LAYER met4 ;
        RECT 1484.205 5007.785 1668.270 5012.435 ;
      LAYER met4 ;
        RECT 1668.670 5007.385 1740.330 5012.835 ;
      LAYER met4 ;
        RECT 1740.730 5007.785 1920.270 5012.435 ;
      LAYER met4 ;
        RECT 1920.670 5007.385 1992.330 5012.835 ;
      LAYER met4 ;
        RECT 1992.730 5007.785 2365.270 5012.435 ;
      LAYER met4 ;
        RECT 2365.670 5007.385 2437.330 5012.835 ;
      LAYER met4 ;
        RECT 2437.730 5007.785 2622.270 5012.435 ;
      LAYER met4 ;
        RECT 2622.670 5007.385 2694.330 5012.835 ;
      LAYER met4 ;
        RECT 2694.730 5007.785 2879.270 5012.435 ;
      LAYER met4 ;
        RECT 2879.670 5007.385 2951.330 5012.835 ;
      LAYER met4 ;
        RECT 2951.730 5007.785 3131.270 5012.435 ;
      LAYER met4 ;
        RECT 3131.670 5007.385 3203.330 5012.835 ;
      LAYER met4 ;
        RECT 3203.730 5007.785 3389.525 5012.435 ;
      LAYER met4 ;
        RECT 3389.925 5011.575 3588.000 5012.835 ;
        RECT 3389.925 5011.310 3444.005 5011.575 ;
        RECT 3389.925 5007.975 3440.725 5011.310 ;
        RECT 3389.925 5007.385 3435.335 5007.975 ;
        RECT 152.665 5006.785 202.745 5007.385 ;
        RECT 381.965 5006.785 455.035 5007.385 ;
        RECT 638.965 5006.785 712.035 5007.385 ;
        RECT 895.965 5006.785 969.035 5007.385 ;
        RECT 1152.240 5006.785 1230.885 5007.385 ;
        RECT 1410.240 5006.785 1488.885 5007.385 ;
        RECT 1667.965 5006.785 1741.035 5007.385 ;
        RECT 1919.965 5006.785 1993.035 5007.385 ;
        RECT 2364.965 5006.785 2438.035 5007.385 ;
        RECT 2621.965 5006.785 2695.035 5007.385 ;
        RECT 2878.965 5006.785 2952.035 5007.385 ;
        RECT 3130.965 5006.785 3204.035 5007.385 ;
        RECT 3388.000 5006.785 3435.335 5007.385 ;
        RECT 152.665 5002.535 202.345 5006.785 ;
      LAYER met4 ;
        RECT 202.745 5002.935 381.965 5006.385 ;
      LAYER met4 ;
        RECT 382.365 5002.535 454.635 5006.785 ;
      LAYER met4 ;
        RECT 455.035 5002.935 638.965 5006.385 ;
      LAYER met4 ;
        RECT 639.365 5002.535 711.635 5006.785 ;
      LAYER met4 ;
        RECT 712.035 5002.935 895.965 5006.385 ;
      LAYER met4 ;
        RECT 896.365 5002.535 968.635 5006.785 ;
      LAYER met4 ;
        RECT 969.035 5002.935 1152.715 5006.385 ;
      LAYER met4 ;
        RECT 1153.115 5002.535 1225.805 5006.785 ;
      LAYER met4 ;
        RECT 1226.205 5002.935 1410.715 5006.385 ;
      LAYER met4 ;
        RECT 1411.115 5002.535 1483.805 5006.785 ;
      LAYER met4 ;
        RECT 1484.205 5002.935 1667.965 5006.385 ;
      LAYER met4 ;
        RECT 1668.365 5002.535 1740.635 5006.785 ;
      LAYER met4 ;
        RECT 1741.035 5002.935 1909.000 5006.385 ;
        RECT 1914.000 5002.935 1919.965 5006.385 ;
      LAYER met4 ;
        RECT 1920.365 5002.535 1992.635 5006.785 ;
      LAYER met4 ;
        RECT 1993.035 5002.935 2364.965 5006.385 ;
      LAYER met4 ;
        RECT 2365.365 5002.535 2437.635 5006.785 ;
      LAYER met4 ;
        RECT 2438.035 5002.935 2621.965 5006.385 ;
      LAYER met4 ;
        RECT 2622.365 5002.535 2694.635 5006.785 ;
      LAYER met4 ;
        RECT 2695.035 5002.935 2878.965 5006.385 ;
      LAYER met4 ;
        RECT 2879.365 5002.535 2951.635 5006.785 ;
      LAYER met4 ;
        RECT 2952.035 5002.935 3130.965 5006.385 ;
      LAYER met4 ;
        RECT 3131.365 5002.535 3203.635 5006.785 ;
      LAYER met4 ;
        RECT 3204.035 5002.935 3389.470 5006.385 ;
      LAYER met4 ;
        RECT 3389.870 5002.535 3435.335 5006.785 ;
        RECT 152.665 5001.935 202.745 5002.535 ;
        RECT 381.965 5001.935 455.035 5002.535 ;
        RECT 638.965 5001.935 712.035 5002.535 ;
        RECT 895.965 5001.935 969.035 5002.535 ;
        RECT 1152.240 5001.935 1230.885 5002.535 ;
        RECT 1410.240 5001.935 1488.885 5002.535 ;
        RECT 1667.965 5001.935 1741.035 5002.535 ;
        RECT 1919.965 5001.935 1993.035 5002.535 ;
        RECT 2364.965 5001.935 2438.035 5002.535 ;
        RECT 2621.965 5001.935 2695.035 5002.535 ;
        RECT 2878.965 5001.935 2952.035 5002.535 ;
        RECT 3130.965 5001.935 3204.035 5002.535 ;
        RECT 3388.000 5001.935 3435.335 5002.535 ;
        RECT 152.665 4996.485 202.330 5001.935 ;
      LAYER met4 ;
        RECT 202.730 4996.885 382.270 5001.535 ;
      LAYER met4 ;
        RECT 382.670 4996.485 454.330 5001.935 ;
      LAYER met4 ;
        RECT 454.730 4996.885 639.270 5001.535 ;
      LAYER met4 ;
        RECT 639.670 4996.485 711.330 5001.935 ;
      LAYER met4 ;
        RECT 711.730 4996.885 896.270 5001.535 ;
      LAYER met4 ;
        RECT 896.670 4996.485 968.330 5001.935 ;
      LAYER met4 ;
        RECT 968.730 4996.885 1152.715 5001.535 ;
      LAYER met4 ;
        RECT 1153.115 4996.485 1230.485 5001.935 ;
      LAYER met4 ;
        RECT 1230.885 4996.885 1410.715 5001.535 ;
      LAYER met4 ;
        RECT 1411.115 4996.485 1488.485 5001.935 ;
      LAYER met4 ;
        RECT 1488.885 4996.885 1668.270 5001.535 ;
      LAYER met4 ;
        RECT 1668.670 4996.485 1740.330 5001.935 ;
      LAYER met4 ;
        RECT 1740.730 4996.885 1914.000 5001.535 ;
        RECT 1919.000 4996.885 1920.270 5001.535 ;
      LAYER met4 ;
        RECT 1920.670 4996.485 1992.330 5001.935 ;
      LAYER met4 ;
        RECT 1992.730 4996.885 2365.270 5001.535 ;
      LAYER met4 ;
        RECT 2365.670 4996.485 2437.330 5001.935 ;
      LAYER met4 ;
        RECT 2437.730 4996.885 2622.270 5001.535 ;
      LAYER met4 ;
        RECT 2622.670 4996.485 2694.330 5001.935 ;
      LAYER met4 ;
        RECT 2694.730 4996.885 2879.270 5001.535 ;
      LAYER met4 ;
        RECT 2879.670 4996.485 2951.330 5001.935 ;
      LAYER met4 ;
        RECT 2951.730 4996.885 3131.270 5001.535 ;
      LAYER met4 ;
        RECT 3131.670 4996.485 3203.330 5001.935 ;
      LAYER met4 ;
        RECT 3203.730 4996.885 3391.785 5001.535 ;
      LAYER met4 ;
        RECT 3392.185 4996.485 3435.335 5001.935 ;
        RECT 152.665 4995.885 202.745 4996.485 ;
        RECT 381.965 4995.885 455.035 4996.485 ;
        RECT 638.965 4995.885 712.035 4996.485 ;
        RECT 895.965 4995.885 969.035 4996.485 ;
        RECT 1152.240 4995.885 1230.885 4996.485 ;
        RECT 1410.240 4995.885 1488.885 4996.485 ;
        RECT 1667.965 4995.885 1741.035 4996.485 ;
        RECT 1919.965 4995.885 1993.035 4996.485 ;
        RECT 2364.965 4995.885 2438.035 4996.485 ;
        RECT 2621.965 4995.885 2695.035 4996.485 ;
        RECT 2878.965 4995.885 2952.035 4996.485 ;
        RECT 3130.965 4995.885 3204.035 4996.485 ;
        RECT 3388.000 4995.885 3435.335 4996.485 ;
        RECT 152.665 4992.185 202.330 4995.885 ;
        RECT 152.665 4990.000 186.065 4992.185 ;
        RECT 152.665 4989.875 169.115 4990.000 ;
        RECT 152.665 4988.000 153.365 4989.875 ;
        RECT 158.815 4989.785 169.115 4989.875 ;
        RECT 158.815 4989.735 164.265 4989.785 ;
        RECT 152.665 4844.330 153.365 4845.035 ;
      LAYER met4 ;
        RECT 153.765 4844.730 158.415 4989.475 ;
      LAYER met4 ;
        RECT 158.815 4988.000 159.415 4989.735 ;
        RECT 158.815 4844.330 159.415 4845.035 ;
      LAYER met4 ;
        RECT 159.815 4844.730 163.265 4989.335 ;
      LAYER met4 ;
        RECT 163.665 4988.000 164.265 4989.735 ;
        RECT 163.665 4844.330 164.265 4845.035 ;
      LAYER met4 ;
        RECT 164.665 4844.730 168.115 4989.385 ;
      LAYER met4 ;
        RECT 168.515 4988.000 169.115 4989.785 ;
        RECT 174.565 4989.925 186.065 4990.000 ;
        RECT 168.515 4844.330 169.115 4845.035 ;
      LAYER met4 ;
        RECT 169.515 4844.730 174.165 4989.600 ;
      LAYER met4 ;
        RECT 174.565 4988.000 175.165 4989.925 ;
        RECT 180.615 4989.870 186.065 4989.925 ;
        RECT 174.565 4844.330 175.165 4845.035 ;
      LAYER met4 ;
        RECT 175.565 4844.730 180.215 4989.525 ;
      LAYER met4 ;
        RECT 180.615 4988.000 181.215 4989.870 ;
      LAYER met4 ;
        RECT 181.615 4845.035 185.065 4989.470 ;
      LAYER met4 ;
        RECT 185.465 4988.000 186.065 4989.870 ;
        RECT 180.615 4844.635 181.215 4845.035 ;
        RECT 185.465 4844.635 186.065 4845.035 ;
      LAYER met4 ;
        RECT 186.465 4844.730 191.115 4991.785 ;
      LAYER met4 ;
        RECT 191.515 4990.750 202.330 4992.185 ;
        RECT 191.515 4988.000 192.115 4990.750 ;
        RECT 180.615 4844.330 186.065 4844.635 ;
        RECT 191.515 4844.330 192.115 4845.035 ;
      LAYER met4 ;
        RECT 192.515 4844.730 197.965 4990.350 ;
      LAYER met4 ;
        RECT 198.365 4989.635 202.330 4990.750 ;
      LAYER met4 ;
        RECT 202.730 4990.035 382.270 4995.485 ;
      LAYER met4 ;
        RECT 382.670 4990.035 454.330 4995.885 ;
      LAYER met4 ;
        RECT 454.730 4990.035 639.270 4995.485 ;
      LAYER met4 ;
        RECT 639.670 4990.035 711.330 4995.885 ;
      LAYER met4 ;
        RECT 711.730 4990.035 896.270 4995.485 ;
      LAYER met4 ;
        RECT 896.670 4990.035 968.330 4995.885 ;
      LAYER met4 ;
        RECT 968.730 4990.035 1152.715 4995.485 ;
      LAYER met4 ;
        RECT 1153.115 4990.035 1230.485 4995.885 ;
      LAYER met4 ;
        RECT 1230.885 4990.035 1410.715 4995.485 ;
      LAYER met4 ;
        RECT 1411.115 4990.035 1488.485 4995.885 ;
      LAYER met4 ;
        RECT 1488.885 4990.035 1668.270 4995.485 ;
      LAYER met4 ;
        RECT 1668.670 4990.035 1740.330 4995.885 ;
      LAYER met4 ;
        RECT 1740.730 4990.035 1920.270 4995.485 ;
      LAYER met4 ;
        RECT 1920.670 4990.035 1992.330 4995.885 ;
      LAYER met4 ;
        RECT 1992.730 4990.035 2365.270 4995.485 ;
      LAYER met4 ;
        RECT 2365.670 4990.035 2437.330 4995.885 ;
      LAYER met4 ;
        RECT 2437.730 4990.035 2622.270 4995.485 ;
      LAYER met4 ;
        RECT 2622.670 4990.035 2694.330 4995.885 ;
      LAYER met4 ;
        RECT 2694.730 4990.035 2879.270 4995.485 ;
      LAYER met4 ;
        RECT 2879.670 4990.035 2951.330 4995.885 ;
      LAYER met4 ;
        RECT 2951.730 4990.035 3131.270 4995.485 ;
      LAYER met4 ;
        RECT 3131.670 4990.035 3203.330 4995.885 ;
      LAYER met4 ;
        RECT 3203.730 4990.035 3390.350 4995.485 ;
      LAYER met4 ;
        RECT 3390.750 4989.635 3435.335 4995.885 ;
        RECT 198.365 4988.000 202.745 4989.635 ;
        RECT 3388.000 4985.670 3435.335 4989.635 ;
        RECT 3388.000 4985.255 3389.635 4985.670 ;
        RECT 152.665 4772.670 197.965 4844.330 ;
      LAYER met4 ;
        RECT 3390.035 4837.285 3395.485 4985.270 ;
      LAYER met4 ;
        RECT 3395.885 4985.255 3396.485 4985.670 ;
        RECT 3401.935 4985.655 3407.385 4985.670 ;
        RECT 3395.885 4836.885 3396.485 4837.760 ;
      LAYER met4 ;
        RECT 3396.885 4837.285 3401.535 4985.270 ;
      LAYER met4 ;
        RECT 3401.935 4985.255 3402.535 4985.655 ;
        RECT 3406.785 4985.255 3407.385 4985.655 ;
        RECT 3401.935 4836.885 3402.535 4837.760 ;
      LAYER met4 ;
        RECT 3402.935 4837.285 3406.385 4985.255 ;
      LAYER met4 ;
        RECT 3406.785 4836.885 3407.385 4837.760 ;
      LAYER met4 ;
        RECT 3407.785 4837.285 3412.435 4985.270 ;
      LAYER met4 ;
        RECT 3412.835 4985.255 3413.435 4985.670 ;
        RECT 3412.835 4836.885 3413.435 4837.760 ;
      LAYER met4 ;
        RECT 3413.835 4837.285 3418.485 4985.270 ;
      LAYER met4 ;
        RECT 3418.885 4985.255 3419.485 4985.670 ;
        RECT 3418.885 4836.885 3419.485 4837.760 ;
      LAYER met4 ;
        RECT 3419.885 4837.285 3423.335 4985.270 ;
      LAYER met4 ;
        RECT 3423.735 4985.255 3424.335 4985.670 ;
        RECT 3423.735 4836.885 3424.335 4837.760 ;
      LAYER met4 ;
        RECT 3424.735 4837.285 3428.185 4985.270 ;
      LAYER met4 ;
        RECT 3428.585 4985.255 3429.185 4985.670 ;
        RECT 3428.585 4837.350 3429.185 4837.760 ;
      LAYER met4 ;
        RECT 3429.585 4837.750 3434.235 4985.270 ;
      LAYER met4 ;
        RECT 3434.635 4985.255 3435.335 4985.670 ;
        RECT 3434.635 4837.350 3435.335 4837.760 ;
        RECT 3428.585 4836.885 3435.335 4837.350 ;
        RECT 152.665 4771.965 153.365 4772.670 ;
        RECT 152.665 4633.330 153.365 4635.000 ;
      LAYER met4 ;
        RECT 153.765 4633.730 158.415 4772.270 ;
      LAYER met4 ;
        RECT 158.815 4771.965 159.415 4772.670 ;
        RECT 158.815 4633.330 159.415 4635.000 ;
      LAYER met4 ;
        RECT 159.815 4633.730 163.265 4772.270 ;
      LAYER met4 ;
        RECT 163.665 4771.965 164.265 4772.670 ;
        RECT 163.665 4633.330 164.265 4635.000 ;
      LAYER met4 ;
        RECT 164.665 4633.730 168.115 4772.270 ;
      LAYER met4 ;
        RECT 168.515 4771.965 169.115 4772.670 ;
        RECT 168.515 4633.330 169.115 4635.000 ;
      LAYER met4 ;
        RECT 169.515 4633.730 174.165 4772.270 ;
      LAYER met4 ;
        RECT 174.565 4771.965 175.165 4772.670 ;
        RECT 180.615 4772.365 186.065 4772.670 ;
        RECT 174.165 4634.935 174.200 4645.935 ;
        RECT 174.565 4633.330 175.165 4635.000 ;
      LAYER met4 ;
        RECT 175.565 4633.730 180.215 4772.270 ;
      LAYER met4 ;
        RECT 180.615 4771.965 181.215 4772.365 ;
        RECT 185.465 4771.965 186.065 4772.365 ;
        RECT 180.615 4633.635 181.215 4635.000 ;
      LAYER met4 ;
        RECT 181.615 4634.035 185.065 4771.965 ;
      LAYER met4 ;
        RECT 185.465 4633.635 186.065 4635.000 ;
      LAYER met4 ;
        RECT 186.465 4633.730 191.115 4772.270 ;
      LAYER met4 ;
        RECT 191.515 4771.965 192.115 4772.670 ;
        RECT 180.615 4633.330 186.065 4633.635 ;
        RECT 191.515 4633.330 192.115 4635.000 ;
      LAYER met4 ;
        RECT 192.515 4633.730 197.965 4772.270 ;
      LAYER met4 ;
        RECT 3390.035 4764.195 3435.335 4836.885 ;
        RECT 3390.035 4759.515 3402.535 4764.195 ;
        RECT 3395.885 4759.115 3396.485 4759.515 ;
        RECT 3401.935 4759.115 3402.535 4759.515 ;
        RECT 152.665 4561.670 197.965 4633.330 ;
      LAYER met4 ;
        RECT 3390.035 4611.730 3395.485 4759.115 ;
      LAYER met4 ;
        RECT 3395.885 4611.330 3396.485 4613.000 ;
      LAYER met4 ;
        RECT 3396.885 4611.730 3401.535 4759.115 ;
      LAYER met4 ;
        RECT 3401.935 4611.635 3402.535 4613.000 ;
      LAYER met4 ;
        RECT 3402.935 4612.035 3406.385 4763.795 ;
      LAYER met4 ;
        RECT 3406.785 4759.115 3407.385 4764.195 ;
        RECT 3406.785 4611.635 3407.385 4613.000 ;
      LAYER met4 ;
        RECT 3407.785 4611.730 3412.435 4763.795 ;
      LAYER met4 ;
        RECT 3412.835 4759.515 3435.335 4764.195 ;
        RECT 3412.835 4759.115 3413.435 4759.515 ;
        RECT 3418.885 4759.115 3419.485 4759.515 ;
        RECT 3423.735 4759.115 3424.335 4759.515 ;
        RECT 3428.585 4759.115 3429.185 4759.515 ;
        RECT 3434.635 4759.115 3435.335 4759.515 ;
        RECT 3401.935 4611.330 3407.385 4611.635 ;
        RECT 3412.835 4611.330 3413.435 4613.000 ;
      LAYER met4 ;
        RECT 3413.835 4611.730 3418.485 4759.115 ;
      LAYER met4 ;
        RECT 3418.885 4611.330 3419.485 4613.000 ;
      LAYER met4 ;
        RECT 3419.885 4611.730 3423.335 4759.115 ;
      LAYER met4 ;
        RECT 3423.735 4611.330 3424.335 4613.000 ;
      LAYER met4 ;
        RECT 3424.735 4611.730 3428.185 4759.115 ;
      LAYER met4 ;
        RECT 3428.585 4611.330 3429.185 4613.000 ;
        RECT 3429.550 4612.930 3429.585 4623.975 ;
      LAYER met4 ;
        RECT 3429.585 4611.730 3434.235 4759.115 ;
      LAYER met4 ;
        RECT 3434.635 4611.330 3435.335 4613.000 ;
        RECT 152.665 4560.000 153.365 4561.670 ;
        RECT 152.665 4422.330 153.365 4423.035 ;
      LAYER met4 ;
        RECT 153.765 4422.730 158.415 4561.270 ;
      LAYER met4 ;
        RECT 158.415 4549.025 158.450 4560.070 ;
        RECT 158.815 4560.000 159.415 4561.670 ;
        RECT 158.815 4422.330 159.415 4423.035 ;
      LAYER met4 ;
        RECT 159.815 4422.730 163.265 4561.270 ;
      LAYER met4 ;
        RECT 163.665 4560.000 164.265 4561.670 ;
        RECT 163.665 4422.330 164.265 4423.035 ;
      LAYER met4 ;
        RECT 164.665 4422.730 168.115 4561.270 ;
      LAYER met4 ;
        RECT 168.515 4560.000 169.115 4561.670 ;
        RECT 168.515 4422.330 169.115 4423.035 ;
      LAYER met4 ;
        RECT 169.515 4422.730 174.165 4561.270 ;
      LAYER met4 ;
        RECT 174.565 4560.000 175.165 4561.670 ;
        RECT 180.615 4561.365 186.065 4561.670 ;
        RECT 174.565 4422.330 175.165 4423.035 ;
      LAYER met4 ;
        RECT 175.565 4422.730 180.215 4561.270 ;
      LAYER met4 ;
        RECT 180.615 4560.000 181.215 4561.365 ;
      LAYER met4 ;
        RECT 181.615 4423.035 185.065 4560.965 ;
      LAYER met4 ;
        RECT 185.465 4560.000 186.065 4561.365 ;
        RECT 180.615 4422.635 181.215 4423.035 ;
        RECT 185.465 4422.635 186.065 4423.035 ;
      LAYER met4 ;
        RECT 186.465 4422.730 191.115 4561.270 ;
      LAYER met4 ;
        RECT 191.515 4560.000 192.115 4561.670 ;
        RECT 180.615 4422.330 186.065 4422.635 ;
        RECT 191.515 4422.330 192.115 4423.035 ;
      LAYER met4 ;
        RECT 192.515 4422.730 197.965 4561.270 ;
      LAYER met4 ;
        RECT 3390.035 4539.670 3435.335 4611.330 ;
        RECT 152.665 4350.670 197.965 4422.330 ;
        RECT 3388.535 4390.330 3389.635 4391.035 ;
      LAYER met4 ;
        RECT 3390.035 4390.730 3395.485 4539.270 ;
      LAYER met4 ;
        RECT 3395.885 4538.000 3396.485 4539.670 ;
        RECT 3401.935 4539.365 3407.385 4539.670 ;
        RECT 3395.885 4390.330 3396.485 4391.035 ;
      LAYER met4 ;
        RECT 3396.885 4390.730 3401.535 4539.270 ;
      LAYER met4 ;
        RECT 3401.935 4538.000 3402.535 4539.365 ;
      LAYER met4 ;
        RECT 3402.935 4391.035 3406.385 4538.965 ;
      LAYER met4 ;
        RECT 3406.785 4538.000 3407.385 4539.365 ;
        RECT 3401.935 4390.635 3402.535 4391.035 ;
        RECT 3406.785 4390.635 3407.385 4391.035 ;
      LAYER met4 ;
        RECT 3407.785 4390.730 3412.435 4539.270 ;
      LAYER met4 ;
        RECT 3412.835 4538.000 3413.435 4539.670 ;
        RECT 3413.800 4527.065 3413.835 4538.065 ;
        RECT 3401.935 4390.330 3407.385 4390.635 ;
        RECT 3412.835 4390.330 3413.435 4391.035 ;
      LAYER met4 ;
        RECT 3413.835 4390.730 3418.485 4539.270 ;
      LAYER met4 ;
        RECT 3418.885 4538.000 3419.485 4539.670 ;
        RECT 3418.885 4390.330 3419.485 4391.035 ;
      LAYER met4 ;
        RECT 3419.885 4390.730 3423.335 4539.270 ;
      LAYER met4 ;
        RECT 3423.735 4538.000 3424.335 4539.670 ;
        RECT 3423.735 4390.330 3424.335 4391.035 ;
      LAYER met4 ;
        RECT 3424.735 4390.730 3428.185 4539.270 ;
      LAYER met4 ;
        RECT 3428.585 4538.000 3429.185 4539.670 ;
        RECT 3428.585 4390.330 3429.185 4391.035 ;
      LAYER met4 ;
        RECT 3429.585 4390.730 3434.235 4539.270 ;
      LAYER met4 ;
        RECT 3434.635 4538.000 3435.335 4539.670 ;
        RECT 3434.635 4390.330 3435.335 4391.035 ;
        RECT 3388.535 4388.990 3435.335 4390.330 ;
      LAYER met4 ;
        RECT 3435.735 4389.390 3436.065 5007.575 ;
      LAYER met4 ;
        RECT 3436.465 5005.955 3440.725 5007.975 ;
        RECT 3436.465 5005.275 3439.245 5005.955 ;
        RECT 152.665 4349.965 153.365 4350.670 ;
        RECT 152.665 4211.330 153.365 4212.035 ;
      LAYER met4 ;
        RECT 153.765 4211.730 158.415 4350.270 ;
      LAYER met4 ;
        RECT 158.815 4349.965 159.415 4350.670 ;
        RECT 158.815 4211.330 159.415 4212.035 ;
      LAYER met4 ;
        RECT 159.815 4211.730 163.265 4350.270 ;
      LAYER met4 ;
        RECT 163.665 4349.965 164.265 4350.670 ;
        RECT 163.665 4211.330 164.265 4212.035 ;
      LAYER met4 ;
        RECT 164.665 4211.730 168.115 4350.270 ;
      LAYER met4 ;
        RECT 168.515 4349.965 169.115 4350.670 ;
        RECT 168.515 4211.330 169.115 4212.035 ;
      LAYER met4 ;
        RECT 169.515 4211.730 174.165 4350.270 ;
      LAYER met4 ;
        RECT 174.565 4349.965 175.165 4350.670 ;
        RECT 180.615 4350.365 186.065 4350.670 ;
        RECT 174.565 4211.330 175.165 4212.035 ;
      LAYER met4 ;
        RECT 175.565 4211.730 180.215 4350.270 ;
      LAYER met4 ;
        RECT 180.615 4349.965 181.215 4350.365 ;
        RECT 185.465 4349.965 186.065 4350.365 ;
      LAYER met4 ;
        RECT 181.615 4212.035 185.065 4349.965 ;
      LAYER met4 ;
        RECT 180.615 4211.635 181.215 4212.035 ;
        RECT 185.465 4211.635 186.065 4212.035 ;
      LAYER met4 ;
        RECT 186.465 4211.730 191.115 4350.270 ;
      LAYER met4 ;
        RECT 191.515 4349.965 192.115 4350.670 ;
        RECT 180.615 4211.330 186.065 4211.635 ;
        RECT 191.515 4211.330 192.115 4212.035 ;
      LAYER met4 ;
        RECT 192.515 4211.730 197.965 4350.270 ;
      LAYER met4 ;
        RECT 3388.535 4345.310 3435.965 4388.990 ;
        RECT 3388.535 4313.670 3435.335 4345.310 ;
        RECT 3388.535 4313.030 3389.635 4313.670 ;
        RECT 152.035 4139.670 197.965 4211.330 ;
      LAYER met4 ;
        RECT 3390.035 4165.730 3395.485 4313.270 ;
      LAYER met4 ;
        RECT 3395.885 4313.030 3396.485 4313.670 ;
        RECT 3401.935 4313.430 3407.385 4313.670 ;
        RECT 3395.885 4165.330 3396.485 4166.035 ;
      LAYER met4 ;
        RECT 3396.885 4165.730 3401.535 4313.270 ;
      LAYER met4 ;
        RECT 3401.935 4313.030 3402.535 4313.430 ;
        RECT 3406.785 4313.030 3407.385 4313.430 ;
      LAYER met4 ;
        RECT 3402.935 4166.035 3406.385 4313.030 ;
      LAYER met4 ;
        RECT 3401.935 4165.635 3402.535 4166.035 ;
        RECT 3406.785 4165.635 3407.385 4166.035 ;
      LAYER met4 ;
        RECT 3407.785 4165.730 3412.435 4313.270 ;
      LAYER met4 ;
        RECT 3412.835 4313.030 3413.435 4313.670 ;
        RECT 3401.935 4165.330 3407.385 4165.635 ;
        RECT 3412.835 4165.330 3413.435 4166.035 ;
      LAYER met4 ;
        RECT 3413.835 4165.730 3418.485 4313.270 ;
      LAYER met4 ;
        RECT 3418.885 4313.030 3419.485 4313.670 ;
        RECT 3418.885 4165.330 3419.485 4166.035 ;
      LAYER met4 ;
        RECT 3419.885 4165.730 3423.335 4313.270 ;
      LAYER met4 ;
        RECT 3423.735 4313.030 3424.335 4313.670 ;
        RECT 3423.735 4165.330 3424.335 4166.035 ;
      LAYER met4 ;
        RECT 3424.735 4165.730 3428.185 4313.270 ;
      LAYER met4 ;
        RECT 3428.585 4313.030 3429.185 4313.670 ;
        RECT 3428.585 4165.330 3429.185 4166.035 ;
      LAYER met4 ;
        RECT 3429.585 4165.730 3434.235 4313.270 ;
      LAYER met4 ;
        RECT 3434.635 4313.030 3435.335 4313.670 ;
        RECT 3434.635 4165.330 3435.335 4166.035 ;
        RECT 147.275 3974.545 151.535 3976.065 ;
        RECT 147.275 3960.360 148.255 3974.545 ;
        RECT 0.000 3958.840 148.255 3960.360 ;
        RECT 0.000 3925.010 143.495 3958.840 ;
        RECT 0.000 3923.670 142.865 3925.010 ;
      LAYER met4 ;
        RECT 0.000 3922.000 24.215 3923.270 ;
      LAYER met4 ;
        RECT 24.615 3922.965 104.600 3923.670 ;
        RECT 0.000 3786.000 104.600 3922.000 ;
      LAYER met4 ;
        RECT 0.000 3784.730 24.215 3786.000 ;
      LAYER met4 ;
        RECT 24.615 3784.330 104.600 3784.970 ;
      LAYER met4 ;
        RECT 105.000 3784.730 129.965 3923.270 ;
      LAYER met4 ;
        RECT 130.365 3922.965 131.065 3923.670 ;
        RECT 130.365 3786.000 131.065 3922.000 ;
        RECT 130.365 3784.330 131.065 3784.970 ;
      LAYER met4 ;
        RECT 131.465 3784.730 135.915 3923.270 ;
      LAYER met4 ;
        RECT 136.315 3922.965 136.915 3923.670 ;
        RECT 136.315 3786.000 136.915 3922.000 ;
        RECT 136.315 3784.330 136.915 3784.970 ;
      LAYER met4 ;
        RECT 137.315 3784.730 141.765 3923.270 ;
      LAYER met4 ;
        RECT 142.165 3922.965 142.865 3923.670 ;
        RECT 142.165 3786.000 142.865 3922.000 ;
        RECT 142.165 3784.330 142.865 3784.970 ;
        RECT 0.000 3752.690 142.865 3784.330 ;
      LAYER met4 ;
        RECT 143.265 3753.090 143.595 3924.610 ;
      LAYER met4 ;
        RECT 0.000 3744.360 143.495 3752.690 ;
      LAYER met4 ;
        RECT 143.895 3744.760 146.875 3958.440 ;
      LAYER met4 ;
        RECT 147.275 3923.670 148.255 3958.840 ;
      LAYER met4 ;
        RECT 147.175 3922.000 148.355 3923.270 ;
      LAYER met4 ;
        RECT 147.175 3786.000 148.355 3922.000 ;
      LAYER met4 ;
        RECT 147.175 3784.730 148.355 3786.000 ;
      LAYER met4 ;
        RECT 147.275 3760.065 148.255 3784.330 ;
      LAYER met4 ;
        RECT 148.655 3760.465 151.635 3974.145 ;
        RECT 151.935 3969.090 152.265 4139.270 ;
      LAYER met4 ;
        RECT 152.665 4138.965 153.365 4139.670 ;
        RECT 152.665 4000.330 153.365 4000.970 ;
      LAYER met4 ;
        RECT 153.765 4000.730 158.415 4139.270 ;
      LAYER met4 ;
        RECT 158.815 4138.965 159.415 4139.670 ;
        RECT 158.815 4000.330 159.415 4000.970 ;
      LAYER met4 ;
        RECT 159.815 4000.730 163.265 4139.270 ;
      LAYER met4 ;
        RECT 163.665 4138.965 164.265 4139.670 ;
        RECT 163.665 4000.330 164.265 4000.970 ;
      LAYER met4 ;
        RECT 164.665 4000.730 168.115 4139.270 ;
      LAYER met4 ;
        RECT 168.515 4138.965 169.115 4139.670 ;
        RECT 168.515 4000.330 169.115 4000.970 ;
      LAYER met4 ;
        RECT 169.515 4000.730 174.165 4139.270 ;
      LAYER met4 ;
        RECT 174.565 4138.965 175.165 4139.670 ;
        RECT 180.615 4139.365 186.065 4139.670 ;
        RECT 174.565 4000.330 175.165 4000.970 ;
      LAYER met4 ;
        RECT 175.565 4000.730 180.215 4139.270 ;
      LAYER met4 ;
        RECT 180.615 4138.965 181.215 4139.365 ;
        RECT 185.465 4138.965 186.065 4139.365 ;
      LAYER met4 ;
        RECT 181.615 4000.970 185.065 4138.965 ;
      LAYER met4 ;
        RECT 180.615 4000.570 181.215 4000.970 ;
        RECT 185.465 4000.570 186.065 4000.970 ;
      LAYER met4 ;
        RECT 186.465 4000.730 191.115 4139.270 ;
      LAYER met4 ;
        RECT 191.515 4138.965 192.115 4139.670 ;
        RECT 180.615 4000.330 186.065 4000.570 ;
        RECT 191.515 4000.330 192.115 4000.970 ;
      LAYER met4 ;
        RECT 192.515 4000.730 197.965 4139.270 ;
      LAYER met4 ;
        RECT 3390.035 4093.670 3435.335 4165.330 ;
        RECT 198.365 4000.330 199.465 4000.970 ;
        RECT 152.665 3968.690 199.465 4000.330 ;
        RECT 152.035 3925.010 199.465 3968.690 ;
        RECT 147.275 3758.545 151.535 3760.065 ;
        RECT 147.275 3744.360 148.255 3758.545 ;
        RECT 0.000 3742.840 148.255 3744.360 ;
        RECT 0.000 3709.010 143.495 3742.840 ;
        RECT 0.000 3707.670 142.865 3709.010 ;
      LAYER met4 ;
        RECT 0.000 3706.000 24.215 3707.270 ;
      LAYER met4 ;
        RECT 24.615 3706.965 104.600 3707.670 ;
        RECT 0.000 3570.000 104.600 3706.000 ;
      LAYER met4 ;
        RECT 0.000 3568.730 24.215 3570.000 ;
      LAYER met4 ;
        RECT 24.615 3568.330 104.600 3568.970 ;
      LAYER met4 ;
        RECT 105.000 3568.730 129.965 3707.270 ;
      LAYER met4 ;
        RECT 130.365 3706.965 131.065 3707.670 ;
        RECT 130.365 3570.000 131.065 3706.000 ;
        RECT 130.365 3568.330 131.065 3568.970 ;
      LAYER met4 ;
        RECT 131.465 3568.730 135.915 3707.270 ;
      LAYER met4 ;
        RECT 136.315 3706.965 136.915 3707.670 ;
        RECT 136.315 3570.000 136.915 3706.000 ;
        RECT 136.315 3568.330 136.915 3568.970 ;
      LAYER met4 ;
        RECT 137.315 3568.730 141.765 3707.270 ;
      LAYER met4 ;
        RECT 142.165 3706.965 142.865 3707.670 ;
        RECT 142.165 3570.000 142.865 3706.000 ;
        RECT 142.165 3568.330 142.865 3568.970 ;
        RECT 0.000 3536.690 142.865 3568.330 ;
      LAYER met4 ;
        RECT 143.265 3537.090 143.595 3708.610 ;
      LAYER met4 ;
        RECT 0.000 3528.360 143.495 3536.690 ;
      LAYER met4 ;
        RECT 143.895 3528.760 146.875 3742.440 ;
      LAYER met4 ;
        RECT 147.275 3707.670 148.255 3742.840 ;
      LAYER met4 ;
        RECT 147.175 3706.000 148.355 3707.270 ;
      LAYER met4 ;
        RECT 147.175 3570.000 148.355 3706.000 ;
      LAYER met4 ;
        RECT 147.175 3568.730 148.355 3570.000 ;
      LAYER met4 ;
        RECT 147.275 3544.065 148.255 3568.330 ;
      LAYER met4 ;
        RECT 148.655 3544.465 151.635 3758.145 ;
        RECT 151.935 3753.090 152.265 3924.610 ;
      LAYER met4 ;
        RECT 152.665 3923.670 199.465 3925.010 ;
        RECT 152.665 3922.965 153.365 3923.670 ;
        RECT 152.665 3784.330 153.365 3784.970 ;
      LAYER met4 ;
        RECT 153.765 3784.730 158.415 3923.270 ;
      LAYER met4 ;
        RECT 158.815 3922.965 159.415 3923.670 ;
        RECT 158.815 3784.330 159.415 3784.970 ;
      LAYER met4 ;
        RECT 159.815 3784.730 163.265 3923.270 ;
      LAYER met4 ;
        RECT 163.665 3922.965 164.265 3923.670 ;
        RECT 163.665 3784.330 164.265 3784.970 ;
      LAYER met4 ;
        RECT 164.665 3784.730 168.115 3923.270 ;
      LAYER met4 ;
        RECT 168.515 3922.965 169.115 3923.670 ;
        RECT 168.515 3784.330 169.115 3784.970 ;
      LAYER met4 ;
        RECT 169.515 3784.730 174.165 3923.270 ;
      LAYER met4 ;
        RECT 174.565 3922.965 175.165 3923.670 ;
        RECT 180.615 3923.365 186.065 3923.670 ;
        RECT 174.565 3784.330 175.165 3784.970 ;
      LAYER met4 ;
        RECT 175.565 3784.730 180.215 3923.270 ;
      LAYER met4 ;
        RECT 180.615 3922.965 181.215 3923.365 ;
        RECT 185.465 3922.965 186.065 3923.365 ;
      LAYER met4 ;
        RECT 181.615 3784.970 185.065 3922.965 ;
      LAYER met4 ;
        RECT 180.615 3784.570 181.215 3784.970 ;
        RECT 185.465 3784.570 186.065 3784.970 ;
      LAYER met4 ;
        RECT 186.465 3784.730 191.115 3923.270 ;
      LAYER met4 ;
        RECT 191.515 3922.965 192.115 3923.670 ;
        RECT 180.615 3784.330 186.065 3784.570 ;
        RECT 191.515 3784.330 192.115 3784.970 ;
      LAYER met4 ;
        RECT 192.515 3784.730 197.965 3923.270 ;
      LAYER met4 ;
        RECT 198.365 3922.965 199.465 3923.670 ;
        RECT 3388.535 3944.330 3389.635 3945.035 ;
      LAYER met4 ;
        RECT 3390.035 3944.730 3395.485 4093.270 ;
      LAYER met4 ;
        RECT 3395.885 4092.965 3396.485 4093.670 ;
        RECT 3401.935 4093.365 3407.385 4093.670 ;
        RECT 3395.885 3944.330 3396.485 3945.035 ;
      LAYER met4 ;
        RECT 3396.885 3944.730 3401.535 4093.270 ;
      LAYER met4 ;
        RECT 3401.935 4092.965 3402.535 4093.365 ;
        RECT 3406.785 4092.965 3407.385 4093.365 ;
      LAYER met4 ;
        RECT 3402.935 3945.035 3406.385 4092.965 ;
      LAYER met4 ;
        RECT 3401.935 3944.635 3402.535 3945.035 ;
        RECT 3406.785 3944.635 3407.385 3945.035 ;
      LAYER met4 ;
        RECT 3407.785 3944.730 3412.435 4093.270 ;
      LAYER met4 ;
        RECT 3412.835 4092.965 3413.435 4093.670 ;
        RECT 3401.935 3944.330 3407.385 3944.635 ;
        RECT 3412.835 3944.330 3413.435 3945.035 ;
      LAYER met4 ;
        RECT 3413.835 3944.730 3418.485 4093.270 ;
      LAYER met4 ;
        RECT 3418.885 4092.965 3419.485 4093.670 ;
        RECT 3418.885 3944.330 3419.485 3945.035 ;
      LAYER met4 ;
        RECT 3419.885 3944.730 3423.335 4093.270 ;
      LAYER met4 ;
        RECT 3423.735 4092.965 3424.335 4093.670 ;
        RECT 3423.735 3944.330 3424.335 3945.035 ;
      LAYER met4 ;
        RECT 3424.735 3944.730 3428.185 4093.270 ;
      LAYER met4 ;
        RECT 3428.585 4092.965 3429.185 4093.670 ;
        RECT 3428.585 3944.330 3429.185 3945.035 ;
      LAYER met4 ;
        RECT 3429.585 3944.730 3434.235 4093.270 ;
      LAYER met4 ;
        RECT 3434.635 4092.965 3435.335 4093.670 ;
        RECT 3434.635 3944.330 3435.335 3945.035 ;
        RECT 3388.535 3942.990 3435.335 3944.330 ;
      LAYER met4 ;
        RECT 3435.735 3943.390 3436.065 4344.910 ;
        RECT 3436.365 4339.855 3439.345 5004.875 ;
        RECT 3439.645 4984.000 3440.825 5005.555 ;
      LAYER met4 ;
        RECT 3439.645 4885.000 3440.825 4984.000 ;
      LAYER met4 ;
        RECT 3439.645 4837.760 3440.825 4885.000 ;
      LAYER met4 ;
        RECT 3439.745 4759.515 3440.725 4837.360 ;
      LAYER met4 ;
        RECT 3439.645 4716.000 3440.825 4759.115 ;
      LAYER met4 ;
        RECT 3439.645 4613.000 3440.825 4716.000 ;
      LAYER met4 ;
        RECT 3439.645 4611.730 3440.825 4613.000 ;
      LAYER met4 ;
        RECT 3439.745 4539.670 3440.725 4611.330 ;
      LAYER met4 ;
        RECT 3439.645 4538.000 3440.825 4539.270 ;
      LAYER met4 ;
        RECT 3439.645 4392.000 3440.825 4538.000 ;
      LAYER met4 ;
        RECT 3439.645 4390.730 3440.825 4392.000 ;
      LAYER met4 ;
        RECT 3439.745 4355.160 3440.725 4390.330 ;
      LAYER met4 ;
        RECT 3441.125 4355.560 3444.105 5010.910 ;
        RECT 3444.405 4389.390 3444.735 5011.175 ;
      LAYER met4 ;
        RECT 3445.135 4986.255 3588.000 5011.575 ;
        RECT 3445.135 4985.670 3457.635 4986.255 ;
        RECT 3445.135 4985.255 3445.835 4985.670 ;
        RECT 3445.135 4885.000 3445.835 4984.000 ;
        RECT 3445.135 4836.885 3445.835 4837.760 ;
      LAYER met4 ;
        RECT 3446.235 4837.285 3450.685 4985.270 ;
      LAYER met4 ;
        RECT 3451.085 4985.255 3451.685 4985.670 ;
        RECT 3451.085 4885.000 3451.685 4984.000 ;
        RECT 3451.085 4836.885 3451.685 4837.760 ;
      LAYER met4 ;
        RECT 3452.085 4837.285 3456.535 4985.270 ;
      LAYER met4 ;
        RECT 3456.935 4985.255 3457.635 4985.670 ;
        RECT 3456.935 4885.000 3457.635 4984.000 ;
        RECT 3456.935 4836.885 3457.635 4837.760 ;
      LAYER met4 ;
        RECT 3458.035 4837.285 3483.000 4985.855 ;
      LAYER met4 ;
        RECT 3483.400 4985.670 3588.000 4986.255 ;
        RECT 3483.400 4985.255 3563.385 4985.670 ;
      LAYER met4 ;
        RECT 3563.785 4984.000 3588.000 4985.270 ;
      LAYER met4 ;
        RECT 3483.400 4885.000 3588.000 4984.000 ;
        RECT 3483.400 4836.885 3563.385 4837.760 ;
        RECT 3445.135 4836.395 3563.385 4836.885 ;
      LAYER met4 ;
        RECT 3563.785 4836.795 3588.000 4885.000 ;
      LAYER met4 ;
        RECT 3445.135 4759.515 3588.000 4836.395 ;
        RECT 3445.135 4759.115 3445.835 4759.515 ;
        RECT 3451.085 4759.115 3451.685 4759.515 ;
        RECT 3456.935 4759.115 3457.635 4759.515 ;
        RECT 3483.400 4759.115 3563.385 4759.515 ;
        RECT 3445.135 4611.330 3445.835 4716.000 ;
      LAYER met4 ;
        RECT 3446.235 4611.730 3450.685 4759.115 ;
      LAYER met4 ;
        RECT 3451.085 4611.330 3451.685 4716.000 ;
      LAYER met4 ;
        RECT 3452.085 4611.730 3456.535 4759.115 ;
      LAYER met4 ;
        RECT 3456.935 4611.330 3457.635 4716.000 ;
      LAYER met4 ;
        RECT 3458.035 4611.730 3483.000 4759.115 ;
        RECT 3563.785 4716.000 3588.000 4759.115 ;
      LAYER met4 ;
        RECT 3483.400 4613.000 3588.000 4716.000 ;
        RECT 3483.400 4611.330 3563.385 4613.000 ;
      LAYER met4 ;
        RECT 3563.785 4611.730 3588.000 4613.000 ;
      LAYER met4 ;
        RECT 3445.135 4539.670 3588.000 4611.330 ;
        RECT 3445.135 4392.000 3445.835 4539.670 ;
        RECT 3445.135 4390.330 3445.835 4391.035 ;
      LAYER met4 ;
        RECT 3446.235 4390.730 3450.685 4539.270 ;
      LAYER met4 ;
        RECT 3451.085 4392.000 3451.685 4539.670 ;
        RECT 3451.085 4390.330 3451.685 4391.035 ;
      LAYER met4 ;
        RECT 3452.085 4390.730 3456.535 4539.270 ;
      LAYER met4 ;
        RECT 3456.935 4392.000 3457.635 4539.670 ;
        RECT 3456.935 4390.330 3457.635 4391.035 ;
      LAYER met4 ;
        RECT 3458.035 4390.730 3483.000 4539.270 ;
      LAYER met4 ;
        RECT 3483.400 4538.000 3563.385 4539.670 ;
        RECT 3563.750 4538.000 3563.785 4538.215 ;
      LAYER met4 ;
        RECT 3563.785 4538.000 3588.000 4539.270 ;
      LAYER met4 ;
        RECT 3483.400 4392.000 3588.000 4538.000 ;
        RECT 3483.400 4390.330 3563.385 4391.035 ;
      LAYER met4 ;
        RECT 3563.785 4390.730 3588.000 4392.000 ;
      LAYER met4 ;
        RECT 3445.135 4388.990 3588.000 4390.330 ;
        RECT 3444.505 4355.160 3588.000 4388.990 ;
        RECT 3439.745 4353.640 3588.000 4355.160 ;
        RECT 3439.745 4339.455 3440.725 4353.640 ;
        RECT 3436.465 4337.935 3440.725 4339.455 ;
        RECT 3388.535 3899.310 3435.965 3942.990 ;
        RECT 3388.535 3867.670 3435.335 3899.310 ;
        RECT 3388.535 3867.030 3389.635 3867.670 ;
        RECT 198.365 3784.330 199.465 3784.970 ;
        RECT 152.665 3752.690 199.465 3784.330 ;
        RECT 152.035 3709.010 199.465 3752.690 ;
        RECT 147.275 3542.545 151.535 3544.065 ;
        RECT 147.275 3528.360 148.255 3542.545 ;
        RECT 0.000 3526.840 148.255 3528.360 ;
        RECT 0.000 3493.010 143.495 3526.840 ;
        RECT 0.000 3491.670 142.865 3493.010 ;
      LAYER met4 ;
        RECT 0.000 3490.000 24.215 3491.270 ;
      LAYER met4 ;
        RECT 24.615 3490.965 104.600 3491.670 ;
        RECT 0.000 3354.000 104.600 3490.000 ;
      LAYER met4 ;
        RECT 0.000 3352.730 24.215 3354.000 ;
      LAYER met4 ;
        RECT 24.615 3352.330 104.600 3352.970 ;
      LAYER met4 ;
        RECT 105.000 3352.730 129.965 3491.270 ;
      LAYER met4 ;
        RECT 130.365 3490.965 131.065 3491.670 ;
        RECT 130.365 3354.000 131.065 3490.000 ;
        RECT 130.365 3352.330 131.065 3352.970 ;
      LAYER met4 ;
        RECT 131.465 3352.730 135.915 3491.270 ;
      LAYER met4 ;
        RECT 136.315 3490.965 136.915 3491.670 ;
        RECT 136.315 3354.000 136.915 3490.000 ;
        RECT 136.315 3352.330 136.915 3352.970 ;
      LAYER met4 ;
        RECT 137.315 3352.730 141.765 3491.270 ;
      LAYER met4 ;
        RECT 142.165 3490.965 142.865 3491.670 ;
        RECT 142.165 3354.000 142.865 3490.000 ;
        RECT 142.165 3352.330 142.865 3352.970 ;
        RECT 0.000 3320.690 142.865 3352.330 ;
      LAYER met4 ;
        RECT 143.265 3321.090 143.595 3492.610 ;
      LAYER met4 ;
        RECT 0.000 3312.360 143.495 3320.690 ;
      LAYER met4 ;
        RECT 143.895 3312.760 146.875 3526.440 ;
      LAYER met4 ;
        RECT 147.275 3491.670 148.255 3526.840 ;
      LAYER met4 ;
        RECT 147.175 3490.000 148.355 3491.270 ;
      LAYER met4 ;
        RECT 147.175 3354.000 148.355 3490.000 ;
      LAYER met4 ;
        RECT 147.175 3352.730 148.355 3354.000 ;
      LAYER met4 ;
        RECT 147.275 3328.065 148.255 3352.330 ;
      LAYER met4 ;
        RECT 148.655 3328.465 151.635 3542.145 ;
        RECT 151.935 3537.090 152.265 3708.610 ;
      LAYER met4 ;
        RECT 152.665 3707.670 199.465 3709.010 ;
        RECT 152.665 3706.965 153.365 3707.670 ;
        RECT 152.665 3568.330 153.365 3568.970 ;
      LAYER met4 ;
        RECT 153.765 3568.730 158.415 3707.270 ;
      LAYER met4 ;
        RECT 158.815 3706.965 159.415 3707.670 ;
        RECT 158.815 3568.330 159.415 3568.970 ;
      LAYER met4 ;
        RECT 159.815 3568.730 163.265 3707.270 ;
      LAYER met4 ;
        RECT 163.665 3706.965 164.265 3707.670 ;
        RECT 163.665 3568.330 164.265 3568.970 ;
      LAYER met4 ;
        RECT 164.665 3568.730 168.115 3707.270 ;
      LAYER met4 ;
        RECT 168.515 3706.965 169.115 3707.670 ;
        RECT 168.515 3568.330 169.115 3568.970 ;
      LAYER met4 ;
        RECT 169.515 3568.730 174.165 3707.270 ;
      LAYER met4 ;
        RECT 174.565 3706.965 175.165 3707.670 ;
        RECT 180.615 3707.365 186.065 3707.670 ;
        RECT 174.565 3568.330 175.165 3568.970 ;
      LAYER met4 ;
        RECT 175.565 3568.730 180.215 3707.270 ;
      LAYER met4 ;
        RECT 180.615 3706.965 181.215 3707.365 ;
        RECT 185.465 3706.965 186.065 3707.365 ;
      LAYER met4 ;
        RECT 181.615 3568.970 185.065 3706.965 ;
      LAYER met4 ;
        RECT 180.615 3568.570 181.215 3568.970 ;
        RECT 185.465 3568.570 186.065 3568.970 ;
      LAYER met4 ;
        RECT 186.465 3568.730 191.115 3707.270 ;
      LAYER met4 ;
        RECT 191.515 3706.965 192.115 3707.670 ;
        RECT 180.615 3568.330 186.065 3568.570 ;
        RECT 191.515 3568.330 192.115 3568.970 ;
      LAYER met4 ;
        RECT 192.515 3568.730 197.965 3707.270 ;
      LAYER met4 ;
        RECT 198.365 3706.965 199.465 3707.670 ;
        RECT 3388.535 3719.330 3389.635 3720.035 ;
      LAYER met4 ;
        RECT 3390.035 3719.730 3395.485 3867.270 ;
      LAYER met4 ;
        RECT 3395.885 3867.030 3396.485 3867.670 ;
        RECT 3401.935 3867.430 3407.385 3867.670 ;
        RECT 3395.885 3719.330 3396.485 3720.035 ;
      LAYER met4 ;
        RECT 3396.885 3719.730 3401.535 3867.270 ;
      LAYER met4 ;
        RECT 3401.935 3867.030 3402.535 3867.430 ;
        RECT 3406.785 3867.030 3407.385 3867.430 ;
      LAYER met4 ;
        RECT 3402.935 3720.035 3406.385 3867.030 ;
      LAYER met4 ;
        RECT 3401.935 3719.635 3402.535 3720.035 ;
        RECT 3406.785 3719.635 3407.385 3720.035 ;
      LAYER met4 ;
        RECT 3407.785 3719.730 3412.435 3867.270 ;
      LAYER met4 ;
        RECT 3412.835 3867.030 3413.435 3867.670 ;
        RECT 3401.935 3719.330 3407.385 3719.635 ;
        RECT 3412.835 3719.330 3413.435 3720.035 ;
      LAYER met4 ;
        RECT 3413.835 3719.730 3418.485 3867.270 ;
      LAYER met4 ;
        RECT 3418.885 3867.030 3419.485 3867.670 ;
        RECT 3418.885 3719.330 3419.485 3720.035 ;
      LAYER met4 ;
        RECT 3419.885 3719.730 3423.335 3867.270 ;
      LAYER met4 ;
        RECT 3423.735 3867.030 3424.335 3867.670 ;
        RECT 3423.735 3719.330 3424.335 3720.035 ;
      LAYER met4 ;
        RECT 3424.735 3719.730 3428.185 3867.270 ;
      LAYER met4 ;
        RECT 3428.585 3867.030 3429.185 3867.670 ;
        RECT 3428.585 3719.330 3429.185 3720.035 ;
      LAYER met4 ;
        RECT 3429.585 3719.730 3434.235 3867.270 ;
      LAYER met4 ;
        RECT 3434.635 3867.030 3435.335 3867.670 ;
        RECT 3434.635 3719.330 3435.335 3720.035 ;
        RECT 3388.535 3717.990 3435.335 3719.330 ;
      LAYER met4 ;
        RECT 3435.735 3718.390 3436.065 3898.910 ;
        RECT 3436.365 3893.855 3439.345 4337.535 ;
      LAYER met4 ;
        RECT 3439.745 4313.670 3440.725 4337.935 ;
      LAYER met4 ;
        RECT 3439.645 4312.000 3440.825 4313.270 ;
      LAYER met4 ;
        RECT 3439.645 4167.000 3440.825 4312.000 ;
      LAYER met4 ;
        RECT 3439.645 4165.730 3440.825 4167.000 ;
      LAYER met4 ;
        RECT 3439.745 4093.670 3440.725 4165.330 ;
      LAYER met4 ;
        RECT 3439.645 4092.000 3440.825 4093.270 ;
      LAYER met4 ;
        RECT 3439.645 3946.000 3440.825 4092.000 ;
      LAYER met4 ;
        RECT 3439.645 3944.730 3440.825 3946.000 ;
      LAYER met4 ;
        RECT 3439.745 3909.160 3440.725 3944.330 ;
      LAYER met4 ;
        RECT 3441.125 3909.560 3444.105 4353.240 ;
      LAYER met4 ;
        RECT 3444.505 4345.310 3588.000 4353.640 ;
      LAYER met4 ;
        RECT 3444.405 3943.390 3444.735 4344.910 ;
      LAYER met4 ;
        RECT 3445.135 4313.670 3588.000 4345.310 ;
        RECT 3445.135 4313.030 3445.835 4313.670 ;
        RECT 3445.135 4167.000 3445.835 4312.000 ;
        RECT 3445.135 4165.330 3445.835 4166.035 ;
      LAYER met4 ;
        RECT 3446.235 4165.730 3450.685 4313.270 ;
      LAYER met4 ;
        RECT 3451.085 4313.030 3451.685 4313.670 ;
        RECT 3451.085 4167.000 3451.685 4312.000 ;
        RECT 3451.085 4165.330 3451.685 4166.035 ;
      LAYER met4 ;
        RECT 3452.085 4165.730 3456.535 4313.270 ;
      LAYER met4 ;
        RECT 3456.935 4313.030 3457.635 4313.670 ;
        RECT 3456.935 4167.000 3457.635 4312.000 ;
        RECT 3456.935 4165.330 3457.635 4166.035 ;
      LAYER met4 ;
        RECT 3458.035 4165.730 3483.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.400 4313.030 3563.385 4313.670 ;
      LAYER met4 ;
        RECT 3563.785 4312.000 3588.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.400 4167.000 3588.000 4312.000 ;
        RECT 3483.400 4165.330 3563.385 4166.035 ;
      LAYER met4 ;
        RECT 3563.785 4165.730 3588.000 4167.000 ;
      LAYER met4 ;
        RECT 3445.135 4093.670 3588.000 4165.330 ;
        RECT 3445.135 4092.965 3445.835 4093.670 ;
        RECT 3445.135 3946.000 3445.835 4092.000 ;
        RECT 3445.135 3944.330 3445.835 3945.035 ;
      LAYER met4 ;
        RECT 3446.235 3944.730 3450.685 4093.270 ;
      LAYER met4 ;
        RECT 3451.085 4092.965 3451.685 4093.670 ;
        RECT 3451.085 3946.000 3451.685 4092.000 ;
        RECT 3451.085 3944.330 3451.685 3945.035 ;
      LAYER met4 ;
        RECT 3452.085 3944.730 3456.535 4093.270 ;
      LAYER met4 ;
        RECT 3456.935 4092.965 3457.635 4093.670 ;
        RECT 3456.935 3946.000 3457.635 4092.000 ;
        RECT 3456.935 3944.330 3457.635 3945.035 ;
      LAYER met4 ;
        RECT 3458.035 3944.730 3483.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.400 4092.965 3563.385 4093.670 ;
      LAYER met4 ;
        RECT 3563.785 4092.000 3588.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.400 3946.000 3588.000 4092.000 ;
        RECT 3483.400 3944.330 3563.385 3945.035 ;
      LAYER met4 ;
        RECT 3563.785 3944.730 3588.000 3946.000 ;
      LAYER met4 ;
        RECT 3445.135 3942.990 3588.000 3944.330 ;
        RECT 3444.505 3909.160 3588.000 3942.990 ;
        RECT 3439.745 3907.640 3588.000 3909.160 ;
        RECT 3439.745 3893.455 3440.725 3907.640 ;
        RECT 3436.465 3891.935 3440.725 3893.455 ;
        RECT 3388.535 3674.310 3435.965 3717.990 ;
        RECT 3388.535 3642.670 3435.335 3674.310 ;
        RECT 3388.535 3642.030 3389.635 3642.670 ;
        RECT 198.365 3568.330 199.465 3568.970 ;
        RECT 152.665 3536.690 199.465 3568.330 ;
        RECT 152.035 3493.010 199.465 3536.690 ;
        RECT 147.275 3326.545 151.535 3328.065 ;
        RECT 147.275 3312.360 148.255 3326.545 ;
        RECT 0.000 3310.840 148.255 3312.360 ;
        RECT 0.000 3277.010 143.495 3310.840 ;
        RECT 0.000 3275.670 142.865 3277.010 ;
      LAYER met4 ;
        RECT 0.000 3274.000 24.215 3275.270 ;
      LAYER met4 ;
        RECT 24.615 3274.965 104.600 3275.670 ;
        RECT 0.000 3138.000 104.600 3274.000 ;
      LAYER met4 ;
        RECT 0.000 3136.730 24.215 3138.000 ;
      LAYER met4 ;
        RECT 24.615 3136.330 104.600 3136.970 ;
      LAYER met4 ;
        RECT 105.000 3136.730 129.965 3275.270 ;
      LAYER met4 ;
        RECT 130.365 3274.965 131.065 3275.670 ;
        RECT 130.365 3138.000 131.065 3274.000 ;
        RECT 130.365 3136.330 131.065 3136.970 ;
      LAYER met4 ;
        RECT 131.465 3136.730 135.915 3275.270 ;
      LAYER met4 ;
        RECT 136.315 3274.965 136.915 3275.670 ;
        RECT 136.315 3138.000 136.915 3274.000 ;
        RECT 136.315 3136.330 136.915 3136.970 ;
      LAYER met4 ;
        RECT 137.315 3136.730 141.765 3275.270 ;
      LAYER met4 ;
        RECT 142.165 3274.965 142.865 3275.670 ;
        RECT 142.165 3138.000 142.865 3274.000 ;
        RECT 142.165 3136.330 142.865 3136.970 ;
        RECT 0.000 3104.690 142.865 3136.330 ;
      LAYER met4 ;
        RECT 143.265 3105.090 143.595 3276.610 ;
      LAYER met4 ;
        RECT 0.000 3096.360 143.495 3104.690 ;
      LAYER met4 ;
        RECT 143.895 3096.760 146.875 3310.440 ;
      LAYER met4 ;
        RECT 147.275 3275.670 148.255 3310.840 ;
      LAYER met4 ;
        RECT 147.175 3274.000 148.355 3275.270 ;
      LAYER met4 ;
        RECT 147.175 3138.000 148.355 3274.000 ;
      LAYER met4 ;
        RECT 147.175 3136.730 148.355 3138.000 ;
      LAYER met4 ;
        RECT 147.275 3112.065 148.255 3136.330 ;
      LAYER met4 ;
        RECT 148.655 3112.465 151.635 3326.145 ;
        RECT 151.935 3321.090 152.265 3492.610 ;
      LAYER met4 ;
        RECT 152.665 3491.670 199.465 3493.010 ;
        RECT 152.665 3490.965 153.365 3491.670 ;
        RECT 152.665 3352.330 153.365 3352.970 ;
      LAYER met4 ;
        RECT 153.765 3352.730 158.415 3491.270 ;
      LAYER met4 ;
        RECT 158.815 3490.965 159.415 3491.670 ;
        RECT 158.815 3352.330 159.415 3352.970 ;
      LAYER met4 ;
        RECT 159.815 3352.730 163.265 3491.270 ;
      LAYER met4 ;
        RECT 163.665 3490.965 164.265 3491.670 ;
        RECT 163.665 3352.330 164.265 3352.970 ;
      LAYER met4 ;
        RECT 164.665 3352.730 168.115 3491.270 ;
      LAYER met4 ;
        RECT 168.515 3490.965 169.115 3491.670 ;
        RECT 168.515 3352.330 169.115 3352.970 ;
      LAYER met4 ;
        RECT 169.515 3352.730 174.165 3491.270 ;
      LAYER met4 ;
        RECT 174.565 3490.965 175.165 3491.670 ;
        RECT 180.615 3491.365 186.065 3491.670 ;
        RECT 174.565 3352.330 175.165 3352.970 ;
      LAYER met4 ;
        RECT 175.565 3352.730 180.215 3491.270 ;
      LAYER met4 ;
        RECT 180.615 3490.965 181.215 3491.365 ;
        RECT 185.465 3490.965 186.065 3491.365 ;
      LAYER met4 ;
        RECT 181.615 3352.970 185.065 3490.965 ;
      LAYER met4 ;
        RECT 180.615 3352.570 181.215 3352.970 ;
        RECT 185.465 3352.570 186.065 3352.970 ;
      LAYER met4 ;
        RECT 186.465 3352.730 191.115 3491.270 ;
      LAYER met4 ;
        RECT 191.515 3490.965 192.115 3491.670 ;
        RECT 180.615 3352.330 186.065 3352.570 ;
        RECT 191.515 3352.330 192.115 3352.970 ;
      LAYER met4 ;
        RECT 192.515 3352.730 197.965 3491.270 ;
      LAYER met4 ;
        RECT 198.365 3490.965 199.465 3491.670 ;
        RECT 3388.535 3494.330 3389.635 3495.035 ;
      LAYER met4 ;
        RECT 3390.035 3494.730 3395.485 3642.270 ;
      LAYER met4 ;
        RECT 3395.885 3642.030 3396.485 3642.670 ;
        RECT 3401.935 3642.430 3407.385 3642.670 ;
        RECT 3395.885 3494.330 3396.485 3495.035 ;
      LAYER met4 ;
        RECT 3396.885 3494.730 3401.535 3642.270 ;
      LAYER met4 ;
        RECT 3401.935 3642.030 3402.535 3642.430 ;
        RECT 3406.785 3642.030 3407.385 3642.430 ;
      LAYER met4 ;
        RECT 3402.935 3495.035 3406.385 3642.030 ;
      LAYER met4 ;
        RECT 3401.935 3494.635 3402.535 3495.035 ;
        RECT 3406.785 3494.635 3407.385 3495.035 ;
      LAYER met4 ;
        RECT 3407.785 3494.730 3412.435 3642.270 ;
      LAYER met4 ;
        RECT 3412.835 3642.030 3413.435 3642.670 ;
        RECT 3401.935 3494.330 3407.385 3494.635 ;
        RECT 3412.835 3494.330 3413.435 3495.035 ;
      LAYER met4 ;
        RECT 3413.835 3494.730 3418.485 3642.270 ;
      LAYER met4 ;
        RECT 3418.885 3642.030 3419.485 3642.670 ;
        RECT 3418.885 3494.330 3419.485 3495.035 ;
      LAYER met4 ;
        RECT 3419.885 3494.730 3423.335 3642.270 ;
      LAYER met4 ;
        RECT 3423.735 3642.030 3424.335 3642.670 ;
        RECT 3423.735 3494.330 3424.335 3495.035 ;
      LAYER met4 ;
        RECT 3424.735 3494.730 3428.185 3642.270 ;
      LAYER met4 ;
        RECT 3428.585 3642.030 3429.185 3642.670 ;
        RECT 3428.585 3494.330 3429.185 3495.035 ;
      LAYER met4 ;
        RECT 3429.585 3494.730 3434.235 3642.270 ;
      LAYER met4 ;
        RECT 3434.635 3642.030 3435.335 3642.670 ;
        RECT 3434.635 3494.330 3435.335 3495.035 ;
        RECT 3388.535 3492.990 3435.335 3494.330 ;
      LAYER met4 ;
        RECT 3435.735 3493.390 3436.065 3673.910 ;
        RECT 3436.365 3668.855 3439.345 3891.535 ;
      LAYER met4 ;
        RECT 3439.745 3867.670 3440.725 3891.935 ;
      LAYER met4 ;
        RECT 3439.645 3866.000 3440.825 3867.270 ;
      LAYER met4 ;
        RECT 3439.645 3721.000 3440.825 3866.000 ;
      LAYER met4 ;
        RECT 3439.645 3719.730 3440.825 3721.000 ;
      LAYER met4 ;
        RECT 3439.745 3684.160 3440.725 3719.330 ;
      LAYER met4 ;
        RECT 3441.125 3684.560 3444.105 3907.240 ;
      LAYER met4 ;
        RECT 3444.505 3899.310 3588.000 3907.640 ;
      LAYER met4 ;
        RECT 3444.405 3718.390 3444.735 3898.910 ;
      LAYER met4 ;
        RECT 3445.135 3867.670 3588.000 3899.310 ;
        RECT 3445.135 3867.030 3445.835 3867.670 ;
        RECT 3445.135 3721.000 3445.835 3866.000 ;
        RECT 3445.135 3719.330 3445.835 3720.035 ;
      LAYER met4 ;
        RECT 3446.235 3719.730 3450.685 3867.270 ;
      LAYER met4 ;
        RECT 3451.085 3867.030 3451.685 3867.670 ;
        RECT 3451.085 3721.000 3451.685 3866.000 ;
        RECT 3451.085 3719.330 3451.685 3720.035 ;
      LAYER met4 ;
        RECT 3452.085 3719.730 3456.535 3867.270 ;
      LAYER met4 ;
        RECT 3456.935 3867.030 3457.635 3867.670 ;
        RECT 3456.935 3721.000 3457.635 3866.000 ;
        RECT 3456.935 3719.330 3457.635 3720.035 ;
      LAYER met4 ;
        RECT 3458.035 3719.730 3483.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.400 3867.030 3563.385 3867.670 ;
      LAYER met4 ;
        RECT 3563.785 3866.000 3588.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.400 3721.000 3588.000 3866.000 ;
        RECT 3483.400 3719.330 3563.385 3720.035 ;
      LAYER met4 ;
        RECT 3563.785 3719.730 3588.000 3721.000 ;
      LAYER met4 ;
        RECT 3445.135 3717.990 3588.000 3719.330 ;
        RECT 3444.505 3684.160 3588.000 3717.990 ;
        RECT 3439.745 3682.640 3588.000 3684.160 ;
        RECT 3439.745 3668.455 3440.725 3682.640 ;
        RECT 3436.465 3666.935 3440.725 3668.455 ;
        RECT 3388.535 3449.310 3435.965 3492.990 ;
        RECT 3388.535 3417.670 3435.335 3449.310 ;
        RECT 3388.535 3417.030 3389.635 3417.670 ;
        RECT 198.365 3352.330 199.465 3352.970 ;
        RECT 152.665 3320.690 199.465 3352.330 ;
        RECT 152.035 3277.010 199.465 3320.690 ;
        RECT 147.275 3110.545 151.535 3112.065 ;
        RECT 147.275 3096.360 148.255 3110.545 ;
        RECT 0.000 3094.840 148.255 3096.360 ;
        RECT 0.000 3061.010 143.495 3094.840 ;
        RECT 0.000 3059.670 142.865 3061.010 ;
      LAYER met4 ;
        RECT 0.000 3058.000 24.215 3059.270 ;
      LAYER met4 ;
        RECT 24.615 3058.965 104.600 3059.670 ;
        RECT 0.000 2922.000 104.600 3058.000 ;
      LAYER met4 ;
        RECT 0.000 2920.730 24.215 2922.000 ;
      LAYER met4 ;
        RECT 24.615 2920.330 104.600 2920.970 ;
      LAYER met4 ;
        RECT 105.000 2920.730 129.965 3059.270 ;
      LAYER met4 ;
        RECT 130.365 3058.965 131.065 3059.670 ;
        RECT 130.365 2922.000 131.065 3058.000 ;
        RECT 130.365 2920.330 131.065 2920.970 ;
      LAYER met4 ;
        RECT 131.465 2920.730 135.915 3059.270 ;
      LAYER met4 ;
        RECT 136.315 3058.965 136.915 3059.670 ;
        RECT 136.315 2922.000 136.915 3058.000 ;
        RECT 136.315 2920.330 136.915 2920.970 ;
      LAYER met4 ;
        RECT 137.315 2920.730 141.765 3059.270 ;
      LAYER met4 ;
        RECT 142.165 3058.965 142.865 3059.670 ;
        RECT 142.165 2922.000 142.865 3058.000 ;
        RECT 142.165 2920.330 142.865 2920.970 ;
        RECT 0.000 2888.690 142.865 2920.330 ;
      LAYER met4 ;
        RECT 143.265 2889.090 143.595 3060.610 ;
      LAYER met4 ;
        RECT 0.000 2880.360 143.495 2888.690 ;
      LAYER met4 ;
        RECT 143.895 2880.760 146.875 3094.440 ;
      LAYER met4 ;
        RECT 147.275 3059.670 148.255 3094.840 ;
      LAYER met4 ;
        RECT 147.175 3058.000 148.355 3059.270 ;
      LAYER met4 ;
        RECT 147.175 2922.000 148.355 3058.000 ;
      LAYER met4 ;
        RECT 147.175 2920.730 148.355 2922.000 ;
      LAYER met4 ;
        RECT 147.275 2896.065 148.255 2920.330 ;
      LAYER met4 ;
        RECT 148.655 2896.465 151.635 3110.145 ;
        RECT 151.935 3105.090 152.265 3276.610 ;
      LAYER met4 ;
        RECT 152.665 3275.670 199.465 3277.010 ;
        RECT 152.665 3274.965 153.365 3275.670 ;
        RECT 152.665 3136.330 153.365 3136.970 ;
      LAYER met4 ;
        RECT 153.765 3136.730 158.415 3275.270 ;
      LAYER met4 ;
        RECT 158.815 3274.965 159.415 3275.670 ;
        RECT 158.815 3136.330 159.415 3136.970 ;
      LAYER met4 ;
        RECT 159.815 3136.730 163.265 3275.270 ;
      LAYER met4 ;
        RECT 163.665 3274.965 164.265 3275.670 ;
        RECT 163.665 3136.330 164.265 3136.970 ;
      LAYER met4 ;
        RECT 164.665 3136.730 168.115 3275.270 ;
      LAYER met4 ;
        RECT 168.515 3274.965 169.115 3275.670 ;
        RECT 168.515 3136.330 169.115 3136.970 ;
      LAYER met4 ;
        RECT 169.515 3136.730 174.165 3275.270 ;
      LAYER met4 ;
        RECT 174.565 3274.965 175.165 3275.670 ;
        RECT 180.615 3275.365 186.065 3275.670 ;
        RECT 174.565 3136.330 175.165 3136.970 ;
      LAYER met4 ;
        RECT 175.565 3136.730 180.215 3275.270 ;
      LAYER met4 ;
        RECT 180.615 3274.965 181.215 3275.365 ;
        RECT 185.465 3274.965 186.065 3275.365 ;
      LAYER met4 ;
        RECT 181.615 3136.970 185.065 3274.965 ;
      LAYER met4 ;
        RECT 180.615 3136.570 181.215 3136.970 ;
        RECT 185.465 3136.570 186.065 3136.970 ;
      LAYER met4 ;
        RECT 186.465 3136.730 191.115 3275.270 ;
      LAYER met4 ;
        RECT 191.515 3274.965 192.115 3275.670 ;
        RECT 180.615 3136.330 186.065 3136.570 ;
        RECT 191.515 3136.330 192.115 3136.970 ;
      LAYER met4 ;
        RECT 192.515 3136.730 197.965 3275.270 ;
      LAYER met4 ;
        RECT 198.365 3274.965 199.465 3275.670 ;
        RECT 3388.535 3268.330 3389.635 3269.035 ;
      LAYER met4 ;
        RECT 3390.035 3268.730 3395.485 3417.270 ;
      LAYER met4 ;
        RECT 3395.885 3417.030 3396.485 3417.670 ;
        RECT 3401.935 3417.430 3407.385 3417.670 ;
        RECT 3395.885 3268.330 3396.485 3269.035 ;
      LAYER met4 ;
        RECT 3396.885 3268.730 3401.535 3417.270 ;
      LAYER met4 ;
        RECT 3401.935 3417.030 3402.535 3417.430 ;
        RECT 3406.785 3417.030 3407.385 3417.430 ;
      LAYER met4 ;
        RECT 3402.935 3269.035 3406.385 3417.030 ;
      LAYER met4 ;
        RECT 3401.935 3268.635 3402.535 3269.035 ;
        RECT 3406.785 3268.635 3407.385 3269.035 ;
      LAYER met4 ;
        RECT 3407.785 3268.730 3412.435 3417.270 ;
      LAYER met4 ;
        RECT 3412.835 3417.030 3413.435 3417.670 ;
        RECT 3401.935 3268.330 3407.385 3268.635 ;
        RECT 3412.835 3268.330 3413.435 3269.035 ;
      LAYER met4 ;
        RECT 3413.835 3268.730 3418.485 3417.270 ;
      LAYER met4 ;
        RECT 3418.885 3417.030 3419.485 3417.670 ;
        RECT 3418.885 3268.330 3419.485 3269.035 ;
      LAYER met4 ;
        RECT 3419.885 3268.730 3423.335 3417.270 ;
      LAYER met4 ;
        RECT 3423.735 3417.030 3424.335 3417.670 ;
        RECT 3423.735 3268.330 3424.335 3269.035 ;
      LAYER met4 ;
        RECT 3424.735 3268.730 3428.185 3417.270 ;
      LAYER met4 ;
        RECT 3428.585 3417.030 3429.185 3417.670 ;
        RECT 3428.585 3268.330 3429.185 3269.035 ;
      LAYER met4 ;
        RECT 3429.585 3268.730 3434.235 3417.270 ;
      LAYER met4 ;
        RECT 3434.635 3417.030 3435.335 3417.670 ;
        RECT 3434.635 3268.330 3435.335 3269.035 ;
        RECT 3388.535 3266.990 3435.335 3268.330 ;
      LAYER met4 ;
        RECT 3435.735 3267.390 3436.065 3448.910 ;
        RECT 3436.365 3443.855 3439.345 3666.535 ;
      LAYER met4 ;
        RECT 3439.745 3642.670 3440.725 3666.935 ;
      LAYER met4 ;
        RECT 3439.645 3641.000 3440.825 3642.270 ;
      LAYER met4 ;
        RECT 3439.645 3496.000 3440.825 3641.000 ;
      LAYER met4 ;
        RECT 3439.645 3494.730 3440.825 3496.000 ;
      LAYER met4 ;
        RECT 3439.745 3459.160 3440.725 3494.330 ;
      LAYER met4 ;
        RECT 3441.125 3459.560 3444.105 3682.240 ;
      LAYER met4 ;
        RECT 3444.505 3674.310 3588.000 3682.640 ;
      LAYER met4 ;
        RECT 3444.405 3493.390 3444.735 3673.910 ;
      LAYER met4 ;
        RECT 3445.135 3642.670 3588.000 3674.310 ;
        RECT 3445.135 3642.030 3445.835 3642.670 ;
        RECT 3445.135 3496.000 3445.835 3641.000 ;
        RECT 3445.135 3494.330 3445.835 3495.035 ;
      LAYER met4 ;
        RECT 3446.235 3494.730 3450.685 3642.270 ;
      LAYER met4 ;
        RECT 3451.085 3642.030 3451.685 3642.670 ;
        RECT 3451.085 3496.000 3451.685 3641.000 ;
        RECT 3451.085 3494.330 3451.685 3495.035 ;
      LAYER met4 ;
        RECT 3452.085 3494.730 3456.535 3642.270 ;
      LAYER met4 ;
        RECT 3456.935 3642.030 3457.635 3642.670 ;
        RECT 3456.935 3496.000 3457.635 3641.000 ;
        RECT 3456.935 3494.330 3457.635 3495.035 ;
      LAYER met4 ;
        RECT 3458.035 3494.730 3483.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.400 3642.030 3563.385 3642.670 ;
      LAYER met4 ;
        RECT 3563.785 3641.000 3588.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.400 3496.000 3588.000 3641.000 ;
        RECT 3483.400 3494.330 3563.385 3495.035 ;
      LAYER met4 ;
        RECT 3563.785 3494.730 3588.000 3496.000 ;
      LAYER met4 ;
        RECT 3445.135 3492.990 3588.000 3494.330 ;
        RECT 3444.505 3459.160 3588.000 3492.990 ;
        RECT 3439.745 3457.640 3588.000 3459.160 ;
        RECT 3439.745 3443.455 3440.725 3457.640 ;
        RECT 3436.465 3441.935 3440.725 3443.455 ;
        RECT 3388.535 3223.310 3435.965 3266.990 ;
        RECT 3388.535 3191.670 3435.335 3223.310 ;
        RECT 3388.535 3191.030 3389.635 3191.670 ;
        RECT 198.365 3136.330 199.465 3136.970 ;
        RECT 152.665 3104.690 199.465 3136.330 ;
        RECT 152.035 3061.010 199.465 3104.690 ;
        RECT 147.275 2894.545 151.535 2896.065 ;
        RECT 147.275 2880.360 148.255 2894.545 ;
        RECT 0.000 2878.840 148.255 2880.360 ;
        RECT 0.000 2845.010 143.495 2878.840 ;
        RECT 0.000 2843.670 142.865 2845.010 ;
      LAYER met4 ;
        RECT 0.000 2842.000 24.215 2843.270 ;
      LAYER met4 ;
        RECT 24.615 2842.965 104.600 2843.670 ;
        RECT 0.000 2706.000 104.600 2842.000 ;
      LAYER met4 ;
        RECT 0.000 2704.730 24.215 2706.000 ;
      LAYER met4 ;
        RECT 24.615 2704.330 104.600 2704.970 ;
      LAYER met4 ;
        RECT 105.000 2704.730 129.965 2843.270 ;
      LAYER met4 ;
        RECT 130.365 2842.965 131.065 2843.670 ;
        RECT 130.365 2706.000 131.065 2842.000 ;
        RECT 130.365 2704.330 131.065 2704.970 ;
      LAYER met4 ;
        RECT 131.465 2704.730 135.915 2843.270 ;
      LAYER met4 ;
        RECT 136.315 2842.965 136.915 2843.670 ;
        RECT 136.315 2706.000 136.915 2842.000 ;
        RECT 136.315 2704.330 136.915 2704.970 ;
      LAYER met4 ;
        RECT 137.315 2704.730 141.765 2843.270 ;
      LAYER met4 ;
        RECT 142.165 2842.965 142.865 2843.670 ;
        RECT 142.165 2706.000 142.865 2842.000 ;
        RECT 142.165 2704.330 142.865 2704.970 ;
        RECT 0.000 2672.690 142.865 2704.330 ;
      LAYER met4 ;
        RECT 143.265 2673.090 143.595 2844.610 ;
      LAYER met4 ;
        RECT 0.000 2664.360 143.495 2672.690 ;
      LAYER met4 ;
        RECT 143.895 2664.760 146.875 2878.440 ;
      LAYER met4 ;
        RECT 147.275 2843.670 148.255 2878.840 ;
      LAYER met4 ;
        RECT 147.175 2842.000 148.355 2843.270 ;
      LAYER met4 ;
        RECT 147.175 2706.000 148.355 2842.000 ;
      LAYER met4 ;
        RECT 147.175 2704.730 148.355 2706.000 ;
      LAYER met4 ;
        RECT 147.275 2680.065 148.255 2704.330 ;
      LAYER met4 ;
        RECT 148.655 2680.465 151.635 2894.145 ;
        RECT 151.935 2889.090 152.265 3060.610 ;
      LAYER met4 ;
        RECT 152.665 3059.670 199.465 3061.010 ;
        RECT 152.665 3058.965 153.365 3059.670 ;
        RECT 152.665 2920.330 153.365 2920.970 ;
      LAYER met4 ;
        RECT 153.765 2920.730 158.415 3059.270 ;
      LAYER met4 ;
        RECT 158.815 3058.965 159.415 3059.670 ;
        RECT 158.815 2920.330 159.415 2920.970 ;
      LAYER met4 ;
        RECT 159.815 2920.730 163.265 3059.270 ;
      LAYER met4 ;
        RECT 163.665 3058.965 164.265 3059.670 ;
        RECT 163.665 2920.330 164.265 2920.970 ;
      LAYER met4 ;
        RECT 164.665 2920.730 168.115 3059.270 ;
      LAYER met4 ;
        RECT 168.515 3058.965 169.115 3059.670 ;
        RECT 168.515 2920.330 169.115 2920.970 ;
      LAYER met4 ;
        RECT 169.515 2920.730 174.165 3059.270 ;
      LAYER met4 ;
        RECT 174.565 3058.965 175.165 3059.670 ;
        RECT 180.615 3059.365 186.065 3059.670 ;
        RECT 174.565 2920.330 175.165 2920.970 ;
      LAYER met4 ;
        RECT 175.565 2920.730 180.215 3059.270 ;
      LAYER met4 ;
        RECT 180.615 3058.965 181.215 3059.365 ;
        RECT 185.465 3058.965 186.065 3059.365 ;
      LAYER met4 ;
        RECT 181.615 2920.970 185.065 3058.965 ;
      LAYER met4 ;
        RECT 180.615 2920.570 181.215 2920.970 ;
        RECT 185.465 2920.570 186.065 2920.970 ;
      LAYER met4 ;
        RECT 186.465 2920.730 191.115 3059.270 ;
      LAYER met4 ;
        RECT 191.515 3058.965 192.115 3059.670 ;
        RECT 180.615 2920.330 186.065 2920.570 ;
        RECT 191.515 2920.330 192.115 2920.970 ;
      LAYER met4 ;
        RECT 192.515 2920.730 197.965 3059.270 ;
      LAYER met4 ;
        RECT 198.365 3058.965 199.465 3059.670 ;
        RECT 3388.535 3043.330 3389.635 3044.035 ;
      LAYER met4 ;
        RECT 3390.035 3043.730 3395.485 3191.270 ;
      LAYER met4 ;
        RECT 3395.885 3191.030 3396.485 3191.670 ;
        RECT 3401.935 3191.430 3407.385 3191.670 ;
        RECT 3395.885 3043.330 3396.485 3044.035 ;
      LAYER met4 ;
        RECT 3396.885 3043.730 3401.535 3191.270 ;
      LAYER met4 ;
        RECT 3401.935 3191.030 3402.535 3191.430 ;
        RECT 3406.785 3191.030 3407.385 3191.430 ;
      LAYER met4 ;
        RECT 3402.935 3044.035 3406.385 3191.030 ;
      LAYER met4 ;
        RECT 3401.935 3043.635 3402.535 3044.035 ;
        RECT 3406.785 3043.635 3407.385 3044.035 ;
      LAYER met4 ;
        RECT 3407.785 3043.730 3412.435 3191.270 ;
      LAYER met4 ;
        RECT 3412.835 3191.030 3413.435 3191.670 ;
        RECT 3401.935 3043.330 3407.385 3043.635 ;
        RECT 3412.835 3043.330 3413.435 3044.035 ;
      LAYER met4 ;
        RECT 3413.835 3043.730 3418.485 3191.270 ;
      LAYER met4 ;
        RECT 3418.885 3191.030 3419.485 3191.670 ;
        RECT 3418.885 3043.330 3419.485 3044.035 ;
      LAYER met4 ;
        RECT 3419.885 3043.730 3423.335 3191.270 ;
      LAYER met4 ;
        RECT 3423.735 3191.030 3424.335 3191.670 ;
        RECT 3423.735 3043.330 3424.335 3044.035 ;
      LAYER met4 ;
        RECT 3424.735 3043.730 3428.185 3191.270 ;
      LAYER met4 ;
        RECT 3428.585 3191.030 3429.185 3191.670 ;
        RECT 3428.585 3043.330 3429.185 3044.035 ;
      LAYER met4 ;
        RECT 3429.585 3043.730 3434.235 3191.270 ;
      LAYER met4 ;
        RECT 3434.635 3191.030 3435.335 3191.670 ;
        RECT 3434.635 3043.330 3435.335 3044.035 ;
        RECT 3388.535 3041.990 3435.335 3043.330 ;
      LAYER met4 ;
        RECT 3435.735 3042.390 3436.065 3222.910 ;
        RECT 3436.365 3217.855 3439.345 3441.535 ;
      LAYER met4 ;
        RECT 3439.745 3417.670 3440.725 3441.935 ;
      LAYER met4 ;
        RECT 3439.645 3416.000 3440.825 3417.270 ;
      LAYER met4 ;
        RECT 3439.645 3270.000 3440.825 3416.000 ;
      LAYER met4 ;
        RECT 3439.645 3268.730 3440.825 3270.000 ;
      LAYER met4 ;
        RECT 3439.745 3233.160 3440.725 3268.330 ;
      LAYER met4 ;
        RECT 3441.125 3233.560 3444.105 3457.240 ;
      LAYER met4 ;
        RECT 3444.505 3449.310 3588.000 3457.640 ;
      LAYER met4 ;
        RECT 3444.405 3267.390 3444.735 3448.910 ;
      LAYER met4 ;
        RECT 3445.135 3417.670 3588.000 3449.310 ;
        RECT 3445.135 3417.030 3445.835 3417.670 ;
        RECT 3445.135 3270.000 3445.835 3416.000 ;
        RECT 3445.135 3268.330 3445.835 3269.035 ;
      LAYER met4 ;
        RECT 3446.235 3268.730 3450.685 3417.270 ;
      LAYER met4 ;
        RECT 3451.085 3417.030 3451.685 3417.670 ;
        RECT 3451.085 3270.000 3451.685 3416.000 ;
        RECT 3451.085 3268.330 3451.685 3269.035 ;
      LAYER met4 ;
        RECT 3452.085 3268.730 3456.535 3417.270 ;
      LAYER met4 ;
        RECT 3456.935 3417.030 3457.635 3417.670 ;
        RECT 3456.935 3270.000 3457.635 3416.000 ;
        RECT 3456.935 3268.330 3457.635 3269.035 ;
      LAYER met4 ;
        RECT 3458.035 3268.730 3483.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.400 3417.030 3563.385 3417.670 ;
      LAYER met4 ;
        RECT 3563.785 3416.000 3588.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.400 3270.000 3588.000 3416.000 ;
        RECT 3483.400 3268.330 3563.385 3269.035 ;
      LAYER met4 ;
        RECT 3563.785 3268.730 3588.000 3270.000 ;
      LAYER met4 ;
        RECT 3445.135 3266.990 3588.000 3268.330 ;
        RECT 3444.505 3233.160 3588.000 3266.990 ;
        RECT 3439.745 3231.640 3588.000 3233.160 ;
        RECT 3439.745 3217.455 3440.725 3231.640 ;
        RECT 3436.465 3215.935 3440.725 3217.455 ;
        RECT 3388.535 2998.310 3435.965 3041.990 ;
        RECT 3388.535 2966.670 3435.335 2998.310 ;
        RECT 3388.535 2966.030 3389.635 2966.670 ;
        RECT 198.365 2920.330 199.465 2920.970 ;
        RECT 152.665 2888.690 199.465 2920.330 ;
        RECT 152.035 2845.010 199.465 2888.690 ;
        RECT 147.275 2678.545 151.535 2680.065 ;
        RECT 147.275 2664.360 148.255 2678.545 ;
        RECT 0.000 2662.840 148.255 2664.360 ;
        RECT 0.000 2629.010 143.495 2662.840 ;
        RECT 0.000 2627.670 142.865 2629.010 ;
      LAYER met4 ;
        RECT 0.000 2626.000 24.215 2627.270 ;
      LAYER met4 ;
        RECT 24.615 2626.965 104.600 2627.670 ;
        RECT 0.000 2490.000 104.600 2626.000 ;
      LAYER met4 ;
        RECT 0.000 2488.730 24.215 2490.000 ;
      LAYER met4 ;
        RECT 24.615 2488.330 104.600 2489.035 ;
      LAYER met4 ;
        RECT 105.000 2488.730 129.965 2627.270 ;
      LAYER met4 ;
        RECT 130.365 2626.965 131.065 2627.670 ;
        RECT 130.365 2490.000 131.065 2626.000 ;
        RECT 130.365 2488.330 131.065 2489.035 ;
      LAYER met4 ;
        RECT 131.465 2488.730 135.915 2627.270 ;
      LAYER met4 ;
        RECT 136.315 2626.965 136.915 2627.670 ;
        RECT 136.315 2490.000 136.915 2626.000 ;
        RECT 136.315 2488.330 136.915 2489.035 ;
      LAYER met4 ;
        RECT 137.315 2488.730 141.765 2627.270 ;
      LAYER met4 ;
        RECT 142.165 2626.965 142.865 2627.670 ;
        RECT 142.165 2490.000 142.865 2626.000 ;
        RECT 142.165 2488.330 142.865 2489.035 ;
        RECT 0.000 2416.670 142.865 2488.330 ;
      LAYER met4 ;
        RECT 0.000 2415.000 24.215 2416.270 ;
      LAYER met4 ;
        RECT 24.615 2415.965 104.600 2416.670 ;
        RECT 0.000 2280.465 104.600 2415.000 ;
        RECT 0.000 2279.000 0.035 2280.465 ;
        RECT 24.215 2279.000 104.600 2280.465 ;
        RECT 24.215 2278.785 24.250 2279.000 ;
        RECT 24.615 2277.330 104.600 2279.000 ;
      LAYER met4 ;
        RECT 105.000 2277.730 129.965 2416.270 ;
      LAYER met4 ;
        RECT 130.365 2415.965 131.065 2416.670 ;
        RECT 130.365 2277.330 131.065 2415.000 ;
      LAYER met4 ;
        RECT 131.465 2277.730 135.915 2416.270 ;
      LAYER met4 ;
        RECT 136.315 2415.965 136.915 2416.670 ;
        RECT 136.315 2277.330 136.915 2415.000 ;
      LAYER met4 ;
        RECT 137.315 2277.730 141.765 2416.270 ;
      LAYER met4 ;
        RECT 142.165 2415.965 142.865 2416.670 ;
        RECT 142.165 2277.330 142.865 2415.000 ;
        RECT 0.000 2205.670 142.865 2277.330 ;
      LAYER met4 ;
        RECT 0.000 2204.000 24.215 2205.270 ;
      LAYER met4 ;
        RECT 24.615 2204.000 104.600 2205.670 ;
        RECT 0.000 2068.000 104.600 2204.000 ;
      LAYER met4 ;
        RECT 0.000 2066.730 24.215 2068.000 ;
      LAYER met4 ;
        RECT 24.615 2066.330 104.600 2066.970 ;
      LAYER met4 ;
        RECT 105.000 2066.730 129.965 2205.270 ;
      LAYER met4 ;
        RECT 130.365 2068.000 131.065 2205.670 ;
        RECT 130.365 2066.330 131.065 2066.970 ;
      LAYER met4 ;
        RECT 131.465 2066.730 135.915 2205.270 ;
      LAYER met4 ;
        RECT 136.315 2068.000 136.915 2205.670 ;
        RECT 136.315 2066.330 136.915 2066.970 ;
      LAYER met4 ;
        RECT 137.315 2066.730 141.765 2205.270 ;
      LAYER met4 ;
        RECT 142.165 2068.000 142.865 2205.670 ;
        RECT 142.165 2066.330 142.865 2066.970 ;
        RECT 0.000 2034.690 142.865 2066.330 ;
        RECT 0.000 2026.360 143.495 2034.690 ;
      LAYER met4 ;
        RECT 143.895 2026.760 146.875 2662.440 ;
      LAYER met4 ;
        RECT 147.275 2627.670 148.255 2662.840 ;
      LAYER met4 ;
        RECT 147.175 2626.000 148.355 2627.270 ;
      LAYER met4 ;
        RECT 147.175 2490.000 148.355 2626.000 ;
      LAYER met4 ;
        RECT 147.175 2488.730 148.355 2490.000 ;
      LAYER met4 ;
        RECT 147.275 2416.670 148.255 2488.330 ;
      LAYER met4 ;
        RECT 147.175 2415.000 148.355 2416.270 ;
      LAYER met4 ;
        RECT 147.175 2279.000 148.355 2415.000 ;
      LAYER met4 ;
        RECT 147.175 2277.730 148.355 2279.000 ;
      LAYER met4 ;
        RECT 147.275 2205.670 148.255 2277.330 ;
      LAYER met4 ;
        RECT 147.175 2204.000 148.355 2205.270 ;
      LAYER met4 ;
        RECT 147.175 2068.000 148.355 2204.000 ;
      LAYER met4 ;
        RECT 147.175 2066.730 148.355 2068.000 ;
      LAYER met4 ;
        RECT 147.275 2042.065 148.255 2066.330 ;
      LAYER met4 ;
        RECT 148.655 2042.465 151.635 2678.145 ;
        RECT 151.935 2673.090 152.265 2844.610 ;
      LAYER met4 ;
        RECT 152.665 2843.670 199.465 2845.010 ;
        RECT 152.665 2842.965 153.365 2843.670 ;
        RECT 152.665 2704.330 153.365 2704.970 ;
      LAYER met4 ;
        RECT 153.765 2704.730 158.415 2843.270 ;
      LAYER met4 ;
        RECT 158.815 2842.965 159.415 2843.670 ;
        RECT 158.815 2704.330 159.415 2704.970 ;
      LAYER met4 ;
        RECT 159.815 2704.730 163.265 2843.270 ;
      LAYER met4 ;
        RECT 163.665 2842.965 164.265 2843.670 ;
        RECT 163.665 2704.330 164.265 2704.970 ;
      LAYER met4 ;
        RECT 164.665 2704.730 168.115 2843.270 ;
      LAYER met4 ;
        RECT 168.515 2842.965 169.115 2843.670 ;
        RECT 168.515 2704.330 169.115 2704.970 ;
      LAYER met4 ;
        RECT 169.515 2704.730 174.165 2843.270 ;
      LAYER met4 ;
        RECT 174.565 2842.965 175.165 2843.670 ;
        RECT 180.615 2843.365 186.065 2843.670 ;
        RECT 174.565 2704.330 175.165 2704.970 ;
      LAYER met4 ;
        RECT 175.565 2704.730 180.215 2843.270 ;
      LAYER met4 ;
        RECT 180.615 2842.965 181.215 2843.365 ;
        RECT 185.465 2842.965 186.065 2843.365 ;
      LAYER met4 ;
        RECT 181.615 2704.970 185.065 2842.965 ;
      LAYER met4 ;
        RECT 180.615 2704.570 181.215 2704.970 ;
        RECT 185.465 2704.570 186.065 2704.970 ;
      LAYER met4 ;
        RECT 186.465 2704.730 191.115 2843.270 ;
      LAYER met4 ;
        RECT 191.515 2842.965 192.115 2843.670 ;
        RECT 180.615 2704.330 186.065 2704.570 ;
        RECT 191.515 2704.330 192.115 2704.970 ;
      LAYER met4 ;
        RECT 192.515 2704.730 197.965 2843.270 ;
      LAYER met4 ;
        RECT 198.365 2842.965 199.465 2843.670 ;
        RECT 3388.535 2817.330 3389.635 2818.035 ;
      LAYER met4 ;
        RECT 3390.035 2817.730 3395.485 2966.270 ;
      LAYER met4 ;
        RECT 3395.885 2966.030 3396.485 2966.670 ;
        RECT 3401.935 2966.430 3407.385 2966.670 ;
        RECT 3395.885 2817.330 3396.485 2818.035 ;
      LAYER met4 ;
        RECT 3396.885 2817.730 3401.535 2966.270 ;
      LAYER met4 ;
        RECT 3401.935 2966.030 3402.535 2966.430 ;
        RECT 3406.785 2966.030 3407.385 2966.430 ;
      LAYER met4 ;
        RECT 3402.935 2818.035 3406.385 2966.030 ;
      LAYER met4 ;
        RECT 3401.935 2817.635 3402.535 2818.035 ;
        RECT 3406.785 2817.635 3407.385 2818.035 ;
      LAYER met4 ;
        RECT 3407.785 2817.730 3412.435 2966.270 ;
      LAYER met4 ;
        RECT 3412.835 2966.030 3413.435 2966.670 ;
        RECT 3401.935 2817.330 3407.385 2817.635 ;
        RECT 3412.835 2817.330 3413.435 2818.035 ;
      LAYER met4 ;
        RECT 3413.835 2817.730 3418.485 2966.270 ;
      LAYER met4 ;
        RECT 3418.885 2966.030 3419.485 2966.670 ;
        RECT 3418.885 2817.330 3419.485 2818.035 ;
      LAYER met4 ;
        RECT 3419.885 2817.730 3423.335 2966.270 ;
      LAYER met4 ;
        RECT 3423.735 2966.030 3424.335 2966.670 ;
        RECT 3423.735 2817.330 3424.335 2818.035 ;
      LAYER met4 ;
        RECT 3424.735 2817.730 3428.185 2966.270 ;
      LAYER met4 ;
        RECT 3428.585 2966.030 3429.185 2966.670 ;
        RECT 3428.585 2817.330 3429.185 2818.035 ;
      LAYER met4 ;
        RECT 3429.585 2817.730 3434.235 2966.270 ;
      LAYER met4 ;
        RECT 3434.635 2966.030 3435.335 2966.670 ;
        RECT 3434.635 2817.330 3435.335 2818.035 ;
        RECT 3388.535 2815.990 3435.335 2817.330 ;
      LAYER met4 ;
        RECT 3435.735 2816.390 3436.065 2997.910 ;
        RECT 3436.365 2992.855 3439.345 3215.535 ;
      LAYER met4 ;
        RECT 3439.745 3191.670 3440.725 3215.935 ;
      LAYER met4 ;
        RECT 3439.645 3190.000 3440.825 3191.270 ;
      LAYER met4 ;
        RECT 3439.645 3045.000 3440.825 3190.000 ;
      LAYER met4 ;
        RECT 3439.645 3043.730 3440.825 3045.000 ;
      LAYER met4 ;
        RECT 3439.745 3008.160 3440.725 3043.330 ;
      LAYER met4 ;
        RECT 3441.125 3008.560 3444.105 3231.240 ;
      LAYER met4 ;
        RECT 3444.505 3223.310 3588.000 3231.640 ;
      LAYER met4 ;
        RECT 3444.405 3042.390 3444.735 3222.910 ;
      LAYER met4 ;
        RECT 3445.135 3191.670 3588.000 3223.310 ;
        RECT 3445.135 3191.030 3445.835 3191.670 ;
        RECT 3445.135 3045.000 3445.835 3190.000 ;
        RECT 3445.135 3043.330 3445.835 3044.035 ;
      LAYER met4 ;
        RECT 3446.235 3043.730 3450.685 3191.270 ;
      LAYER met4 ;
        RECT 3451.085 3191.030 3451.685 3191.670 ;
        RECT 3451.085 3045.000 3451.685 3190.000 ;
        RECT 3451.085 3043.330 3451.685 3044.035 ;
      LAYER met4 ;
        RECT 3452.085 3043.730 3456.535 3191.270 ;
      LAYER met4 ;
        RECT 3456.935 3191.030 3457.635 3191.670 ;
        RECT 3456.935 3045.000 3457.635 3190.000 ;
        RECT 3456.935 3043.330 3457.635 3044.035 ;
      LAYER met4 ;
        RECT 3458.035 3043.730 3483.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.400 3191.030 3563.385 3191.670 ;
      LAYER met4 ;
        RECT 3563.785 3190.000 3588.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.400 3045.000 3588.000 3190.000 ;
        RECT 3483.400 3043.330 3563.385 3044.035 ;
      LAYER met4 ;
        RECT 3563.785 3043.730 3588.000 3045.000 ;
      LAYER met4 ;
        RECT 3445.135 3041.990 3588.000 3043.330 ;
        RECT 3444.505 3008.160 3588.000 3041.990 ;
        RECT 3439.745 3006.640 3588.000 3008.160 ;
        RECT 3439.745 2992.455 3440.725 3006.640 ;
        RECT 3436.465 2990.935 3440.725 2992.455 ;
        RECT 3388.535 2772.310 3435.965 2815.990 ;
        RECT 3388.535 2740.670 3435.335 2772.310 ;
        RECT 3388.535 2740.030 3389.635 2740.670 ;
        RECT 198.365 2704.330 199.465 2704.970 ;
        RECT 152.665 2672.690 199.465 2704.330 ;
        RECT 152.035 2629.010 199.465 2672.690 ;
        RECT 147.275 2040.545 151.535 2042.065 ;
        RECT 147.275 2026.360 148.255 2040.545 ;
        RECT 0.000 2024.840 148.255 2026.360 ;
        RECT 0.000 1991.010 143.495 2024.840 ;
        RECT 0.000 1989.670 142.865 1991.010 ;
      LAYER met4 ;
        RECT 0.000 1988.000 24.215 1989.270 ;
      LAYER met4 ;
        RECT 24.615 1988.965 104.600 1989.670 ;
        RECT 0.000 1852.000 104.600 1988.000 ;
      LAYER met4 ;
        RECT 0.000 1850.730 24.215 1852.000 ;
      LAYER met4 ;
        RECT 24.615 1850.330 104.600 1850.970 ;
      LAYER met4 ;
        RECT 105.000 1850.730 129.965 1989.270 ;
      LAYER met4 ;
        RECT 130.365 1988.965 131.065 1989.670 ;
        RECT 130.365 1852.000 131.065 1988.000 ;
        RECT 130.365 1850.330 131.065 1850.970 ;
      LAYER met4 ;
        RECT 131.465 1850.730 135.915 1989.270 ;
      LAYER met4 ;
        RECT 136.315 1988.965 136.915 1989.670 ;
        RECT 136.315 1852.000 136.915 1988.000 ;
        RECT 136.315 1850.330 136.915 1850.970 ;
      LAYER met4 ;
        RECT 137.315 1850.730 141.765 1989.270 ;
      LAYER met4 ;
        RECT 142.165 1988.965 142.865 1989.670 ;
        RECT 142.165 1852.000 142.865 1988.000 ;
        RECT 142.165 1850.330 142.865 1850.970 ;
        RECT 0.000 1818.690 142.865 1850.330 ;
      LAYER met4 ;
        RECT 143.265 1819.090 143.595 1990.610 ;
      LAYER met4 ;
        RECT 0.000 1810.360 143.495 1818.690 ;
      LAYER met4 ;
        RECT 143.895 1810.760 146.875 2024.440 ;
      LAYER met4 ;
        RECT 147.275 1989.670 148.255 2024.840 ;
      LAYER met4 ;
        RECT 147.175 1988.000 148.355 1989.270 ;
      LAYER met4 ;
        RECT 147.175 1852.000 148.355 1988.000 ;
      LAYER met4 ;
        RECT 147.175 1850.730 148.355 1852.000 ;
      LAYER met4 ;
        RECT 147.275 1826.065 148.255 1850.330 ;
      LAYER met4 ;
        RECT 148.655 1826.465 151.635 2040.145 ;
        RECT 151.935 2035.090 152.265 2628.610 ;
      LAYER met4 ;
        RECT 152.665 2627.670 199.465 2629.010 ;
        RECT 152.665 2626.965 153.365 2627.670 ;
        RECT 152.665 2488.330 153.365 2489.035 ;
      LAYER met4 ;
        RECT 153.765 2488.730 158.415 2627.270 ;
      LAYER met4 ;
        RECT 158.815 2626.965 159.415 2627.670 ;
        RECT 158.815 2488.330 159.415 2489.035 ;
      LAYER met4 ;
        RECT 159.815 2488.730 163.265 2627.270 ;
      LAYER met4 ;
        RECT 163.665 2626.965 164.265 2627.670 ;
        RECT 163.665 2488.330 164.265 2489.035 ;
      LAYER met4 ;
        RECT 164.665 2488.730 168.115 2627.270 ;
      LAYER met4 ;
        RECT 168.515 2626.965 169.115 2627.670 ;
        RECT 168.515 2488.330 169.115 2489.035 ;
      LAYER met4 ;
        RECT 169.515 2488.730 174.165 2627.270 ;
      LAYER met4 ;
        RECT 174.565 2626.965 175.165 2627.670 ;
        RECT 180.615 2627.365 186.065 2627.670 ;
        RECT 174.565 2488.330 175.165 2489.035 ;
      LAYER met4 ;
        RECT 175.565 2488.730 180.215 2627.270 ;
      LAYER met4 ;
        RECT 180.615 2626.965 181.215 2627.365 ;
        RECT 185.465 2626.965 186.065 2627.365 ;
      LAYER met4 ;
        RECT 181.615 2489.035 185.065 2626.965 ;
      LAYER met4 ;
        RECT 180.615 2488.635 181.215 2489.035 ;
        RECT 185.465 2488.635 186.065 2489.035 ;
      LAYER met4 ;
        RECT 186.465 2488.730 191.115 2627.270 ;
      LAYER met4 ;
        RECT 191.515 2626.965 192.115 2627.670 ;
        RECT 180.615 2488.330 186.065 2488.635 ;
        RECT 191.515 2488.330 192.115 2489.035 ;
      LAYER met4 ;
        RECT 192.515 2488.730 197.965 2627.270 ;
      LAYER met4 ;
        RECT 198.365 2626.965 199.465 2627.670 ;
      LAYER met4 ;
        RECT 3390.035 2592.730 3395.485 2740.270 ;
      LAYER met4 ;
        RECT 3395.885 2740.030 3396.485 2740.670 ;
        RECT 3401.935 2740.430 3407.385 2740.670 ;
        RECT 3395.885 2592.330 3396.485 2593.035 ;
      LAYER met4 ;
        RECT 3396.885 2592.730 3401.535 2740.270 ;
      LAYER met4 ;
        RECT 3401.935 2740.030 3402.535 2740.430 ;
        RECT 3406.785 2740.030 3407.385 2740.430 ;
      LAYER met4 ;
        RECT 3402.935 2593.035 3406.385 2740.030 ;
      LAYER met4 ;
        RECT 3401.935 2592.635 3402.535 2593.035 ;
        RECT 3406.785 2592.635 3407.385 2593.035 ;
      LAYER met4 ;
        RECT 3407.785 2592.730 3412.435 2740.270 ;
      LAYER met4 ;
        RECT 3412.835 2740.030 3413.435 2740.670 ;
        RECT 3401.935 2592.330 3407.385 2592.635 ;
        RECT 3412.835 2592.330 3413.435 2593.035 ;
      LAYER met4 ;
        RECT 3413.835 2592.730 3418.485 2740.270 ;
      LAYER met4 ;
        RECT 3418.885 2740.030 3419.485 2740.670 ;
        RECT 3418.885 2592.330 3419.485 2593.035 ;
      LAYER met4 ;
        RECT 3419.885 2592.730 3423.335 2740.270 ;
      LAYER met4 ;
        RECT 3423.735 2740.030 3424.335 2740.670 ;
        RECT 3423.735 2592.330 3424.335 2593.035 ;
      LAYER met4 ;
        RECT 3424.735 2592.730 3428.185 2740.270 ;
      LAYER met4 ;
        RECT 3428.585 2740.030 3429.185 2740.670 ;
        RECT 3428.585 2592.330 3429.185 2593.035 ;
      LAYER met4 ;
        RECT 3429.585 2592.730 3434.235 2740.270 ;
      LAYER met4 ;
        RECT 3434.635 2740.030 3435.335 2740.670 ;
        RECT 3434.635 2592.330 3435.335 2593.035 ;
        RECT 3390.035 2520.670 3435.335 2592.330 ;
        RECT 152.665 2416.670 197.965 2488.330 ;
        RECT 152.665 2415.965 153.365 2416.670 ;
        RECT 152.665 2277.330 153.365 2279.000 ;
      LAYER met4 ;
        RECT 153.765 2277.730 158.415 2416.270 ;
      LAYER met4 ;
        RECT 158.815 2415.965 159.415 2416.670 ;
        RECT 158.815 2277.330 159.415 2279.000 ;
      LAYER met4 ;
        RECT 159.815 2277.730 163.265 2416.270 ;
      LAYER met4 ;
        RECT 163.665 2415.965 164.265 2416.670 ;
        RECT 168.515 2415.965 169.115 2416.670 ;
        RECT 163.665 2277.330 164.265 2279.000 ;
        RECT 168.515 2277.330 169.115 2279.000 ;
      LAYER met4 ;
        RECT 169.515 2277.730 174.165 2416.270 ;
      LAYER met4 ;
        RECT 174.565 2415.965 175.165 2416.670 ;
        RECT 180.615 2416.365 186.065 2416.670 ;
        RECT 174.165 2278.935 174.200 2289.935 ;
        RECT 174.565 2277.330 175.165 2279.000 ;
      LAYER met4 ;
        RECT 175.565 2277.730 180.215 2416.270 ;
      LAYER met4 ;
        RECT 180.615 2415.965 181.215 2416.365 ;
        RECT 185.465 2415.965 186.065 2416.365 ;
        RECT 191.515 2415.965 192.115 2416.670 ;
      LAYER met4 ;
        RECT 3390.035 2372.730 3395.485 2520.270 ;
      LAYER met4 ;
        RECT 3395.885 2519.965 3396.485 2520.670 ;
        RECT 3401.935 2520.365 3407.385 2520.670 ;
        RECT 3395.885 2372.330 3396.485 2374.000 ;
      LAYER met4 ;
        RECT 3396.885 2372.730 3401.535 2520.270 ;
      LAYER met4 ;
        RECT 3401.935 2519.965 3402.535 2520.365 ;
        RECT 3406.785 2519.965 3407.385 2520.365 ;
        RECT 3401.935 2372.635 3402.535 2374.000 ;
      LAYER met4 ;
        RECT 3402.935 2373.035 3406.385 2519.965 ;
      LAYER met4 ;
        RECT 3406.785 2372.635 3407.385 2374.000 ;
      LAYER met4 ;
        RECT 3407.785 2372.730 3412.435 2520.270 ;
      LAYER met4 ;
        RECT 3412.835 2519.965 3413.435 2520.670 ;
        RECT 3401.935 2372.330 3407.385 2372.635 ;
        RECT 3412.835 2372.330 3413.435 2374.000 ;
      LAYER met4 ;
        RECT 3413.835 2372.730 3418.485 2520.270 ;
      LAYER met4 ;
        RECT 3418.885 2519.965 3419.485 2520.670 ;
        RECT 3418.885 2372.330 3419.485 2374.000 ;
      LAYER met4 ;
        RECT 3419.885 2372.730 3423.335 2520.270 ;
      LAYER met4 ;
        RECT 3423.735 2519.965 3424.335 2520.670 ;
        RECT 3423.735 2372.330 3424.335 2374.000 ;
      LAYER met4 ;
        RECT 3424.735 2372.730 3428.185 2520.270 ;
      LAYER met4 ;
        RECT 3428.585 2519.965 3429.185 2520.670 ;
        RECT 3428.585 2372.330 3429.185 2374.000 ;
        RECT 3429.550 2373.930 3429.585 2384.975 ;
      LAYER met4 ;
        RECT 3429.585 2372.730 3434.235 2520.270 ;
      LAYER met4 ;
        RECT 3434.635 2519.965 3435.335 2520.670 ;
        RECT 3434.635 2372.330 3435.335 2374.000 ;
        RECT 3390.035 2300.670 3435.335 2372.330 ;
        RECT 180.615 2277.635 181.215 2279.000 ;
        RECT 185.465 2277.635 186.065 2279.000 ;
        RECT 180.615 2277.330 186.065 2277.635 ;
        RECT 191.515 2277.330 192.115 2279.000 ;
        RECT 152.665 2205.670 197.965 2277.330 ;
        RECT 152.665 2204.000 153.365 2205.670 ;
        RECT 152.665 2066.330 153.365 2066.970 ;
      LAYER met4 ;
        RECT 153.765 2066.730 158.415 2205.270 ;
      LAYER met4 ;
        RECT 158.415 2193.025 158.450 2204.070 ;
        RECT 158.815 2204.000 159.415 2205.670 ;
        RECT 158.815 2066.330 159.415 2066.970 ;
      LAYER met4 ;
        RECT 159.815 2066.730 163.265 2205.270 ;
      LAYER met4 ;
        RECT 163.665 2204.000 164.265 2205.670 ;
        RECT 163.665 2066.330 164.265 2066.970 ;
      LAYER met4 ;
        RECT 164.665 2066.730 168.115 2205.270 ;
      LAYER met4 ;
        RECT 168.515 2204.000 169.115 2205.670 ;
        RECT 168.515 2066.330 169.115 2066.970 ;
      LAYER met4 ;
        RECT 169.515 2066.730 174.165 2205.270 ;
      LAYER met4 ;
        RECT 174.565 2204.000 175.165 2205.670 ;
        RECT 180.615 2205.365 186.065 2205.670 ;
        RECT 174.565 2066.330 175.165 2066.970 ;
      LAYER met4 ;
        RECT 175.565 2066.730 180.215 2205.270 ;
      LAYER met4 ;
        RECT 180.615 2204.000 181.215 2205.365 ;
      LAYER met4 ;
        RECT 181.615 2066.970 185.065 2204.965 ;
      LAYER met4 ;
        RECT 185.465 2204.000 186.065 2205.365 ;
        RECT 180.615 2066.570 181.215 2066.970 ;
        RECT 185.465 2066.570 186.065 2066.970 ;
      LAYER met4 ;
        RECT 186.465 2066.730 191.115 2205.270 ;
      LAYER met4 ;
        RECT 191.515 2204.000 192.115 2205.670 ;
        RECT 180.615 2066.330 186.065 2066.570 ;
        RECT 191.515 2066.330 192.115 2066.970 ;
      LAYER met4 ;
        RECT 192.515 2066.730 197.965 2205.270 ;
        RECT 3390.035 2151.730 3395.485 2300.270 ;
      LAYER met4 ;
        RECT 3395.885 2299.000 3396.485 2300.670 ;
        RECT 3401.935 2300.365 3407.385 2300.670 ;
        RECT 3401.935 2299.000 3402.535 2300.365 ;
        RECT 3406.785 2299.000 3407.385 2300.365 ;
        RECT 3395.885 2151.330 3396.485 2152.035 ;
        RECT 3401.935 2151.635 3402.535 2152.035 ;
        RECT 3406.785 2151.635 3407.385 2152.035 ;
      LAYER met4 ;
        RECT 3407.785 2151.730 3412.435 2300.270 ;
      LAYER met4 ;
        RECT 3412.835 2299.000 3413.435 2300.670 ;
        RECT 3413.800 2288.065 3413.835 2299.065 ;
        RECT 3401.935 2151.330 3407.385 2151.635 ;
        RECT 3412.835 2151.330 3413.435 2152.035 ;
      LAYER met4 ;
        RECT 3413.835 2151.730 3418.485 2300.270 ;
      LAYER met4 ;
        RECT 3418.885 2299.000 3419.485 2300.670 ;
        RECT 3418.885 2151.330 3419.485 2152.035 ;
      LAYER met4 ;
        RECT 3419.885 2151.730 3423.335 2300.270 ;
      LAYER met4 ;
        RECT 3423.735 2299.000 3424.335 2300.670 ;
        RECT 3423.735 2151.330 3424.335 2152.035 ;
      LAYER met4 ;
        RECT 3424.735 2151.730 3428.185 2300.270 ;
      LAYER met4 ;
        RECT 3428.585 2299.000 3429.185 2300.670 ;
        RECT 3428.585 2151.330 3429.185 2152.035 ;
      LAYER met4 ;
        RECT 3429.585 2151.730 3434.235 2300.270 ;
      LAYER met4 ;
        RECT 3434.635 2299.000 3435.335 2300.670 ;
        RECT 3434.635 2151.330 3435.335 2152.035 ;
      LAYER met4 ;
        RECT 3435.735 2151.730 3436.065 2771.910 ;
        RECT 3436.365 2766.855 3439.345 2990.535 ;
      LAYER met4 ;
        RECT 3439.745 2966.670 3440.725 2990.935 ;
      LAYER met4 ;
        RECT 3439.645 2965.000 3440.825 2966.270 ;
      LAYER met4 ;
        RECT 3439.645 2819.000 3440.825 2965.000 ;
      LAYER met4 ;
        RECT 3439.645 2817.730 3440.825 2819.000 ;
      LAYER met4 ;
        RECT 3439.745 2782.160 3440.725 2817.330 ;
      LAYER met4 ;
        RECT 3441.125 2782.560 3444.105 3006.240 ;
      LAYER met4 ;
        RECT 3444.505 2998.310 3588.000 3006.640 ;
      LAYER met4 ;
        RECT 3444.405 2816.390 3444.735 2997.910 ;
      LAYER met4 ;
        RECT 3445.135 2966.670 3588.000 2998.310 ;
        RECT 3445.135 2966.030 3445.835 2966.670 ;
        RECT 3445.135 2819.000 3445.835 2965.000 ;
        RECT 3445.135 2817.330 3445.835 2818.035 ;
      LAYER met4 ;
        RECT 3446.235 2817.730 3450.685 2966.270 ;
      LAYER met4 ;
        RECT 3451.085 2966.030 3451.685 2966.670 ;
        RECT 3451.085 2819.000 3451.685 2965.000 ;
        RECT 3451.085 2817.330 3451.685 2818.035 ;
      LAYER met4 ;
        RECT 3452.085 2817.730 3456.535 2966.270 ;
      LAYER met4 ;
        RECT 3456.935 2966.030 3457.635 2966.670 ;
        RECT 3456.935 2819.000 3457.635 2965.000 ;
        RECT 3456.935 2817.330 3457.635 2818.035 ;
      LAYER met4 ;
        RECT 3458.035 2817.730 3483.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.400 2966.030 3563.385 2966.670 ;
      LAYER met4 ;
        RECT 3563.785 2965.000 3588.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.400 2819.000 3588.000 2965.000 ;
        RECT 3483.400 2817.330 3563.385 2818.035 ;
      LAYER met4 ;
        RECT 3563.785 2817.730 3588.000 2819.000 ;
      LAYER met4 ;
        RECT 3445.135 2815.990 3588.000 2817.330 ;
        RECT 3444.505 2782.160 3588.000 2815.990 ;
        RECT 3439.745 2780.640 3588.000 2782.160 ;
        RECT 3439.745 2766.455 3440.725 2780.640 ;
        RECT 3436.465 2764.935 3440.725 2766.455 ;
        RECT 3390.035 2079.670 3435.965 2151.330 ;
        RECT 198.365 2066.330 199.465 2066.970 ;
        RECT 152.665 2034.690 199.465 2066.330 ;
        RECT 152.035 1991.010 199.465 2034.690 ;
        RECT 147.275 1824.545 151.535 1826.065 ;
        RECT 147.275 1810.360 148.255 1824.545 ;
        RECT 0.000 1808.840 148.255 1810.360 ;
        RECT 0.000 1775.010 143.495 1808.840 ;
        RECT 0.000 1773.670 142.865 1775.010 ;
      LAYER met4 ;
        RECT 0.000 1772.000 24.215 1773.270 ;
      LAYER met4 ;
        RECT 24.615 1772.965 104.600 1773.670 ;
        RECT 0.000 1636.000 104.600 1772.000 ;
      LAYER met4 ;
        RECT 0.000 1634.730 24.215 1636.000 ;
      LAYER met4 ;
        RECT 24.615 1634.330 104.600 1634.970 ;
      LAYER met4 ;
        RECT 105.000 1634.730 129.965 1773.270 ;
      LAYER met4 ;
        RECT 130.365 1772.965 131.065 1773.670 ;
        RECT 130.365 1636.000 131.065 1772.000 ;
        RECT 130.365 1634.330 131.065 1634.970 ;
      LAYER met4 ;
        RECT 131.465 1634.730 135.915 1773.270 ;
      LAYER met4 ;
        RECT 136.315 1772.965 136.915 1773.670 ;
        RECT 136.315 1636.000 136.915 1772.000 ;
        RECT 136.315 1634.330 136.915 1634.970 ;
      LAYER met4 ;
        RECT 137.315 1634.730 141.765 1773.270 ;
      LAYER met4 ;
        RECT 142.165 1772.965 142.865 1773.670 ;
        RECT 142.165 1636.000 142.865 1772.000 ;
        RECT 142.165 1634.330 142.865 1634.970 ;
        RECT 0.000 1602.690 142.865 1634.330 ;
      LAYER met4 ;
        RECT 143.265 1603.090 143.595 1774.610 ;
      LAYER met4 ;
        RECT 0.000 1594.360 143.495 1602.690 ;
      LAYER met4 ;
        RECT 143.895 1594.760 146.875 1808.440 ;
      LAYER met4 ;
        RECT 147.275 1773.670 148.255 1808.840 ;
      LAYER met4 ;
        RECT 147.175 1772.000 148.355 1773.270 ;
      LAYER met4 ;
        RECT 147.175 1636.000 148.355 1772.000 ;
      LAYER met4 ;
        RECT 147.175 1634.730 148.355 1636.000 ;
      LAYER met4 ;
        RECT 147.275 1610.065 148.255 1634.330 ;
      LAYER met4 ;
        RECT 148.655 1610.465 151.635 1824.145 ;
        RECT 151.935 1819.090 152.265 1990.610 ;
      LAYER met4 ;
        RECT 152.665 1989.670 199.465 1991.010 ;
        RECT 152.665 1988.965 153.365 1989.670 ;
        RECT 152.665 1850.330 153.365 1850.970 ;
      LAYER met4 ;
        RECT 153.765 1850.730 158.415 1989.270 ;
      LAYER met4 ;
        RECT 158.815 1988.965 159.415 1989.670 ;
        RECT 158.815 1850.330 159.415 1850.970 ;
      LAYER met4 ;
        RECT 159.815 1850.730 163.265 1989.270 ;
      LAYER met4 ;
        RECT 163.665 1988.965 164.265 1989.670 ;
        RECT 163.665 1850.330 164.265 1850.970 ;
      LAYER met4 ;
        RECT 164.665 1850.730 168.115 1989.270 ;
      LAYER met4 ;
        RECT 168.515 1988.965 169.115 1989.670 ;
        RECT 168.515 1850.330 169.115 1850.970 ;
      LAYER met4 ;
        RECT 169.515 1850.730 174.165 1989.270 ;
      LAYER met4 ;
        RECT 174.565 1988.965 175.165 1989.670 ;
        RECT 180.615 1989.365 186.065 1989.670 ;
        RECT 174.565 1850.330 175.165 1850.970 ;
      LAYER met4 ;
        RECT 175.565 1850.730 180.215 1989.270 ;
      LAYER met4 ;
        RECT 180.615 1988.965 181.215 1989.365 ;
        RECT 185.465 1988.965 186.065 1989.365 ;
      LAYER met4 ;
        RECT 181.615 1850.970 185.065 1988.965 ;
      LAYER met4 ;
        RECT 180.615 1850.570 181.215 1850.970 ;
        RECT 185.465 1850.570 186.065 1850.970 ;
      LAYER met4 ;
        RECT 186.465 1850.730 191.115 1989.270 ;
      LAYER met4 ;
        RECT 191.515 1988.965 192.115 1989.670 ;
        RECT 180.615 1850.330 186.065 1850.570 ;
        RECT 191.515 1850.330 192.115 1850.970 ;
      LAYER met4 ;
        RECT 192.515 1850.730 197.965 1989.270 ;
      LAYER met4 ;
        RECT 198.365 1988.965 199.465 1989.670 ;
        RECT 3388.535 1931.330 3389.635 1932.035 ;
      LAYER met4 ;
        RECT 3390.035 1931.730 3395.485 2079.270 ;
      LAYER met4 ;
        RECT 3395.885 2078.965 3396.485 2079.670 ;
        RECT 3401.935 2079.365 3407.385 2079.670 ;
        RECT 3395.885 1931.330 3396.485 1932.035 ;
      LAYER met4 ;
        RECT 3396.885 1931.730 3401.535 2079.270 ;
      LAYER met4 ;
        RECT 3401.935 2078.965 3402.535 2079.365 ;
        RECT 3406.785 2078.965 3407.385 2079.365 ;
      LAYER met4 ;
        RECT 3402.935 1932.035 3406.385 2078.965 ;
      LAYER met4 ;
        RECT 3401.935 1931.635 3402.535 1932.035 ;
        RECT 3406.785 1931.635 3407.385 1932.035 ;
      LAYER met4 ;
        RECT 3407.785 1931.730 3412.435 2079.270 ;
      LAYER met4 ;
        RECT 3412.835 2078.965 3413.435 2079.670 ;
        RECT 3401.935 1931.330 3407.385 1931.635 ;
        RECT 3412.835 1931.330 3413.435 1932.035 ;
      LAYER met4 ;
        RECT 3413.835 1931.730 3418.485 2079.270 ;
      LAYER met4 ;
        RECT 3418.885 2078.965 3419.485 2079.670 ;
        RECT 3418.885 1931.330 3419.485 1932.035 ;
      LAYER met4 ;
        RECT 3419.885 1931.730 3423.335 2079.270 ;
      LAYER met4 ;
        RECT 3423.735 2078.965 3424.335 2079.670 ;
        RECT 3423.735 1931.330 3424.335 1932.035 ;
      LAYER met4 ;
        RECT 3424.735 1931.730 3428.185 2079.270 ;
      LAYER met4 ;
        RECT 3428.585 2078.965 3429.185 2079.670 ;
        RECT 3428.585 1931.330 3429.185 1932.035 ;
      LAYER met4 ;
        RECT 3429.585 1931.730 3434.235 2079.270 ;
      LAYER met4 ;
        RECT 3434.635 2078.965 3435.335 2079.670 ;
        RECT 3434.635 1931.330 3435.335 1932.035 ;
        RECT 3388.535 1929.990 3435.335 1931.330 ;
      LAYER met4 ;
        RECT 3435.735 1930.390 3436.065 2079.270 ;
      LAYER met4 ;
        RECT 3388.535 1886.310 3435.965 1929.990 ;
        RECT 3388.535 1854.670 3435.335 1886.310 ;
        RECT 3388.535 1854.030 3389.635 1854.670 ;
        RECT 198.365 1850.330 199.465 1850.970 ;
        RECT 152.665 1818.690 199.465 1850.330 ;
        RECT 152.035 1775.010 199.465 1818.690 ;
        RECT 147.275 1608.545 151.535 1610.065 ;
        RECT 147.275 1594.360 148.255 1608.545 ;
        RECT 0.000 1592.840 148.255 1594.360 ;
        RECT 0.000 1559.010 143.495 1592.840 ;
        RECT 0.000 1557.670 142.865 1559.010 ;
      LAYER met4 ;
        RECT 0.000 1556.000 24.215 1557.270 ;
      LAYER met4 ;
        RECT 24.615 1556.965 104.600 1557.670 ;
        RECT 0.000 1420.000 104.600 1556.000 ;
      LAYER met4 ;
        RECT 0.000 1418.730 24.215 1420.000 ;
      LAYER met4 ;
        RECT 24.615 1418.330 104.600 1418.970 ;
      LAYER met4 ;
        RECT 105.000 1418.730 129.965 1557.270 ;
      LAYER met4 ;
        RECT 130.365 1556.965 131.065 1557.670 ;
        RECT 130.365 1420.000 131.065 1556.000 ;
        RECT 130.365 1418.330 131.065 1418.970 ;
      LAYER met4 ;
        RECT 131.465 1418.730 135.915 1557.270 ;
      LAYER met4 ;
        RECT 136.315 1556.965 136.915 1557.670 ;
        RECT 136.315 1420.000 136.915 1556.000 ;
        RECT 136.315 1418.330 136.915 1418.970 ;
      LAYER met4 ;
        RECT 137.315 1418.730 141.765 1557.270 ;
      LAYER met4 ;
        RECT 142.165 1556.965 142.865 1557.670 ;
        RECT 142.165 1420.000 142.865 1556.000 ;
        RECT 142.165 1418.330 142.865 1418.970 ;
        RECT 0.000 1386.690 142.865 1418.330 ;
      LAYER met4 ;
        RECT 143.265 1387.090 143.595 1558.610 ;
      LAYER met4 ;
        RECT 0.000 1378.360 143.495 1386.690 ;
      LAYER met4 ;
        RECT 143.895 1378.760 146.875 1592.440 ;
      LAYER met4 ;
        RECT 147.275 1557.670 148.255 1592.840 ;
      LAYER met4 ;
        RECT 147.175 1556.000 148.355 1557.270 ;
      LAYER met4 ;
        RECT 147.175 1420.000 148.355 1556.000 ;
      LAYER met4 ;
        RECT 147.175 1418.730 148.355 1420.000 ;
      LAYER met4 ;
        RECT 147.275 1394.065 148.255 1418.330 ;
      LAYER met4 ;
        RECT 148.655 1394.465 151.635 1608.145 ;
        RECT 151.935 1603.090 152.265 1774.610 ;
      LAYER met4 ;
        RECT 152.665 1773.670 199.465 1775.010 ;
        RECT 152.665 1772.965 153.365 1773.670 ;
        RECT 152.665 1634.330 153.365 1634.970 ;
      LAYER met4 ;
        RECT 153.765 1634.730 158.415 1773.270 ;
      LAYER met4 ;
        RECT 158.815 1772.965 159.415 1773.670 ;
        RECT 158.815 1634.330 159.415 1634.970 ;
      LAYER met4 ;
        RECT 159.815 1634.730 163.265 1773.270 ;
      LAYER met4 ;
        RECT 163.665 1772.965 164.265 1773.670 ;
        RECT 163.665 1634.330 164.265 1634.970 ;
      LAYER met4 ;
        RECT 164.665 1634.730 168.115 1773.270 ;
      LAYER met4 ;
        RECT 168.515 1772.965 169.115 1773.670 ;
        RECT 168.515 1634.330 169.115 1634.970 ;
      LAYER met4 ;
        RECT 169.515 1634.730 174.165 1773.270 ;
      LAYER met4 ;
        RECT 174.565 1772.965 175.165 1773.670 ;
        RECT 180.615 1773.365 186.065 1773.670 ;
        RECT 174.565 1634.330 175.165 1634.970 ;
      LAYER met4 ;
        RECT 175.565 1634.730 180.215 1773.270 ;
      LAYER met4 ;
        RECT 180.615 1772.965 181.215 1773.365 ;
        RECT 185.465 1772.965 186.065 1773.365 ;
      LAYER met4 ;
        RECT 181.615 1634.970 185.065 1772.965 ;
      LAYER met4 ;
        RECT 180.615 1634.570 181.215 1634.970 ;
        RECT 185.465 1634.570 186.065 1634.970 ;
      LAYER met4 ;
        RECT 186.465 1634.730 191.115 1773.270 ;
      LAYER met4 ;
        RECT 191.515 1772.965 192.115 1773.670 ;
        RECT 180.615 1634.330 186.065 1634.570 ;
        RECT 191.515 1634.330 192.115 1634.970 ;
      LAYER met4 ;
        RECT 192.515 1634.730 197.965 1773.270 ;
      LAYER met4 ;
        RECT 198.365 1772.965 199.465 1773.670 ;
        RECT 3388.535 1705.330 3389.635 1706.035 ;
      LAYER met4 ;
        RECT 3390.035 1705.730 3395.485 1854.270 ;
      LAYER met4 ;
        RECT 3395.885 1854.030 3396.485 1854.670 ;
        RECT 3401.935 1854.430 3407.385 1854.670 ;
        RECT 3395.885 1705.330 3396.485 1706.035 ;
      LAYER met4 ;
        RECT 3396.885 1705.730 3401.535 1854.270 ;
      LAYER met4 ;
        RECT 3401.935 1854.030 3402.535 1854.430 ;
        RECT 3406.785 1854.030 3407.385 1854.430 ;
      LAYER met4 ;
        RECT 3402.935 1706.035 3406.385 1854.030 ;
      LAYER met4 ;
        RECT 3401.935 1705.635 3402.535 1706.035 ;
        RECT 3406.785 1705.635 3407.385 1706.035 ;
      LAYER met4 ;
        RECT 3407.785 1705.730 3412.435 1854.270 ;
      LAYER met4 ;
        RECT 3412.835 1854.030 3413.435 1854.670 ;
        RECT 3401.935 1705.330 3407.385 1705.635 ;
        RECT 3412.835 1705.330 3413.435 1706.035 ;
      LAYER met4 ;
        RECT 3413.835 1705.730 3418.485 1854.270 ;
      LAYER met4 ;
        RECT 3418.885 1854.030 3419.485 1854.670 ;
        RECT 3418.885 1705.330 3419.485 1706.035 ;
      LAYER met4 ;
        RECT 3419.885 1705.730 3423.335 1854.270 ;
      LAYER met4 ;
        RECT 3423.735 1854.030 3424.335 1854.670 ;
        RECT 3423.735 1705.330 3424.335 1706.035 ;
      LAYER met4 ;
        RECT 3424.735 1705.730 3428.185 1854.270 ;
      LAYER met4 ;
        RECT 3428.585 1854.030 3429.185 1854.670 ;
        RECT 3428.585 1705.330 3429.185 1706.035 ;
      LAYER met4 ;
        RECT 3429.585 1705.730 3434.235 1854.270 ;
      LAYER met4 ;
        RECT 3434.635 1854.030 3435.335 1854.670 ;
        RECT 3434.635 1705.330 3435.335 1706.035 ;
        RECT 3388.535 1703.990 3435.335 1705.330 ;
      LAYER met4 ;
        RECT 3435.735 1704.390 3436.065 1885.910 ;
        RECT 3436.365 1880.855 3439.345 2764.535 ;
      LAYER met4 ;
        RECT 3439.745 2740.670 3440.725 2764.935 ;
      LAYER met4 ;
        RECT 3439.645 2739.000 3440.825 2740.270 ;
      LAYER met4 ;
        RECT 3439.645 2594.000 3440.825 2739.000 ;
      LAYER met4 ;
        RECT 3439.645 2592.730 3440.825 2594.000 ;
      LAYER met4 ;
        RECT 3439.745 2520.670 3440.725 2592.330 ;
      LAYER met4 ;
        RECT 3439.645 2519.000 3440.825 2520.270 ;
      LAYER met4 ;
        RECT 3439.645 2374.000 3440.825 2519.000 ;
      LAYER met4 ;
        RECT 3439.645 2372.730 3440.825 2374.000 ;
      LAYER met4 ;
        RECT 3439.745 2300.670 3440.725 2372.330 ;
      LAYER met4 ;
        RECT 3439.645 2299.000 3440.825 2300.270 ;
      LAYER met4 ;
        RECT 3439.645 2153.000 3440.825 2299.000 ;
      LAYER met4 ;
        RECT 3439.645 2151.730 3440.825 2153.000 ;
      LAYER met4 ;
        RECT 3439.745 2079.670 3440.725 2151.330 ;
      LAYER met4 ;
        RECT 3439.645 2078.000 3440.825 2079.270 ;
      LAYER met4 ;
        RECT 3439.645 1933.000 3440.825 2078.000 ;
      LAYER met4 ;
        RECT 3439.645 1931.730 3440.825 1933.000 ;
      LAYER met4 ;
        RECT 3439.745 1896.160 3440.725 1931.330 ;
      LAYER met4 ;
        RECT 3441.125 1896.560 3444.105 2780.240 ;
      LAYER met4 ;
        RECT 3444.505 2772.310 3588.000 2780.640 ;
        RECT 3445.135 2740.670 3588.000 2772.310 ;
        RECT 3445.135 2740.030 3445.835 2740.670 ;
        RECT 3445.135 2594.000 3445.835 2739.000 ;
        RECT 3445.135 2592.330 3445.835 2593.035 ;
      LAYER met4 ;
        RECT 3446.235 2592.730 3450.685 2740.270 ;
      LAYER met4 ;
        RECT 3451.085 2740.030 3451.685 2740.670 ;
        RECT 3451.085 2594.000 3451.685 2739.000 ;
        RECT 3451.085 2592.330 3451.685 2593.035 ;
      LAYER met4 ;
        RECT 3452.085 2592.730 3456.535 2740.270 ;
      LAYER met4 ;
        RECT 3456.935 2740.030 3457.635 2740.670 ;
        RECT 3456.935 2594.000 3457.635 2739.000 ;
        RECT 3456.935 2592.330 3457.635 2593.035 ;
      LAYER met4 ;
        RECT 3458.035 2592.730 3483.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.400 2740.030 3563.385 2740.670 ;
      LAYER met4 ;
        RECT 3563.785 2739.000 3588.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.400 2594.000 3588.000 2739.000 ;
        RECT 3483.400 2592.330 3563.385 2593.035 ;
      LAYER met4 ;
        RECT 3563.785 2592.730 3588.000 2594.000 ;
      LAYER met4 ;
        RECT 3445.135 2520.670 3588.000 2592.330 ;
        RECT 3445.135 2519.965 3445.835 2520.670 ;
        RECT 3445.135 2372.330 3445.835 2519.000 ;
      LAYER met4 ;
        RECT 3446.235 2372.730 3450.685 2520.270 ;
      LAYER met4 ;
        RECT 3451.085 2519.965 3451.685 2520.670 ;
        RECT 3451.085 2372.330 3451.685 2519.000 ;
      LAYER met4 ;
        RECT 3452.085 2372.730 3456.535 2520.270 ;
      LAYER met4 ;
        RECT 3456.935 2519.965 3457.635 2520.670 ;
        RECT 3456.935 2372.330 3457.635 2519.000 ;
      LAYER met4 ;
        RECT 3458.035 2372.730 3483.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.400 2519.965 3563.385 2520.670 ;
      LAYER met4 ;
        RECT 3563.785 2519.000 3588.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.400 2374.000 3588.000 2519.000 ;
        RECT 3483.400 2372.330 3563.385 2374.000 ;
      LAYER met4 ;
        RECT 3563.785 2372.730 3588.000 2374.000 ;
      LAYER met4 ;
        RECT 3445.135 2300.670 3588.000 2372.330 ;
        RECT 3445.135 2153.000 3445.835 2300.670 ;
        RECT 3445.135 2151.330 3445.835 2152.035 ;
      LAYER met4 ;
        RECT 3446.235 2151.730 3450.685 2300.270 ;
      LAYER met4 ;
        RECT 3451.085 2153.000 3451.685 2300.670 ;
        RECT 3451.085 2151.330 3451.685 2152.035 ;
      LAYER met4 ;
        RECT 3452.085 2151.730 3456.535 2300.270 ;
      LAYER met4 ;
        RECT 3456.935 2153.000 3457.635 2300.670 ;
        RECT 3456.935 2151.330 3457.635 2152.035 ;
      LAYER met4 ;
        RECT 3458.035 2151.730 3483.000 2300.270 ;
      LAYER met4 ;
        RECT 3483.400 2299.000 3563.385 2300.670 ;
        RECT 3563.750 2299.000 3563.785 2299.215 ;
      LAYER met4 ;
        RECT 3563.785 2299.000 3588.000 2300.270 ;
      LAYER met4 ;
        RECT 3483.400 2153.000 3588.000 2299.000 ;
        RECT 3483.400 2151.330 3563.385 2152.035 ;
      LAYER met4 ;
        RECT 3563.785 2151.730 3588.000 2153.000 ;
      LAYER met4 ;
        RECT 3444.505 2079.670 3588.000 2151.330 ;
      LAYER met4 ;
        RECT 3444.405 1930.390 3444.735 2079.270 ;
      LAYER met4 ;
        RECT 3445.135 2078.965 3445.835 2079.670 ;
        RECT 3445.135 1933.000 3445.835 2078.000 ;
        RECT 3445.135 1931.330 3445.835 1932.035 ;
      LAYER met4 ;
        RECT 3446.235 1931.730 3450.685 2079.270 ;
      LAYER met4 ;
        RECT 3451.085 2078.965 3451.685 2079.670 ;
        RECT 3451.085 1933.000 3451.685 2078.000 ;
        RECT 3451.085 1931.330 3451.685 1932.035 ;
      LAYER met4 ;
        RECT 3452.085 1931.730 3456.535 2079.270 ;
      LAYER met4 ;
        RECT 3456.935 2078.965 3457.635 2079.670 ;
        RECT 3456.935 1933.000 3457.635 2078.000 ;
        RECT 3456.935 1931.330 3457.635 1932.035 ;
      LAYER met4 ;
        RECT 3458.035 1931.730 3483.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.400 2078.965 3563.385 2079.670 ;
      LAYER met4 ;
        RECT 3563.785 2078.000 3588.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.400 1933.000 3588.000 2078.000 ;
        RECT 3483.400 1931.330 3563.385 1932.035 ;
      LAYER met4 ;
        RECT 3563.785 1931.730 3588.000 1933.000 ;
      LAYER met4 ;
        RECT 3445.135 1929.990 3588.000 1931.330 ;
        RECT 3444.505 1896.160 3588.000 1929.990 ;
        RECT 3439.745 1894.640 3588.000 1896.160 ;
        RECT 3439.745 1880.455 3440.725 1894.640 ;
        RECT 3436.465 1878.935 3440.725 1880.455 ;
        RECT 3388.535 1660.310 3435.965 1703.990 ;
        RECT 198.365 1634.330 199.465 1634.970 ;
        RECT 152.665 1602.690 199.465 1634.330 ;
        RECT 3388.535 1628.670 3435.335 1660.310 ;
        RECT 3388.535 1628.030 3389.635 1628.670 ;
        RECT 152.035 1559.010 199.465 1602.690 ;
        RECT 147.275 1392.545 151.535 1394.065 ;
        RECT 147.275 1378.360 148.255 1392.545 ;
        RECT 0.000 1376.840 148.255 1378.360 ;
        RECT 0.000 1343.010 143.495 1376.840 ;
        RECT 0.000 1341.670 142.865 1343.010 ;
      LAYER met4 ;
        RECT 0.000 1340.000 24.215 1341.270 ;
      LAYER met4 ;
        RECT 24.615 1340.965 104.600 1341.670 ;
        RECT 0.000 1204.000 104.600 1340.000 ;
      LAYER met4 ;
        RECT 0.000 1202.730 24.215 1204.000 ;
      LAYER met4 ;
        RECT 24.615 1202.330 104.600 1202.970 ;
      LAYER met4 ;
        RECT 105.000 1202.730 129.965 1341.270 ;
      LAYER met4 ;
        RECT 130.365 1340.965 131.065 1341.670 ;
        RECT 130.365 1204.000 131.065 1340.000 ;
        RECT 130.365 1202.330 131.065 1202.970 ;
      LAYER met4 ;
        RECT 131.465 1202.730 135.915 1341.270 ;
      LAYER met4 ;
        RECT 136.315 1340.965 136.915 1341.670 ;
        RECT 136.315 1204.000 136.915 1340.000 ;
        RECT 136.315 1202.330 136.915 1202.970 ;
      LAYER met4 ;
        RECT 137.315 1202.730 141.765 1341.270 ;
      LAYER met4 ;
        RECT 142.165 1340.965 142.865 1341.670 ;
        RECT 142.165 1204.000 142.865 1340.000 ;
        RECT 142.165 1202.330 142.865 1202.970 ;
        RECT 0.000 1170.690 142.865 1202.330 ;
      LAYER met4 ;
        RECT 143.265 1171.090 143.595 1342.610 ;
      LAYER met4 ;
        RECT 0.000 1162.360 143.495 1170.690 ;
      LAYER met4 ;
        RECT 143.895 1162.760 146.875 1376.440 ;
      LAYER met4 ;
        RECT 147.275 1341.670 148.255 1376.840 ;
      LAYER met4 ;
        RECT 147.175 1340.000 148.355 1341.270 ;
      LAYER met4 ;
        RECT 147.175 1204.000 148.355 1340.000 ;
      LAYER met4 ;
        RECT 147.175 1202.730 148.355 1204.000 ;
      LAYER met4 ;
        RECT 147.275 1178.065 148.255 1202.330 ;
      LAYER met4 ;
        RECT 148.655 1178.465 151.635 1392.145 ;
        RECT 151.935 1387.090 152.265 1558.610 ;
      LAYER met4 ;
        RECT 152.665 1557.670 199.465 1559.010 ;
        RECT 152.665 1556.965 153.365 1557.670 ;
        RECT 152.665 1418.330 153.365 1418.970 ;
      LAYER met4 ;
        RECT 153.765 1418.730 158.415 1557.270 ;
      LAYER met4 ;
        RECT 158.815 1556.965 159.415 1557.670 ;
        RECT 158.815 1418.330 159.415 1418.970 ;
      LAYER met4 ;
        RECT 159.815 1418.730 163.265 1557.270 ;
      LAYER met4 ;
        RECT 163.665 1556.965 164.265 1557.670 ;
        RECT 163.665 1418.330 164.265 1418.970 ;
      LAYER met4 ;
        RECT 164.665 1418.730 168.115 1557.270 ;
      LAYER met4 ;
        RECT 168.515 1556.965 169.115 1557.670 ;
        RECT 168.515 1418.330 169.115 1418.970 ;
      LAYER met4 ;
        RECT 169.515 1418.730 174.165 1557.270 ;
      LAYER met4 ;
        RECT 174.565 1556.965 175.165 1557.670 ;
        RECT 180.615 1557.365 186.065 1557.670 ;
        RECT 174.565 1418.330 175.165 1418.970 ;
      LAYER met4 ;
        RECT 175.565 1418.730 180.215 1557.270 ;
      LAYER met4 ;
        RECT 180.615 1556.965 181.215 1557.365 ;
        RECT 185.465 1556.965 186.065 1557.365 ;
      LAYER met4 ;
        RECT 181.615 1418.970 185.065 1556.965 ;
      LAYER met4 ;
        RECT 180.615 1418.570 181.215 1418.970 ;
        RECT 185.465 1418.570 186.065 1418.970 ;
      LAYER met4 ;
        RECT 186.465 1418.730 191.115 1557.270 ;
      LAYER met4 ;
        RECT 191.515 1556.965 192.115 1557.670 ;
        RECT 180.615 1418.330 186.065 1418.570 ;
        RECT 191.515 1418.330 192.115 1418.970 ;
      LAYER met4 ;
        RECT 192.515 1418.730 197.965 1557.270 ;
      LAYER met4 ;
        RECT 198.365 1556.965 199.465 1557.670 ;
        RECT 3388.535 1480.330 3389.635 1481.035 ;
      LAYER met4 ;
        RECT 3390.035 1480.730 3395.485 1628.270 ;
      LAYER met4 ;
        RECT 3395.885 1628.030 3396.485 1628.670 ;
        RECT 3401.935 1628.430 3407.385 1628.670 ;
        RECT 3395.885 1480.330 3396.485 1481.035 ;
      LAYER met4 ;
        RECT 3396.885 1480.730 3401.535 1628.270 ;
      LAYER met4 ;
        RECT 3401.935 1628.030 3402.535 1628.430 ;
        RECT 3406.785 1628.030 3407.385 1628.430 ;
      LAYER met4 ;
        RECT 3402.935 1481.035 3406.385 1628.030 ;
      LAYER met4 ;
        RECT 3401.935 1480.635 3402.535 1481.035 ;
        RECT 3406.785 1480.635 3407.385 1481.035 ;
      LAYER met4 ;
        RECT 3407.785 1480.730 3412.435 1628.270 ;
      LAYER met4 ;
        RECT 3412.835 1628.030 3413.435 1628.670 ;
        RECT 3401.935 1480.330 3407.385 1480.635 ;
        RECT 3412.835 1480.330 3413.435 1481.035 ;
      LAYER met4 ;
        RECT 3413.835 1480.730 3418.485 1628.270 ;
      LAYER met4 ;
        RECT 3418.885 1628.030 3419.485 1628.670 ;
        RECT 3418.885 1480.330 3419.485 1481.035 ;
      LAYER met4 ;
        RECT 3419.885 1480.730 3423.335 1628.270 ;
      LAYER met4 ;
        RECT 3423.735 1628.030 3424.335 1628.670 ;
        RECT 3423.735 1480.330 3424.335 1481.035 ;
      LAYER met4 ;
        RECT 3424.735 1480.730 3428.185 1628.270 ;
      LAYER met4 ;
        RECT 3428.585 1628.030 3429.185 1628.670 ;
        RECT 3428.585 1480.330 3429.185 1481.035 ;
      LAYER met4 ;
        RECT 3429.585 1480.730 3434.235 1628.270 ;
      LAYER met4 ;
        RECT 3434.635 1628.030 3435.335 1628.670 ;
        RECT 3434.635 1480.330 3435.335 1481.035 ;
        RECT 3388.535 1478.990 3435.335 1480.330 ;
      LAYER met4 ;
        RECT 3435.735 1479.390 3436.065 1659.910 ;
        RECT 3436.365 1654.855 3439.345 1878.535 ;
      LAYER met4 ;
        RECT 3439.745 1854.670 3440.725 1878.935 ;
      LAYER met4 ;
        RECT 3439.645 1853.000 3440.825 1854.270 ;
      LAYER met4 ;
        RECT 3439.645 1707.000 3440.825 1853.000 ;
      LAYER met4 ;
        RECT 3439.645 1705.730 3440.825 1707.000 ;
      LAYER met4 ;
        RECT 3439.745 1670.160 3440.725 1705.330 ;
      LAYER met4 ;
        RECT 3441.125 1670.560 3444.105 1894.240 ;
      LAYER met4 ;
        RECT 3444.505 1886.310 3588.000 1894.640 ;
      LAYER met4 ;
        RECT 3444.405 1704.390 3444.735 1885.910 ;
      LAYER met4 ;
        RECT 3445.135 1854.670 3588.000 1886.310 ;
        RECT 3445.135 1854.030 3445.835 1854.670 ;
        RECT 3445.135 1707.000 3445.835 1853.000 ;
        RECT 3445.135 1705.330 3445.835 1706.035 ;
      LAYER met4 ;
        RECT 3446.235 1705.730 3450.685 1854.270 ;
      LAYER met4 ;
        RECT 3451.085 1854.030 3451.685 1854.670 ;
        RECT 3451.085 1707.000 3451.685 1853.000 ;
        RECT 3451.085 1705.330 3451.685 1706.035 ;
      LAYER met4 ;
        RECT 3452.085 1705.730 3456.535 1854.270 ;
      LAYER met4 ;
        RECT 3456.935 1854.030 3457.635 1854.670 ;
        RECT 3456.935 1707.000 3457.635 1853.000 ;
        RECT 3456.935 1705.330 3457.635 1706.035 ;
      LAYER met4 ;
        RECT 3458.035 1705.730 3483.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.400 1854.030 3563.385 1854.670 ;
      LAYER met4 ;
        RECT 3563.785 1853.000 3588.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.400 1707.000 3588.000 1853.000 ;
        RECT 3483.400 1705.330 3563.385 1706.035 ;
      LAYER met4 ;
        RECT 3563.785 1705.730 3588.000 1707.000 ;
      LAYER met4 ;
        RECT 3445.135 1703.990 3588.000 1705.330 ;
        RECT 3444.505 1670.160 3588.000 1703.990 ;
        RECT 3439.745 1668.640 3588.000 1670.160 ;
        RECT 3439.745 1654.455 3440.725 1668.640 ;
        RECT 3436.465 1652.935 3440.725 1654.455 ;
        RECT 3388.535 1435.310 3435.965 1478.990 ;
        RECT 198.365 1418.330 199.465 1418.970 ;
        RECT 152.665 1386.690 199.465 1418.330 ;
        RECT 3388.535 1403.670 3435.335 1435.310 ;
        RECT 3388.535 1403.030 3389.635 1403.670 ;
        RECT 152.035 1343.010 199.465 1386.690 ;
        RECT 147.275 1176.545 151.535 1178.065 ;
        RECT 147.275 1162.360 148.255 1176.545 ;
        RECT 0.000 1160.840 148.255 1162.360 ;
        RECT 0.000 1127.010 143.495 1160.840 ;
        RECT 0.000 1125.670 142.865 1127.010 ;
      LAYER met4 ;
        RECT 0.000 1124.000 24.215 1125.270 ;
      LAYER met4 ;
        RECT 24.615 1124.965 104.600 1125.670 ;
        RECT 0.000 988.000 104.600 1124.000 ;
      LAYER met4 ;
        RECT 0.000 986.730 24.215 988.000 ;
      LAYER met4 ;
        RECT 24.615 986.330 104.600 986.970 ;
      LAYER met4 ;
        RECT 105.000 986.730 129.965 1125.270 ;
      LAYER met4 ;
        RECT 130.365 1124.965 131.065 1125.670 ;
        RECT 130.365 988.000 131.065 1124.000 ;
        RECT 130.365 986.330 131.065 986.970 ;
      LAYER met4 ;
        RECT 131.465 986.730 135.915 1125.270 ;
      LAYER met4 ;
        RECT 136.315 1124.965 136.915 1125.670 ;
        RECT 136.315 988.000 136.915 1124.000 ;
        RECT 136.315 986.330 136.915 986.970 ;
      LAYER met4 ;
        RECT 137.315 986.730 141.765 1125.270 ;
      LAYER met4 ;
        RECT 142.165 1124.965 142.865 1125.670 ;
        RECT 142.165 988.000 142.865 1124.000 ;
        RECT 142.165 986.330 142.865 986.970 ;
        RECT 0.000 954.690 142.865 986.330 ;
      LAYER met4 ;
        RECT 143.265 955.090 143.595 1126.610 ;
      LAYER met4 ;
        RECT 0.000 946.360 143.495 954.690 ;
      LAYER met4 ;
        RECT 143.895 946.760 146.875 1160.440 ;
      LAYER met4 ;
        RECT 147.275 1125.670 148.255 1160.840 ;
      LAYER met4 ;
        RECT 147.175 1124.000 148.355 1125.270 ;
      LAYER met4 ;
        RECT 147.175 988.000 148.355 1124.000 ;
      LAYER met4 ;
        RECT 147.175 986.730 148.355 988.000 ;
      LAYER met4 ;
        RECT 147.275 962.065 148.255 986.330 ;
      LAYER met4 ;
        RECT 148.655 962.465 151.635 1176.145 ;
        RECT 151.935 1171.090 152.265 1342.610 ;
      LAYER met4 ;
        RECT 152.665 1341.670 199.465 1343.010 ;
        RECT 152.665 1340.965 153.365 1341.670 ;
        RECT 152.665 1202.330 153.365 1202.970 ;
      LAYER met4 ;
        RECT 153.765 1202.730 158.415 1341.270 ;
      LAYER met4 ;
        RECT 158.815 1340.965 159.415 1341.670 ;
        RECT 158.815 1202.330 159.415 1202.970 ;
      LAYER met4 ;
        RECT 159.815 1202.730 163.265 1341.270 ;
      LAYER met4 ;
        RECT 163.665 1340.965 164.265 1341.670 ;
        RECT 163.665 1202.330 164.265 1202.970 ;
      LAYER met4 ;
        RECT 164.665 1202.730 168.115 1341.270 ;
      LAYER met4 ;
        RECT 168.515 1340.965 169.115 1341.670 ;
        RECT 168.515 1202.330 169.115 1202.970 ;
      LAYER met4 ;
        RECT 169.515 1202.730 174.165 1341.270 ;
      LAYER met4 ;
        RECT 174.565 1340.965 175.165 1341.670 ;
        RECT 180.615 1341.365 186.065 1341.670 ;
        RECT 174.565 1202.330 175.165 1202.970 ;
      LAYER met4 ;
        RECT 175.565 1202.730 180.215 1341.270 ;
      LAYER met4 ;
        RECT 180.615 1340.965 181.215 1341.365 ;
        RECT 185.465 1340.965 186.065 1341.365 ;
      LAYER met4 ;
        RECT 181.615 1202.970 185.065 1340.965 ;
      LAYER met4 ;
        RECT 180.615 1202.570 181.215 1202.970 ;
        RECT 185.465 1202.570 186.065 1202.970 ;
      LAYER met4 ;
        RECT 186.465 1202.730 191.115 1341.270 ;
      LAYER met4 ;
        RECT 191.515 1340.965 192.115 1341.670 ;
        RECT 180.615 1202.330 186.065 1202.570 ;
        RECT 191.515 1202.330 192.115 1202.970 ;
      LAYER met4 ;
        RECT 192.515 1202.730 197.965 1341.270 ;
      LAYER met4 ;
        RECT 198.365 1340.965 199.465 1341.670 ;
        RECT 3388.535 1255.330 3389.635 1256.035 ;
      LAYER met4 ;
        RECT 3390.035 1255.730 3395.485 1403.270 ;
      LAYER met4 ;
        RECT 3395.885 1403.030 3396.485 1403.670 ;
        RECT 3401.935 1403.430 3407.385 1403.670 ;
        RECT 3395.885 1255.330 3396.485 1256.035 ;
      LAYER met4 ;
        RECT 3396.885 1255.730 3401.535 1403.270 ;
      LAYER met4 ;
        RECT 3401.935 1403.030 3402.535 1403.430 ;
        RECT 3406.785 1403.030 3407.385 1403.430 ;
      LAYER met4 ;
        RECT 3402.935 1256.035 3406.385 1403.030 ;
      LAYER met4 ;
        RECT 3401.935 1255.635 3402.535 1256.035 ;
        RECT 3406.785 1255.635 3407.385 1256.035 ;
      LAYER met4 ;
        RECT 3407.785 1255.730 3412.435 1403.270 ;
      LAYER met4 ;
        RECT 3412.835 1403.030 3413.435 1403.670 ;
        RECT 3401.935 1255.330 3407.385 1255.635 ;
        RECT 3412.835 1255.330 3413.435 1256.035 ;
      LAYER met4 ;
        RECT 3413.835 1255.730 3418.485 1403.270 ;
      LAYER met4 ;
        RECT 3418.885 1403.030 3419.485 1403.670 ;
        RECT 3418.885 1255.330 3419.485 1256.035 ;
      LAYER met4 ;
        RECT 3419.885 1255.730 3423.335 1403.270 ;
      LAYER met4 ;
        RECT 3423.735 1403.030 3424.335 1403.670 ;
        RECT 3423.735 1255.330 3424.335 1256.035 ;
      LAYER met4 ;
        RECT 3424.735 1255.730 3428.185 1403.270 ;
      LAYER met4 ;
        RECT 3428.585 1403.030 3429.185 1403.670 ;
        RECT 3428.585 1255.330 3429.185 1256.035 ;
      LAYER met4 ;
        RECT 3429.585 1255.730 3434.235 1403.270 ;
      LAYER met4 ;
        RECT 3434.635 1403.030 3435.335 1403.670 ;
        RECT 3434.635 1255.330 3435.335 1256.035 ;
        RECT 3388.535 1253.990 3435.335 1255.330 ;
      LAYER met4 ;
        RECT 3435.735 1254.390 3436.065 1434.910 ;
        RECT 3436.365 1429.855 3439.345 1652.535 ;
      LAYER met4 ;
        RECT 3439.745 1628.670 3440.725 1652.935 ;
      LAYER met4 ;
        RECT 3439.645 1627.000 3440.825 1628.270 ;
      LAYER met4 ;
        RECT 3439.645 1482.000 3440.825 1627.000 ;
      LAYER met4 ;
        RECT 3439.645 1480.730 3440.825 1482.000 ;
      LAYER met4 ;
        RECT 3439.745 1445.160 3440.725 1480.330 ;
      LAYER met4 ;
        RECT 3441.125 1445.560 3444.105 1668.240 ;
      LAYER met4 ;
        RECT 3444.505 1660.310 3588.000 1668.640 ;
      LAYER met4 ;
        RECT 3444.405 1479.390 3444.735 1659.910 ;
      LAYER met4 ;
        RECT 3445.135 1628.670 3588.000 1660.310 ;
        RECT 3445.135 1628.030 3445.835 1628.670 ;
        RECT 3445.135 1482.000 3445.835 1627.000 ;
        RECT 3445.135 1480.330 3445.835 1481.035 ;
      LAYER met4 ;
        RECT 3446.235 1480.730 3450.685 1628.270 ;
      LAYER met4 ;
        RECT 3451.085 1628.030 3451.685 1628.670 ;
        RECT 3451.085 1482.000 3451.685 1627.000 ;
        RECT 3451.085 1480.330 3451.685 1481.035 ;
      LAYER met4 ;
        RECT 3452.085 1480.730 3456.535 1628.270 ;
      LAYER met4 ;
        RECT 3456.935 1628.030 3457.635 1628.670 ;
        RECT 3456.935 1482.000 3457.635 1627.000 ;
        RECT 3456.935 1480.330 3457.635 1481.035 ;
      LAYER met4 ;
        RECT 3458.035 1480.730 3483.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.400 1628.030 3563.385 1628.670 ;
      LAYER met4 ;
        RECT 3563.785 1627.000 3588.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.400 1482.000 3588.000 1627.000 ;
        RECT 3483.400 1480.330 3563.385 1481.035 ;
      LAYER met4 ;
        RECT 3563.785 1480.730 3588.000 1482.000 ;
      LAYER met4 ;
        RECT 3445.135 1478.990 3588.000 1480.330 ;
        RECT 3444.505 1445.160 3588.000 1478.990 ;
        RECT 3439.745 1443.640 3588.000 1445.160 ;
        RECT 3439.745 1429.455 3440.725 1443.640 ;
        RECT 3436.465 1427.935 3440.725 1429.455 ;
        RECT 3388.535 1210.310 3435.965 1253.990 ;
        RECT 198.365 1202.330 199.465 1202.970 ;
        RECT 152.665 1170.690 199.465 1202.330 ;
        RECT 3388.535 1178.670 3435.335 1210.310 ;
        RECT 3388.535 1178.030 3389.635 1178.670 ;
        RECT 152.035 1127.010 199.465 1170.690 ;
        RECT 147.275 960.545 151.535 962.065 ;
        RECT 147.275 946.360 148.255 960.545 ;
        RECT 0.000 944.840 148.255 946.360 ;
        RECT 0.000 911.010 143.495 944.840 ;
        RECT 0.000 909.670 142.865 911.010 ;
      LAYER met4 ;
        RECT 0.000 908.000 24.215 909.270 ;
      LAYER met4 ;
        RECT 24.615 908.965 104.600 909.670 ;
        RECT 0.000 631.000 104.600 908.000 ;
        RECT 0.000 626.000 24.215 631.000 ;
      LAYER met4 ;
        RECT 0.000 624.730 24.215 626.000 ;
      LAYER met4 ;
        RECT 24.615 624.330 104.600 625.035 ;
      LAYER met4 ;
        RECT 105.000 624.730 129.965 909.270 ;
      LAYER met4 ;
        RECT 130.365 908.965 131.065 909.670 ;
        RECT 130.365 631.000 131.065 908.000 ;
        RECT 130.365 624.330 131.065 625.035 ;
      LAYER met4 ;
        RECT 131.465 624.730 135.915 909.270 ;
      LAYER met4 ;
        RECT 136.315 908.965 136.915 909.670 ;
        RECT 136.315 631.000 136.915 908.000 ;
        RECT 136.315 624.330 136.915 625.035 ;
      LAYER met4 ;
        RECT 137.315 624.730 141.765 909.270 ;
      LAYER met4 ;
        RECT 142.165 908.965 142.865 909.670 ;
        RECT 142.165 631.000 142.865 908.000 ;
      LAYER met4 ;
        RECT 143.265 631.000 143.595 910.610 ;
      LAYER met4 ;
        RECT 142.165 624.330 142.865 625.035 ;
        RECT 0.000 552.670 142.865 624.330 ;
      LAYER met4 ;
        RECT 0.000 551.000 24.215 552.270 ;
      LAYER met4 ;
        RECT 24.615 551.965 104.600 552.670 ;
        RECT 0.000 415.000 104.600 551.000 ;
      LAYER met4 ;
        RECT 0.000 413.730 24.215 415.000 ;
      LAYER met4 ;
        RECT 24.615 413.330 104.600 415.000 ;
      LAYER met4 ;
        RECT 105.000 413.730 129.965 552.270 ;
      LAYER met4 ;
        RECT 130.365 551.965 131.065 552.670 ;
        RECT 130.365 413.330 131.065 551.000 ;
      LAYER met4 ;
        RECT 131.465 413.730 135.915 552.270 ;
      LAYER met4 ;
        RECT 136.315 551.965 136.915 552.670 ;
        RECT 136.315 413.330 136.915 551.000 ;
      LAYER met4 ;
        RECT 137.315 413.730 141.765 552.270 ;
      LAYER met4 ;
        RECT 142.165 551.965 142.865 552.670 ;
        RECT 142.165 413.330 142.865 551.000 ;
        RECT 0.000 341.670 142.865 413.330 ;
      LAYER met4 ;
        RECT 0.000 340.000 24.215 341.270 ;
      LAYER met4 ;
        RECT 24.615 340.965 104.600 341.670 ;
        RECT 0.000 204.000 104.600 340.000 ;
      LAYER met4 ;
        RECT 0.000 202.730 24.215 204.000 ;
      LAYER met4 ;
        RECT 24.615 202.330 104.600 202.745 ;
        RECT 0.000 201.745 104.600 202.330 ;
      LAYER met4 ;
        RECT 105.000 202.145 129.965 341.270 ;
      LAYER met4 ;
        RECT 130.365 340.965 131.065 341.670 ;
        RECT 130.365 204.000 131.065 340.000 ;
        RECT 130.365 202.330 131.065 202.745 ;
      LAYER met4 ;
        RECT 131.465 202.730 135.915 341.270 ;
      LAYER met4 ;
        RECT 136.315 340.965 136.915 341.670 ;
        RECT 136.315 204.000 136.915 340.000 ;
        RECT 136.315 202.330 136.915 202.745 ;
      LAYER met4 ;
        RECT 137.315 202.730 141.765 341.270 ;
      LAYER met4 ;
        RECT 142.165 340.965 142.865 341.670 ;
        RECT 142.165 204.000 142.865 340.000 ;
        RECT 142.165 202.330 142.865 202.745 ;
        RECT 130.365 201.745 142.865 202.330 ;
        RECT 0.000 176.425 142.865 201.745 ;
      LAYER met4 ;
        RECT 143.265 176.825 143.595 626.000 ;
        RECT 143.895 177.090 146.875 944.440 ;
      LAYER met4 ;
        RECT 147.275 909.670 148.255 944.840 ;
      LAYER met4 ;
        RECT 147.175 908.000 148.355 909.270 ;
      LAYER met4 ;
        RECT 147.175 631.000 148.355 908.000 ;
      LAYER met4 ;
        RECT 147.175 624.730 148.355 626.000 ;
      LAYER met4 ;
        RECT 147.275 552.670 148.255 624.330 ;
      LAYER met4 ;
        RECT 147.175 551.000 148.355 552.270 ;
      LAYER met4 ;
        RECT 147.175 415.000 148.355 551.000 ;
      LAYER met4 ;
        RECT 147.175 413.730 148.355 415.000 ;
      LAYER met4 ;
        RECT 147.275 341.670 148.255 413.330 ;
      LAYER met4 ;
        RECT 147.175 340.000 148.355 341.270 ;
      LAYER met4 ;
        RECT 147.175 204.000 148.355 340.000 ;
      LAYER met4 ;
        RECT 147.175 182.445 148.355 204.000 ;
        RECT 148.655 183.125 151.635 960.145 ;
        RECT 151.935 955.090 152.265 1126.610 ;
      LAYER met4 ;
        RECT 152.665 1125.670 199.465 1127.010 ;
        RECT 152.665 1124.965 153.365 1125.670 ;
        RECT 152.665 986.330 153.365 986.970 ;
      LAYER met4 ;
        RECT 153.765 986.730 158.415 1125.270 ;
      LAYER met4 ;
        RECT 158.815 1124.965 159.415 1125.670 ;
        RECT 158.815 986.330 159.415 986.970 ;
      LAYER met4 ;
        RECT 159.815 986.730 163.265 1125.270 ;
      LAYER met4 ;
        RECT 163.665 1124.965 164.265 1125.670 ;
        RECT 163.665 986.330 164.265 986.970 ;
      LAYER met4 ;
        RECT 164.665 986.730 168.115 1125.270 ;
      LAYER met4 ;
        RECT 168.515 1124.965 169.115 1125.670 ;
        RECT 168.515 986.330 169.115 986.970 ;
      LAYER met4 ;
        RECT 169.515 986.730 174.165 1125.270 ;
      LAYER met4 ;
        RECT 174.565 1124.965 175.165 1125.670 ;
        RECT 180.615 1125.365 186.065 1125.670 ;
        RECT 174.565 986.330 175.165 986.970 ;
      LAYER met4 ;
        RECT 175.565 986.730 180.215 1125.270 ;
      LAYER met4 ;
        RECT 180.615 1124.965 181.215 1125.365 ;
        RECT 185.465 1124.965 186.065 1125.365 ;
      LAYER met4 ;
        RECT 181.615 986.970 185.065 1124.965 ;
      LAYER met4 ;
        RECT 180.615 986.570 181.215 986.970 ;
        RECT 185.465 986.570 186.065 986.970 ;
      LAYER met4 ;
        RECT 186.465 986.730 191.115 1125.270 ;
      LAYER met4 ;
        RECT 191.515 1124.965 192.115 1125.670 ;
        RECT 180.615 986.330 186.065 986.570 ;
        RECT 191.515 986.330 192.115 986.970 ;
      LAYER met4 ;
        RECT 192.515 986.730 197.965 1125.270 ;
      LAYER met4 ;
        RECT 198.365 1124.965 199.465 1125.670 ;
        RECT 3388.535 1029.330 3389.635 1030.035 ;
      LAYER met4 ;
        RECT 3390.035 1029.730 3395.485 1178.270 ;
      LAYER met4 ;
        RECT 3395.885 1178.030 3396.485 1178.670 ;
        RECT 3401.935 1178.430 3407.385 1178.670 ;
        RECT 3395.885 1029.330 3396.485 1030.035 ;
      LAYER met4 ;
        RECT 3396.885 1029.730 3401.535 1178.270 ;
      LAYER met4 ;
        RECT 3401.935 1178.030 3402.535 1178.430 ;
        RECT 3406.785 1178.030 3407.385 1178.430 ;
      LAYER met4 ;
        RECT 3402.935 1030.035 3406.385 1178.030 ;
      LAYER met4 ;
        RECT 3401.935 1029.635 3402.535 1030.035 ;
        RECT 3406.785 1029.635 3407.385 1030.035 ;
      LAYER met4 ;
        RECT 3407.785 1029.730 3412.435 1178.270 ;
      LAYER met4 ;
        RECT 3412.835 1178.030 3413.435 1178.670 ;
        RECT 3401.935 1029.330 3407.385 1029.635 ;
        RECT 3412.835 1029.330 3413.435 1030.035 ;
      LAYER met4 ;
        RECT 3413.835 1029.730 3418.485 1178.270 ;
      LAYER met4 ;
        RECT 3418.885 1178.030 3419.485 1178.670 ;
        RECT 3418.885 1029.330 3419.485 1030.035 ;
      LAYER met4 ;
        RECT 3419.885 1029.730 3423.335 1178.270 ;
      LAYER met4 ;
        RECT 3423.735 1178.030 3424.335 1178.670 ;
        RECT 3423.735 1029.330 3424.335 1030.035 ;
      LAYER met4 ;
        RECT 3424.735 1029.730 3428.185 1178.270 ;
      LAYER met4 ;
        RECT 3428.585 1178.030 3429.185 1178.670 ;
        RECT 3428.585 1029.330 3429.185 1030.035 ;
      LAYER met4 ;
        RECT 3429.585 1029.730 3434.235 1178.270 ;
      LAYER met4 ;
        RECT 3434.635 1178.030 3435.335 1178.670 ;
        RECT 3434.635 1029.330 3435.335 1030.035 ;
        RECT 3388.535 1027.990 3435.335 1029.330 ;
      LAYER met4 ;
        RECT 3435.735 1028.390 3436.065 1209.910 ;
        RECT 3436.365 1204.855 3439.345 1427.535 ;
      LAYER met4 ;
        RECT 3439.745 1403.670 3440.725 1427.935 ;
      LAYER met4 ;
        RECT 3439.645 1402.000 3440.825 1403.270 ;
      LAYER met4 ;
        RECT 3439.645 1257.000 3440.825 1402.000 ;
      LAYER met4 ;
        RECT 3439.645 1255.730 3440.825 1257.000 ;
      LAYER met4 ;
        RECT 3439.745 1220.160 3440.725 1255.330 ;
      LAYER met4 ;
        RECT 3441.125 1220.560 3444.105 1443.240 ;
      LAYER met4 ;
        RECT 3444.505 1435.310 3588.000 1443.640 ;
      LAYER met4 ;
        RECT 3444.405 1254.390 3444.735 1434.910 ;
      LAYER met4 ;
        RECT 3445.135 1403.670 3588.000 1435.310 ;
        RECT 3445.135 1403.030 3445.835 1403.670 ;
        RECT 3445.135 1257.000 3445.835 1402.000 ;
        RECT 3445.135 1255.330 3445.835 1256.035 ;
      LAYER met4 ;
        RECT 3446.235 1255.730 3450.685 1403.270 ;
      LAYER met4 ;
        RECT 3451.085 1403.030 3451.685 1403.670 ;
        RECT 3451.085 1257.000 3451.685 1402.000 ;
        RECT 3451.085 1255.330 3451.685 1256.035 ;
      LAYER met4 ;
        RECT 3452.085 1255.730 3456.535 1403.270 ;
      LAYER met4 ;
        RECT 3456.935 1403.030 3457.635 1403.670 ;
        RECT 3456.935 1257.000 3457.635 1402.000 ;
        RECT 3456.935 1255.330 3457.635 1256.035 ;
      LAYER met4 ;
        RECT 3458.035 1255.730 3483.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.400 1403.030 3563.385 1403.670 ;
      LAYER met4 ;
        RECT 3563.785 1402.000 3588.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.400 1257.000 3588.000 1402.000 ;
        RECT 3483.400 1255.330 3563.385 1256.035 ;
      LAYER met4 ;
        RECT 3563.785 1255.730 3588.000 1257.000 ;
      LAYER met4 ;
        RECT 3445.135 1253.990 3588.000 1255.330 ;
        RECT 3444.505 1220.160 3588.000 1253.990 ;
        RECT 3439.745 1218.640 3588.000 1220.160 ;
        RECT 3439.745 1204.455 3440.725 1218.640 ;
        RECT 3436.465 1202.935 3440.725 1204.455 ;
        RECT 198.365 986.330 199.465 986.970 ;
        RECT 152.665 954.690 199.465 986.330 ;
        RECT 152.035 911.010 199.465 954.690 ;
        RECT 3388.535 984.310 3435.965 1027.990 ;
        RECT 3388.535 952.670 3435.335 984.310 ;
        RECT 3388.535 952.030 3389.635 952.670 ;
      LAYER met4 ;
        RECT 151.935 631.000 152.265 910.610 ;
      LAYER met4 ;
        RECT 152.665 909.670 199.465 911.010 ;
        RECT 152.665 908.965 153.365 909.670 ;
      LAYER met4 ;
        RECT 153.765 636.000 158.415 909.270 ;
      LAYER met4 ;
        RECT 158.815 908.965 159.415 909.670 ;
      LAYER met4 ;
        RECT 159.815 631.000 163.265 909.270 ;
      LAYER met4 ;
        RECT 163.665 908.965 164.265 909.670 ;
        RECT 148.755 182.045 151.535 182.725 ;
        RECT 147.275 180.025 151.535 182.045 ;
      LAYER met4 ;
        RECT 151.935 180.425 152.265 626.000 ;
      LAYER met4 ;
        RECT 152.665 624.330 153.365 625.035 ;
      LAYER met4 ;
        RECT 153.765 624.730 158.415 631.000 ;
      LAYER met4 ;
        RECT 158.815 624.330 159.415 625.035 ;
      LAYER met4 ;
        RECT 159.815 624.730 163.265 626.000 ;
      LAYER met4 ;
        RECT 163.665 624.330 164.265 625.035 ;
      LAYER met4 ;
        RECT 164.665 624.730 168.115 909.270 ;
      LAYER met4 ;
        RECT 168.515 908.965 169.115 909.670 ;
        RECT 168.515 624.330 169.115 625.035 ;
      LAYER met4 ;
        RECT 169.515 624.730 174.165 909.270 ;
      LAYER met4 ;
        RECT 174.565 908.965 175.165 909.670 ;
        RECT 180.615 909.365 186.065 909.670 ;
        RECT 174.565 624.330 175.165 625.035 ;
      LAYER met4 ;
        RECT 175.565 624.730 180.215 909.270 ;
      LAYER met4 ;
        RECT 180.615 908.965 181.215 909.365 ;
        RECT 185.465 908.965 186.065 909.365 ;
      LAYER met4 ;
        RECT 181.615 631.000 185.065 908.965 ;
        RECT 186.465 636.000 191.115 909.270 ;
      LAYER met4 ;
        RECT 191.515 908.965 192.115 909.670 ;
      LAYER met4 ;
        RECT 181.615 625.035 185.065 626.000 ;
      LAYER met4 ;
        RECT 180.615 624.635 181.215 625.035 ;
        RECT 185.465 624.635 186.065 625.035 ;
      LAYER met4 ;
        RECT 186.465 624.730 191.115 631.000 ;
      LAYER met4 ;
        RECT 180.615 624.330 186.065 624.635 ;
        RECT 191.515 624.330 192.115 625.035 ;
      LAYER met4 ;
        RECT 192.515 624.730 197.965 909.270 ;
      LAYER met4 ;
        RECT 198.365 908.965 199.465 909.670 ;
        RECT 3388.535 804.330 3389.635 805.035 ;
      LAYER met4 ;
        RECT 3390.035 804.730 3395.485 952.270 ;
      LAYER met4 ;
        RECT 3395.885 952.030 3396.485 952.670 ;
        RECT 3401.935 952.430 3407.385 952.670 ;
        RECT 3395.885 804.330 3396.485 805.035 ;
      LAYER met4 ;
        RECT 3396.885 804.730 3401.535 952.270 ;
      LAYER met4 ;
        RECT 3401.935 952.030 3402.535 952.430 ;
        RECT 3406.785 952.030 3407.385 952.430 ;
      LAYER met4 ;
        RECT 3402.935 805.035 3406.385 952.030 ;
      LAYER met4 ;
        RECT 3401.935 804.635 3402.535 805.035 ;
        RECT 3406.785 804.635 3407.385 805.035 ;
      LAYER met4 ;
        RECT 3407.785 804.730 3412.435 952.270 ;
      LAYER met4 ;
        RECT 3412.835 952.030 3413.435 952.670 ;
        RECT 3401.935 804.330 3407.385 804.635 ;
        RECT 3412.835 804.330 3413.435 805.035 ;
      LAYER met4 ;
        RECT 3413.835 804.730 3418.485 952.270 ;
      LAYER met4 ;
        RECT 3418.885 952.030 3419.485 952.670 ;
        RECT 3418.885 804.330 3419.485 805.035 ;
      LAYER met4 ;
        RECT 3419.885 804.730 3423.335 952.270 ;
      LAYER met4 ;
        RECT 3423.735 952.030 3424.335 952.670 ;
        RECT 3423.735 804.330 3424.335 805.035 ;
      LAYER met4 ;
        RECT 3424.735 804.730 3428.185 952.270 ;
      LAYER met4 ;
        RECT 3428.585 952.030 3429.185 952.670 ;
        RECT 3428.585 804.330 3429.185 805.035 ;
      LAYER met4 ;
        RECT 3429.585 804.730 3434.235 952.270 ;
      LAYER met4 ;
        RECT 3434.635 952.030 3435.335 952.670 ;
        RECT 3434.635 804.330 3435.335 805.035 ;
        RECT 3388.535 802.990 3435.335 804.330 ;
      LAYER met4 ;
        RECT 3435.735 803.390 3436.065 983.910 ;
        RECT 3436.365 978.855 3439.345 1202.535 ;
      LAYER met4 ;
        RECT 3439.745 1178.670 3440.725 1202.935 ;
      LAYER met4 ;
        RECT 3439.645 1177.000 3440.825 1178.270 ;
      LAYER met4 ;
        RECT 3439.645 1031.000 3440.825 1177.000 ;
      LAYER met4 ;
        RECT 3439.645 1029.730 3440.825 1031.000 ;
      LAYER met4 ;
        RECT 3439.745 994.160 3440.725 1029.330 ;
      LAYER met4 ;
        RECT 3441.125 994.560 3444.105 1218.240 ;
      LAYER met4 ;
        RECT 3444.505 1210.310 3588.000 1218.640 ;
      LAYER met4 ;
        RECT 3444.405 1028.390 3444.735 1209.910 ;
      LAYER met4 ;
        RECT 3445.135 1178.670 3588.000 1210.310 ;
        RECT 3445.135 1178.030 3445.835 1178.670 ;
        RECT 3445.135 1031.000 3445.835 1177.000 ;
        RECT 3445.135 1029.330 3445.835 1030.035 ;
      LAYER met4 ;
        RECT 3446.235 1029.730 3450.685 1178.270 ;
      LAYER met4 ;
        RECT 3451.085 1178.030 3451.685 1178.670 ;
        RECT 3451.085 1031.000 3451.685 1177.000 ;
        RECT 3451.085 1029.330 3451.685 1030.035 ;
      LAYER met4 ;
        RECT 3452.085 1029.730 3456.535 1178.270 ;
      LAYER met4 ;
        RECT 3456.935 1178.030 3457.635 1178.670 ;
        RECT 3456.935 1031.000 3457.635 1177.000 ;
        RECT 3456.935 1029.330 3457.635 1030.035 ;
      LAYER met4 ;
        RECT 3458.035 1029.730 3483.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.400 1178.030 3563.385 1178.670 ;
      LAYER met4 ;
        RECT 3563.785 1177.000 3588.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.400 1031.000 3588.000 1177.000 ;
        RECT 3483.400 1029.330 3563.385 1030.035 ;
      LAYER met4 ;
        RECT 3563.785 1029.730 3588.000 1031.000 ;
      LAYER met4 ;
        RECT 3445.135 1027.990 3588.000 1029.330 ;
        RECT 3444.505 994.160 3588.000 1027.990 ;
        RECT 3439.745 992.640 3588.000 994.160 ;
        RECT 3439.745 978.455 3440.725 992.640 ;
        RECT 3436.465 976.935 3440.725 978.455 ;
        RECT 3388.535 759.310 3435.965 802.990 ;
        RECT 3388.535 727.670 3435.335 759.310 ;
        RECT 3388.535 727.030 3389.635 727.670 ;
        RECT 152.665 552.670 197.965 624.330 ;
        RECT 3388.535 578.330 3389.635 579.035 ;
      LAYER met4 ;
        RECT 3390.035 578.730 3395.485 727.270 ;
      LAYER met4 ;
        RECT 3395.885 727.030 3396.485 727.670 ;
        RECT 3401.935 727.430 3407.385 727.670 ;
        RECT 3395.885 578.330 3396.485 579.035 ;
      LAYER met4 ;
        RECT 3396.885 578.730 3401.535 727.270 ;
      LAYER met4 ;
        RECT 3401.935 727.030 3402.535 727.430 ;
        RECT 3406.785 727.030 3407.385 727.430 ;
      LAYER met4 ;
        RECT 3402.935 579.035 3406.385 727.030 ;
      LAYER met4 ;
        RECT 3401.935 578.635 3402.535 579.035 ;
        RECT 3406.785 578.635 3407.385 579.035 ;
      LAYER met4 ;
        RECT 3407.785 578.730 3412.435 727.270 ;
      LAYER met4 ;
        RECT 3412.835 727.030 3413.435 727.670 ;
        RECT 3401.935 578.330 3407.385 578.635 ;
        RECT 3412.835 578.330 3413.435 579.035 ;
      LAYER met4 ;
        RECT 3413.835 578.730 3418.485 727.270 ;
      LAYER met4 ;
        RECT 3418.885 727.030 3419.485 727.670 ;
        RECT 3418.885 578.330 3419.485 579.035 ;
      LAYER met4 ;
        RECT 3419.885 578.730 3423.335 727.270 ;
      LAYER met4 ;
        RECT 3423.735 727.030 3424.335 727.670 ;
        RECT 3423.735 578.330 3424.335 579.035 ;
      LAYER met4 ;
        RECT 3424.735 578.730 3428.185 727.270 ;
      LAYER met4 ;
        RECT 3428.585 727.030 3429.185 727.670 ;
        RECT 3428.585 578.330 3429.185 579.035 ;
      LAYER met4 ;
        RECT 3429.585 578.730 3434.235 727.270 ;
      LAYER met4 ;
        RECT 3434.635 727.030 3435.335 727.670 ;
        RECT 3434.635 578.330 3435.335 579.035 ;
        RECT 3388.535 576.990 3435.335 578.330 ;
      LAYER met4 ;
        RECT 3435.735 577.390 3436.065 758.910 ;
        RECT 3436.365 753.855 3439.345 976.535 ;
      LAYER met4 ;
        RECT 3439.745 952.670 3440.725 976.935 ;
      LAYER met4 ;
        RECT 3439.645 951.000 3440.825 952.270 ;
      LAYER met4 ;
        RECT 3439.645 806.000 3440.825 951.000 ;
      LAYER met4 ;
        RECT 3439.645 804.730 3440.825 806.000 ;
      LAYER met4 ;
        RECT 3439.745 769.160 3440.725 804.330 ;
      LAYER met4 ;
        RECT 3441.125 769.560 3444.105 992.240 ;
      LAYER met4 ;
        RECT 3444.505 984.310 3588.000 992.640 ;
      LAYER met4 ;
        RECT 3444.405 803.390 3444.735 983.910 ;
      LAYER met4 ;
        RECT 3445.135 952.670 3588.000 984.310 ;
        RECT 3445.135 952.030 3445.835 952.670 ;
        RECT 3445.135 806.000 3445.835 951.000 ;
        RECT 3445.135 804.330 3445.835 805.035 ;
      LAYER met4 ;
        RECT 3446.235 804.730 3450.685 952.270 ;
      LAYER met4 ;
        RECT 3451.085 952.030 3451.685 952.670 ;
        RECT 3451.085 806.000 3451.685 951.000 ;
        RECT 3451.085 804.330 3451.685 805.035 ;
      LAYER met4 ;
        RECT 3452.085 804.730 3456.535 952.270 ;
      LAYER met4 ;
        RECT 3456.935 952.030 3457.635 952.670 ;
        RECT 3456.935 806.000 3457.635 951.000 ;
        RECT 3456.935 804.330 3457.635 805.035 ;
      LAYER met4 ;
        RECT 3458.035 804.730 3483.000 952.270 ;
      LAYER met4 ;
        RECT 3483.400 952.030 3563.385 952.670 ;
      LAYER met4 ;
        RECT 3563.785 951.000 3588.000 952.270 ;
      LAYER met4 ;
        RECT 3483.400 806.000 3588.000 951.000 ;
        RECT 3483.400 804.330 3563.385 805.035 ;
      LAYER met4 ;
        RECT 3563.785 804.730 3588.000 806.000 ;
      LAYER met4 ;
        RECT 3445.135 802.990 3588.000 804.330 ;
        RECT 3444.505 769.160 3588.000 802.990 ;
        RECT 3439.745 767.640 3588.000 769.160 ;
        RECT 3439.745 753.455 3440.725 767.640 ;
        RECT 3436.465 751.935 3440.725 753.455 ;
        RECT 152.665 551.965 153.365 552.670 ;
        RECT 152.665 413.330 153.365 415.000 ;
      LAYER met4 ;
        RECT 153.765 413.730 158.415 552.270 ;
      LAYER met4 ;
        RECT 158.815 551.965 159.415 552.670 ;
        RECT 158.815 413.330 159.415 415.000 ;
      LAYER met4 ;
        RECT 159.815 413.730 163.265 552.270 ;
      LAYER met4 ;
        RECT 163.665 551.965 164.265 552.670 ;
        RECT 163.665 413.330 164.265 415.000 ;
      LAYER met4 ;
        RECT 164.665 413.730 168.115 552.270 ;
      LAYER met4 ;
        RECT 168.515 551.965 169.115 552.670 ;
        RECT 168.515 413.330 169.115 415.000 ;
      LAYER met4 ;
        RECT 169.515 413.730 174.165 552.270 ;
      LAYER met4 ;
        RECT 174.565 551.965 175.165 552.670 ;
        RECT 180.615 552.365 186.065 552.670 ;
        RECT 174.565 413.330 175.165 415.000 ;
      LAYER met4 ;
        RECT 175.565 413.730 180.215 552.270 ;
      LAYER met4 ;
        RECT 180.615 551.965 181.215 552.365 ;
        RECT 185.465 551.965 186.065 552.365 ;
        RECT 180.615 413.635 181.215 415.000 ;
      LAYER met4 ;
        RECT 181.615 414.035 185.065 551.965 ;
      LAYER met4 ;
        RECT 185.465 413.635 186.065 415.000 ;
      LAYER met4 ;
        RECT 186.465 413.730 191.115 552.270 ;
      LAYER met4 ;
        RECT 191.515 551.965 192.115 552.670 ;
        RECT 180.615 413.330 186.065 413.635 ;
        RECT 191.515 413.330 192.115 415.000 ;
      LAYER met4 ;
        RECT 192.515 413.730 197.965 552.270 ;
      LAYER met4 ;
        RECT 3388.535 533.310 3435.965 576.990 ;
        RECT 3388.535 501.670 3435.335 533.310 ;
        RECT 3388.535 501.030 3389.635 501.670 ;
        RECT 152.665 341.670 197.965 413.330 ;
        RECT 152.665 340.965 153.365 341.670 ;
        RECT 152.665 202.330 153.365 202.745 ;
      LAYER met4 ;
        RECT 153.765 202.730 158.415 341.270 ;
      LAYER met4 ;
        RECT 158.815 340.965 159.415 341.670 ;
        RECT 158.815 202.330 159.415 202.745 ;
      LAYER met4 ;
        RECT 159.815 202.730 163.265 341.270 ;
      LAYER met4 ;
        RECT 163.665 340.965 164.265 341.670 ;
        RECT 163.665 202.330 164.265 202.745 ;
      LAYER met4 ;
        RECT 164.665 202.730 168.115 341.270 ;
      LAYER met4 ;
        RECT 168.515 340.965 169.115 341.670 ;
        RECT 168.515 202.330 169.115 202.745 ;
      LAYER met4 ;
        RECT 169.515 202.730 174.165 341.270 ;
      LAYER met4 ;
        RECT 174.565 340.965 175.165 341.670 ;
        RECT 180.615 341.365 186.065 341.670 ;
        RECT 174.565 202.330 175.165 202.745 ;
      LAYER met4 ;
        RECT 175.565 202.730 180.215 341.270 ;
      LAYER met4 ;
        RECT 180.615 340.965 181.215 341.365 ;
        RECT 185.465 340.965 186.065 341.365 ;
      LAYER met4 ;
        RECT 181.615 202.745 185.065 340.965 ;
      LAYER met4 ;
        RECT 180.615 202.345 181.215 202.745 ;
        RECT 185.465 202.345 186.065 202.745 ;
      LAYER met4 ;
        RECT 186.465 202.730 191.115 341.270 ;
      LAYER met4 ;
        RECT 191.515 340.965 192.115 341.670 ;
        RECT 180.615 202.330 186.065 202.345 ;
        RECT 191.515 202.330 192.115 202.745 ;
      LAYER met4 ;
        RECT 192.515 202.730 197.965 341.270 ;
      LAYER met4 ;
        RECT 198.365 202.330 200.000 202.745 ;
        RECT 152.665 198.365 200.000 202.330 ;
        RECT 933.030 198.365 1011.035 199.465 ;
        RECT 1476.030 198.365 1554.035 199.465 ;
        RECT 1750.030 198.365 1828.035 199.465 ;
        RECT 2024.030 198.365 2102.035 199.465 ;
        RECT 2298.030 198.365 2376.035 199.465 ;
        RECT 2572.030 198.365 2650.035 199.465 ;
        RECT 3385.255 198.365 3389.635 200.000 ;
        RECT 152.665 192.115 197.250 198.365 ;
      LAYER met4 ;
        RECT 197.650 192.515 395.270 197.965 ;
      LAYER met4 ;
        RECT 395.670 192.115 467.330 197.965 ;
      LAYER met4 ;
        RECT 467.730 192.515 664.270 197.965 ;
      LAYER met4 ;
        RECT 664.670 192.115 736.330 197.965 ;
      LAYER met4 ;
        RECT 736.730 192.515 933.270 197.965 ;
      LAYER met4 ;
        RECT 933.670 192.115 1010.330 198.365 ;
      LAYER met4 ;
        RECT 1010.730 192.515 1207.270 197.965 ;
      LAYER met4 ;
        RECT 1207.670 192.115 1279.330 197.965 ;
      LAYER met4 ;
        RECT 1279.730 192.515 1476.270 197.965 ;
      LAYER met4 ;
        RECT 1476.670 192.115 1553.330 198.365 ;
      LAYER met4 ;
        RECT 1553.730 192.515 1750.270 197.965 ;
      LAYER met4 ;
        RECT 1750.670 192.115 1827.330 198.365 ;
      LAYER met4 ;
        RECT 1827.730 192.515 2024.270 197.965 ;
      LAYER met4 ;
        RECT 2024.670 192.115 2101.330 198.365 ;
      LAYER met4 ;
        RECT 2101.730 192.515 2298.270 197.965 ;
      LAYER met4 ;
        RECT 2298.670 192.115 2375.330 198.365 ;
      LAYER met4 ;
        RECT 2375.730 192.515 2572.270 197.965 ;
      LAYER met4 ;
        RECT 2572.670 192.115 2649.330 198.365 ;
      LAYER met4 ;
        RECT 2649.730 192.515 2846.270 197.965 ;
      LAYER met4 ;
        RECT 2846.670 192.115 2918.330 197.965 ;
      LAYER met4 ;
        RECT 2918.730 192.515 3115.270 197.965 ;
      LAYER met4 ;
        RECT 3115.670 192.115 3187.330 197.965 ;
      LAYER met4 ;
        RECT 3187.730 192.515 3385.270 197.965 ;
      LAYER met4 ;
        RECT 3385.670 197.250 3389.635 198.365 ;
      LAYER met4 ;
        RECT 3390.035 197.650 3395.485 501.270 ;
      LAYER met4 ;
        RECT 3395.885 501.030 3396.485 501.670 ;
        RECT 3401.935 501.430 3407.385 501.670 ;
      LAYER met4 ;
        RECT 3396.885 355.000 3401.535 501.270 ;
      LAYER met4 ;
        RECT 3401.935 501.030 3402.535 501.430 ;
        RECT 3406.785 501.030 3407.385 501.430 ;
      LAYER met4 ;
        RECT 3402.935 350.000 3406.385 501.030 ;
      LAYER met4 ;
        RECT 3395.885 197.250 3396.485 200.000 ;
        RECT 3385.670 195.815 3396.485 197.250 ;
      LAYER met4 ;
        RECT 3396.885 196.215 3401.535 350.000 ;
      LAYER met4 ;
        RECT 3401.935 198.130 3402.535 200.000 ;
      LAYER met4 ;
        RECT 3402.935 198.530 3406.385 345.000 ;
      LAYER met4 ;
        RECT 3406.785 198.130 3407.385 200.000 ;
      LAYER met4 ;
        RECT 3407.785 198.475 3412.435 501.270 ;
      LAYER met4 ;
        RECT 3412.835 501.030 3413.435 501.670 ;
        RECT 3401.935 198.075 3407.385 198.130 ;
        RECT 3412.835 198.075 3413.435 200.000 ;
      LAYER met4 ;
        RECT 3413.835 198.400 3418.485 501.270 ;
      LAYER met4 ;
        RECT 3418.885 501.030 3419.485 501.670 ;
        RECT 3401.935 198.000 3413.435 198.075 ;
        RECT 3418.885 198.215 3419.485 200.000 ;
      LAYER met4 ;
        RECT 3419.885 198.615 3423.335 501.270 ;
      LAYER met4 ;
        RECT 3423.735 501.030 3424.335 501.670 ;
      LAYER met4 ;
        RECT 3424.735 350.000 3428.185 501.270 ;
      LAYER met4 ;
        RECT 3428.585 501.030 3429.185 501.670 ;
      LAYER met4 ;
        RECT 3429.585 355.000 3434.235 501.270 ;
      LAYER met4 ;
        RECT 3434.635 501.030 3435.335 501.670 ;
      LAYER met4 ;
        RECT 3435.735 350.000 3436.065 532.910 ;
        RECT 3436.365 527.855 3439.345 751.535 ;
      LAYER met4 ;
        RECT 3439.745 727.670 3440.725 751.935 ;
      LAYER met4 ;
        RECT 3439.645 726.000 3440.825 727.270 ;
      LAYER met4 ;
        RECT 3439.645 580.000 3440.825 726.000 ;
      LAYER met4 ;
        RECT 3439.645 578.730 3440.825 580.000 ;
      LAYER met4 ;
        RECT 3439.745 543.160 3440.725 578.330 ;
      LAYER met4 ;
        RECT 3441.125 543.560 3444.105 767.240 ;
      LAYER met4 ;
        RECT 3444.505 759.310 3588.000 767.640 ;
      LAYER met4 ;
        RECT 3444.405 577.390 3444.735 758.910 ;
      LAYER met4 ;
        RECT 3445.135 727.670 3588.000 759.310 ;
        RECT 3445.135 727.030 3445.835 727.670 ;
        RECT 3445.135 580.000 3445.835 726.000 ;
        RECT 3445.135 578.330 3445.835 579.035 ;
      LAYER met4 ;
        RECT 3446.235 578.730 3450.685 727.270 ;
      LAYER met4 ;
        RECT 3451.085 727.030 3451.685 727.670 ;
        RECT 3451.085 580.000 3451.685 726.000 ;
        RECT 3451.085 578.330 3451.685 579.035 ;
      LAYER met4 ;
        RECT 3452.085 578.730 3456.535 727.270 ;
      LAYER met4 ;
        RECT 3456.935 727.030 3457.635 727.670 ;
        RECT 3456.935 580.000 3457.635 726.000 ;
        RECT 3456.935 578.330 3457.635 579.035 ;
      LAYER met4 ;
        RECT 3458.035 578.730 3483.000 727.270 ;
      LAYER met4 ;
        RECT 3483.400 727.030 3563.385 727.670 ;
      LAYER met4 ;
        RECT 3563.785 726.000 3588.000 727.270 ;
      LAYER met4 ;
        RECT 3483.400 580.000 3588.000 726.000 ;
        RECT 3483.400 578.330 3563.385 579.035 ;
      LAYER met4 ;
        RECT 3563.785 578.730 3588.000 580.000 ;
      LAYER met4 ;
        RECT 3445.135 576.990 3588.000 578.330 ;
        RECT 3444.505 543.160 3588.000 576.990 ;
        RECT 3439.745 541.640 3588.000 543.160 ;
        RECT 3439.745 527.455 3440.725 541.640 ;
        RECT 3436.465 525.935 3440.725 527.455 ;
        RECT 3423.735 198.265 3424.335 200.000 ;
      LAYER met4 ;
        RECT 3424.735 198.665 3428.185 345.000 ;
      LAYER met4 ;
        RECT 3428.585 198.265 3429.185 200.000 ;
      LAYER met4 ;
        RECT 3429.585 198.525 3434.235 350.000 ;
      LAYER met4 ;
        RECT 3423.735 198.215 3429.185 198.265 ;
        RECT 3418.885 198.125 3429.185 198.215 ;
        RECT 3434.635 198.125 3435.335 200.000 ;
        RECT 3418.885 198.000 3435.335 198.125 ;
        RECT 3401.935 195.815 3435.335 198.000 ;
        RECT 3385.670 192.115 3435.335 195.815 ;
        RECT 152.665 191.515 200.000 192.115 ;
        RECT 394.965 191.515 468.035 192.115 ;
        RECT 663.965 191.515 737.035 192.115 ;
        RECT 933.030 191.515 1011.035 192.115 ;
        RECT 1206.000 191.515 1280.035 192.115 ;
        RECT 1476.030 191.515 1554.035 192.115 ;
        RECT 1750.030 191.515 1828.035 192.115 ;
        RECT 2024.030 191.515 2102.035 192.115 ;
        RECT 2298.030 191.515 2376.035 192.115 ;
        RECT 2572.030 191.515 2650.035 192.115 ;
        RECT 2845.965 191.515 2919.035 192.115 ;
        RECT 3114.965 191.515 3188.035 192.115 ;
        RECT 3385.255 191.515 3435.335 192.115 ;
        RECT 152.665 186.065 195.815 191.515 ;
      LAYER met4 ;
        RECT 196.215 186.465 395.270 191.115 ;
      LAYER met4 ;
        RECT 395.670 186.065 467.330 191.515 ;
      LAYER met4 ;
        RECT 467.730 186.465 664.270 191.115 ;
      LAYER met4 ;
        RECT 664.670 186.065 736.330 191.515 ;
      LAYER met4 ;
        RECT 736.730 186.465 933.270 191.115 ;
      LAYER met4 ;
        RECT 933.670 186.065 1010.330 191.515 ;
      LAYER met4 ;
        RECT 1010.730 186.465 1207.270 191.115 ;
      LAYER met4 ;
        RECT 1207.670 186.065 1279.330 191.515 ;
      LAYER met4 ;
        RECT 1279.730 186.465 1476.270 191.115 ;
      LAYER met4 ;
        RECT 1476.670 186.065 1553.330 191.515 ;
      LAYER met4 ;
        RECT 1553.730 186.465 1750.270 191.115 ;
      LAYER met4 ;
        RECT 1750.670 186.065 1827.330 191.515 ;
      LAYER met4 ;
        RECT 1827.730 186.465 2024.270 191.115 ;
      LAYER met4 ;
        RECT 2024.670 186.065 2101.330 191.515 ;
      LAYER met4 ;
        RECT 2101.730 186.465 2298.270 191.115 ;
      LAYER met4 ;
        RECT 2298.670 186.065 2375.330 191.515 ;
      LAYER met4 ;
        RECT 2375.730 186.465 2572.270 191.115 ;
      LAYER met4 ;
        RECT 2572.670 186.065 2649.330 191.515 ;
      LAYER met4 ;
        RECT 2649.730 186.465 2846.270 191.115 ;
      LAYER met4 ;
        RECT 2846.670 186.065 2918.330 191.515 ;
      LAYER met4 ;
        RECT 2918.730 186.465 3115.270 191.115 ;
      LAYER met4 ;
        RECT 3115.670 186.065 3187.330 191.515 ;
      LAYER met4 ;
        RECT 3187.730 186.465 3385.270 191.115 ;
      LAYER met4 ;
        RECT 3385.670 186.065 3435.335 191.515 ;
        RECT 152.665 185.465 200.000 186.065 ;
        RECT 394.965 185.465 468.035 186.065 ;
        RECT 663.965 185.465 737.035 186.065 ;
        RECT 933.030 185.465 1011.035 186.065 ;
        RECT 1206.000 185.465 1280.035 186.065 ;
        RECT 1476.030 185.465 1554.035 186.065 ;
        RECT 1750.030 185.465 1828.035 186.065 ;
        RECT 2024.030 185.465 2102.035 186.065 ;
        RECT 2298.030 185.465 2376.035 186.065 ;
        RECT 2572.030 185.465 2650.035 186.065 ;
        RECT 2845.965 185.465 2919.035 186.065 ;
        RECT 3114.965 185.465 3188.035 186.065 ;
        RECT 3385.255 185.465 3435.335 186.065 ;
        RECT 152.665 181.215 198.130 185.465 ;
      LAYER met4 ;
        RECT 198.530 181.615 394.965 185.065 ;
      LAYER met4 ;
        RECT 395.365 181.215 467.635 185.465 ;
        RECT 664.365 181.215 736.635 185.465 ;
      LAYER met4 ;
        RECT 737.035 181.615 933.030 185.065 ;
      LAYER met4 ;
        RECT 933.430 181.215 1010.635 185.465 ;
      LAYER met4 ;
        RECT 1011.035 181.615 1206.965 185.065 ;
      LAYER met4 ;
        RECT 1207.365 181.215 1279.635 185.465 ;
      LAYER met4 ;
        RECT 1280.035 181.615 1476.030 185.065 ;
      LAYER met4 ;
        RECT 1476.430 181.215 1553.635 185.465 ;
      LAYER met4 ;
        RECT 1554.035 181.615 1750.030 185.065 ;
      LAYER met4 ;
        RECT 1750.430 181.215 1827.635 185.465 ;
      LAYER met4 ;
        RECT 1828.035 181.615 2024.030 185.065 ;
      LAYER met4 ;
        RECT 2024.430 181.215 2101.635 185.465 ;
      LAYER met4 ;
        RECT 2102.035 181.615 2298.030 185.065 ;
      LAYER met4 ;
        RECT 2298.430 181.215 2375.635 185.465 ;
      LAYER met4 ;
        RECT 2376.035 181.615 2572.030 185.065 ;
      LAYER met4 ;
        RECT 2572.430 181.215 2649.635 185.465 ;
      LAYER met4 ;
        RECT 2650.035 181.615 2845.965 185.065 ;
      LAYER met4 ;
        RECT 2846.365 181.215 2918.635 185.465 ;
      LAYER met4 ;
        RECT 2919.035 181.615 3114.965 185.065 ;
      LAYER met4 ;
        RECT 3115.365 181.215 3187.635 185.465 ;
      LAYER met4 ;
        RECT 3188.035 181.615 3385.255 185.065 ;
      LAYER met4 ;
        RECT 3385.655 181.215 3435.335 185.465 ;
        RECT 152.665 180.615 200.000 181.215 ;
        RECT 394.965 180.615 468.035 181.215 ;
        RECT 663.965 180.615 737.035 181.215 ;
        RECT 933.030 180.615 1011.035 181.215 ;
        RECT 1206.000 180.615 1280.035 181.215 ;
        RECT 1476.030 180.615 1554.035 181.215 ;
        RECT 1750.030 180.615 1828.035 181.215 ;
        RECT 2024.030 180.615 2102.035 181.215 ;
        RECT 2298.030 180.615 2376.035 181.215 ;
        RECT 2572.030 180.615 2650.035 181.215 ;
        RECT 2845.965 180.615 2919.035 181.215 ;
        RECT 3114.965 180.615 3188.035 181.215 ;
        RECT 3385.255 180.615 3435.335 181.215 ;
        RECT 152.665 180.025 198.075 180.615 ;
        RECT 147.275 176.690 198.075 180.025 ;
        RECT 143.995 176.425 198.075 176.690 ;
        RECT 0.000 175.165 198.075 176.425 ;
      LAYER met4 ;
        RECT 198.475 175.565 395.270 180.215 ;
      LAYER met4 ;
        RECT 395.670 175.165 467.330 180.615 ;
      LAYER met4 ;
        RECT 467.730 175.565 664.270 180.215 ;
      LAYER met4 ;
        RECT 664.670 175.165 736.330 180.615 ;
      LAYER met4 ;
        RECT 736.730 175.565 933.270 180.215 ;
      LAYER met4 ;
        RECT 933.670 175.165 1010.330 180.615 ;
      LAYER met4 ;
        RECT 1010.730 175.565 1207.270 180.215 ;
      LAYER met4 ;
        RECT 1207.670 175.165 1279.330 180.615 ;
      LAYER met4 ;
        RECT 1279.730 175.565 1476.270 180.215 ;
      LAYER met4 ;
        RECT 1476.670 175.165 1553.330 180.615 ;
      LAYER met4 ;
        RECT 1553.730 175.565 1750.270 180.215 ;
      LAYER met4 ;
        RECT 1750.670 175.165 1827.330 180.615 ;
      LAYER met4 ;
        RECT 1827.730 175.565 2024.270 180.215 ;
      LAYER met4 ;
        RECT 2024.670 175.165 2101.330 180.615 ;
      LAYER met4 ;
        RECT 2101.730 175.565 2298.270 180.215 ;
      LAYER met4 ;
        RECT 2298.670 175.165 2375.330 180.615 ;
      LAYER met4 ;
        RECT 2375.730 175.565 2572.270 180.215 ;
      LAYER met4 ;
        RECT 2572.670 175.165 2649.330 180.615 ;
      LAYER met4 ;
        RECT 2649.730 175.565 2846.270 180.215 ;
      LAYER met4 ;
        RECT 2846.670 175.165 2918.330 180.615 ;
      LAYER met4 ;
        RECT 2918.730 175.565 3115.270 180.215 ;
      LAYER met4 ;
        RECT 3115.670 175.165 3187.330 180.615 ;
      LAYER met4 ;
        RECT 3187.730 175.565 3385.270 180.215 ;
      LAYER met4 ;
        RECT 3385.670 180.025 3435.335 180.615 ;
      LAYER met4 ;
        RECT 3435.735 180.425 3436.065 345.000 ;
      LAYER met4 ;
        RECT 3385.670 178.665 3435.965 180.025 ;
      LAYER met4 ;
        RECT 3436.365 179.065 3439.345 525.535 ;
      LAYER met4 ;
        RECT 3439.745 501.670 3440.725 525.935 ;
      LAYER met4 ;
        RECT 3439.645 500.000 3440.825 501.270 ;
      LAYER met4 ;
        RECT 3439.645 350.000 3440.825 500.000 ;
        RECT 3439.645 200.000 3440.825 345.000 ;
        RECT 3385.670 178.050 3439.245 178.665 ;
      LAYER met4 ;
        RECT 3439.645 178.450 3440.825 200.000 ;
      LAYER met4 ;
        RECT 3385.670 176.690 3440.725 178.050 ;
      LAYER met4 ;
        RECT 3441.125 177.090 3444.105 541.240 ;
      LAYER met4 ;
        RECT 3444.505 533.310 3588.000 541.640 ;
      LAYER met4 ;
        RECT 3444.405 350.000 3444.735 532.910 ;
      LAYER met4 ;
        RECT 3445.135 501.670 3588.000 533.310 ;
        RECT 3445.135 501.030 3445.835 501.670 ;
        RECT 3445.135 350.000 3445.835 500.000 ;
      LAYER met4 ;
        RECT 3444.405 176.825 3444.735 345.000 ;
      LAYER met4 ;
        RECT 3445.135 197.975 3445.835 345.000 ;
      LAYER met4 ;
        RECT 3446.235 198.375 3450.685 501.270 ;
      LAYER met4 ;
        RECT 3451.085 501.030 3451.685 501.670 ;
        RECT 3451.085 350.000 3451.685 500.000 ;
        RECT 3451.085 198.120 3451.685 345.000 ;
      LAYER met4 ;
        RECT 3452.085 198.520 3456.535 501.270 ;
      LAYER met4 ;
        RECT 3456.935 501.030 3457.635 501.670 ;
        RECT 3456.935 350.000 3457.635 500.000 ;
        RECT 3456.935 198.120 3457.635 345.000 ;
        RECT 3451.085 197.975 3457.635 198.120 ;
        RECT 3445.135 196.955 3457.635 197.975 ;
      LAYER met4 ;
        RECT 3458.035 197.355 3483.000 501.270 ;
      LAYER met4 ;
        RECT 3483.400 501.030 3563.385 501.670 ;
      LAYER met4 ;
        RECT 3563.785 500.000 3588.000 501.270 ;
      LAYER met4 ;
        RECT 3483.400 350.000 3588.000 500.000 ;
        RECT 3563.785 345.000 3588.000 350.000 ;
        RECT 3483.400 200.000 3588.000 345.000 ;
        RECT 3483.400 198.165 3563.385 200.000 ;
      LAYER met4 ;
        RECT 3563.785 198.565 3588.000 200.000 ;
      LAYER met4 ;
        RECT 3483.400 196.955 3588.000 198.165 ;
        RECT 3385.670 176.425 3444.005 176.690 ;
        RECT 3445.135 176.425 3588.000 196.955 ;
        RECT 3385.670 175.165 3588.000 176.425 ;
        RECT 0.000 174.565 200.000 175.165 ;
        RECT 394.965 174.565 468.035 175.165 ;
        RECT 663.965 174.565 737.035 175.165 ;
        RECT 933.030 174.565 1011.035 175.165 ;
        RECT 1206.000 174.565 1280.035 175.165 ;
        RECT 1476.030 174.565 1554.035 175.165 ;
        RECT 1750.030 174.565 1828.035 175.165 ;
        RECT 2024.030 174.565 2102.035 175.165 ;
        RECT 2298.030 174.565 2376.035 175.165 ;
        RECT 2572.030 174.565 2650.035 175.165 ;
        RECT 2845.965 174.565 2919.035 175.165 ;
        RECT 3114.965 174.565 3188.035 175.165 ;
        RECT 3385.255 174.565 3588.000 175.165 ;
        RECT 0.000 169.115 198.000 174.565 ;
      LAYER met4 ;
        RECT 198.400 169.515 395.270 174.165 ;
      LAYER met4 ;
        RECT 395.670 169.115 467.330 174.565 ;
      LAYER met4 ;
        RECT 467.730 169.515 664.270 174.165 ;
      LAYER met4 ;
        RECT 664.670 169.115 736.330 174.565 ;
      LAYER met4 ;
        RECT 736.730 169.515 933.270 174.165 ;
      LAYER met4 ;
        RECT 933.670 169.115 1010.330 174.565 ;
      LAYER met4 ;
        RECT 1010.730 169.515 1207.270 174.165 ;
      LAYER met4 ;
        RECT 1207.670 169.115 1279.330 174.565 ;
      LAYER met4 ;
        RECT 1279.730 169.515 1476.270 174.165 ;
      LAYER met4 ;
        RECT 1476.670 169.115 1553.330 174.565 ;
      LAYER met4 ;
        RECT 1553.730 169.515 1750.270 174.165 ;
      LAYER met4 ;
        RECT 1750.670 169.115 1827.330 174.565 ;
      LAYER met4 ;
        RECT 1827.730 169.515 2024.270 174.165 ;
      LAYER met4 ;
        RECT 2024.670 169.115 2101.330 174.565 ;
      LAYER met4 ;
        RECT 2101.730 169.515 2298.270 174.165 ;
      LAYER met4 ;
        RECT 2298.670 169.115 2375.330 174.565 ;
      LAYER met4 ;
        RECT 2375.730 169.515 2572.270 174.165 ;
      LAYER met4 ;
        RECT 2572.670 169.115 2649.330 174.565 ;
      LAYER met4 ;
        RECT 2649.730 169.515 2846.270 174.165 ;
      LAYER met4 ;
        RECT 2846.670 169.115 2918.330 174.565 ;
      LAYER met4 ;
        RECT 2918.730 169.515 3115.270 174.165 ;
      LAYER met4 ;
        RECT 3115.670 169.115 3187.330 174.565 ;
      LAYER met4 ;
        RECT 3187.730 169.515 3385.270 174.165 ;
      LAYER met4 ;
        RECT 3385.670 169.115 3588.000 174.565 ;
        RECT 0.000 168.515 200.000 169.115 ;
        RECT 394.965 168.515 468.035 169.115 ;
        RECT 663.965 168.515 737.035 169.115 ;
        RECT 933.030 168.515 1011.035 169.115 ;
        RECT 1206.000 168.515 1280.035 169.115 ;
        RECT 1476.030 168.515 1554.035 169.115 ;
        RECT 1750.030 168.515 1828.035 169.115 ;
        RECT 2024.030 168.515 2102.035 169.115 ;
        RECT 2298.030 168.515 2376.035 169.115 ;
        RECT 2572.030 168.515 2650.035 169.115 ;
        RECT 2845.965 168.515 2919.035 169.115 ;
        RECT 3114.965 168.515 3188.035 169.115 ;
        RECT 3385.255 168.515 3588.000 169.115 ;
        RECT 0.000 164.265 198.215 168.515 ;
      LAYER met4 ;
        RECT 198.615 164.665 395.270 168.115 ;
      LAYER met4 ;
        RECT 395.670 164.265 467.330 168.515 ;
      LAYER met4 ;
        RECT 467.730 164.665 664.270 168.115 ;
      LAYER met4 ;
        RECT 664.670 164.265 736.330 168.515 ;
      LAYER met4 ;
        RECT 736.730 164.665 933.270 168.115 ;
      LAYER met4 ;
        RECT 933.670 164.265 1010.330 168.515 ;
      LAYER met4 ;
        RECT 1010.730 164.665 1207.270 168.115 ;
      LAYER met4 ;
        RECT 1207.670 164.265 1279.330 168.515 ;
      LAYER met4 ;
        RECT 1279.730 164.665 1476.270 168.115 ;
      LAYER met4 ;
        RECT 1476.670 164.265 1553.330 168.515 ;
      LAYER met4 ;
        RECT 1553.730 164.665 1750.270 168.115 ;
      LAYER met4 ;
        RECT 1750.670 164.265 1827.330 168.515 ;
      LAYER met4 ;
        RECT 1827.730 164.665 2024.270 168.115 ;
      LAYER met4 ;
        RECT 2024.670 164.265 2101.330 168.515 ;
      LAYER met4 ;
        RECT 2101.730 164.665 2298.270 168.115 ;
      LAYER met4 ;
        RECT 2298.670 164.265 2375.330 168.515 ;
      LAYER met4 ;
        RECT 2375.730 164.665 2572.270 168.115 ;
      LAYER met4 ;
        RECT 2572.670 164.265 2649.330 168.515 ;
      LAYER met4 ;
        RECT 2649.730 164.665 2846.270 168.115 ;
      LAYER met4 ;
        RECT 2846.670 164.265 2918.330 168.515 ;
      LAYER met4 ;
        RECT 2918.730 164.665 3115.270 168.115 ;
      LAYER met4 ;
        RECT 3115.670 164.265 3187.330 168.515 ;
      LAYER met4 ;
        RECT 3187.730 164.665 3385.270 168.115 ;
      LAYER met4 ;
        RECT 3385.670 164.265 3588.000 168.515 ;
        RECT 0.000 163.665 200.000 164.265 ;
        RECT 394.965 163.665 468.035 164.265 ;
        RECT 663.965 163.665 737.035 164.265 ;
        RECT 933.030 163.665 1011.035 164.265 ;
        RECT 1206.000 163.665 1280.035 164.265 ;
        RECT 1476.030 163.665 1554.035 164.265 ;
        RECT 1750.030 163.665 1828.035 164.265 ;
        RECT 2024.030 163.665 2102.035 164.265 ;
        RECT 2298.030 163.665 2376.035 164.265 ;
        RECT 2572.030 163.665 2650.035 164.265 ;
        RECT 2845.965 163.665 2919.035 164.265 ;
        RECT 3114.965 163.665 3188.035 164.265 ;
        RECT 3385.255 163.665 3588.000 164.265 ;
        RECT 0.000 159.415 198.265 163.665 ;
      LAYER met4 ;
        RECT 198.665 159.815 395.270 163.265 ;
      LAYER met4 ;
        RECT 395.670 159.415 467.330 163.665 ;
      LAYER met4 ;
        RECT 467.730 159.815 664.270 163.265 ;
      LAYER met4 ;
        RECT 664.670 159.415 736.330 163.665 ;
      LAYER met4 ;
        RECT 736.730 159.815 933.270 163.265 ;
      LAYER met4 ;
        RECT 933.670 159.415 1010.330 163.665 ;
      LAYER met4 ;
        RECT 1010.730 159.815 1207.270 163.265 ;
      LAYER met4 ;
        RECT 1207.670 159.415 1279.330 163.665 ;
      LAYER met4 ;
        RECT 1279.730 159.815 1476.270 163.265 ;
      LAYER met4 ;
        RECT 1476.670 159.415 1553.330 163.665 ;
      LAYER met4 ;
        RECT 1553.730 159.815 1750.270 163.265 ;
      LAYER met4 ;
        RECT 1750.670 159.415 1827.330 163.665 ;
      LAYER met4 ;
        RECT 1827.730 159.815 2024.270 163.265 ;
      LAYER met4 ;
        RECT 2024.670 159.415 2101.330 163.665 ;
      LAYER met4 ;
        RECT 2101.730 159.815 2298.270 163.265 ;
      LAYER met4 ;
        RECT 2298.670 159.415 2375.330 163.665 ;
      LAYER met4 ;
        RECT 2375.730 159.815 2572.270 163.265 ;
      LAYER met4 ;
        RECT 2572.670 159.415 2649.330 163.665 ;
      LAYER met4 ;
        RECT 2649.730 159.815 2846.270 163.265 ;
      LAYER met4 ;
        RECT 2846.670 159.415 2918.330 163.665 ;
      LAYER met4 ;
        RECT 2918.730 159.815 3115.270 163.265 ;
      LAYER met4 ;
        RECT 3115.670 159.415 3187.330 163.665 ;
      LAYER met4 ;
        RECT 3187.730 159.815 3385.270 163.265 ;
      LAYER met4 ;
        RECT 3385.670 159.415 3588.000 163.665 ;
        RECT 0.000 158.815 200.000 159.415 ;
        RECT 394.965 158.815 468.035 159.415 ;
        RECT 663.965 158.815 737.035 159.415 ;
        RECT 933.030 158.815 1011.035 159.415 ;
        RECT 1206.000 158.815 1280.035 159.415 ;
        RECT 1476.030 158.815 1554.035 159.415 ;
        RECT 1750.030 158.815 1828.035 159.415 ;
        RECT 2024.030 158.815 2102.035 159.415 ;
        RECT 2298.030 158.815 2376.035 159.415 ;
        RECT 2572.030 158.815 2650.035 159.415 ;
        RECT 2845.965 158.815 2919.035 159.415 ;
        RECT 3114.965 158.815 3188.035 159.415 ;
        RECT 3385.255 158.815 3588.000 159.415 ;
        RECT 0.000 153.365 198.125 158.815 ;
      LAYER met4 ;
        RECT 198.525 153.765 395.270 158.415 ;
      LAYER met4 ;
        RECT 395.670 153.365 467.330 158.815 ;
        RECT 664.670 158.770 736.330 158.815 ;
        RECT 664.745 153.410 736.330 158.770 ;
      LAYER met4 ;
        RECT 736.730 153.765 933.270 158.415 ;
      LAYER met4 ;
        RECT 664.670 153.365 736.330 153.410 ;
        RECT 933.670 153.365 1010.330 158.815 ;
      LAYER met4 ;
        RECT 1010.730 153.765 1207.270 158.415 ;
      LAYER met4 ;
        RECT 1207.670 153.365 1279.330 158.815 ;
      LAYER met4 ;
        RECT 1279.730 153.765 1476.270 158.415 ;
      LAYER met4 ;
        RECT 1476.670 153.365 1553.330 158.815 ;
      LAYER met4 ;
        RECT 1553.730 153.765 1750.270 158.415 ;
      LAYER met4 ;
        RECT 1750.670 153.365 1827.330 158.815 ;
      LAYER met4 ;
        RECT 1827.730 153.765 2024.270 158.415 ;
      LAYER met4 ;
        RECT 2024.670 153.365 2101.330 158.815 ;
      LAYER met4 ;
        RECT 2101.730 153.765 2298.270 158.415 ;
      LAYER met4 ;
        RECT 2298.670 153.365 2375.330 158.815 ;
      LAYER met4 ;
        RECT 2375.730 153.765 2572.270 158.415 ;
      LAYER met4 ;
        RECT 2572.670 153.365 2649.330 158.815 ;
      LAYER met4 ;
        RECT 2649.730 153.765 2846.270 158.415 ;
      LAYER met4 ;
        RECT 2846.670 153.365 2918.330 158.815 ;
      LAYER met4 ;
        RECT 2918.730 153.765 3115.270 158.415 ;
      LAYER met4 ;
        RECT 3115.670 153.365 3187.330 158.815 ;
      LAYER met4 ;
        RECT 3187.730 153.765 3385.270 158.415 ;
      LAYER met4 ;
        RECT 3385.670 153.365 3588.000 158.815 ;
        RECT 0.000 152.665 200.000 153.365 ;
        RECT 394.965 152.665 468.035 153.365 ;
        RECT 663.965 152.665 737.035 153.365 ;
        RECT 933.030 152.665 1011.035 153.365 ;
        RECT 1206.000 152.665 1280.035 153.365 ;
        RECT 1476.030 152.665 1554.035 153.365 ;
        RECT 1750.030 152.665 1828.035 153.365 ;
        RECT 2024.030 152.665 2102.035 153.365 ;
        RECT 2298.030 152.665 2376.035 153.365 ;
        RECT 2572.030 152.665 2650.035 153.365 ;
        RECT 2845.965 152.665 2919.035 153.365 ;
        RECT 3114.965 152.665 3188.035 153.365 ;
        RECT 3385.255 152.665 3588.000 153.365 ;
        RECT 0.000 152.035 180.025 152.665 ;
        RECT 0.000 148.755 178.665 152.035 ;
      LAYER met4 ;
        RECT 180.425 151.935 395.270 152.265 ;
      LAYER met4 ;
        RECT 395.670 152.035 467.330 152.665 ;
      LAYER met4 ;
        RECT 467.730 151.935 964.910 152.265 ;
      LAYER met4 ;
        RECT 965.310 152.035 1008.990 152.665 ;
      LAYER met4 ;
        RECT 1009.390 151.935 1507.910 152.265 ;
      LAYER met4 ;
        RECT 1508.310 152.035 1551.990 152.665 ;
      LAYER met4 ;
        RECT 1552.390 151.935 1781.910 152.265 ;
      LAYER met4 ;
        RECT 1782.310 152.035 1825.990 152.665 ;
      LAYER met4 ;
        RECT 1826.390 151.935 2055.910 152.265 ;
      LAYER met4 ;
        RECT 2056.310 152.035 2099.990 152.665 ;
      LAYER met4 ;
        RECT 2100.390 151.935 2329.910 152.265 ;
      LAYER met4 ;
        RECT 2330.310 152.035 2373.990 152.665 ;
      LAYER met4 ;
        RECT 2374.390 151.935 2603.910 152.265 ;
      LAYER met4 ;
        RECT 2604.310 152.035 2647.990 152.665 ;
      LAYER met4 ;
        RECT 2648.390 151.935 3407.575 152.265 ;
      LAYER met4 ;
        RECT 0.000 147.275 178.050 148.755 ;
      LAYER met4 ;
        RECT 179.065 148.655 957.535 151.635 ;
      LAYER met4 ;
        RECT 0.000 143.995 176.690 147.275 ;
      LAYER met4 ;
        RECT 178.450 147.175 200.000 148.355 ;
      LAYER met4 ;
        RECT 200.000 147.175 394.000 148.355 ;
      LAYER met4 ;
        RECT 394.000 147.175 395.270 148.355 ;
      LAYER met4 ;
        RECT 395.670 147.275 467.330 148.255 ;
      LAYER met4 ;
        RECT 467.730 147.175 469.000 148.355 ;
      LAYER met4 ;
        RECT 469.000 147.175 663.000 148.355 ;
      LAYER met4 ;
        RECT 663.000 147.175 664.270 148.355 ;
      LAYER met4 ;
        RECT 664.670 147.275 736.330 148.255 ;
      LAYER met4 ;
        RECT 736.730 147.175 738.000 148.355 ;
      LAYER met4 ;
        RECT 738.000 147.175 932.000 148.355 ;
      LAYER met4 ;
        RECT 932.000 147.175 933.270 148.355 ;
      LAYER met4 ;
        RECT 957.935 148.255 959.455 151.535 ;
      LAYER met4 ;
        RECT 959.855 148.655 1500.535 151.635 ;
      LAYER met4 ;
        RECT 933.670 147.275 1010.330 148.255 ;
        RECT 0.000 142.865 176.425 143.995 ;
      LAYER met4 ;
        RECT 177.090 143.895 973.240 146.875 ;
        RECT 176.825 143.265 395.270 143.595 ;
      LAYER met4 ;
        RECT 973.640 143.495 975.160 147.275 ;
      LAYER met4 ;
        RECT 1010.730 147.175 1012.000 148.355 ;
      LAYER met4 ;
        RECT 1012.000 147.175 1206.000 148.355 ;
      LAYER met4 ;
        RECT 1206.000 147.175 1207.270 148.355 ;
      LAYER met4 ;
        RECT 1207.670 147.275 1279.330 148.255 ;
      LAYER met4 ;
        RECT 1279.730 147.175 1281.000 148.355 ;
      LAYER met4 ;
        RECT 1281.000 147.175 1475.000 148.355 ;
      LAYER met4 ;
        RECT 1475.000 147.175 1476.270 148.355 ;
      LAYER met4 ;
        RECT 1500.935 148.255 1502.455 151.535 ;
      LAYER met4 ;
        RECT 1502.855 148.655 1774.535 151.635 ;
      LAYER met4 ;
        RECT 1476.670 147.275 1553.330 148.255 ;
      LAYER met4 ;
        RECT 975.560 143.895 1516.240 146.875 ;
      LAYER met4 ;
        RECT 395.670 142.865 467.330 143.495 ;
        RECT 965.310 142.865 1008.990 143.495 ;
      LAYER met4 ;
        RECT 1009.390 143.265 1507.910 143.595 ;
      LAYER met4 ;
        RECT 1516.640 143.495 1518.160 147.275 ;
      LAYER met4 ;
        RECT 1553.730 147.175 1555.000 148.355 ;
      LAYER met4 ;
        RECT 1555.000 147.175 1749.000 148.355 ;
      LAYER met4 ;
        RECT 1749.000 147.175 1750.270 148.355 ;
      LAYER met4 ;
        RECT 1774.935 148.255 1776.455 151.535 ;
      LAYER met4 ;
        RECT 1776.855 148.655 2048.535 151.635 ;
      LAYER met4 ;
        RECT 1750.670 147.275 1827.330 148.255 ;
      LAYER met4 ;
        RECT 1518.560 143.895 1790.240 146.875 ;
      LAYER met4 ;
        RECT 1508.310 142.865 1551.990 143.495 ;
      LAYER met4 ;
        RECT 1552.390 143.265 1781.910 143.595 ;
      LAYER met4 ;
        RECT 1790.640 143.495 1792.160 147.275 ;
      LAYER met4 ;
        RECT 1827.730 147.175 1829.000 148.355 ;
      LAYER met4 ;
        RECT 1829.000 147.175 2023.000 148.355 ;
      LAYER met4 ;
        RECT 2023.000 147.175 2024.270 148.355 ;
      LAYER met4 ;
        RECT 2048.935 148.255 2050.455 151.535 ;
      LAYER met4 ;
        RECT 2050.855 148.655 2322.535 151.635 ;
      LAYER met4 ;
        RECT 2024.670 147.275 2101.330 148.255 ;
      LAYER met4 ;
        RECT 1792.560 143.895 2064.240 146.875 ;
      LAYER met4 ;
        RECT 1782.310 142.865 1825.990 143.495 ;
      LAYER met4 ;
        RECT 1826.390 143.265 2055.910 143.595 ;
      LAYER met4 ;
        RECT 2064.640 143.495 2066.160 147.275 ;
      LAYER met4 ;
        RECT 2101.730 147.175 2103.000 148.355 ;
      LAYER met4 ;
        RECT 2103.000 147.175 2297.000 148.355 ;
      LAYER met4 ;
        RECT 2297.000 147.175 2298.270 148.355 ;
      LAYER met4 ;
        RECT 2322.935 148.255 2324.455 151.535 ;
      LAYER met4 ;
        RECT 2324.855 148.655 2596.535 151.635 ;
      LAYER met4 ;
        RECT 2298.670 147.275 2375.330 148.255 ;
      LAYER met4 ;
        RECT 2066.560 143.895 2338.240 146.875 ;
      LAYER met4 ;
        RECT 2056.310 142.865 2099.990 143.495 ;
      LAYER met4 ;
        RECT 2100.390 143.265 2329.910 143.595 ;
      LAYER met4 ;
        RECT 2338.640 143.495 2340.160 147.275 ;
      LAYER met4 ;
        RECT 2375.730 147.175 2377.000 148.355 ;
      LAYER met4 ;
        RECT 2377.000 147.175 2571.000 148.355 ;
      LAYER met4 ;
        RECT 2571.000 147.175 2572.270 148.355 ;
      LAYER met4 ;
        RECT 2596.935 148.255 2598.455 151.535 ;
      LAYER met4 ;
        RECT 2598.855 148.655 3404.875 151.635 ;
      LAYER met4 ;
        RECT 3407.975 151.535 3588.000 152.665 ;
        RECT 3405.275 148.755 3588.000 151.535 ;
        RECT 2572.670 147.275 2649.330 148.255 ;
      LAYER met4 ;
        RECT 2340.560 143.895 2612.240 146.875 ;
      LAYER met4 ;
        RECT 2330.310 142.865 2373.990 143.495 ;
      LAYER met4 ;
        RECT 2374.390 143.265 2603.910 143.595 ;
      LAYER met4 ;
        RECT 2612.640 143.495 2614.160 147.275 ;
      LAYER met4 ;
        RECT 2649.730 147.175 2651.000 148.355 ;
      LAYER met4 ;
        RECT 2651.000 147.175 2845.000 148.355 ;
      LAYER met4 ;
        RECT 2845.000 147.175 2846.270 148.355 ;
      LAYER met4 ;
        RECT 2846.670 147.275 2918.330 148.255 ;
      LAYER met4 ;
        RECT 2918.730 147.175 2920.000 148.355 ;
      LAYER met4 ;
        RECT 2920.000 147.175 3114.000 148.355 ;
      LAYER met4 ;
        RECT 3114.000 147.175 3115.270 148.355 ;
      LAYER met4 ;
        RECT 3115.670 147.275 3187.330 148.255 ;
      LAYER met4 ;
        RECT 3187.730 147.175 3189.000 148.355 ;
      LAYER met4 ;
        RECT 3189.000 147.175 3384.000 148.355 ;
      LAYER met4 ;
        RECT 3384.000 147.175 3405.555 148.355 ;
      LAYER met4 ;
        RECT 3405.955 147.275 3588.000 148.755 ;
      LAYER met4 ;
        RECT 2614.560 143.895 3410.910 146.875 ;
      LAYER met4 ;
        RECT 3411.310 143.995 3588.000 147.275 ;
        RECT 2604.310 142.865 2647.990 143.495 ;
      LAYER met4 ;
        RECT 2648.390 143.265 3411.175 143.595 ;
      LAYER met4 ;
        RECT 3411.575 142.865 3588.000 143.995 ;
        RECT 0.000 142.165 394.000 142.865 ;
        RECT 394.965 142.165 468.035 142.865 ;
        RECT 469.000 142.165 663.000 142.865 ;
        RECT 663.965 142.165 737.035 142.865 ;
        RECT 738.000 142.165 932.000 142.865 ;
        RECT 933.030 142.165 1011.035 142.865 ;
        RECT 1012.000 142.165 1280.035 142.865 ;
        RECT 1281.000 142.165 1475.000 142.865 ;
        RECT 1476.030 142.165 1554.035 142.865 ;
        RECT 1555.000 142.165 1749.000 142.865 ;
        RECT 1750.030 142.165 1828.035 142.865 ;
        RECT 1829.000 142.165 2023.000 142.865 ;
        RECT 2024.030 142.165 2102.035 142.865 ;
        RECT 2103.000 142.165 2297.000 142.865 ;
        RECT 2298.030 142.165 2376.035 142.865 ;
        RECT 2377.000 142.165 2571.000 142.865 ;
        RECT 2572.030 142.165 2650.035 142.865 ;
        RECT 2651.000 142.165 2845.000 142.865 ;
        RECT 2845.965 142.165 2919.035 142.865 ;
        RECT 2920.000 142.165 3114.000 142.865 ;
        RECT 3114.965 142.165 3188.035 142.865 ;
        RECT 3189.000 142.165 3384.000 142.865 ;
        RECT 3385.255 142.165 3588.000 142.865 ;
        RECT 0.000 136.915 197.975 142.165 ;
      LAYER met4 ;
        RECT 198.375 137.315 395.270 141.765 ;
      LAYER met4 ;
        RECT 395.670 136.915 467.330 142.165 ;
      LAYER met4 ;
        RECT 467.730 137.315 664.270 141.765 ;
      LAYER met4 ;
        RECT 664.670 136.915 736.330 142.165 ;
      LAYER met4 ;
        RECT 736.730 137.315 933.270 141.765 ;
      LAYER met4 ;
        RECT 933.670 136.915 1010.330 142.165 ;
      LAYER met4 ;
        RECT 1010.730 137.315 1207.270 141.765 ;
      LAYER met4 ;
        RECT 1207.670 136.915 1279.330 142.165 ;
      LAYER met4 ;
        RECT 1279.730 137.315 1476.270 141.765 ;
      LAYER met4 ;
        RECT 1476.670 136.915 1553.330 142.165 ;
      LAYER met4 ;
        RECT 1553.730 137.315 1750.270 141.765 ;
      LAYER met4 ;
        RECT 1750.670 136.915 1827.330 142.165 ;
      LAYER met4 ;
        RECT 1827.730 137.315 2024.270 141.765 ;
      LAYER met4 ;
        RECT 2024.670 136.915 2101.330 142.165 ;
      LAYER met4 ;
        RECT 2101.730 137.315 2298.270 141.765 ;
      LAYER met4 ;
        RECT 2298.670 136.915 2375.330 142.165 ;
      LAYER met4 ;
        RECT 2375.730 137.315 2572.270 141.765 ;
      LAYER met4 ;
        RECT 2572.670 136.915 2649.330 142.165 ;
      LAYER met4 ;
        RECT 2649.730 137.315 2846.270 141.765 ;
      LAYER met4 ;
        RECT 2846.670 136.915 2918.330 142.165 ;
      LAYER met4 ;
        RECT 2918.730 137.315 3115.270 141.765 ;
      LAYER met4 ;
        RECT 3115.670 136.915 3187.330 142.165 ;
      LAYER met4 ;
        RECT 3187.730 137.315 3385.270 141.765 ;
      LAYER met4 ;
        RECT 3385.670 136.915 3588.000 142.165 ;
        RECT 0.000 136.315 394.000 136.915 ;
        RECT 394.965 136.315 468.035 136.915 ;
        RECT 469.000 136.315 663.000 136.915 ;
        RECT 663.965 136.315 737.035 136.915 ;
        RECT 738.000 136.315 932.000 136.915 ;
        RECT 933.030 136.315 1011.035 136.915 ;
        RECT 1012.000 136.315 1280.035 136.915 ;
        RECT 1281.000 136.315 1475.000 136.915 ;
        RECT 1476.030 136.315 1554.035 136.915 ;
        RECT 1555.000 136.315 1749.000 136.915 ;
        RECT 1750.030 136.315 1828.035 136.915 ;
        RECT 1829.000 136.315 2023.000 136.915 ;
        RECT 2024.030 136.315 2102.035 136.915 ;
        RECT 2103.000 136.315 2297.000 136.915 ;
        RECT 2298.030 136.315 2376.035 136.915 ;
        RECT 2377.000 136.315 2571.000 136.915 ;
        RECT 2572.030 136.315 2650.035 136.915 ;
        RECT 2651.000 136.315 2845.000 136.915 ;
        RECT 2845.965 136.315 2919.035 136.915 ;
        RECT 2920.000 136.315 3114.000 136.915 ;
        RECT 3114.965 136.315 3188.035 136.915 ;
        RECT 3189.000 136.315 3384.000 136.915 ;
        RECT 3385.255 136.315 3588.000 136.915 ;
        RECT 0.000 131.065 198.120 136.315 ;
      LAYER met4 ;
        RECT 198.520 131.465 395.270 135.915 ;
      LAYER met4 ;
        RECT 395.670 131.065 467.330 136.315 ;
      LAYER met4 ;
        RECT 467.730 131.465 664.270 135.915 ;
      LAYER met4 ;
        RECT 664.670 131.065 736.330 136.315 ;
      LAYER met4 ;
        RECT 736.730 131.465 933.270 135.915 ;
      LAYER met4 ;
        RECT 933.670 131.065 1010.330 136.315 ;
      LAYER met4 ;
        RECT 1010.730 131.465 1207.270 135.915 ;
      LAYER met4 ;
        RECT 1207.670 131.065 1279.330 136.315 ;
      LAYER met4 ;
        RECT 1279.730 131.465 1476.270 135.915 ;
      LAYER met4 ;
        RECT 1476.670 131.065 1553.330 136.315 ;
      LAYER met4 ;
        RECT 1553.730 131.465 1750.270 135.915 ;
      LAYER met4 ;
        RECT 1750.670 131.065 1827.330 136.315 ;
      LAYER met4 ;
        RECT 1827.730 131.465 2024.270 135.915 ;
      LAYER met4 ;
        RECT 2024.670 131.065 2101.330 136.315 ;
      LAYER met4 ;
        RECT 2101.730 131.465 2298.270 135.915 ;
      LAYER met4 ;
        RECT 2298.670 131.065 2375.330 136.315 ;
      LAYER met4 ;
        RECT 2375.730 131.465 2572.270 135.915 ;
      LAYER met4 ;
        RECT 2572.670 131.065 2649.330 136.315 ;
      LAYER met4 ;
        RECT 2649.730 131.465 2846.270 135.915 ;
      LAYER met4 ;
        RECT 2846.670 131.065 2918.330 136.315 ;
      LAYER met4 ;
        RECT 2918.730 131.465 3115.270 135.915 ;
      LAYER met4 ;
        RECT 3115.670 131.065 3187.330 136.315 ;
      LAYER met4 ;
        RECT 3187.730 131.465 3385.270 135.915 ;
      LAYER met4 ;
        RECT 3385.670 131.065 3588.000 136.315 ;
        RECT 0.000 130.365 394.000 131.065 ;
        RECT 394.965 130.365 468.035 131.065 ;
        RECT 469.000 130.365 663.000 131.065 ;
        RECT 663.965 130.365 737.035 131.065 ;
        RECT 738.000 130.365 932.000 131.065 ;
        RECT 933.030 130.365 1011.035 131.065 ;
        RECT 1012.000 130.365 1280.035 131.065 ;
        RECT 1281.000 130.365 1475.000 131.065 ;
        RECT 1476.030 130.365 1554.035 131.065 ;
        RECT 1555.000 130.365 1749.000 131.065 ;
        RECT 1750.030 130.365 1828.035 131.065 ;
        RECT 1829.000 130.365 2023.000 131.065 ;
        RECT 2024.030 130.365 2102.035 131.065 ;
        RECT 2103.000 130.365 2297.000 131.065 ;
        RECT 2298.030 130.365 2376.035 131.065 ;
        RECT 2377.000 130.365 2571.000 131.065 ;
        RECT 2572.030 130.365 2650.035 131.065 ;
        RECT 2651.000 130.365 2845.000 131.065 ;
        RECT 2845.965 130.365 2919.035 131.065 ;
        RECT 2920.000 130.365 3114.000 131.065 ;
        RECT 3114.965 130.365 3188.035 131.065 ;
        RECT 3189.000 130.365 3384.000 131.065 ;
        RECT 3385.255 130.365 3588.000 131.065 ;
        RECT 0.000 104.600 196.955 130.365 ;
      LAYER met4 ;
        RECT 197.355 105.000 395.270 129.965 ;
      LAYER met4 ;
        RECT 395.670 104.600 467.330 130.365 ;
      LAYER met4 ;
        RECT 467.730 105.000 664.270 129.965 ;
      LAYER met4 ;
        RECT 664.670 104.600 736.330 130.365 ;
      LAYER met4 ;
        RECT 736.730 105.000 933.270 129.965 ;
      LAYER met4 ;
        RECT 933.670 104.600 1010.330 130.365 ;
      LAYER met4 ;
        RECT 1010.730 105.000 1207.270 129.965 ;
      LAYER met4 ;
        RECT 1207.670 104.600 1279.330 130.365 ;
      LAYER met4 ;
        RECT 1279.730 105.000 1476.270 129.965 ;
      LAYER met4 ;
        RECT 1476.670 104.600 1553.330 130.365 ;
      LAYER met4 ;
        RECT 1553.730 105.000 1750.270 129.965 ;
      LAYER met4 ;
        RECT 1750.670 104.600 1827.330 130.365 ;
      LAYER met4 ;
        RECT 1827.730 105.000 2024.270 129.965 ;
      LAYER met4 ;
        RECT 2024.670 104.600 2101.330 130.365 ;
      LAYER met4 ;
        RECT 2101.730 105.000 2298.270 129.965 ;
      LAYER met4 ;
        RECT 2298.670 104.600 2375.330 130.365 ;
      LAYER met4 ;
        RECT 2375.730 105.000 2572.270 129.965 ;
      LAYER met4 ;
        RECT 2572.670 104.600 2649.330 130.365 ;
      LAYER met4 ;
        RECT 2649.730 105.000 2846.270 129.965 ;
      LAYER met4 ;
        RECT 2846.670 104.600 2918.330 130.365 ;
      LAYER met4 ;
        RECT 2918.730 105.000 3115.270 129.965 ;
      LAYER met4 ;
        RECT 3115.670 104.600 3187.330 130.365 ;
      LAYER met4 ;
        RECT 3187.730 105.000 3385.855 129.965 ;
      LAYER met4 ;
        RECT 3386.255 104.600 3588.000 130.365 ;
        RECT 0.000 24.615 394.000 104.600 ;
        RECT 394.965 24.615 468.035 104.600 ;
        RECT 0.000 0.000 198.165 24.615 ;
      LAYER met4 ;
        RECT 198.565 0.000 200.000 24.215 ;
      LAYER met4 ;
        RECT 200.000 0.000 394.000 24.615 ;
      LAYER met4 ;
        RECT 394.000 0.000 395.270 24.215 ;
      LAYER met4 ;
        RECT 395.670 0.000 467.330 24.615 ;
      LAYER met4 ;
        RECT 467.730 0.000 469.000 24.215 ;
      LAYER met4 ;
        RECT 469.000 0.000 663.000 104.600 ;
        RECT 663.965 24.615 737.035 104.600 ;
      LAYER met4 ;
        RECT 663.000 0.000 664.270 24.215 ;
      LAYER met4 ;
        RECT 664.670 0.000 736.330 24.615 ;
      LAYER met4 ;
        RECT 736.730 0.000 738.000 24.215 ;
      LAYER met4 ;
        RECT 738.000 0.000 932.000 104.600 ;
        RECT 933.030 24.615 1011.035 104.600 ;
        RECT 1012.000 24.615 1280.035 104.600 ;
      LAYER met4 ;
        RECT 932.000 0.000 933.270 24.215 ;
      LAYER met4 ;
        RECT 933.670 0.000 1010.330 24.615 ;
      LAYER met4 ;
        RECT 1010.730 0.000 1012.000 24.215 ;
      LAYER met4 ;
        RECT 1012.000 0.000 1206.000 24.615 ;
      LAYER met4 ;
        RECT 1206.000 0.000 1207.270 24.215 ;
      LAYER met4 ;
        RECT 1207.670 0.000 1279.330 24.615 ;
      LAYER met4 ;
        RECT 1279.730 0.000 1281.000 24.215 ;
      LAYER met4 ;
        RECT 1281.000 0.000 1475.000 104.600 ;
        RECT 1476.030 24.615 1554.035 104.600 ;
      LAYER met4 ;
        RECT 1475.000 0.000 1476.270 24.215 ;
      LAYER met4 ;
        RECT 1476.670 0.000 1553.330 24.615 ;
      LAYER met4 ;
        RECT 1553.730 0.000 1555.000 24.215 ;
      LAYER met4 ;
        RECT 1555.000 0.000 1749.000 104.600 ;
        RECT 1750.030 24.615 1828.035 104.600 ;
      LAYER met4 ;
        RECT 1749.000 0.000 1750.270 24.215 ;
      LAYER met4 ;
        RECT 1750.670 0.000 1827.330 24.615 ;
      LAYER met4 ;
        RECT 1827.730 0.000 1829.000 24.215 ;
      LAYER met4 ;
        RECT 1829.000 0.000 2023.000 104.600 ;
        RECT 2024.030 24.615 2102.035 104.600 ;
      LAYER met4 ;
        RECT 2023.000 0.000 2024.270 24.215 ;
      LAYER met4 ;
        RECT 2024.670 0.000 2101.330 24.615 ;
      LAYER met4 ;
        RECT 2101.730 0.000 2103.000 24.215 ;
      LAYER met4 ;
        RECT 2103.000 0.000 2297.000 104.600 ;
        RECT 2298.030 24.615 2376.035 104.600 ;
      LAYER met4 ;
        RECT 2297.000 0.000 2298.270 24.215 ;
      LAYER met4 ;
        RECT 2298.670 0.000 2375.330 24.615 ;
      LAYER met4 ;
        RECT 2375.730 0.000 2377.000 24.215 ;
      LAYER met4 ;
        RECT 2377.000 0.000 2571.000 104.600 ;
        RECT 2572.030 24.615 2650.035 104.600 ;
      LAYER met4 ;
        RECT 2571.000 0.000 2572.270 24.215 ;
      LAYER met4 ;
        RECT 2572.670 0.000 2649.330 24.615 ;
      LAYER met4 ;
        RECT 2649.730 0.000 2651.000 24.215 ;
      LAYER met4 ;
        RECT 2651.000 0.000 2845.000 104.600 ;
        RECT 2845.965 24.615 2919.035 104.600 ;
      LAYER met4 ;
        RECT 2845.000 0.000 2846.270 24.215 ;
      LAYER met4 ;
        RECT 2846.670 0.000 2918.330 24.615 ;
      LAYER met4 ;
        RECT 2918.730 0.000 2920.000 24.215 ;
      LAYER met4 ;
        RECT 2920.000 0.000 3114.000 104.600 ;
        RECT 3114.965 24.615 3188.035 104.600 ;
      LAYER met4 ;
        RECT 3114.000 0.000 3115.270 24.215 ;
      LAYER met4 ;
        RECT 3115.670 0.000 3187.330 24.615 ;
      LAYER met4 ;
        RECT 3187.730 0.000 3189.000 24.215 ;
      LAYER met4 ;
        RECT 3189.000 0.000 3384.000 104.600 ;
        RECT 3385.255 24.615 3588.000 104.600 ;
      LAYER met4 ;
        RECT 3384.000 0.000 3385.270 24.215 ;
      LAYER met4 ;
        RECT 3385.670 0.000 3588.000 24.615 ;
      LAYER met5 ;
        RECT 0.000 5084.585 204.000 5188.000 ;
      LAYER met5 ;
        RECT 204.000 5163.785 382.270 5188.000 ;
      LAYER met5 ;
        RECT 383.870 5162.185 453.130 5188.000 ;
      LAYER met5 ;
        RECT 454.730 5163.785 639.270 5188.000 ;
      LAYER met5 ;
        RECT 640.870 5162.185 710.130 5188.000 ;
      LAYER met5 ;
        RECT 711.730 5163.785 896.270 5188.000 ;
      LAYER met5 ;
        RECT 897.870 5162.185 967.130 5188.000 ;
      LAYER met5 ;
        RECT 968.730 5163.785 1105.000 5188.000 ;
      LAYER met5 ;
        RECT 381.000 5155.545 456.000 5162.185 ;
        RECT 381.000 5091.520 386.450 5155.545 ;
        RECT 450.490 5091.520 456.000 5155.545 ;
        RECT 381.000 5084.585 456.000 5091.520 ;
        RECT 638.000 5155.545 713.000 5162.185 ;
        RECT 638.000 5091.520 643.450 5155.545 ;
        RECT 707.490 5091.520 713.000 5155.545 ;
        RECT 638.000 5084.585 713.000 5091.520 ;
        RECT 895.000 5155.545 970.000 5162.185 ;
        RECT 895.000 5091.520 900.450 5155.545 ;
        RECT 964.490 5091.520 970.000 5155.545 ;
        RECT 895.000 5084.585 970.000 5091.520 ;
        RECT 1105.000 5155.545 1274.000 5188.000 ;
      LAYER met5 ;
        RECT 1274.000 5163.785 1363.000 5188.000 ;
      LAYER met5 ;
        RECT 1105.000 5091.520 1157.450 5155.545 ;
        RECT 1221.490 5091.520 1274.000 5155.545 ;
        RECT 1105.000 5084.585 1274.000 5091.520 ;
        RECT 1363.000 5155.545 1532.000 5188.000 ;
      LAYER met5 ;
        RECT 1532.000 5163.785 1667.000 5188.000 ;
      LAYER met5 ;
        RECT 1363.000 5091.520 1415.450 5155.545 ;
        RECT 1479.490 5091.520 1532.000 5155.545 ;
        RECT 1363.000 5084.585 1532.000 5091.520 ;
        RECT 1667.000 5155.545 1742.000 5188.000 ;
      LAYER met5 ;
        RECT 1742.000 5163.785 1920.270 5188.000 ;
      LAYER met5 ;
        RECT 1921.870 5162.185 1991.130 5188.000 ;
      LAYER met5 ;
        RECT 1992.730 5163.785 2365.270 5188.000 ;
      LAYER met5 ;
        RECT 2366.870 5162.185 2436.130 5188.000 ;
      LAYER met5 ;
        RECT 2437.730 5163.785 2622.270 5188.000 ;
      LAYER met5 ;
        RECT 2623.870 5162.185 2693.130 5188.000 ;
      LAYER met5 ;
        RECT 2694.730 5163.785 2878.000 5188.000 ;
      LAYER met5 ;
        RECT 1667.000 5091.520 1672.450 5155.545 ;
        RECT 1736.490 5091.520 1742.000 5155.545 ;
        RECT 1667.000 5084.585 1742.000 5091.520 ;
        RECT 1919.000 5155.545 1994.000 5162.185 ;
        RECT 1919.000 5091.520 1924.450 5155.545 ;
        RECT 1988.490 5091.520 1994.000 5155.545 ;
        RECT 1919.000 5084.585 1994.000 5091.520 ;
        RECT 2364.000 5155.545 2439.000 5162.185 ;
        RECT 2364.000 5091.520 2369.450 5155.545 ;
        RECT 2433.490 5091.520 2439.000 5155.545 ;
        RECT 2364.000 5084.585 2439.000 5091.520 ;
        RECT 2621.000 5155.545 2696.000 5162.185 ;
        RECT 2621.000 5091.520 2626.450 5155.545 ;
        RECT 2690.490 5091.520 2696.000 5155.545 ;
        RECT 2621.000 5084.585 2696.000 5091.520 ;
        RECT 2878.000 5155.545 2953.000 5188.000 ;
      LAYER met5 ;
        RECT 2953.000 5163.785 3131.270 5188.000 ;
      LAYER met5 ;
        RECT 3132.870 5162.185 3202.130 5188.000 ;
      LAYER met5 ;
        RECT 3203.730 5163.785 3388.000 5188.000 ;
      LAYER met5 ;
        RECT 2878.000 5091.520 2883.450 5155.545 ;
        RECT 2947.490 5091.520 2953.000 5155.545 ;
        RECT 2878.000 5084.585 2953.000 5091.520 ;
        RECT 3130.000 5155.545 3205.000 5162.185 ;
        RECT 3130.000 5091.520 3135.450 5155.545 ;
        RECT 3199.490 5091.520 3205.000 5155.545 ;
        RECT 3130.000 5084.585 3205.000 5091.520 ;
        RECT 3388.000 5084.585 3588.000 5188.000 ;
        RECT 0.000 5056.435 200.545 5084.585 ;
      LAYER met5 ;
        RECT 202.145 5058.035 382.270 5082.985 ;
      LAYER met5 ;
        RECT 0.000 5046.335 201.130 5056.435 ;
      LAYER met5 ;
        RECT 202.730 5052.185 382.270 5056.435 ;
        RECT 202.730 5046.335 382.270 5050.585 ;
      LAYER met5 ;
        RECT 0.000 5034.135 175.245 5046.335 ;
      LAYER met5 ;
        RECT 176.845 5035.735 382.270 5044.735 ;
      LAYER met5 ;
        RECT 0.000 5012.755 201.130 5034.135 ;
      LAYER met5 ;
        RECT 202.730 5029.685 382.270 5034.135 ;
        RECT 202.730 5024.840 382.270 5028.085 ;
      LAYER met5 ;
        RECT 383.870 5024.840 453.130 5084.585 ;
      LAYER met5 ;
        RECT 454.730 5058.035 639.270 5082.985 ;
        RECT 454.730 5052.185 639.270 5056.435 ;
        RECT 454.730 5046.335 639.270 5050.585 ;
        RECT 454.730 5035.735 639.270 5044.735 ;
        RECT 454.730 5029.685 639.270 5034.135 ;
        RECT 454.730 5024.840 639.270 5028.085 ;
      LAYER met5 ;
        RECT 640.870 5024.840 710.130 5084.585 ;
      LAYER met5 ;
        RECT 711.730 5058.035 896.270 5082.985 ;
        RECT 711.730 5052.185 896.270 5056.435 ;
        RECT 711.730 5046.335 896.270 5050.585 ;
        RECT 711.730 5035.735 896.270 5044.735 ;
        RECT 711.730 5029.685 896.270 5034.135 ;
        RECT 711.730 5024.840 896.270 5028.085 ;
      LAYER met5 ;
        RECT 897.870 5024.840 967.130 5084.585 ;
      LAYER met5 ;
        RECT 968.730 5058.035 1152.715 5082.985 ;
        RECT 968.730 5052.185 1152.715 5056.435 ;
        RECT 968.730 5046.335 1152.715 5050.585 ;
      LAYER met5 ;
        RECT 1154.315 5044.735 1229.285 5084.585 ;
      LAYER met5 ;
        RECT 1230.885 5058.035 1410.715 5082.985 ;
        RECT 1230.885 5052.185 1410.715 5056.435 ;
        RECT 1230.885 5046.335 1410.715 5050.585 ;
      LAYER met5 ;
        RECT 1412.315 5044.735 1487.285 5084.585 ;
      LAYER met5 ;
        RECT 1488.885 5058.035 1668.270 5082.985 ;
        RECT 1488.885 5052.185 1668.270 5056.435 ;
        RECT 1488.885 5046.335 1668.270 5050.585 ;
        RECT 968.730 5035.735 1152.240 5044.735 ;
      LAYER met5 ;
        RECT 1153.840 5035.735 1229.285 5044.735 ;
      LAYER met5 ;
        RECT 1230.885 5035.735 1410.240 5044.735 ;
      LAYER met5 ;
        RECT 1411.840 5035.735 1487.285 5044.735 ;
      LAYER met5 ;
        RECT 1488.885 5035.735 1668.270 5044.735 ;
        RECT 968.730 5029.685 1152.715 5034.135 ;
        RECT 968.730 5024.840 1152.715 5028.085 ;
        RECT 204.000 5024.835 381.000 5024.840 ;
      LAYER met5 ;
        RECT 381.000 5024.835 456.000 5024.840 ;
      LAYER met5 ;
        RECT 456.000 5024.835 638.000 5024.840 ;
      LAYER met5 ;
        RECT 638.000 5024.835 713.000 5024.840 ;
      LAYER met5 ;
        RECT 713.000 5024.835 895.000 5024.840 ;
      LAYER met5 ;
        RECT 895.000 5024.835 970.000 5024.840 ;
      LAYER met5 ;
        RECT 970.000 5024.835 1152.715 5024.840 ;
        RECT 202.730 5019.985 382.270 5023.235 ;
        RECT 202.730 5013.935 382.270 5018.385 ;
      LAYER met5 ;
        RECT 0.000 4992.245 141.665 5012.755 ;
        RECT 0.000 4988.000 103.415 4992.245 ;
        RECT 131.565 4991.225 141.665 4992.245 ;
        RECT 131.565 4991.080 135.815 4991.225 ;
      LAYER met5 ;
        RECT 0.000 4844.730 24.215 4988.000 ;
      LAYER met5 ;
        RECT 25.815 4843.130 103.415 4846.000 ;
      LAYER met5 ;
        RECT 105.015 4844.730 129.965 4990.645 ;
        RECT 131.565 4844.730 135.815 4989.480 ;
        RECT 137.415 4844.730 141.665 4989.625 ;
        RECT 143.265 4844.730 152.265 5011.155 ;
      LAYER met5 ;
        RECT 153.865 5006.285 201.130 5012.755 ;
      LAYER met5 ;
        RECT 202.730 5007.885 382.270 5012.335 ;
      LAYER met5 ;
        RECT 383.870 5006.285 453.130 5024.835 ;
      LAYER met5 ;
        RECT 454.730 5019.985 639.270 5023.235 ;
        RECT 454.730 5013.935 639.270 5018.385 ;
        RECT 454.730 5007.885 639.270 5012.335 ;
      LAYER met5 ;
        RECT 640.870 5006.285 710.130 5024.835 ;
      LAYER met5 ;
        RECT 711.730 5019.985 896.270 5023.235 ;
        RECT 711.730 5013.935 896.270 5018.385 ;
        RECT 711.730 5007.885 896.270 5012.335 ;
      LAYER met5 ;
        RECT 897.870 5006.285 967.130 5024.835 ;
      LAYER met5 ;
        RECT 968.730 5019.985 1152.715 5023.235 ;
        RECT 968.730 5013.935 1152.715 5018.385 ;
        RECT 968.730 5007.885 1152.715 5012.335 ;
      LAYER met5 ;
        RECT 1154.315 5007.885 1229.285 5035.735 ;
      LAYER met5 ;
        RECT 1230.885 5029.685 1410.715 5034.135 ;
        RECT 1230.885 5024.835 1410.715 5028.085 ;
        RECT 1230.885 5019.985 1410.715 5023.235 ;
        RECT 1230.885 5013.935 1410.715 5018.385 ;
        RECT 1230.885 5007.885 1410.715 5012.335 ;
      LAYER met5 ;
        RECT 1412.315 5007.885 1487.285 5035.735 ;
      LAYER met5 ;
        RECT 1488.885 5029.685 1668.270 5034.135 ;
        RECT 1488.885 5024.840 1668.270 5028.085 ;
      LAYER met5 ;
        RECT 1669.870 5024.840 1739.130 5084.585 ;
      LAYER met5 ;
        RECT 1740.730 5058.035 1920.270 5082.985 ;
        RECT 1740.730 5052.185 1920.270 5056.435 ;
        RECT 1740.730 5046.335 1920.270 5050.585 ;
        RECT 1740.730 5035.735 1909.000 5044.735 ;
        RECT 1914.000 5035.735 1920.270 5044.735 ;
        RECT 1740.730 5029.685 1914.000 5034.135 ;
        RECT 1919.000 5029.685 1920.270 5034.135 ;
        RECT 1740.730 5024.840 1909.000 5028.085 ;
        RECT 1488.885 5024.835 1667.000 5024.840 ;
      LAYER met5 ;
        RECT 1667.000 5024.835 1742.000 5024.840 ;
      LAYER met5 ;
        RECT 1742.000 5024.835 1909.000 5024.840 ;
        RECT 1914.000 5024.840 1920.270 5028.085 ;
      LAYER met5 ;
        RECT 1921.870 5024.840 1991.130 5084.585 ;
      LAYER met5 ;
        RECT 1992.730 5058.035 2365.270 5082.985 ;
        RECT 1992.730 5052.185 2365.270 5056.435 ;
        RECT 1992.730 5046.335 2365.270 5050.585 ;
        RECT 1992.730 5035.735 2365.270 5044.735 ;
        RECT 1992.730 5029.685 2365.270 5034.135 ;
        RECT 1992.730 5024.840 2365.270 5028.085 ;
      LAYER met5 ;
        RECT 2366.870 5024.840 2436.130 5084.585 ;
      LAYER met5 ;
        RECT 2437.730 5058.035 2622.270 5082.985 ;
        RECT 2437.730 5052.185 2622.270 5056.435 ;
        RECT 2437.730 5046.335 2622.270 5050.585 ;
        RECT 2437.730 5035.735 2622.270 5044.735 ;
        RECT 2437.730 5029.685 2622.270 5034.135 ;
        RECT 2437.730 5024.840 2622.270 5028.085 ;
      LAYER met5 ;
        RECT 2623.870 5024.840 2693.130 5084.585 ;
      LAYER met5 ;
        RECT 2694.730 5058.035 2879.270 5082.985 ;
        RECT 2694.730 5052.185 2879.270 5056.435 ;
        RECT 2694.730 5046.335 2879.270 5050.585 ;
        RECT 2694.730 5035.735 2879.270 5044.735 ;
        RECT 2694.730 5029.685 2879.270 5034.135 ;
        RECT 2694.730 5024.840 2879.270 5028.085 ;
      LAYER met5 ;
        RECT 2880.870 5024.840 2950.130 5084.585 ;
      LAYER met5 ;
        RECT 2951.730 5058.035 3131.270 5082.985 ;
        RECT 2951.730 5052.185 3131.270 5056.435 ;
        RECT 2951.730 5046.335 3131.270 5050.585 ;
        RECT 2951.730 5035.735 3131.270 5044.735 ;
        RECT 2951.730 5029.685 3131.270 5034.135 ;
        RECT 2951.730 5024.840 3131.270 5028.085 ;
      LAYER met5 ;
        RECT 3132.870 5024.840 3202.130 5084.585 ;
      LAYER met5 ;
        RECT 3203.730 5058.035 3390.645 5082.985 ;
      LAYER met5 ;
        RECT 3392.245 5056.435 3588.000 5084.585 ;
      LAYER met5 ;
        RECT 3203.730 5052.185 3389.480 5056.435 ;
      LAYER met5 ;
        RECT 3391.080 5052.185 3588.000 5056.435 ;
      LAYER met5 ;
        RECT 3203.730 5046.335 3389.625 5050.585 ;
      LAYER met5 ;
        RECT 3391.225 5046.335 3588.000 5052.185 ;
      LAYER met5 ;
        RECT 3203.730 5035.735 3411.155 5044.735 ;
      LAYER met5 ;
        RECT 3412.755 5034.135 3588.000 5046.335 ;
      LAYER met5 ;
        RECT 3203.730 5029.685 3389.475 5034.135 ;
      LAYER met5 ;
        RECT 3391.075 5028.085 3588.000 5034.135 ;
      LAYER met5 ;
        RECT 3203.730 5024.840 3389.335 5028.085 ;
        RECT 1914.000 5024.835 1919.000 5024.840 ;
      LAYER met5 ;
        RECT 1919.000 5024.835 1994.000 5024.840 ;
      LAYER met5 ;
        RECT 1994.000 5024.835 2364.000 5024.840 ;
      LAYER met5 ;
        RECT 2364.000 5024.835 2439.000 5024.840 ;
      LAYER met5 ;
        RECT 2439.000 5024.835 2621.000 5024.840 ;
      LAYER met5 ;
        RECT 2621.000 5024.835 2696.000 5024.840 ;
      LAYER met5 ;
        RECT 2696.000 5024.835 2878.000 5024.840 ;
      LAYER met5 ;
        RECT 2878.000 5024.835 2953.000 5024.840 ;
      LAYER met5 ;
        RECT 2953.000 5024.835 3130.000 5024.840 ;
      LAYER met5 ;
        RECT 3130.000 5024.835 3205.000 5024.840 ;
      LAYER met5 ;
        RECT 3205.000 5024.835 3389.335 5024.840 ;
      LAYER met5 ;
        RECT 3390.935 5024.835 3588.000 5028.085 ;
      LAYER met5 ;
        RECT 1488.885 5019.985 1668.270 5023.235 ;
        RECT 1488.885 5013.935 1668.270 5018.385 ;
        RECT 1488.885 5007.885 1668.270 5012.335 ;
      LAYER met5 ;
        RECT 153.865 5003.035 201.145 5006.285 ;
      LAYER met5 ;
        RECT 202.745 5003.035 381.965 5006.285 ;
      LAYER met5 ;
        RECT 383.565 5003.035 453.435 5006.285 ;
      LAYER met5 ;
        RECT 455.035 5003.035 638.965 5006.285 ;
      LAYER met5 ;
        RECT 640.565 5003.035 710.435 5006.285 ;
      LAYER met5 ;
        RECT 712.035 5003.035 895.965 5006.285 ;
      LAYER met5 ;
        RECT 897.565 5003.035 967.435 5006.285 ;
      LAYER met5 ;
        RECT 969.035 5003.035 1152.715 5006.285 ;
      LAYER met5 ;
        RECT 153.865 4993.385 201.130 5003.035 ;
      LAYER met5 ;
        RECT 202.730 4996.985 382.270 5001.435 ;
      LAYER met5 ;
        RECT 153.865 4991.200 184.965 4993.385 ;
        RECT 192.615 4991.950 201.130 4993.385 ;
        RECT 153.865 4991.075 168.015 4991.200 ;
        RECT 175.665 4991.125 184.965 4991.200 ;
        RECT 159.915 4990.985 168.015 4991.075 ;
        RECT 181.715 4991.070 184.965 4991.125 ;
        RECT 159.915 4990.935 163.165 4990.985 ;
      LAYER met5 ;
        RECT 153.865 4844.730 158.315 4989.475 ;
        RECT 159.915 4846.000 163.165 4989.335 ;
        RECT 159.915 4844.730 163.160 4846.000 ;
      LAYER met5 ;
        RECT 163.160 4843.130 163.165 4846.000 ;
      LAYER met5 ;
        RECT 164.765 4844.730 168.015 4989.385 ;
        RECT 169.615 4844.730 174.065 4989.600 ;
        RECT 175.665 4844.730 180.115 4989.525 ;
        RECT 181.715 4845.035 184.965 4989.470 ;
        RECT 186.565 4844.730 191.015 4991.785 ;
        RECT 192.615 4844.730 197.865 4990.350 ;
      LAYER met5 ;
        RECT 199.465 4988.535 201.130 4991.950 ;
      LAYER met5 ;
        RECT 202.730 4990.135 382.270 4995.385 ;
      LAYER met5 ;
        RECT 383.870 4990.135 453.130 5003.035 ;
      LAYER met5 ;
        RECT 454.730 4996.985 639.270 5001.435 ;
        RECT 454.730 4990.135 639.270 4995.385 ;
      LAYER met5 ;
        RECT 640.870 4990.135 710.130 5003.035 ;
      LAYER met5 ;
        RECT 711.730 4996.985 896.270 5001.435 ;
        RECT 711.730 4990.135 896.270 4995.385 ;
      LAYER met5 ;
        RECT 897.870 4990.135 967.130 5003.035 ;
        RECT 1154.315 5001.435 1224.605 5007.885 ;
      LAYER met5 ;
        RECT 1226.205 5003.035 1410.715 5006.285 ;
      LAYER met5 ;
        RECT 1412.315 5001.435 1482.605 5007.885 ;
        RECT 1669.870 5006.285 1739.130 5024.835 ;
      LAYER met5 ;
        RECT 1740.730 5019.985 1920.270 5023.235 ;
        RECT 1740.730 5013.935 1920.270 5018.385 ;
        RECT 1740.730 5007.885 1920.270 5012.335 ;
      LAYER met5 ;
        RECT 1921.870 5006.285 1991.130 5024.835 ;
      LAYER met5 ;
        RECT 1992.730 5019.985 2365.270 5023.235 ;
        RECT 1992.730 5013.935 2365.270 5018.385 ;
        RECT 1992.730 5007.885 2365.270 5012.335 ;
      LAYER met5 ;
        RECT 2366.870 5006.285 2436.130 5024.835 ;
      LAYER met5 ;
        RECT 2437.730 5019.985 2622.270 5023.235 ;
        RECT 2437.730 5013.935 2622.270 5018.385 ;
        RECT 2437.730 5007.885 2622.270 5012.335 ;
      LAYER met5 ;
        RECT 2623.870 5006.285 2693.130 5024.835 ;
      LAYER met5 ;
        RECT 2694.730 5019.985 2879.270 5023.235 ;
        RECT 2694.730 5013.935 2879.270 5018.385 ;
        RECT 2694.730 5007.885 2879.270 5012.335 ;
      LAYER met5 ;
        RECT 2880.870 5006.285 2950.130 5024.835 ;
      LAYER met5 ;
        RECT 2951.730 5019.985 3131.270 5023.235 ;
        RECT 2951.730 5013.935 3131.270 5018.385 ;
        RECT 2951.730 5007.885 3131.270 5012.335 ;
      LAYER met5 ;
        RECT 3132.870 5006.285 3202.130 5024.835 ;
      LAYER met5 ;
        RECT 3203.730 5019.985 3389.385 5023.235 ;
      LAYER met5 ;
        RECT 3390.985 5019.985 3588.000 5024.835 ;
      LAYER met5 ;
        RECT 3203.730 5013.935 3389.600 5018.385 ;
      LAYER met5 ;
        RECT 3391.200 5012.755 3588.000 5019.985 ;
        RECT 3391.200 5012.335 3434.135 5012.755 ;
      LAYER met5 ;
        RECT 3203.730 5007.885 3389.525 5012.335 ;
      LAYER met5 ;
        RECT 3391.125 5006.285 3434.135 5012.335 ;
      LAYER met5 ;
        RECT 1484.205 5003.035 1667.965 5006.285 ;
      LAYER met5 ;
        RECT 1669.565 5003.035 1739.435 5006.285 ;
      LAYER met5 ;
        RECT 1741.035 5003.035 1909.000 5006.285 ;
        RECT 1914.000 5003.035 1919.965 5006.285 ;
      LAYER met5 ;
        RECT 1921.565 5003.035 1991.435 5006.285 ;
      LAYER met5 ;
        RECT 1993.035 5003.035 2364.965 5006.285 ;
      LAYER met5 ;
        RECT 2366.565 5003.035 2436.435 5006.285 ;
      LAYER met5 ;
        RECT 2438.035 5003.035 2621.965 5006.285 ;
      LAYER met5 ;
        RECT 2623.565 5003.035 2693.435 5006.285 ;
      LAYER met5 ;
        RECT 2695.035 5003.035 2878.965 5006.285 ;
      LAYER met5 ;
        RECT 2880.565 5003.035 2950.435 5006.285 ;
      LAYER met5 ;
        RECT 2952.035 5003.035 3130.965 5006.285 ;
      LAYER met5 ;
        RECT 3132.565 5003.035 3202.435 5006.285 ;
      LAYER met5 ;
        RECT 3204.035 5003.035 3389.470 5006.285 ;
      LAYER met5 ;
        RECT 3391.070 5003.035 3434.135 5006.285 ;
      LAYER met5 ;
        RECT 968.730 4996.985 1152.715 5001.435 ;
        RECT 968.730 4990.135 1152.715 4995.385 ;
      LAYER met5 ;
        RECT 1154.315 4990.135 1229.285 5001.435 ;
      LAYER met5 ;
        RECT 1230.885 4996.985 1410.715 5001.435 ;
        RECT 1230.885 4990.135 1410.715 4995.385 ;
      LAYER met5 ;
        RECT 1412.315 4990.135 1487.285 5001.435 ;
      LAYER met5 ;
        RECT 1488.885 4996.985 1668.270 5001.435 ;
        RECT 1488.885 4990.135 1668.270 4995.385 ;
      LAYER met5 ;
        RECT 1669.870 4990.135 1739.130 5003.035 ;
      LAYER met5 ;
        RECT 1740.730 4996.985 1914.000 5001.435 ;
        RECT 1919.000 4996.985 1920.270 5001.435 ;
        RECT 1740.730 4990.135 1920.270 4995.385 ;
      LAYER met5 ;
        RECT 1921.870 4990.135 1991.130 5003.035 ;
      LAYER met5 ;
        RECT 1992.730 4996.985 2365.270 5001.435 ;
        RECT 1992.730 4990.135 2365.270 4995.385 ;
      LAYER met5 ;
        RECT 2366.870 4990.135 2436.130 5003.035 ;
      LAYER met5 ;
        RECT 2437.730 4996.985 2622.270 5001.435 ;
        RECT 2437.730 4990.135 2622.270 4995.385 ;
      LAYER met5 ;
        RECT 2623.870 4990.135 2693.130 5003.035 ;
      LAYER met5 ;
        RECT 2694.730 4996.985 2879.270 5001.435 ;
        RECT 2694.730 4990.135 2879.270 4995.385 ;
      LAYER met5 ;
        RECT 2880.870 4990.135 2950.130 5003.035 ;
      LAYER met5 ;
        RECT 2951.730 4996.985 3131.270 5001.435 ;
        RECT 2951.730 4990.135 3131.270 4995.385 ;
      LAYER met5 ;
        RECT 3132.870 4990.135 3202.130 5003.035 ;
      LAYER met5 ;
        RECT 3203.730 4996.985 3391.785 5001.435 ;
      LAYER met5 ;
        RECT 3393.385 4995.385 3434.135 5003.035 ;
      LAYER met5 ;
        RECT 3203.730 4990.135 3390.350 4995.385 ;
      LAYER met5 ;
        RECT 3391.950 4988.535 3434.135 4995.385 ;
        RECT 199.465 4988.000 204.000 4988.535 ;
        RECT 3388.000 4986.870 3434.135 4988.535 ;
        RECT 3388.000 4984.000 3388.535 4986.870 ;
        RECT 3403.035 4986.855 3406.285 4986.870 ;
        RECT 181.715 4843.130 184.965 4843.435 ;
        RECT 0.000 4840.490 197.865 4843.130 ;
        RECT 0.000 4776.450 32.455 4840.490 ;
        RECT 96.480 4776.450 197.865 4840.490 ;
      LAYER met5 ;
        RECT 3390.135 4837.285 3395.385 4985.270 ;
        RECT 3396.985 4837.285 3401.435 4985.270 ;
        RECT 3403.035 4837.285 3406.285 4985.255 ;
        RECT 3407.885 4837.285 3412.335 4985.270 ;
        RECT 3413.935 4837.285 3418.385 4985.270 ;
        RECT 3419.985 4837.285 3423.235 4985.270 ;
        RECT 3424.840 4984.000 3428.085 4985.270 ;
        RECT 3424.835 4837.285 3428.085 4984.000 ;
        RECT 3429.685 4837.285 3434.135 4985.270 ;
        RECT 3435.735 4837.760 3444.735 5011.155 ;
      LAYER met5 ;
        RECT 3446.335 4987.455 3588.000 5012.755 ;
        RECT 3446.335 4986.870 3456.435 4987.455 ;
      LAYER met5 ;
        RECT 3446.335 4837.285 3450.585 4985.270 ;
        RECT 3452.185 4837.285 3456.435 4985.270 ;
        RECT 3458.035 4837.285 3482.985 4985.855 ;
      LAYER met5 ;
        RECT 3484.585 4984.000 3588.000 4987.455 ;
      LAYER met5 ;
        RECT 3563.785 4885.000 3588.000 4984.000 ;
      LAYER met5 ;
        RECT 3435.735 4835.685 3444.735 4836.160 ;
        RECT 3484.585 4835.685 3588.000 4885.000 ;
        RECT 0.000 4773.870 197.865 4776.450 ;
        RECT 3390.135 4832.550 3588.000 4835.685 ;
      LAYER met5 ;
        RECT 0.000 4635.000 24.215 4772.270 ;
      LAYER met5 ;
        RECT 25.815 4771.000 103.415 4773.870 ;
        RECT 0.000 4632.130 103.415 4635.000 ;
      LAYER met5 ;
        RECT 105.015 4633.730 129.965 4772.270 ;
        RECT 131.565 4633.730 135.815 4772.270 ;
        RECT 137.415 4633.730 141.665 4772.270 ;
        RECT 143.265 4633.730 152.265 4772.270 ;
        RECT 153.865 4633.730 158.315 4772.270 ;
        RECT 159.915 4771.000 163.160 4772.270 ;
      LAYER met5 ;
        RECT 163.160 4771.000 163.165 4773.870 ;
        RECT 181.715 4773.565 184.965 4773.870 ;
      LAYER met5 ;
        RECT 159.915 4635.000 163.165 4771.000 ;
        RECT 159.915 4633.730 163.160 4635.000 ;
        RECT 164.765 4633.730 168.015 4772.270 ;
        RECT 169.615 4633.730 174.065 4772.270 ;
        RECT 175.665 4633.730 180.115 4772.270 ;
        RECT 181.715 4634.035 184.965 4771.965 ;
        RECT 186.565 4633.730 191.015 4772.270 ;
        RECT 192.615 4633.730 197.865 4772.270 ;
      LAYER met5 ;
        RECT 3390.135 4768.510 3491.520 4832.550 ;
        RECT 3555.545 4768.510 3588.000 4832.550 ;
        RECT 3390.135 4765.395 3588.000 4768.510 ;
        RECT 3390.135 4760.715 3401.435 4765.395 ;
        RECT 181.715 4632.130 184.965 4632.435 ;
        RECT 0.000 4626.270 197.865 4632.130 ;
        RECT 0.000 4568.670 29.235 4626.270 ;
        RECT 99.700 4568.670 197.865 4626.270 ;
      LAYER met5 ;
        RECT 3390.135 4611.730 3395.385 4759.115 ;
        RECT 3396.985 4611.730 3401.435 4759.115 ;
        RECT 3403.035 4612.035 3406.285 4763.795 ;
      LAYER met5 ;
        RECT 3407.885 4760.715 3588.000 4765.395 ;
      LAYER met5 ;
        RECT 3407.885 4611.730 3412.335 4759.115 ;
        RECT 3413.935 4611.730 3418.385 4759.115 ;
        RECT 3419.985 4611.730 3423.235 4759.115 ;
        RECT 3424.835 4613.000 3428.085 4759.115 ;
        RECT 3424.840 4611.730 3428.085 4613.000 ;
        RECT 3429.685 4611.730 3434.135 4759.115 ;
        RECT 3435.735 4611.730 3444.735 4759.115 ;
        RECT 3446.335 4611.730 3450.585 4759.115 ;
        RECT 3452.185 4611.730 3456.435 4759.115 ;
        RECT 3458.035 4611.730 3482.985 4759.115 ;
      LAYER met5 ;
        RECT 3484.585 4716.000 3588.000 4760.715 ;
      LAYER met5 ;
        RECT 3563.785 4613.000 3588.000 4716.000 ;
      LAYER met5 ;
        RECT 3403.035 4610.130 3406.285 4610.435 ;
        RECT 3484.585 4610.130 3588.000 4613.000 ;
        RECT 0.000 4562.870 197.865 4568.670 ;
        RECT 3390.135 4604.330 3588.000 4610.130 ;
        RECT 0.000 4560.000 103.415 4562.870 ;
        RECT 181.715 4562.565 184.965 4562.870 ;
      LAYER met5 ;
        RECT 0.000 4424.000 24.215 4560.000 ;
      LAYER met5 ;
        RECT 0.000 4421.130 103.415 4424.000 ;
      LAYER met5 ;
        RECT 105.015 4422.730 129.965 4561.270 ;
        RECT 131.565 4422.730 135.815 4561.270 ;
        RECT 137.415 4422.730 141.665 4561.270 ;
        RECT 143.265 4422.730 152.265 4561.270 ;
        RECT 153.865 4422.730 158.315 4561.270 ;
        RECT 159.915 4560.000 163.160 4561.270 ;
        RECT 159.915 4424.000 163.165 4560.000 ;
        RECT 159.915 4422.730 163.160 4424.000 ;
      LAYER met5 ;
        RECT 163.160 4421.130 163.165 4424.000 ;
      LAYER met5 ;
        RECT 164.765 4422.730 168.015 4561.270 ;
        RECT 169.615 4422.730 174.065 4561.270 ;
        RECT 175.665 4422.730 180.115 4561.270 ;
        RECT 181.715 4423.035 184.965 4560.965 ;
        RECT 186.565 4422.730 191.015 4561.270 ;
        RECT 192.615 4422.730 197.865 4561.270 ;
      LAYER met5 ;
        RECT 3390.135 4546.730 3488.300 4604.330 ;
        RECT 3558.765 4546.730 3588.000 4604.330 ;
        RECT 3390.135 4540.870 3588.000 4546.730 ;
        RECT 3403.035 4540.565 3406.285 4540.870 ;
        RECT 181.715 4421.130 184.965 4421.435 ;
        RECT 0.000 4418.490 197.865 4421.130 ;
        RECT 0.000 4354.450 32.455 4418.490 ;
        RECT 96.480 4354.450 197.865 4418.490 ;
      LAYER met5 ;
        RECT 3390.135 4390.730 3395.385 4539.270 ;
        RECT 3396.985 4390.730 3401.435 4539.270 ;
        RECT 3403.035 4391.035 3406.285 4538.965 ;
        RECT 3407.885 4390.730 3412.335 4539.270 ;
        RECT 3413.935 4390.730 3418.385 4539.270 ;
        RECT 3419.985 4390.730 3423.235 4539.270 ;
        RECT 3424.840 4538.000 3428.085 4539.270 ;
        RECT 3424.835 4392.000 3428.085 4538.000 ;
        RECT 3424.840 4390.730 3428.085 4392.000 ;
        RECT 3429.685 4390.730 3434.135 4539.270 ;
        RECT 3435.735 4390.730 3444.735 4539.270 ;
        RECT 3446.335 4390.730 3450.585 4539.270 ;
        RECT 3452.185 4390.730 3456.435 4539.270 ;
        RECT 3458.035 4390.730 3482.985 4539.270 ;
      LAYER met5 ;
        RECT 3484.585 4538.000 3588.000 4540.870 ;
      LAYER met5 ;
        RECT 3563.785 4392.000 3588.000 4538.000 ;
      LAYER met5 ;
        RECT 3403.035 4389.130 3406.285 4389.435 ;
        RECT 3484.585 4389.130 3588.000 4392.000 ;
        RECT 0.000 4351.870 197.865 4354.450 ;
        RECT 3390.135 4382.500 3588.000 4389.130 ;
        RECT 0.000 4349.000 103.415 4351.870 ;
      LAYER met5 ;
        RECT 0.000 4213.000 24.215 4349.000 ;
      LAYER met5 ;
        RECT 0.000 4210.130 103.415 4213.000 ;
      LAYER met5 ;
        RECT 105.015 4211.730 129.965 4350.270 ;
        RECT 131.565 4211.730 135.815 4350.270 ;
        RECT 137.415 4211.730 141.665 4350.270 ;
        RECT 143.265 4211.730 152.265 4350.270 ;
        RECT 153.865 4211.730 158.315 4350.270 ;
        RECT 159.915 4349.000 163.160 4350.270 ;
      LAYER met5 ;
        RECT 163.160 4349.000 163.165 4351.870 ;
        RECT 181.715 4351.565 184.965 4351.870 ;
      LAYER met5 ;
        RECT 159.915 4213.000 163.165 4349.000 ;
        RECT 159.915 4211.730 163.160 4213.000 ;
      LAYER met5 ;
        RECT 163.160 4210.130 163.165 4213.000 ;
      LAYER met5 ;
        RECT 164.765 4211.730 168.015 4350.270 ;
        RECT 169.615 4211.730 174.065 4350.270 ;
        RECT 175.665 4211.730 180.115 4350.270 ;
        RECT 181.715 4212.035 184.965 4349.965 ;
        RECT 186.565 4211.730 191.015 4350.270 ;
        RECT 192.615 4211.730 197.865 4350.270 ;
      LAYER met5 ;
        RECT 3390.135 4316.600 3490.960 4382.500 ;
        RECT 3556.610 4316.600 3588.000 4382.500 ;
        RECT 3390.135 4314.870 3588.000 4316.600 ;
        RECT 3403.035 4314.630 3406.285 4314.870 ;
        RECT 181.715 4210.130 184.965 4210.435 ;
        RECT 0.000 4207.490 197.865 4210.130 ;
        RECT 0.000 4143.450 32.455 4207.490 ;
        RECT 96.480 4143.450 197.865 4207.490 ;
      LAYER met5 ;
        RECT 3390.135 4165.730 3395.385 4313.270 ;
        RECT 3396.985 4165.730 3401.435 4313.270 ;
        RECT 3403.035 4166.035 3406.285 4313.030 ;
        RECT 3407.885 4165.730 3412.335 4313.270 ;
        RECT 3413.935 4165.730 3418.385 4313.270 ;
        RECT 3419.985 4165.730 3423.235 4313.270 ;
        RECT 3424.840 4312.000 3428.085 4313.270 ;
        RECT 3424.835 4167.000 3428.085 4312.000 ;
      LAYER met5 ;
        RECT 3403.035 4164.130 3406.285 4164.435 ;
        RECT 3424.835 4164.130 3424.840 4167.000 ;
      LAYER met5 ;
        RECT 3424.840 4165.730 3428.085 4167.000 ;
        RECT 3429.685 4165.730 3434.135 4313.270 ;
        RECT 3435.735 4165.730 3444.735 4313.270 ;
        RECT 3446.335 4165.730 3450.585 4313.270 ;
        RECT 3452.185 4165.730 3456.435 4313.270 ;
        RECT 3458.035 4165.730 3482.985 4313.270 ;
      LAYER met5 ;
        RECT 3484.585 4312.000 3588.000 4314.870 ;
      LAYER met5 ;
        RECT 3563.785 4167.000 3588.000 4312.000 ;
      LAYER met5 ;
        RECT 3484.585 4164.130 3588.000 4167.000 ;
        RECT 0.000 4140.870 197.865 4143.450 ;
        RECT 3390.135 4161.550 3588.000 4164.130 ;
        RECT 0.000 4138.000 103.415 4140.870 ;
      LAYER met5 ;
        RECT 0.000 4002.000 24.215 4138.000 ;
      LAYER met5 ;
        RECT 0.000 3999.130 103.415 4002.000 ;
      LAYER met5 ;
        RECT 105.015 4000.730 129.965 4139.270 ;
        RECT 131.565 4000.730 135.815 4139.270 ;
        RECT 137.415 4000.730 141.665 4139.270 ;
        RECT 143.265 4000.730 152.265 4139.270 ;
        RECT 153.865 4000.730 158.315 4139.270 ;
        RECT 159.915 4138.000 163.160 4139.270 ;
      LAYER met5 ;
        RECT 163.160 4138.000 163.165 4140.870 ;
        RECT 181.715 4140.565 184.965 4140.870 ;
      LAYER met5 ;
        RECT 159.915 4002.000 163.165 4138.000 ;
        RECT 159.915 4000.730 163.160 4002.000 ;
        RECT 164.765 4000.730 168.015 4139.270 ;
        RECT 169.615 4000.730 174.065 4139.270 ;
        RECT 175.665 4000.730 180.115 4139.270 ;
        RECT 181.715 4000.970 184.965 4138.965 ;
        RECT 186.565 4000.730 191.015 4139.270 ;
        RECT 192.615 4000.730 197.865 4139.270 ;
      LAYER met5 ;
        RECT 3390.135 4097.510 3491.520 4161.550 ;
        RECT 3555.545 4097.510 3588.000 4161.550 ;
        RECT 3390.135 4094.870 3588.000 4097.510 ;
        RECT 3403.035 4094.565 3406.285 4094.870 ;
        RECT 181.715 3999.130 184.965 3999.370 ;
        RECT 0.000 3997.400 197.865 3999.130 ;
        RECT 0.000 3931.500 31.390 3997.400 ;
        RECT 97.040 3931.500 197.865 3997.400 ;
      LAYER met5 ;
        RECT 3390.135 3944.730 3395.385 4093.270 ;
        RECT 3396.985 3944.730 3401.435 4093.270 ;
        RECT 3403.035 3945.035 3406.285 4092.965 ;
        RECT 3407.885 3944.730 3412.335 4093.270 ;
        RECT 3413.935 3944.730 3418.385 4093.270 ;
        RECT 3419.985 3944.730 3423.235 4093.270 ;
      LAYER met5 ;
        RECT 3424.835 4092.000 3424.840 4094.870 ;
      LAYER met5 ;
        RECT 3424.840 4092.000 3428.085 4093.270 ;
        RECT 3424.835 3946.000 3428.085 4092.000 ;
        RECT 3424.840 3944.730 3428.085 3946.000 ;
        RECT 3429.685 3944.730 3434.135 4093.270 ;
        RECT 3435.735 3944.730 3444.735 4093.270 ;
        RECT 3446.335 3944.730 3450.585 4093.270 ;
        RECT 3452.185 3944.730 3456.435 4093.270 ;
        RECT 3458.035 3944.730 3482.985 4093.270 ;
      LAYER met5 ;
        RECT 3484.585 4092.000 3588.000 4094.870 ;
      LAYER met5 ;
        RECT 3563.785 3946.000 3588.000 4092.000 ;
      LAYER met5 ;
        RECT 3403.035 3943.130 3406.285 3943.435 ;
        RECT 3484.585 3943.130 3588.000 3946.000 ;
        RECT 0.000 3924.870 197.865 3931.500 ;
        RECT 3390.135 3936.500 3588.000 3943.130 ;
        RECT 0.000 3922.000 103.415 3924.870 ;
        RECT 181.715 3924.565 184.965 3924.870 ;
      LAYER met5 ;
        RECT 0.000 3786.000 24.215 3922.000 ;
      LAYER met5 ;
        RECT 0.000 3783.130 103.415 3786.000 ;
      LAYER met5 ;
        RECT 105.015 3784.730 129.965 3923.270 ;
        RECT 131.565 3784.730 135.815 3923.270 ;
        RECT 137.415 3784.730 141.665 3923.270 ;
        RECT 143.265 3784.730 152.265 3923.270 ;
        RECT 153.865 3784.730 158.315 3923.270 ;
        RECT 159.915 3922.000 163.160 3923.270 ;
        RECT 159.915 3786.000 163.165 3922.000 ;
        RECT 159.915 3784.730 163.160 3786.000 ;
        RECT 164.765 3784.730 168.015 3923.270 ;
        RECT 169.615 3784.730 174.065 3923.270 ;
        RECT 175.665 3784.730 180.115 3923.270 ;
        RECT 181.715 3784.970 184.965 3922.965 ;
        RECT 186.565 3784.730 191.015 3923.270 ;
        RECT 192.615 3784.730 197.865 3923.270 ;
      LAYER met5 ;
        RECT 3390.135 3870.600 3490.960 3936.500 ;
        RECT 3556.610 3870.600 3588.000 3936.500 ;
        RECT 3390.135 3868.870 3588.000 3870.600 ;
        RECT 3403.035 3868.630 3406.285 3868.870 ;
        RECT 181.715 3783.130 184.965 3783.370 ;
        RECT 0.000 3781.400 197.865 3783.130 ;
        RECT 0.000 3715.500 31.390 3781.400 ;
        RECT 97.040 3715.500 197.865 3781.400 ;
      LAYER met5 ;
        RECT 3390.135 3719.730 3395.385 3867.270 ;
        RECT 3396.985 3719.730 3401.435 3867.270 ;
        RECT 3403.035 3720.035 3406.285 3867.030 ;
        RECT 3407.885 3719.730 3412.335 3867.270 ;
        RECT 3413.935 3719.730 3418.385 3867.270 ;
        RECT 3419.985 3719.730 3423.235 3867.270 ;
        RECT 3424.840 3866.000 3428.085 3867.270 ;
        RECT 3424.835 3721.000 3428.085 3866.000 ;
        RECT 3424.840 3719.730 3428.085 3721.000 ;
        RECT 3429.685 3719.730 3434.135 3867.270 ;
        RECT 3435.735 3719.730 3444.735 3867.270 ;
        RECT 3446.335 3719.730 3450.585 3867.270 ;
        RECT 3452.185 3719.730 3456.435 3867.270 ;
        RECT 3458.035 3719.730 3482.985 3867.270 ;
      LAYER met5 ;
        RECT 3484.585 3866.000 3588.000 3868.870 ;
      LAYER met5 ;
        RECT 3563.785 3721.000 3588.000 3866.000 ;
      LAYER met5 ;
        RECT 3403.035 3718.130 3406.285 3718.435 ;
        RECT 3484.585 3718.130 3588.000 3721.000 ;
        RECT 0.000 3708.870 197.865 3715.500 ;
        RECT 3390.135 3711.500 3588.000 3718.130 ;
        RECT 0.000 3706.000 103.415 3708.870 ;
        RECT 181.715 3708.565 184.965 3708.870 ;
      LAYER met5 ;
        RECT 0.000 3570.000 24.215 3706.000 ;
      LAYER met5 ;
        RECT 0.000 3567.130 103.415 3570.000 ;
      LAYER met5 ;
        RECT 105.015 3568.730 129.965 3707.270 ;
        RECT 131.565 3568.730 135.815 3707.270 ;
        RECT 137.415 3568.730 141.665 3707.270 ;
        RECT 143.265 3568.730 152.265 3707.270 ;
        RECT 153.865 3568.730 158.315 3707.270 ;
        RECT 159.915 3706.000 163.160 3707.270 ;
        RECT 159.915 3570.000 163.165 3706.000 ;
        RECT 159.915 3568.730 163.160 3570.000 ;
        RECT 164.765 3568.730 168.015 3707.270 ;
        RECT 169.615 3568.730 174.065 3707.270 ;
        RECT 175.665 3568.730 180.115 3707.270 ;
        RECT 181.715 3568.970 184.965 3706.965 ;
        RECT 186.565 3568.730 191.015 3707.270 ;
        RECT 192.615 3568.730 197.865 3707.270 ;
      LAYER met5 ;
        RECT 3390.135 3645.600 3490.960 3711.500 ;
        RECT 3556.610 3645.600 3588.000 3711.500 ;
        RECT 3390.135 3643.870 3588.000 3645.600 ;
        RECT 3403.035 3643.630 3406.285 3643.870 ;
        RECT 181.715 3567.130 184.965 3567.370 ;
        RECT 0.000 3565.400 197.865 3567.130 ;
        RECT 0.000 3499.500 31.390 3565.400 ;
        RECT 97.040 3499.500 197.865 3565.400 ;
        RECT 0.000 3492.870 197.865 3499.500 ;
      LAYER met5 ;
        RECT 3390.135 3494.730 3395.385 3642.270 ;
        RECT 3396.985 3494.730 3401.435 3642.270 ;
        RECT 3403.035 3495.035 3406.285 3642.030 ;
        RECT 3407.885 3494.730 3412.335 3642.270 ;
        RECT 3413.935 3494.730 3418.385 3642.270 ;
        RECT 3419.985 3494.730 3423.235 3642.270 ;
        RECT 3424.840 3641.000 3428.085 3642.270 ;
        RECT 3424.835 3496.000 3428.085 3641.000 ;
        RECT 3424.840 3494.730 3428.085 3496.000 ;
        RECT 3429.685 3494.730 3434.135 3642.270 ;
        RECT 3435.735 3494.730 3444.735 3642.270 ;
        RECT 3446.335 3494.730 3450.585 3642.270 ;
        RECT 3452.185 3494.730 3456.435 3642.270 ;
        RECT 3458.035 3494.730 3482.985 3642.270 ;
      LAYER met5 ;
        RECT 3484.585 3641.000 3588.000 3643.870 ;
      LAYER met5 ;
        RECT 3563.785 3496.000 3588.000 3641.000 ;
      LAYER met5 ;
        RECT 3403.035 3493.130 3406.285 3493.435 ;
        RECT 3484.585 3493.130 3588.000 3496.000 ;
        RECT 0.000 3490.000 103.415 3492.870 ;
        RECT 181.715 3492.565 184.965 3492.870 ;
      LAYER met5 ;
        RECT 0.000 3354.000 24.215 3490.000 ;
      LAYER met5 ;
        RECT 0.000 3351.130 103.415 3354.000 ;
      LAYER met5 ;
        RECT 105.015 3352.730 129.965 3491.270 ;
        RECT 131.565 3352.730 135.815 3491.270 ;
        RECT 137.415 3352.730 141.665 3491.270 ;
        RECT 143.265 3352.730 152.265 3491.270 ;
        RECT 153.865 3352.730 158.315 3491.270 ;
        RECT 159.915 3490.000 163.160 3491.270 ;
        RECT 159.915 3354.000 163.165 3490.000 ;
        RECT 159.915 3352.730 163.160 3354.000 ;
        RECT 164.765 3352.730 168.015 3491.270 ;
        RECT 169.615 3352.730 174.065 3491.270 ;
        RECT 175.665 3352.730 180.115 3491.270 ;
        RECT 181.715 3352.970 184.965 3490.965 ;
        RECT 186.565 3352.730 191.015 3491.270 ;
        RECT 192.615 3352.730 197.865 3491.270 ;
      LAYER met5 ;
        RECT 3390.135 3486.500 3588.000 3493.130 ;
        RECT 3390.135 3420.600 3490.960 3486.500 ;
        RECT 3556.610 3420.600 3588.000 3486.500 ;
        RECT 3390.135 3418.870 3588.000 3420.600 ;
        RECT 3403.035 3418.630 3406.285 3418.870 ;
        RECT 181.715 3351.130 184.965 3351.370 ;
        RECT 0.000 3349.400 197.865 3351.130 ;
        RECT 0.000 3283.500 31.390 3349.400 ;
        RECT 97.040 3283.500 197.865 3349.400 ;
        RECT 0.000 3276.870 197.865 3283.500 ;
        RECT 0.000 3274.000 103.415 3276.870 ;
        RECT 181.715 3276.565 184.965 3276.870 ;
      LAYER met5 ;
        RECT 0.000 3138.000 24.215 3274.000 ;
      LAYER met5 ;
        RECT 0.000 3135.130 103.415 3138.000 ;
      LAYER met5 ;
        RECT 105.015 3136.730 129.965 3275.270 ;
        RECT 131.565 3136.730 135.815 3275.270 ;
        RECT 137.415 3136.730 141.665 3275.270 ;
        RECT 143.265 3136.730 152.265 3275.270 ;
        RECT 153.865 3136.730 158.315 3275.270 ;
        RECT 159.915 3274.000 163.160 3275.270 ;
        RECT 159.915 3138.000 163.165 3274.000 ;
        RECT 159.915 3136.730 163.160 3138.000 ;
        RECT 164.765 3136.730 168.015 3275.270 ;
        RECT 169.615 3136.730 174.065 3275.270 ;
        RECT 175.665 3136.730 180.115 3275.270 ;
        RECT 181.715 3136.970 184.965 3274.965 ;
        RECT 186.565 3136.730 191.015 3275.270 ;
        RECT 192.615 3136.730 197.865 3275.270 ;
        RECT 3390.135 3268.730 3395.385 3417.270 ;
        RECT 3396.985 3268.730 3401.435 3417.270 ;
        RECT 3403.035 3269.035 3406.285 3417.030 ;
        RECT 3407.885 3268.730 3412.335 3417.270 ;
        RECT 3413.935 3268.730 3418.385 3417.270 ;
        RECT 3419.985 3268.730 3423.235 3417.270 ;
        RECT 3424.840 3416.000 3428.085 3417.270 ;
        RECT 3424.835 3270.000 3428.085 3416.000 ;
        RECT 3424.840 3268.730 3428.085 3270.000 ;
        RECT 3429.685 3268.730 3434.135 3417.270 ;
        RECT 3435.735 3268.730 3444.735 3417.270 ;
        RECT 3446.335 3268.730 3450.585 3417.270 ;
        RECT 3452.185 3268.730 3456.435 3417.270 ;
        RECT 3458.035 3268.730 3482.985 3417.270 ;
      LAYER met5 ;
        RECT 3484.585 3416.000 3588.000 3418.870 ;
      LAYER met5 ;
        RECT 3563.785 3270.000 3588.000 3416.000 ;
      LAYER met5 ;
        RECT 3403.035 3267.130 3406.285 3267.435 ;
        RECT 3484.585 3267.130 3588.000 3270.000 ;
        RECT 3390.135 3260.500 3588.000 3267.130 ;
        RECT 3390.135 3194.600 3490.960 3260.500 ;
        RECT 3556.610 3194.600 3588.000 3260.500 ;
        RECT 3390.135 3192.870 3588.000 3194.600 ;
        RECT 3403.035 3192.630 3406.285 3192.870 ;
        RECT 181.715 3135.130 184.965 3135.370 ;
        RECT 0.000 3133.400 197.865 3135.130 ;
        RECT 0.000 3067.500 31.390 3133.400 ;
        RECT 97.040 3067.500 197.865 3133.400 ;
        RECT 0.000 3060.870 197.865 3067.500 ;
        RECT 0.000 3058.000 103.415 3060.870 ;
        RECT 181.715 3060.565 184.965 3060.870 ;
      LAYER met5 ;
        RECT 0.000 2922.000 24.215 3058.000 ;
      LAYER met5 ;
        RECT 0.000 2919.130 103.415 2922.000 ;
      LAYER met5 ;
        RECT 105.015 2920.730 129.965 3059.270 ;
        RECT 131.565 2920.730 135.815 3059.270 ;
        RECT 137.415 2920.730 141.665 3059.270 ;
        RECT 143.265 2920.730 152.265 3059.270 ;
        RECT 153.865 2920.730 158.315 3059.270 ;
        RECT 159.915 3058.000 163.160 3059.270 ;
        RECT 159.915 2922.000 163.165 3058.000 ;
        RECT 159.915 2920.730 163.160 2922.000 ;
        RECT 164.765 2920.730 168.015 3059.270 ;
        RECT 169.615 2920.730 174.065 3059.270 ;
        RECT 175.665 2920.730 180.115 3059.270 ;
        RECT 181.715 2920.970 184.965 3058.965 ;
        RECT 186.565 2920.730 191.015 3059.270 ;
        RECT 192.615 2920.730 197.865 3059.270 ;
        RECT 3390.135 3043.730 3395.385 3191.270 ;
        RECT 3396.985 3043.730 3401.435 3191.270 ;
        RECT 3403.035 3044.035 3406.285 3191.030 ;
        RECT 3407.885 3043.730 3412.335 3191.270 ;
        RECT 3413.935 3043.730 3418.385 3191.270 ;
        RECT 3419.985 3043.730 3423.235 3191.270 ;
        RECT 3424.840 3190.000 3428.085 3191.270 ;
        RECT 3424.835 3045.000 3428.085 3190.000 ;
        RECT 3424.840 3043.730 3428.085 3045.000 ;
        RECT 3429.685 3043.730 3434.135 3191.270 ;
        RECT 3435.735 3043.730 3444.735 3191.270 ;
        RECT 3446.335 3043.730 3450.585 3191.270 ;
        RECT 3452.185 3043.730 3456.435 3191.270 ;
        RECT 3458.035 3043.730 3482.985 3191.270 ;
      LAYER met5 ;
        RECT 3484.585 3190.000 3588.000 3192.870 ;
      LAYER met5 ;
        RECT 3563.785 3045.000 3588.000 3190.000 ;
      LAYER met5 ;
        RECT 3403.035 3042.130 3406.285 3042.435 ;
        RECT 3484.585 3042.130 3588.000 3045.000 ;
        RECT 3390.135 3035.500 3588.000 3042.130 ;
        RECT 3390.135 2969.600 3490.960 3035.500 ;
        RECT 3556.610 2969.600 3588.000 3035.500 ;
        RECT 3390.135 2967.870 3588.000 2969.600 ;
        RECT 3403.035 2967.630 3406.285 2967.870 ;
        RECT 181.715 2919.130 184.965 2919.370 ;
        RECT 0.000 2917.400 197.865 2919.130 ;
        RECT 0.000 2851.500 31.390 2917.400 ;
        RECT 97.040 2851.500 197.865 2917.400 ;
        RECT 0.000 2844.870 197.865 2851.500 ;
        RECT 0.000 2842.000 103.415 2844.870 ;
        RECT 181.715 2844.565 184.965 2844.870 ;
      LAYER met5 ;
        RECT 0.000 2706.000 24.215 2842.000 ;
      LAYER met5 ;
        RECT 0.000 2703.130 103.415 2706.000 ;
      LAYER met5 ;
        RECT 105.015 2704.730 129.965 2843.270 ;
        RECT 131.565 2704.730 135.815 2843.270 ;
        RECT 137.415 2704.730 141.665 2843.270 ;
        RECT 143.265 2704.730 152.265 2843.270 ;
        RECT 153.865 2704.730 158.315 2843.270 ;
        RECT 159.915 2842.000 163.160 2843.270 ;
        RECT 159.915 2706.000 163.165 2842.000 ;
        RECT 159.915 2704.730 163.160 2706.000 ;
        RECT 164.765 2704.730 168.015 2843.270 ;
        RECT 169.615 2704.730 174.065 2843.270 ;
        RECT 175.665 2704.730 180.115 2843.270 ;
        RECT 181.715 2704.970 184.965 2842.965 ;
        RECT 186.565 2704.730 191.015 2843.270 ;
        RECT 192.615 2704.730 197.865 2843.270 ;
        RECT 3390.135 2817.730 3395.385 2966.270 ;
        RECT 3396.985 2817.730 3401.435 2966.270 ;
        RECT 3403.035 2818.035 3406.285 2966.030 ;
        RECT 3407.885 2817.730 3412.335 2966.270 ;
        RECT 3413.935 2817.730 3418.385 2966.270 ;
        RECT 3419.985 2817.730 3423.235 2966.270 ;
        RECT 3424.840 2965.000 3428.085 2966.270 ;
        RECT 3424.835 2819.000 3428.085 2965.000 ;
        RECT 3424.840 2817.730 3428.085 2819.000 ;
        RECT 3429.685 2817.730 3434.135 2966.270 ;
        RECT 3435.735 2817.730 3444.735 2966.270 ;
        RECT 3446.335 2817.730 3450.585 2966.270 ;
        RECT 3452.185 2817.730 3456.435 2966.270 ;
        RECT 3458.035 2817.730 3482.985 2966.270 ;
      LAYER met5 ;
        RECT 3484.585 2965.000 3588.000 2967.870 ;
      LAYER met5 ;
        RECT 3563.785 2819.000 3588.000 2965.000 ;
      LAYER met5 ;
        RECT 3403.035 2816.130 3406.285 2816.435 ;
        RECT 3484.585 2816.130 3588.000 2819.000 ;
        RECT 3390.135 2809.500 3588.000 2816.130 ;
        RECT 3390.135 2743.600 3490.960 2809.500 ;
        RECT 3556.610 2743.600 3588.000 2809.500 ;
        RECT 3390.135 2741.870 3588.000 2743.600 ;
        RECT 3403.035 2741.630 3406.285 2741.870 ;
        RECT 181.715 2703.130 184.965 2703.370 ;
        RECT 0.000 2701.400 197.865 2703.130 ;
        RECT 0.000 2635.500 31.390 2701.400 ;
        RECT 97.040 2635.500 197.865 2701.400 ;
        RECT 0.000 2628.870 197.865 2635.500 ;
        RECT 0.000 2626.000 103.415 2628.870 ;
        RECT 181.715 2628.565 184.965 2628.870 ;
      LAYER met5 ;
        RECT 0.000 2490.000 24.215 2626.000 ;
      LAYER met5 ;
        RECT 0.000 2487.130 103.415 2490.000 ;
      LAYER met5 ;
        RECT 105.015 2488.730 129.965 2627.270 ;
        RECT 131.565 2488.730 135.815 2627.270 ;
        RECT 137.415 2488.730 141.665 2627.270 ;
        RECT 143.265 2488.730 152.265 2627.270 ;
        RECT 153.865 2488.730 158.315 2627.270 ;
        RECT 159.915 2626.000 163.160 2627.270 ;
        RECT 159.915 2490.000 163.165 2626.000 ;
        RECT 159.915 2488.730 163.160 2490.000 ;
      LAYER met5 ;
        RECT 163.160 2487.130 163.165 2490.000 ;
      LAYER met5 ;
        RECT 164.765 2488.730 168.015 2627.270 ;
        RECT 169.615 2488.730 174.065 2627.270 ;
        RECT 175.665 2488.730 180.115 2627.270 ;
        RECT 181.715 2489.035 184.965 2626.965 ;
        RECT 186.565 2488.730 191.015 2627.270 ;
        RECT 192.615 2488.730 197.865 2627.270 ;
        RECT 3390.135 2592.730 3395.385 2740.270 ;
        RECT 3396.985 2592.730 3401.435 2740.270 ;
        RECT 3403.035 2593.035 3406.285 2740.030 ;
        RECT 3407.885 2592.730 3412.335 2740.270 ;
        RECT 3413.935 2592.730 3418.385 2740.270 ;
        RECT 3419.985 2592.730 3423.235 2740.270 ;
        RECT 3424.840 2739.000 3428.085 2740.270 ;
        RECT 3424.835 2594.000 3428.085 2739.000 ;
      LAYER met5 ;
        RECT 3403.035 2591.130 3406.285 2591.435 ;
        RECT 3424.835 2591.130 3424.840 2594.000 ;
      LAYER met5 ;
        RECT 3424.840 2592.730 3428.085 2594.000 ;
        RECT 3429.685 2592.730 3434.135 2740.270 ;
        RECT 3435.735 2592.730 3444.735 2740.270 ;
        RECT 3446.335 2592.730 3450.585 2740.270 ;
        RECT 3452.185 2592.730 3456.435 2740.270 ;
        RECT 3458.035 2592.730 3482.985 2740.270 ;
      LAYER met5 ;
        RECT 3484.585 2739.000 3588.000 2741.870 ;
      LAYER met5 ;
        RECT 3563.785 2594.000 3588.000 2739.000 ;
      LAYER met5 ;
        RECT 3484.585 2591.130 3588.000 2594.000 ;
        RECT 3390.135 2588.550 3588.000 2591.130 ;
        RECT 3390.135 2524.510 3491.520 2588.550 ;
        RECT 3555.545 2524.510 3588.000 2588.550 ;
        RECT 3390.135 2521.870 3588.000 2524.510 ;
        RECT 3403.035 2521.565 3406.285 2521.870 ;
        RECT 181.715 2487.130 184.965 2487.435 ;
        RECT 0.000 2484.490 197.865 2487.130 ;
        RECT 0.000 2420.450 32.455 2484.490 ;
        RECT 96.480 2420.450 197.865 2484.490 ;
        RECT 0.000 2417.870 197.865 2420.450 ;
        RECT 0.000 2415.000 103.415 2417.870 ;
      LAYER met5 ;
        RECT 0.000 2279.000 24.215 2415.000 ;
      LAYER met5 ;
        RECT 0.000 2276.130 103.415 2279.000 ;
      LAYER met5 ;
        RECT 105.015 2277.730 129.965 2416.270 ;
        RECT 131.565 2277.730 135.815 2416.270 ;
        RECT 137.415 2277.730 141.665 2416.270 ;
        RECT 143.265 2277.730 152.265 2416.270 ;
        RECT 153.865 2277.730 158.315 2416.270 ;
        RECT 159.915 2415.000 163.160 2416.270 ;
      LAYER met5 ;
        RECT 163.160 2415.000 163.165 2417.870 ;
        RECT 181.715 2417.565 184.965 2417.870 ;
      LAYER met5 ;
        RECT 159.915 2279.000 163.165 2415.000 ;
        RECT 159.915 2277.730 163.160 2279.000 ;
        RECT 164.765 2277.730 168.015 2416.270 ;
        RECT 169.615 2277.730 174.065 2416.270 ;
        RECT 175.665 2277.730 180.115 2416.270 ;
        RECT 181.715 2278.035 184.965 2415.965 ;
        RECT 186.565 2277.730 191.015 2416.270 ;
        RECT 192.615 2277.730 197.865 2416.270 ;
        RECT 3390.135 2372.730 3395.385 2520.270 ;
        RECT 3396.985 2372.730 3401.435 2520.270 ;
        RECT 3403.035 2373.035 3406.285 2519.965 ;
        RECT 3407.885 2372.730 3412.335 2520.270 ;
        RECT 3413.935 2372.730 3418.385 2520.270 ;
        RECT 3419.985 2372.730 3423.235 2520.270 ;
      LAYER met5 ;
        RECT 3424.835 2519.000 3424.840 2521.870 ;
      LAYER met5 ;
        RECT 3424.840 2519.000 3428.085 2520.270 ;
        RECT 3424.835 2374.000 3428.085 2519.000 ;
        RECT 3424.840 2372.730 3428.085 2374.000 ;
        RECT 3429.685 2372.730 3434.135 2520.270 ;
        RECT 3435.735 2372.730 3444.735 2520.270 ;
        RECT 3446.335 2372.730 3450.585 2520.270 ;
        RECT 3452.185 2372.730 3456.435 2520.270 ;
        RECT 3458.035 2372.730 3482.985 2520.270 ;
      LAYER met5 ;
        RECT 3484.585 2519.000 3588.000 2521.870 ;
      LAYER met5 ;
        RECT 3563.785 2374.000 3588.000 2519.000 ;
      LAYER met5 ;
        RECT 3403.035 2371.130 3406.285 2371.435 ;
        RECT 3484.585 2371.130 3588.000 2374.000 ;
        RECT 3390.135 2365.330 3588.000 2371.130 ;
        RECT 3390.135 2307.730 3488.300 2365.330 ;
        RECT 3558.765 2307.730 3588.000 2365.330 ;
        RECT 3390.135 2301.870 3588.000 2307.730 ;
        RECT 3403.035 2301.565 3406.285 2301.870 ;
        RECT 181.715 2276.130 184.965 2276.435 ;
        RECT 0.000 2270.270 197.865 2276.130 ;
        RECT 0.000 2212.670 29.235 2270.270 ;
        RECT 99.700 2212.670 197.865 2270.270 ;
        RECT 0.000 2206.870 197.865 2212.670 ;
        RECT 0.000 2204.000 103.415 2206.870 ;
        RECT 181.715 2206.565 184.965 2206.870 ;
      LAYER met5 ;
        RECT 0.000 2068.000 24.215 2204.000 ;
      LAYER met5 ;
        RECT 0.000 2065.130 103.415 2068.000 ;
      LAYER met5 ;
        RECT 105.015 2066.730 129.965 2205.270 ;
        RECT 131.565 2066.730 135.815 2205.270 ;
        RECT 137.415 2066.730 141.665 2205.270 ;
        RECT 143.265 2066.730 152.265 2205.270 ;
        RECT 153.865 2066.730 158.315 2205.270 ;
        RECT 159.915 2204.000 163.160 2205.270 ;
        RECT 159.915 2068.000 163.165 2204.000 ;
        RECT 159.915 2066.730 163.160 2068.000 ;
        RECT 164.765 2066.730 168.015 2205.270 ;
        RECT 169.615 2066.730 174.065 2205.270 ;
        RECT 175.665 2066.730 180.115 2205.270 ;
        RECT 181.715 2066.970 184.965 2204.965 ;
        RECT 186.565 2066.730 191.015 2205.270 ;
        RECT 192.615 2066.730 197.865 2205.270 ;
        RECT 3390.135 2151.730 3395.385 2300.270 ;
        RECT 3396.985 2151.730 3401.435 2300.270 ;
        RECT 3403.035 2152.035 3406.285 2299.965 ;
        RECT 3407.885 2151.730 3412.335 2300.270 ;
        RECT 3413.935 2151.730 3418.385 2300.270 ;
        RECT 3419.985 2151.730 3423.235 2300.270 ;
        RECT 3424.840 2299.000 3428.085 2300.270 ;
        RECT 3424.835 2153.000 3428.085 2299.000 ;
      LAYER met5 ;
        RECT 3403.035 2150.130 3406.285 2150.435 ;
        RECT 3424.835 2150.130 3424.840 2153.000 ;
      LAYER met5 ;
        RECT 3424.840 2151.730 3428.085 2153.000 ;
        RECT 3429.685 2151.730 3434.135 2300.270 ;
        RECT 3435.735 2151.730 3444.735 2300.270 ;
        RECT 3446.335 2151.730 3450.585 2300.270 ;
        RECT 3452.185 2151.730 3456.435 2300.270 ;
        RECT 3458.035 2151.730 3482.985 2300.270 ;
      LAYER met5 ;
        RECT 3484.585 2299.000 3588.000 2301.870 ;
      LAYER met5 ;
        RECT 3563.785 2153.000 3588.000 2299.000 ;
      LAYER met5 ;
        RECT 3484.585 2150.130 3588.000 2153.000 ;
        RECT 3390.135 2147.550 3588.000 2150.130 ;
        RECT 3390.135 2083.510 3491.520 2147.550 ;
        RECT 3555.545 2083.510 3588.000 2147.550 ;
        RECT 3390.135 2080.870 3588.000 2083.510 ;
        RECT 3403.035 2080.565 3406.285 2080.870 ;
        RECT 181.715 2065.130 184.965 2065.370 ;
        RECT 0.000 2063.400 197.865 2065.130 ;
        RECT 0.000 1997.500 31.390 2063.400 ;
        RECT 97.040 1997.500 197.865 2063.400 ;
        RECT 0.000 1990.870 197.865 1997.500 ;
        RECT 0.000 1988.000 103.415 1990.870 ;
        RECT 181.715 1990.565 184.965 1990.870 ;
      LAYER met5 ;
        RECT 0.000 1852.000 24.215 1988.000 ;
      LAYER met5 ;
        RECT 0.000 1849.130 103.415 1852.000 ;
      LAYER met5 ;
        RECT 105.015 1850.730 129.965 1989.270 ;
        RECT 131.565 1850.730 135.815 1989.270 ;
        RECT 137.415 1850.730 141.665 1989.270 ;
        RECT 143.265 1850.730 152.265 1989.270 ;
        RECT 153.865 1850.730 158.315 1989.270 ;
        RECT 159.915 1988.000 163.160 1989.270 ;
        RECT 159.915 1852.000 163.165 1988.000 ;
        RECT 159.915 1850.730 163.160 1852.000 ;
        RECT 164.765 1850.730 168.015 1989.270 ;
        RECT 169.615 1850.730 174.065 1989.270 ;
        RECT 175.665 1850.730 180.115 1989.270 ;
        RECT 181.715 1850.970 184.965 1988.965 ;
        RECT 186.565 1850.730 191.015 1989.270 ;
        RECT 192.615 1850.730 197.865 1989.270 ;
        RECT 3390.135 1931.730 3395.385 2079.270 ;
        RECT 3396.985 1931.730 3401.435 2079.270 ;
        RECT 3403.035 1932.035 3406.285 2078.965 ;
        RECT 3407.885 1931.730 3412.335 2079.270 ;
        RECT 3413.935 1931.730 3418.385 2079.270 ;
        RECT 3419.985 1931.730 3423.235 2079.270 ;
      LAYER met5 ;
        RECT 3424.835 2078.000 3424.840 2080.870 ;
      LAYER met5 ;
        RECT 3424.840 2078.000 3428.085 2079.270 ;
        RECT 3424.835 1933.000 3428.085 2078.000 ;
        RECT 3424.840 1931.730 3428.085 1933.000 ;
        RECT 3429.685 1931.730 3434.135 2079.270 ;
        RECT 3435.735 1931.730 3444.735 2079.270 ;
        RECT 3446.335 1931.730 3450.585 2079.270 ;
        RECT 3452.185 1931.730 3456.435 2079.270 ;
        RECT 3458.035 1931.730 3482.985 2079.270 ;
      LAYER met5 ;
        RECT 3484.585 2078.000 3588.000 2080.870 ;
      LAYER met5 ;
        RECT 3563.785 1933.000 3588.000 2078.000 ;
      LAYER met5 ;
        RECT 3403.035 1930.130 3406.285 1930.435 ;
        RECT 3484.585 1930.130 3588.000 1933.000 ;
        RECT 3390.135 1923.500 3588.000 1930.130 ;
        RECT 3390.135 1857.600 3490.960 1923.500 ;
        RECT 3556.610 1857.600 3588.000 1923.500 ;
        RECT 3390.135 1855.870 3588.000 1857.600 ;
        RECT 3403.035 1855.630 3406.285 1855.870 ;
        RECT 181.715 1849.130 184.965 1849.370 ;
        RECT 0.000 1847.400 197.865 1849.130 ;
        RECT 0.000 1781.500 31.390 1847.400 ;
        RECT 97.040 1781.500 197.865 1847.400 ;
        RECT 0.000 1774.870 197.865 1781.500 ;
        RECT 0.000 1772.000 103.415 1774.870 ;
        RECT 181.715 1774.565 184.965 1774.870 ;
      LAYER met5 ;
        RECT 0.000 1636.000 24.215 1772.000 ;
      LAYER met5 ;
        RECT 0.000 1633.130 103.415 1636.000 ;
      LAYER met5 ;
        RECT 105.015 1634.730 129.965 1773.270 ;
        RECT 131.565 1634.730 135.815 1773.270 ;
        RECT 137.415 1634.730 141.665 1773.270 ;
        RECT 143.265 1634.730 152.265 1773.270 ;
        RECT 153.865 1634.730 158.315 1773.270 ;
        RECT 159.915 1772.000 163.160 1773.270 ;
        RECT 159.915 1636.000 163.165 1772.000 ;
        RECT 159.915 1634.730 163.160 1636.000 ;
        RECT 164.765 1634.730 168.015 1773.270 ;
        RECT 169.615 1634.730 174.065 1773.270 ;
        RECT 175.665 1634.730 180.115 1773.270 ;
        RECT 181.715 1634.970 184.965 1772.965 ;
        RECT 186.565 1634.730 191.015 1773.270 ;
        RECT 192.615 1634.730 197.865 1773.270 ;
        RECT 3390.135 1705.730 3395.385 1854.270 ;
        RECT 3396.985 1705.730 3401.435 1854.270 ;
        RECT 3403.035 1706.035 3406.285 1854.030 ;
        RECT 3407.885 1705.730 3412.335 1854.270 ;
        RECT 3413.935 1705.730 3418.385 1854.270 ;
        RECT 3419.985 1705.730 3423.235 1854.270 ;
        RECT 3424.840 1853.000 3428.085 1854.270 ;
        RECT 3424.835 1707.000 3428.085 1853.000 ;
        RECT 3424.840 1705.730 3428.085 1707.000 ;
        RECT 3429.685 1705.730 3434.135 1854.270 ;
        RECT 3435.735 1705.730 3444.735 1854.270 ;
        RECT 3446.335 1705.730 3450.585 1854.270 ;
        RECT 3452.185 1705.730 3456.435 1854.270 ;
        RECT 3458.035 1705.730 3482.985 1854.270 ;
      LAYER met5 ;
        RECT 3484.585 1853.000 3588.000 1855.870 ;
      LAYER met5 ;
        RECT 3563.785 1707.000 3588.000 1853.000 ;
      LAYER met5 ;
        RECT 3403.035 1704.130 3406.285 1704.435 ;
        RECT 3484.585 1704.130 3588.000 1707.000 ;
        RECT 3390.135 1697.500 3588.000 1704.130 ;
        RECT 181.715 1633.130 184.965 1633.370 ;
        RECT 0.000 1631.400 197.865 1633.130 ;
        RECT 0.000 1565.500 31.390 1631.400 ;
        RECT 97.040 1565.500 197.865 1631.400 ;
        RECT 3390.135 1631.600 3490.960 1697.500 ;
        RECT 3556.610 1631.600 3588.000 1697.500 ;
        RECT 3390.135 1629.870 3588.000 1631.600 ;
        RECT 3403.035 1629.630 3406.285 1629.870 ;
        RECT 0.000 1558.870 197.865 1565.500 ;
        RECT 0.000 1556.000 103.415 1558.870 ;
        RECT 181.715 1558.565 184.965 1558.870 ;
      LAYER met5 ;
        RECT 0.000 1420.000 24.215 1556.000 ;
      LAYER met5 ;
        RECT 0.000 1417.130 103.415 1420.000 ;
      LAYER met5 ;
        RECT 105.015 1418.730 129.965 1557.270 ;
        RECT 131.565 1418.730 135.815 1557.270 ;
        RECT 137.415 1418.730 141.665 1557.270 ;
        RECT 143.265 1418.730 152.265 1557.270 ;
        RECT 153.865 1418.730 158.315 1557.270 ;
        RECT 159.915 1556.000 163.160 1557.270 ;
        RECT 159.915 1420.000 163.165 1556.000 ;
        RECT 159.915 1418.730 163.160 1420.000 ;
        RECT 164.765 1418.730 168.015 1557.270 ;
        RECT 169.615 1418.730 174.065 1557.270 ;
        RECT 175.665 1418.730 180.115 1557.270 ;
        RECT 181.715 1418.970 184.965 1556.965 ;
        RECT 186.565 1418.730 191.015 1557.270 ;
        RECT 192.615 1418.730 197.865 1557.270 ;
        RECT 3390.135 1480.730 3395.385 1628.270 ;
        RECT 3396.985 1480.730 3401.435 1628.270 ;
        RECT 3403.035 1481.035 3406.285 1628.030 ;
        RECT 3407.885 1480.730 3412.335 1628.270 ;
        RECT 3413.935 1480.730 3418.385 1628.270 ;
        RECT 3419.985 1480.730 3423.235 1628.270 ;
        RECT 3424.840 1627.000 3428.085 1628.270 ;
        RECT 3424.835 1482.000 3428.085 1627.000 ;
        RECT 3424.840 1480.730 3428.085 1482.000 ;
        RECT 3429.685 1480.730 3434.135 1628.270 ;
        RECT 3435.735 1480.730 3444.735 1628.270 ;
        RECT 3446.335 1480.730 3450.585 1628.270 ;
        RECT 3452.185 1480.730 3456.435 1628.270 ;
        RECT 3458.035 1480.730 3482.985 1628.270 ;
      LAYER met5 ;
        RECT 3484.585 1627.000 3588.000 1629.870 ;
      LAYER met5 ;
        RECT 3563.785 1482.000 3588.000 1627.000 ;
      LAYER met5 ;
        RECT 3403.035 1479.130 3406.285 1479.435 ;
        RECT 3484.585 1479.130 3588.000 1482.000 ;
        RECT 3390.135 1472.500 3588.000 1479.130 ;
        RECT 181.715 1417.130 184.965 1417.370 ;
        RECT 0.000 1415.400 197.865 1417.130 ;
        RECT 0.000 1349.500 31.390 1415.400 ;
        RECT 97.040 1349.500 197.865 1415.400 ;
        RECT 3390.135 1406.600 3490.960 1472.500 ;
        RECT 3556.610 1406.600 3588.000 1472.500 ;
        RECT 3390.135 1404.870 3588.000 1406.600 ;
        RECT 3403.035 1404.630 3406.285 1404.870 ;
        RECT 0.000 1342.870 197.865 1349.500 ;
        RECT 0.000 1340.000 103.415 1342.870 ;
        RECT 181.715 1342.565 184.965 1342.870 ;
      LAYER met5 ;
        RECT 0.000 1204.000 24.215 1340.000 ;
      LAYER met5 ;
        RECT 0.000 1201.130 103.415 1204.000 ;
      LAYER met5 ;
        RECT 105.015 1202.730 129.965 1341.270 ;
        RECT 131.565 1202.730 135.815 1341.270 ;
        RECT 137.415 1202.730 141.665 1341.270 ;
        RECT 143.265 1202.730 152.265 1341.270 ;
        RECT 153.865 1202.730 158.315 1341.270 ;
        RECT 159.915 1340.000 163.160 1341.270 ;
        RECT 159.915 1204.000 163.165 1340.000 ;
        RECT 159.915 1202.730 163.160 1204.000 ;
        RECT 164.765 1202.730 168.015 1341.270 ;
        RECT 169.615 1202.730 174.065 1341.270 ;
        RECT 175.665 1202.730 180.115 1341.270 ;
        RECT 181.715 1202.970 184.965 1340.965 ;
        RECT 186.565 1202.730 191.015 1341.270 ;
        RECT 192.615 1202.730 197.865 1341.270 ;
        RECT 3390.135 1255.730 3395.385 1403.270 ;
        RECT 3396.985 1255.730 3401.435 1403.270 ;
        RECT 3403.035 1256.035 3406.285 1403.030 ;
        RECT 3407.885 1255.730 3412.335 1403.270 ;
        RECT 3413.935 1255.730 3418.385 1403.270 ;
        RECT 3419.985 1255.730 3423.235 1403.270 ;
        RECT 3424.840 1402.000 3428.085 1403.270 ;
        RECT 3424.835 1257.000 3428.085 1402.000 ;
        RECT 3424.840 1255.730 3428.085 1257.000 ;
        RECT 3429.685 1255.730 3434.135 1403.270 ;
        RECT 3435.735 1255.730 3444.735 1403.270 ;
        RECT 3446.335 1255.730 3450.585 1403.270 ;
        RECT 3452.185 1255.730 3456.435 1403.270 ;
        RECT 3458.035 1255.730 3482.985 1403.270 ;
      LAYER met5 ;
        RECT 3484.585 1402.000 3588.000 1404.870 ;
      LAYER met5 ;
        RECT 3563.785 1257.000 3588.000 1402.000 ;
      LAYER met5 ;
        RECT 3403.035 1254.130 3406.285 1254.435 ;
        RECT 3484.585 1254.130 3588.000 1257.000 ;
        RECT 3390.135 1247.500 3588.000 1254.130 ;
        RECT 181.715 1201.130 184.965 1201.370 ;
        RECT 0.000 1199.400 197.865 1201.130 ;
        RECT 0.000 1133.500 31.390 1199.400 ;
        RECT 97.040 1133.500 197.865 1199.400 ;
        RECT 3390.135 1181.600 3490.960 1247.500 ;
        RECT 3556.610 1181.600 3588.000 1247.500 ;
        RECT 3390.135 1179.870 3588.000 1181.600 ;
        RECT 3403.035 1179.630 3406.285 1179.870 ;
        RECT 0.000 1126.870 197.865 1133.500 ;
        RECT 0.000 1124.000 103.415 1126.870 ;
        RECT 181.715 1126.565 184.965 1126.870 ;
      LAYER met5 ;
        RECT 0.000 988.000 24.215 1124.000 ;
      LAYER met5 ;
        RECT 0.000 985.130 103.415 988.000 ;
      LAYER met5 ;
        RECT 105.015 986.730 129.965 1125.270 ;
        RECT 131.565 986.730 135.815 1125.270 ;
        RECT 137.415 986.730 141.665 1125.270 ;
        RECT 143.265 986.730 152.265 1125.270 ;
        RECT 153.865 986.730 158.315 1125.270 ;
        RECT 159.915 1124.000 163.160 1125.270 ;
        RECT 159.915 988.000 163.165 1124.000 ;
        RECT 159.915 986.730 163.160 988.000 ;
        RECT 164.765 986.730 168.015 1125.270 ;
        RECT 169.615 986.730 174.065 1125.270 ;
        RECT 175.665 986.730 180.115 1125.270 ;
        RECT 181.715 986.970 184.965 1124.965 ;
        RECT 186.565 986.730 191.015 1125.270 ;
        RECT 192.615 986.730 197.865 1125.270 ;
        RECT 3390.135 1029.730 3395.385 1178.270 ;
        RECT 3396.985 1029.730 3401.435 1178.270 ;
        RECT 3403.035 1030.035 3406.285 1178.030 ;
        RECT 3407.885 1029.730 3412.335 1178.270 ;
        RECT 3413.935 1029.730 3418.385 1178.270 ;
        RECT 3419.985 1029.730 3423.235 1178.270 ;
        RECT 3424.840 1177.000 3428.085 1178.270 ;
        RECT 3424.835 1031.000 3428.085 1177.000 ;
        RECT 3424.840 1029.730 3428.085 1031.000 ;
        RECT 3429.685 1029.730 3434.135 1178.270 ;
        RECT 3435.735 1029.730 3444.735 1178.270 ;
        RECT 3446.335 1029.730 3450.585 1178.270 ;
        RECT 3452.185 1029.730 3456.435 1178.270 ;
        RECT 3458.035 1029.730 3482.985 1178.270 ;
      LAYER met5 ;
        RECT 3484.585 1177.000 3588.000 1179.870 ;
      LAYER met5 ;
        RECT 3563.785 1031.000 3588.000 1177.000 ;
      LAYER met5 ;
        RECT 3403.035 1028.130 3406.285 1028.435 ;
        RECT 3484.585 1028.130 3588.000 1031.000 ;
        RECT 3390.135 1021.500 3588.000 1028.130 ;
        RECT 181.715 985.130 184.965 985.370 ;
        RECT 0.000 983.400 197.865 985.130 ;
        RECT 0.000 917.500 31.390 983.400 ;
        RECT 97.040 917.500 197.865 983.400 ;
        RECT 3390.135 955.600 3490.960 1021.500 ;
        RECT 3556.610 955.600 3588.000 1021.500 ;
        RECT 3390.135 953.870 3588.000 955.600 ;
        RECT 3403.035 953.630 3406.285 953.870 ;
        RECT 0.000 910.870 197.865 917.500 ;
        RECT 0.000 908.000 103.415 910.870 ;
        RECT 181.715 910.565 184.965 910.870 ;
      LAYER met5 ;
        RECT 0.000 626.000 24.215 908.000 ;
      LAYER met5 ;
        RECT 0.000 623.130 103.415 626.000 ;
      LAYER met5 ;
        RECT 105.015 624.730 129.965 909.270 ;
        RECT 131.565 624.730 135.815 909.270 ;
        RECT 137.415 624.730 141.665 909.270 ;
        RECT 143.265 631.000 152.265 909.270 ;
        RECT 153.865 636.000 158.315 909.270 ;
        RECT 159.915 908.000 163.160 909.270 ;
        RECT 159.915 631.000 163.165 908.000 ;
        RECT 143.265 624.730 152.265 626.000 ;
        RECT 153.865 624.730 158.315 631.000 ;
        RECT 159.915 624.730 163.160 626.000 ;
      LAYER met5 ;
        RECT 163.160 623.130 163.165 626.000 ;
      LAYER met5 ;
        RECT 164.765 624.730 168.015 909.270 ;
        RECT 169.615 624.730 174.065 909.270 ;
        RECT 175.665 624.730 180.115 909.270 ;
        RECT 181.715 631.000 184.965 908.965 ;
        RECT 186.565 636.000 191.015 909.270 ;
        RECT 181.715 625.035 184.965 626.000 ;
        RECT 186.565 624.730 191.015 631.000 ;
        RECT 192.615 624.730 197.865 909.270 ;
        RECT 3390.135 804.730 3395.385 952.270 ;
        RECT 3396.985 804.730 3401.435 952.270 ;
        RECT 3403.035 805.035 3406.285 952.030 ;
        RECT 3407.885 804.730 3412.335 952.270 ;
        RECT 3413.935 804.730 3418.385 952.270 ;
        RECT 3419.985 804.730 3423.235 952.270 ;
        RECT 3424.840 951.000 3428.085 952.270 ;
        RECT 3424.835 806.000 3428.085 951.000 ;
        RECT 3424.840 804.730 3428.085 806.000 ;
        RECT 3429.685 804.730 3434.135 952.270 ;
        RECT 3435.735 804.730 3444.735 952.270 ;
        RECT 3446.335 804.730 3450.585 952.270 ;
        RECT 3452.185 804.730 3456.435 952.270 ;
        RECT 3458.035 804.730 3482.985 952.270 ;
      LAYER met5 ;
        RECT 3484.585 951.000 3588.000 953.870 ;
      LAYER met5 ;
        RECT 3563.785 806.000 3588.000 951.000 ;
      LAYER met5 ;
        RECT 3403.035 803.130 3406.285 803.435 ;
        RECT 3484.585 803.130 3588.000 806.000 ;
        RECT 3390.135 796.500 3588.000 803.130 ;
        RECT 3390.135 730.600 3490.960 796.500 ;
        RECT 3556.610 730.600 3588.000 796.500 ;
        RECT 3390.135 728.870 3588.000 730.600 ;
        RECT 3403.035 728.630 3406.285 728.870 ;
        RECT 181.715 623.130 184.965 623.435 ;
        RECT 0.000 620.490 197.865 623.130 ;
        RECT 0.000 556.450 32.455 620.490 ;
        RECT 96.480 556.450 197.865 620.490 ;
      LAYER met5 ;
        RECT 3390.135 578.730 3395.385 727.270 ;
        RECT 3396.985 578.730 3401.435 727.270 ;
        RECT 3403.035 579.035 3406.285 727.030 ;
        RECT 3407.885 578.730 3412.335 727.270 ;
        RECT 3413.935 578.730 3418.385 727.270 ;
        RECT 3419.985 578.730 3423.235 727.270 ;
        RECT 3424.840 726.000 3428.085 727.270 ;
        RECT 3424.835 580.000 3428.085 726.000 ;
        RECT 3424.840 578.730 3428.085 580.000 ;
        RECT 3429.685 578.730 3434.135 727.270 ;
        RECT 3435.735 578.730 3444.735 727.270 ;
        RECT 3446.335 578.730 3450.585 727.270 ;
        RECT 3452.185 578.730 3456.435 727.270 ;
        RECT 3458.035 578.730 3482.985 727.270 ;
      LAYER met5 ;
        RECT 3484.585 726.000 3588.000 728.870 ;
      LAYER met5 ;
        RECT 3563.785 580.000 3588.000 726.000 ;
      LAYER met5 ;
        RECT 3403.035 577.130 3406.285 577.435 ;
        RECT 3484.585 577.130 3588.000 580.000 ;
        RECT 0.000 553.870 197.865 556.450 ;
        RECT 3390.135 570.500 3588.000 577.130 ;
        RECT 0.000 551.000 103.415 553.870 ;
      LAYER met5 ;
        RECT 0.000 415.000 24.215 551.000 ;
      LAYER met5 ;
        RECT 0.000 412.130 103.415 415.000 ;
      LAYER met5 ;
        RECT 105.015 413.730 129.965 552.270 ;
        RECT 131.565 413.730 135.815 552.270 ;
        RECT 137.415 413.730 141.665 552.270 ;
        RECT 143.265 413.730 152.265 552.270 ;
        RECT 153.865 413.730 158.315 552.270 ;
        RECT 159.915 551.000 163.160 552.270 ;
      LAYER met5 ;
        RECT 163.160 551.000 163.165 553.870 ;
        RECT 181.715 553.565 184.965 553.870 ;
      LAYER met5 ;
        RECT 159.915 415.000 163.165 551.000 ;
        RECT 159.915 413.730 163.160 415.000 ;
      LAYER met5 ;
        RECT 163.160 412.130 163.165 415.000 ;
      LAYER met5 ;
        RECT 164.765 413.730 168.015 552.270 ;
        RECT 169.615 413.730 174.065 552.270 ;
        RECT 175.665 413.730 180.115 552.270 ;
        RECT 181.715 414.035 184.965 551.965 ;
        RECT 186.565 413.730 191.015 552.270 ;
        RECT 192.615 413.730 197.865 552.270 ;
      LAYER met5 ;
        RECT 3390.135 504.600 3490.960 570.500 ;
        RECT 3556.610 504.600 3588.000 570.500 ;
        RECT 3390.135 502.870 3588.000 504.600 ;
        RECT 3403.035 502.630 3406.285 502.870 ;
        RECT 181.715 412.130 184.965 412.435 ;
        RECT 0.000 406.270 197.865 412.130 ;
        RECT 0.000 348.670 29.235 406.270 ;
        RECT 99.700 348.670 197.865 406.270 ;
        RECT 0.000 342.870 197.865 348.670 ;
        RECT 0.000 340.000 103.415 342.870 ;
      LAYER met5 ;
        RECT 0.000 204.000 24.215 340.000 ;
      LAYER met5 ;
        RECT 0.000 200.545 103.415 204.000 ;
      LAYER met5 ;
        RECT 105.015 202.145 129.965 341.270 ;
        RECT 131.565 202.730 135.815 341.270 ;
        RECT 137.415 202.730 141.665 341.270 ;
      LAYER met5 ;
        RECT 131.565 200.545 141.665 201.130 ;
        RECT 0.000 175.245 141.665 200.545 ;
      LAYER met5 ;
        RECT 143.265 176.845 152.265 341.270 ;
        RECT 153.865 202.730 158.315 341.270 ;
        RECT 159.915 340.000 163.160 341.270 ;
      LAYER met5 ;
        RECT 163.160 340.000 163.165 342.870 ;
        RECT 181.715 342.565 184.965 342.870 ;
      LAYER met5 ;
        RECT 159.915 204.000 163.165 340.000 ;
        RECT 159.915 202.730 163.160 204.000 ;
        RECT 164.765 202.730 168.015 341.270 ;
        RECT 169.615 202.730 174.065 341.270 ;
        RECT 175.665 202.730 180.115 341.270 ;
        RECT 181.715 202.745 184.965 340.965 ;
        RECT 186.565 202.730 191.015 341.270 ;
        RECT 192.615 202.730 197.865 341.270 ;
      LAYER met5 ;
        RECT 181.715 201.130 184.965 201.145 ;
        RECT 199.465 201.130 200.000 204.000 ;
        RECT 153.865 199.465 200.000 201.130 ;
        RECT 3384.000 199.465 3388.535 200.000 ;
        RECT 153.865 192.615 196.050 199.465 ;
      LAYER met5 ;
        RECT 197.650 192.615 395.270 197.865 ;
      LAYER met5 ;
        RECT 153.865 184.965 194.615 192.615 ;
      LAYER met5 ;
        RECT 237.000 191.015 357.000 192.615 ;
        RECT 196.215 186.565 395.270 191.015 ;
      LAYER met5 ;
        RECT 396.870 184.965 466.130 197.865 ;
      LAYER met5 ;
        RECT 467.730 192.615 664.270 197.865 ;
        RECT 506.000 191.015 626.000 192.615 ;
        RECT 467.730 186.565 664.270 191.015 ;
      LAYER met5 ;
        RECT 665.870 184.965 735.130 197.865 ;
      LAYER met5 ;
        RECT 736.730 192.615 933.270 197.865 ;
        RECT 775.000 191.015 895.000 192.615 ;
        RECT 736.730 186.565 933.270 191.015 ;
      LAYER met5 ;
        RECT 934.870 184.965 1009.130 197.865 ;
      LAYER met5 ;
        RECT 1010.730 192.615 1207.270 197.865 ;
        RECT 1049.000 191.015 1169.000 192.615 ;
        RECT 1010.730 186.565 1207.270 191.015 ;
      LAYER met5 ;
        RECT 1208.870 184.965 1278.130 197.865 ;
      LAYER met5 ;
        RECT 1279.730 192.615 1476.270 197.865 ;
        RECT 1318.000 191.015 1438.000 192.615 ;
        RECT 1279.730 186.565 1476.270 191.015 ;
      LAYER met5 ;
        RECT 1477.870 184.965 1552.130 197.865 ;
      LAYER met5 ;
        RECT 1553.730 192.615 1750.270 197.865 ;
        RECT 1592.000 191.015 1712.000 192.615 ;
        RECT 1553.730 186.565 1750.270 191.015 ;
      LAYER met5 ;
        RECT 1751.870 184.965 1826.130 197.865 ;
      LAYER met5 ;
        RECT 1827.730 192.615 2024.270 197.865 ;
        RECT 1866.000 191.015 1986.000 192.615 ;
        RECT 1827.730 186.565 2024.270 191.015 ;
      LAYER met5 ;
        RECT 2025.870 184.965 2100.130 197.865 ;
      LAYER met5 ;
        RECT 2101.730 192.615 2298.270 197.865 ;
        RECT 2140.000 191.015 2260.000 192.615 ;
        RECT 2101.730 186.565 2298.270 191.015 ;
      LAYER met5 ;
        RECT 2299.870 184.965 2374.130 197.865 ;
      LAYER met5 ;
        RECT 2375.730 192.615 2572.270 197.865 ;
        RECT 2414.000 191.015 2534.000 192.615 ;
        RECT 2375.730 186.565 2572.270 191.015 ;
      LAYER met5 ;
        RECT 2573.870 184.965 2648.130 197.865 ;
      LAYER met5 ;
        RECT 2649.730 192.615 2846.270 197.865 ;
        RECT 2688.000 191.015 2808.000 192.615 ;
        RECT 2649.730 186.565 2846.270 191.015 ;
      LAYER met5 ;
        RECT 2847.870 184.965 2917.130 197.865 ;
      LAYER met5 ;
        RECT 2918.730 192.615 3115.270 197.865 ;
        RECT 2957.000 191.015 3077.000 192.615 ;
        RECT 2918.730 186.565 3115.270 191.015 ;
      LAYER met5 ;
        RECT 3116.870 184.965 3186.130 197.865 ;
      LAYER met5 ;
        RECT 3187.730 192.615 3385.270 197.865 ;
      LAYER met5 ;
        RECT 3386.870 196.050 3388.535 199.465 ;
      LAYER met5 ;
        RECT 3390.135 197.650 3395.385 501.270 ;
        RECT 3396.985 355.000 3401.435 501.270 ;
        RECT 3403.035 350.000 3406.285 501.030 ;
        RECT 3396.985 196.215 3401.435 350.000 ;
        RECT 3403.035 198.530 3406.285 345.000 ;
        RECT 3407.885 198.475 3412.335 501.270 ;
        RECT 3413.935 198.400 3418.385 501.270 ;
        RECT 3419.985 198.615 3423.235 501.270 ;
        RECT 3424.840 500.000 3428.085 501.270 ;
        RECT 3424.835 350.000 3428.085 500.000 ;
        RECT 3429.685 355.000 3434.135 501.270 ;
        RECT 3435.735 350.000 3444.735 501.270 ;
        RECT 3424.835 198.665 3428.085 345.000 ;
        RECT 3429.685 198.525 3434.135 350.000 ;
      LAYER met5 ;
        RECT 3424.835 197.015 3428.085 197.065 ;
        RECT 3403.035 196.875 3406.285 196.930 ;
        RECT 3419.985 196.925 3428.085 197.015 ;
        RECT 3403.035 196.800 3412.335 196.875 ;
        RECT 3419.985 196.800 3434.135 196.925 ;
        RECT 3386.870 194.615 3395.385 196.050 ;
        RECT 3403.035 194.615 3434.135 196.800 ;
      LAYER met5 ;
        RECT 3226.000 191.015 3346.000 192.615 ;
        RECT 3187.730 186.565 3385.270 191.015 ;
      LAYER met5 ;
        RECT 3386.870 184.965 3434.135 194.615 ;
        RECT 153.865 181.715 196.930 184.965 ;
      LAYER met5 ;
        RECT 198.530 181.715 394.965 184.965 ;
      LAYER met5 ;
        RECT 396.565 181.715 466.435 184.965 ;
      LAYER met5 ;
        RECT 468.035 181.715 663.965 184.965 ;
      LAYER met5 ;
        RECT 665.565 181.715 735.435 184.965 ;
      LAYER met5 ;
        RECT 737.035 181.715 933.030 184.965 ;
      LAYER met5 ;
        RECT 934.630 181.715 1009.435 184.965 ;
      LAYER met5 ;
        RECT 1011.035 181.715 1206.965 184.965 ;
      LAYER met5 ;
        RECT 1208.565 181.715 1278.435 184.965 ;
      LAYER met5 ;
        RECT 1280.035 181.715 1476.030 184.965 ;
      LAYER met5 ;
        RECT 1477.630 181.715 1552.435 184.965 ;
      LAYER met5 ;
        RECT 1554.035 181.715 1750.030 184.965 ;
      LAYER met5 ;
        RECT 1751.630 181.715 1826.435 184.965 ;
      LAYER met5 ;
        RECT 1828.035 181.715 2024.030 184.965 ;
      LAYER met5 ;
        RECT 2025.630 181.715 2100.435 184.965 ;
      LAYER met5 ;
        RECT 2102.035 181.715 2298.030 184.965 ;
      LAYER met5 ;
        RECT 2299.630 181.715 2374.435 184.965 ;
      LAYER met5 ;
        RECT 2376.035 181.715 2572.030 184.965 ;
      LAYER met5 ;
        RECT 2573.630 181.715 2648.435 184.965 ;
      LAYER met5 ;
        RECT 2650.035 181.715 2845.965 184.965 ;
      LAYER met5 ;
        RECT 2847.565 181.715 2917.435 184.965 ;
      LAYER met5 ;
        RECT 2919.035 181.715 3114.965 184.965 ;
      LAYER met5 ;
        RECT 3116.565 181.715 3186.435 184.965 ;
      LAYER met5 ;
        RECT 3188.035 181.715 3385.255 184.965 ;
      LAYER met5 ;
        RECT 3386.855 181.715 3434.135 184.965 ;
        RECT 153.865 175.665 196.875 181.715 ;
      LAYER met5 ;
        RECT 198.475 175.665 395.270 180.115 ;
      LAYER met5 ;
        RECT 153.865 175.245 196.800 175.665 ;
        RECT 0.000 168.015 196.800 175.245 ;
      LAYER met5 ;
        RECT 198.400 169.615 395.270 174.065 ;
      LAYER met5 ;
        RECT 0.000 163.165 197.015 168.015 ;
      LAYER met5 ;
        RECT 198.615 164.765 395.270 168.015 ;
      LAYER met5 ;
        RECT 396.870 163.165 466.130 181.715 ;
      LAYER met5 ;
        RECT 467.730 175.665 664.270 180.115 ;
        RECT 467.730 169.615 664.270 174.065 ;
        RECT 467.730 164.765 664.270 168.015 ;
      LAYER met5 ;
        RECT 0.000 159.915 197.065 163.165 ;
      LAYER met5 ;
        RECT 198.665 163.160 394.000 163.165 ;
      LAYER met5 ;
        RECT 394.000 163.160 469.000 163.165 ;
      LAYER met5 ;
        RECT 469.000 163.160 663.000 163.165 ;
        RECT 198.665 159.915 395.270 163.160 ;
      LAYER met5 ;
        RECT 0.000 153.865 196.925 159.915 ;
      LAYER met5 ;
        RECT 198.525 153.865 395.270 158.315 ;
      LAYER met5 ;
        RECT 0.000 141.665 175.245 153.865 ;
      LAYER met5 ;
        RECT 176.845 143.265 395.270 152.265 ;
      LAYER met5 ;
        RECT 0.000 135.815 196.775 141.665 ;
      LAYER met5 ;
        RECT 198.375 137.415 395.270 141.665 ;
      LAYER met5 ;
        RECT 0.000 131.565 196.920 135.815 ;
      LAYER met5 ;
        RECT 198.520 131.565 395.270 135.815 ;
      LAYER met5 ;
        RECT 0.000 103.415 195.755 131.565 ;
      LAYER met5 ;
        RECT 197.355 105.015 395.270 129.965 ;
      LAYER met5 ;
        RECT 396.870 103.415 466.130 163.160 ;
      LAYER met5 ;
        RECT 467.730 159.915 664.270 163.160 ;
        RECT 467.730 153.865 664.270 158.315 ;
        RECT 467.730 143.265 664.270 152.265 ;
        RECT 467.730 137.415 664.270 141.665 ;
        RECT 467.730 131.565 664.270 135.815 ;
        RECT 467.730 105.015 664.270 129.965 ;
      LAYER met5 ;
        RECT 665.870 103.415 735.130 181.715 ;
      LAYER met5 ;
        RECT 736.730 175.665 933.270 180.115 ;
        RECT 736.730 169.615 933.270 174.065 ;
        RECT 736.730 164.765 933.270 168.015 ;
        RECT 738.000 163.160 932.000 163.165 ;
        RECT 736.730 159.915 933.270 163.160 ;
        RECT 736.730 153.865 933.270 158.315 ;
        RECT 736.730 143.265 933.270 152.265 ;
        RECT 736.730 137.415 933.270 141.665 ;
        RECT 736.730 131.565 933.270 135.815 ;
        RECT 736.730 105.015 933.270 129.965 ;
      LAYER met5 ;
        RECT 934.870 103.415 1009.130 181.715 ;
      LAYER met5 ;
        RECT 1010.730 175.665 1207.270 180.115 ;
        RECT 1010.730 169.615 1207.270 174.065 ;
        RECT 1010.730 164.765 1207.270 168.015 ;
      LAYER met5 ;
        RECT 1208.870 163.165 1278.130 181.715 ;
      LAYER met5 ;
        RECT 1279.730 175.665 1476.270 180.115 ;
        RECT 1279.730 169.615 1476.270 174.065 ;
        RECT 1279.730 164.765 1476.270 168.015 ;
        RECT 1012.000 163.160 1206.000 163.165 ;
      LAYER met5 ;
        RECT 1206.000 163.160 1281.000 163.165 ;
      LAYER met5 ;
        RECT 1281.000 163.160 1475.000 163.165 ;
        RECT 1010.730 159.915 1207.270 163.160 ;
        RECT 1010.730 153.865 1207.270 158.315 ;
        RECT 1010.730 143.265 1207.270 152.265 ;
        RECT 1010.730 137.415 1207.270 141.665 ;
        RECT 1010.730 131.565 1207.270 135.815 ;
        RECT 1010.730 105.015 1207.270 129.965 ;
      LAYER met5 ;
        RECT 1208.870 103.415 1278.130 163.160 ;
      LAYER met5 ;
        RECT 1279.730 159.915 1476.270 163.160 ;
        RECT 1279.730 153.865 1476.270 158.315 ;
        RECT 1279.730 143.265 1476.270 152.265 ;
        RECT 1279.730 137.415 1476.270 141.665 ;
        RECT 1279.730 131.565 1476.270 135.815 ;
        RECT 1279.730 105.015 1476.270 129.965 ;
      LAYER met5 ;
        RECT 1477.870 103.415 1552.130 181.715 ;
      LAYER met5 ;
        RECT 1553.730 175.665 1750.270 180.115 ;
        RECT 1553.730 169.615 1750.270 174.065 ;
        RECT 1553.730 164.765 1750.270 168.015 ;
        RECT 1555.000 163.160 1749.000 163.165 ;
        RECT 1553.730 159.915 1750.270 163.160 ;
        RECT 1553.730 153.865 1750.270 158.315 ;
        RECT 1553.730 143.265 1750.270 152.265 ;
        RECT 1553.730 137.415 1750.270 141.665 ;
        RECT 1553.730 131.565 1750.270 135.815 ;
        RECT 1553.730 105.015 1750.270 129.965 ;
      LAYER met5 ;
        RECT 1751.870 103.415 1826.130 181.715 ;
      LAYER met5 ;
        RECT 1827.730 175.665 2024.270 180.115 ;
        RECT 1827.730 169.615 2024.270 174.065 ;
        RECT 1827.730 164.765 2024.270 168.015 ;
        RECT 1829.000 163.160 2023.000 163.165 ;
        RECT 1827.730 159.915 2024.270 163.160 ;
        RECT 1827.730 153.865 2024.270 158.315 ;
        RECT 1827.730 143.265 2024.270 152.265 ;
        RECT 1827.730 137.415 2024.270 141.665 ;
        RECT 1827.730 131.565 2024.270 135.815 ;
        RECT 1827.730 105.015 2024.270 129.965 ;
      LAYER met5 ;
        RECT 2025.870 103.415 2100.130 181.715 ;
      LAYER met5 ;
        RECT 2101.730 175.665 2298.270 180.115 ;
        RECT 2101.730 169.615 2298.270 174.065 ;
        RECT 2101.730 164.765 2298.270 168.015 ;
        RECT 2103.000 163.160 2297.000 163.165 ;
        RECT 2101.730 159.915 2298.270 163.160 ;
        RECT 2101.730 153.865 2298.270 158.315 ;
        RECT 2101.730 143.265 2298.270 152.265 ;
        RECT 2101.730 137.415 2298.270 141.665 ;
        RECT 2101.730 131.565 2298.270 135.815 ;
        RECT 2101.730 105.015 2298.270 129.965 ;
      LAYER met5 ;
        RECT 2299.870 103.415 2374.130 181.715 ;
      LAYER met5 ;
        RECT 2375.730 175.665 2572.270 180.115 ;
        RECT 2375.730 169.615 2572.270 174.065 ;
        RECT 2375.730 164.765 2572.270 168.015 ;
        RECT 2377.000 163.160 2571.000 163.165 ;
        RECT 2375.730 159.915 2572.270 163.160 ;
        RECT 2375.730 153.865 2572.270 158.315 ;
        RECT 2375.730 143.265 2572.270 152.265 ;
        RECT 2375.730 137.415 2572.270 141.665 ;
        RECT 2375.730 131.565 2572.270 135.815 ;
        RECT 2375.730 105.015 2572.270 129.965 ;
      LAYER met5 ;
        RECT 2573.870 103.415 2648.130 181.715 ;
      LAYER met5 ;
        RECT 2649.730 175.665 2846.270 180.115 ;
        RECT 2649.730 169.615 2846.270 174.065 ;
        RECT 2649.730 164.765 2846.270 168.015 ;
      LAYER met5 ;
        RECT 2847.870 163.165 2917.130 181.715 ;
      LAYER met5 ;
        RECT 2918.730 175.665 3115.270 180.115 ;
        RECT 2918.730 169.615 3115.270 174.065 ;
        RECT 2918.730 164.765 3115.270 168.015 ;
      LAYER met5 ;
        RECT 3116.870 163.165 3186.130 181.715 ;
      LAYER met5 ;
        RECT 3187.730 175.665 3385.270 180.115 ;
      LAYER met5 ;
        RECT 3386.870 175.245 3434.135 181.715 ;
      LAYER met5 ;
        RECT 3435.735 176.845 3444.735 345.000 ;
        RECT 3446.335 198.375 3450.585 501.270 ;
        RECT 3452.185 198.520 3456.435 501.270 ;
        RECT 3458.035 197.355 3482.985 501.270 ;
      LAYER met5 ;
        RECT 3484.585 500.000 3588.000 502.870 ;
      LAYER met5 ;
        RECT 3563.785 200.000 3588.000 500.000 ;
      LAYER met5 ;
        RECT 3452.185 196.775 3456.435 196.920 ;
        RECT 3446.335 195.755 3456.435 196.775 ;
        RECT 3484.585 195.755 3588.000 200.000 ;
        RECT 3446.335 175.245 3588.000 195.755 ;
      LAYER met5 ;
        RECT 3187.730 169.615 3385.270 174.065 ;
        RECT 3187.730 164.765 3385.270 168.015 ;
        RECT 2651.000 163.160 2845.000 163.165 ;
      LAYER met5 ;
        RECT 2845.000 163.160 2920.000 163.165 ;
      LAYER met5 ;
        RECT 2920.000 163.160 3114.000 163.165 ;
      LAYER met5 ;
        RECT 3114.000 163.160 3189.000 163.165 ;
      LAYER met5 ;
        RECT 3189.000 163.160 3384.000 163.165 ;
        RECT 2649.730 159.915 2846.270 163.160 ;
        RECT 2649.730 153.865 2846.270 158.315 ;
        RECT 2649.730 143.265 2846.270 152.265 ;
        RECT 2649.730 137.415 2846.270 141.665 ;
        RECT 2649.730 131.565 2846.270 135.815 ;
        RECT 2649.730 105.015 2846.270 129.965 ;
      LAYER met5 ;
        RECT 2847.870 103.415 2917.130 163.160 ;
      LAYER met5 ;
        RECT 2918.730 159.915 3115.270 163.160 ;
        RECT 2918.730 153.865 3115.270 158.315 ;
        RECT 2918.730 143.265 3115.270 152.265 ;
        RECT 2918.730 137.415 3115.270 141.665 ;
        RECT 2918.730 131.565 3115.270 135.815 ;
        RECT 2918.730 105.015 3115.270 129.965 ;
      LAYER met5 ;
        RECT 3116.870 103.415 3186.130 163.160 ;
      LAYER met5 ;
        RECT 3187.730 159.915 3385.270 163.160 ;
        RECT 3187.730 153.865 3385.270 158.315 ;
      LAYER met5 ;
        RECT 3386.870 153.865 3588.000 175.245 ;
      LAYER met5 ;
        RECT 3187.730 143.265 3411.155 152.265 ;
      LAYER met5 ;
        RECT 3412.755 141.665 3588.000 153.865 ;
      LAYER met5 ;
        RECT 3187.730 137.415 3385.270 141.665 ;
        RECT 3187.730 131.565 3385.270 135.815 ;
      LAYER met5 ;
        RECT 3386.870 131.565 3588.000 141.665 ;
      LAYER met5 ;
        RECT 3187.730 105.015 3385.855 129.965 ;
      LAYER met5 ;
        RECT 3387.455 103.415 3588.000 131.565 ;
        RECT 0.000 0.000 200.000 103.415 ;
        RECT 394.000 96.480 469.000 103.415 ;
        RECT 394.000 32.455 399.510 96.480 ;
        RECT 463.550 32.455 469.000 96.480 ;
      LAYER met5 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met5 ;
        RECT 394.000 0.000 469.000 32.455 ;
        RECT 663.000 93.145 738.000 103.415 ;
        RECT 663.000 34.115 681.965 93.145 ;
        RECT 722.350 34.115 738.000 93.145 ;
        RECT 663.000 25.815 738.000 34.115 ;
        RECT 932.000 97.040 1012.000 103.415 ;
        RECT 932.000 31.390 936.600 97.040 ;
        RECT 1002.500 31.390 1012.000 97.040 ;
      LAYER met5 ;
        RECT 469.000 0.000 664.270 24.215 ;
      LAYER met5 ;
        RECT 665.870 0.000 735.130 25.815 ;
      LAYER met5 ;
        RECT 736.730 0.000 932.000 24.215 ;
      LAYER met5 ;
        RECT 932.000 0.000 1012.000 31.390 ;
        RECT 1206.000 99.700 1281.000 103.415 ;
        RECT 1206.000 29.235 1214.730 99.700 ;
        RECT 1272.330 29.235 1281.000 99.700 ;
      LAYER met5 ;
        RECT 1012.000 0.000 1206.000 24.215 ;
      LAYER met5 ;
        RECT 1206.000 0.000 1281.000 29.235 ;
        RECT 1475.000 97.040 1555.000 103.415 ;
        RECT 1475.000 31.390 1479.600 97.040 ;
        RECT 1545.500 31.390 1555.000 97.040 ;
      LAYER met5 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met5 ;
        RECT 1475.000 0.000 1555.000 31.390 ;
        RECT 1749.000 97.040 1829.000 103.415 ;
        RECT 1749.000 31.390 1753.600 97.040 ;
        RECT 1819.500 31.390 1829.000 97.040 ;
      LAYER met5 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met5 ;
        RECT 1749.000 0.000 1829.000 31.390 ;
        RECT 2023.000 97.040 2103.000 103.415 ;
        RECT 2023.000 31.390 2027.600 97.040 ;
        RECT 2093.500 31.390 2103.000 97.040 ;
      LAYER met5 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met5 ;
        RECT 2023.000 0.000 2103.000 31.390 ;
        RECT 2297.000 97.040 2377.000 103.415 ;
        RECT 2297.000 31.390 2301.600 97.040 ;
        RECT 2367.500 31.390 2377.000 97.040 ;
      LAYER met5 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met5 ;
        RECT 2297.000 0.000 2377.000 31.390 ;
        RECT 2571.000 97.040 2651.000 103.415 ;
        RECT 2571.000 31.390 2575.600 97.040 ;
        RECT 2641.500 31.390 2651.000 97.040 ;
      LAYER met5 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met5 ;
        RECT 2571.000 0.000 2651.000 31.390 ;
        RECT 2845.000 96.480 2920.000 103.415 ;
        RECT 2845.000 32.455 2850.510 96.480 ;
        RECT 2914.550 32.455 2920.000 96.480 ;
      LAYER met5 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met5 ;
        RECT 2845.000 0.000 2920.000 32.455 ;
        RECT 3114.000 96.480 3189.000 103.415 ;
        RECT 3114.000 32.455 3119.510 96.480 ;
        RECT 3183.550 32.455 3189.000 96.480 ;
      LAYER met5 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met5 ;
        RECT 3114.000 0.000 3189.000 32.455 ;
      LAYER met5 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met5 ;
        RECT 3384.000 0.000 3588.000 103.415 ;
  END
END chip_io_alt
END LIBRARY

