magic
tech sky130A
magscale 1 2
timestamp 1623348572
<< nwell >>
rect 11772 9130 23593 9434
<< pwell >>
rect 10099 9180 11657 13751
<< obsli1 >>
rect 9522 9400 23971 48932
rect 9522 9206 11631 9400
rect 11807 9377 12009 9400
rect 23346 9377 23536 9400
rect 11807 9187 23536 9377
<< obsm1 >>
rect 9437 9400 23983 48938
rect 10125 9219 11171 9400
rect 11807 9377 12070 9400
tri 12070 9377 12093 9400 sw
tri 23285 9377 23308 9400 se
rect 23308 9377 23536 9400
rect 11807 9187 23536 9377
<< metal2 >>
rect 9499 8993 14279 9404
rect 19478 8993 24258 14125
<< obsm2 >>
rect 9453 14181 24258 48008
rect 9453 9460 19422 14181
rect 14335 9400 19422 9460
rect 14579 8993 14979 9377
<< metal3 >>
rect 0 8993 14279 12130
rect 14579 8993 16779 9538
rect 16978 8993 19178 11259
rect 19478 8993 33800 12130
<< obsm3 >>
rect 0 12210 33800 48993
rect 0 12130 4307 12210
rect 14359 11339 19398 12210
rect 14359 9618 16898 11339
rect 14359 9538 14499 9618
rect 16859 9538 16898 9618
rect 19258 9538 19398 11339
<< metal4 >>
rect 0 44150 9641 48993
rect 25649 44150 33800 48993
rect 0 23000 9543 27993
rect 25177 23000 33800 27993
rect 0 21810 9543 22700
rect 25177 21810 33800 22700
rect 0 20640 9543 21530
rect 25177 20640 33800 21530
rect 0 20274 33800 20340
rect 0 19618 33800 20214
rect 0 19322 9448 19558
rect 25177 19322 33800 19558
rect 0 18666 33800 19262
rect 0 18540 33800 18606
rect 0 17310 9450 18240
rect 25177 17310 33800 18240
rect 0 16340 9543 17030
rect 25177 16340 33800 17030
rect 0 15370 9543 16060
rect 25177 15370 33800 16060
rect 0 14160 9543 15090
rect 25177 14160 33800 15090
rect 0 12950 9543 13880
rect 24241 12950 33800 13880
rect 0 11980 9543 12670
rect 24241 11980 33800 12670
rect 0 10770 9543 11700
rect 25177 10770 33800 11700
rect 0 9400 9543 10490
rect 25177 9400 33800 10490
<< obsm4 >>
rect 9721 44070 25569 48993
rect 9448 28073 25649 44070
rect 9623 22920 25097 28073
rect 9448 22780 25649 22920
rect 9623 21730 25097 22780
rect 9448 21610 25649 21730
rect 9623 20560 25097 21610
rect 9448 20420 25649 20560
rect 9528 19342 25097 19538
rect 9448 18320 25649 18460
rect 9530 17230 25097 18320
rect 9448 17110 25649 17230
rect 9623 16260 25097 17110
rect 9448 16140 25649 16260
rect 9623 15290 25097 16140
rect 9448 15170 25649 15290
rect 9623 14080 25097 15170
rect 9448 13960 25649 14080
rect 9623 12870 24161 13960
rect 9448 12750 25649 12870
rect 9623 11900 24161 12750
rect 9448 11780 25649 11900
rect 9623 10690 25097 11780
rect 9448 10570 25649 10690
rect 9623 9400 25097 10570
<< metal5 >>
rect 10810 30017 22978 42182
rect 0 23000 9543 27990
rect 0 21830 9543 22680
rect 0 20660 9543 21510
rect 25177 23000 33800 27990
rect 25177 21830 33800 22680
rect 25177 20660 33800 21510
rect 0 18540 9448 20340
rect 25177 18540 33800 20340
rect 0 17330 9543 18220
rect 0 16360 9543 17010
rect 0 15390 9543 16040
rect 0 14180 9543 15070
rect 0 12970 9543 13860
rect 25177 17330 33800 18220
rect 25177 16360 33800 17010
rect 25177 15390 33800 16040
rect 25177 14180 33800 15070
rect 25177 12970 33800 13860
rect 0 12000 9543 12650
rect 24241 12000 33800 12650
rect 0 10790 9543 11680
rect 0 9420 9543 10470
rect 25177 10790 33800 11680
rect 25177 9420 33800 10470
<< obsm5 >>
rect 0 42502 33800 48993
rect 0 29697 10490 42502
rect 23298 29697 33800 42502
rect 0 28310 33800 29697
rect 9863 20340 24857 28310
rect 9768 18540 24857 20340
rect 9863 12970 24857 18540
rect 9863 11680 23921 12970
rect 9863 9420 24857 11680
<< labels >>
rlabel metal4 s 0 19618 33800 20214 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 19618 254 20214 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 18666 33800 19262 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal4 s 0 18666 254 19262 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal2 s 19478 8993 24258 14125 6 DRN_HVC
port 3 nsew power bidirectional
rlabel metal3 s 16978 8993 19178 11259 6 DRN_HVC
port 3 nsew power bidirectional
rlabel metal3 s 0 8993 14279 12130 6 P_CORE
port 4 nsew power bidirectional
rlabel metal3 s 19478 8993 33800 12130 6 P_CORE
port 4 nsew power bidirectional
rlabel metal5 s 10810 30017 22978 42182 6 P_PAD
port 5 nsew power bidirectional
rlabel metal2 s 9499 8993 14279 9404 6 SRC_BDY_HVC
port 6 nsew ground bidirectional
rlabel metal3 s 14579 8993 16779 9538 6 SRC_BDY_HVC
port 6 nsew ground bidirectional
rlabel metal5 s 25177 18540 33800 20340 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 25177 16360 33800 17010 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 25177 19322 33800 19558 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 20274 33800 20340 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 18540 33800 18606 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 25177 16340 33800 17030 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 18540 9448 20340 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 16360 9543 17010 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 18540 254 18606 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 19322 9448 19558 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 20274 254 20340 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 16340 9543 17030 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 24241 12000 33800 12650 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 24241 11980 33800 12670 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 12000 9543 12650 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 11980 9543 12670 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 25177 15390 33800 16040 6 VSWITCH
port 9 nsew power bidirectional
rlabel metal4 s 25177 15370 33800 16060 6 VSWITCH
port 9 nsew power bidirectional
rlabel metal5 s 0 15390 9543 16040 6 VSWITCH
port 9 nsew power bidirectional
rlabel metal4 s 0 15370 9543 16060 6 VSWITCH
port 9 nsew power bidirectional
rlabel metal5 s 25177 21830 33800 22680 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 25177 21810 33800 22700 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 0 21830 9543 22680 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 0 21810 9543 22700 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 25177 9420 33800 10470 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 25177 9400 33800 10490 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal5 s 0 9420 9543 10470 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 0 9400 9543 10490 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal5 s 25177 23000 33800 27990 6 VDDIO
port 12 nsew power bidirectional
rlabel metal5 s 25177 12970 33800 13860 6 VDDIO
port 12 nsew power bidirectional
rlabel metal4 s 24241 12950 33800 13880 6 VDDIO
port 12 nsew power bidirectional
rlabel metal4 s 25177 23000 33800 27993 6 VDDIO
port 12 nsew power bidirectional
rlabel metal5 s 0 23000 9543 27990 6 VDDIO
port 12 nsew power bidirectional
rlabel metal5 s 0 12970 9543 13860 6 VDDIO
port 12 nsew power bidirectional
rlabel metal4 s 0 12950 9543 13880 6 VDDIO
port 12 nsew power bidirectional
rlabel metal4 s 0 23000 9543 27993 6 VDDIO
port 12 nsew power bidirectional
rlabel metal5 s 25177 10790 33800 11680 6 VCCD
port 13 nsew power bidirectional
rlabel metal4 s 25177 10770 33800 11700 6 VCCD
port 13 nsew power bidirectional
rlabel metal5 s 0 10790 9543 11680 6 VCCD
port 13 nsew power bidirectional
rlabel metal4 s 0 10770 9543 11700 6 VCCD
port 13 nsew power bidirectional
rlabel metal4 s 25649 44150 33800 48993 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 33672 47313 33674 47315 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal5 s 25177 14180 33800 15070 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 25177 14160 33800 15090 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 33546 44150 33800 48993 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 0 44150 9641 48993 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 126 47313 128 47315 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal5 s 0 14180 9543 15070 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 0 44150 254 48993 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 0 14160 9543 15090 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal5 s 25177 17330 33800 18220 6 VSSD
port 15 nsew ground bidirectional
rlabel metal4 s 25177 17310 33800 18240 6 VSSD
port 15 nsew ground bidirectional
rlabel metal5 s 0 17330 9543 18220 6 VSSD
port 15 nsew ground bidirectional
rlabel metal4 s 0 17310 9450 18240 6 VSSD
port 15 nsew ground bidirectional
rlabel metal5 s 25177 20660 33800 21510 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal4 s 25177 20640 33800 21530 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal5 s 0 20660 9543 21510 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal4 s 0 20640 9543 21530 6 VSSIO_Q
port 16 nsew ground bidirectional
<< properties >>
string LEFclass PAD POWER
string FIXED_BBOX 0 9400 33800 48993
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_END 1824342
string GDS_START 1807708
<< end >>
