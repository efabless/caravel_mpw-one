magic
tech sky130A
magscale 1 2
timestamp 1607567185
<< checkpaint >>
rect -2854 -2865 202770 13745
<< locali >>
rect 94329 9911 94363 10557
rect 143549 9979 143583 10149
rect 143399 9945 143457 9979
rect 153117 9911 153151 10149
rect 153209 9979 153243 10149
rect 157993 9911 158027 10149
rect 103253 8347 103287 8585
rect 101965 7259 101999 7497
rect 157165 7497 157533 7531
rect 130117 7259 130151 7429
rect 110429 6715 110463 6885
rect 110521 6715 110555 6817
rect 157165 6715 157199 7497
rect 161799 7361 162041 7395
rect 181729 7361 182005 7395
rect 181729 7327 181763 7361
rect 107669 6239 107703 6409
rect 74733 6103 74767 6205
rect 118801 6103 118835 6341
rect 96445 5151 96479 5321
rect 99573 5015 99607 5253
rect 87061 4539 87095 4641
rect 106657 4607 106691 4709
rect 119905 4471 119939 4709
rect 144193 4607 144227 4709
rect 124505 4063 124539 4165
rect 114477 3927 114511 4029
rect 130393 3927 130427 4029
rect 121929 3383 121963 3621
rect 138581 3451 138615 3621
rect 4445 2839 4479 3009
rect 156981 2907 157015 3349
rect 157073 2907 157107 3009
rect 157257 2975 157291 3145
rect 157257 2941 157441 2975
rect 157625 2907 157659 2941
rect 157383 2873 157659 2907
rect 162627 2941 162961 2975
rect 161305 2839 161339 2941
rect 164559 2873 164835 2907
rect 156923 2805 157533 2839
rect 164801 2839 164835 2873
rect 152473 1751 152507 1853
rect 163789 1751 163823 1921
rect 193137 1343 193171 1445
rect 140973 1207 141007 1309
rect 144963 969 145021 1003
rect 129841 595 129875 765
rect 133245 663 133279 901
rect 135119 697 135269 731
rect 137569 323 137603 969
rect 140789 391 140823 561
rect 141893 391 141927 833
rect 143733 595 143767 901
rect 145055 765 146033 799
rect 149805 731 149839 901
rect 161857 323 161891 425
rect 161949 323 161983 901
rect 165997 731 166031 969
rect 182189 799 182223 901
rect 166825 255 166859 493
<< viali >>
rect 94329 10557 94363 10591
rect 143549 10149 143583 10183
rect 143365 9945 143399 9979
rect 143457 9945 143491 9979
rect 143549 9945 143583 9979
rect 153117 10149 153151 10183
rect 94329 9877 94363 9911
rect 153209 10149 153243 10183
rect 153209 9945 153243 9979
rect 157993 10149 158027 10183
rect 153117 9877 153151 9911
rect 157993 9877 158027 9911
rect 3065 9673 3099 9707
rect 156705 9605 156739 9639
rect 165261 9605 165295 9639
rect 171333 9605 171367 9639
rect 182741 9605 182775 9639
rect 185593 9605 185627 9639
rect 194149 9605 194183 9639
rect 196633 9605 196667 9639
rect 5457 9537 5491 9571
rect 7941 9537 7975 9571
rect 16497 9537 16531 9571
rect 45017 9537 45051 9571
rect 69857 9537 69891 9571
rect 81449 9537 81483 9571
rect 94329 9537 94363 9571
rect 101045 9537 101079 9571
rect 111441 9537 111475 9571
rect 113925 9537 113959 9571
rect 119629 9537 119663 9571
rect 121009 9537 121043 9571
rect 125517 9537 125551 9571
rect 128553 9537 128587 9571
rect 129565 9537 129599 9571
rect 130577 9537 130611 9571
rect 141985 9537 142019 9571
rect 151277 9537 151311 9571
rect 153853 9537 153887 9571
rect 158821 9537 158855 9571
rect 159833 9537 159867 9571
rect 168113 9537 168147 9571
rect 173817 9537 173851 9571
rect 176945 9537 176979 9571
rect 181269 9537 181303 9571
rect 186881 9537 186915 9571
rect 188353 9537 188387 9571
rect 190929 9537 190963 9571
rect 195161 9537 195195 9571
rect 2973 9469 3007 9503
rect 4445 9469 4479 9503
rect 5549 9469 5583 9503
rect 6929 9469 6963 9503
rect 8033 9469 8067 9503
rect 15485 9469 15519 9503
rect 17049 9469 17083 9503
rect 44005 9469 44039 9503
rect 45109 9469 45143 9503
rect 61301 9469 61335 9503
rect 61485 9469 61519 9503
rect 61669 9469 61703 9503
rect 67557 9469 67591 9503
rect 81357 9469 81391 9503
rect 81817 9469 81851 9503
rect 91293 9469 91327 9503
rect 92857 9469 92891 9503
rect 94421 9469 94455 9503
rect 95617 9469 95651 9503
rect 95709 9469 95743 9503
rect 96077 9469 96111 9503
rect 104909 9469 104943 9503
rect 107485 9469 107519 9503
rect 109969 9469 110003 9503
rect 111533 9469 111567 9503
rect 112453 9469 112487 9503
rect 114017 9469 114051 9503
rect 118157 9469 118191 9503
rect 119721 9469 119755 9503
rect 122757 9469 122791 9503
rect 124137 9469 124171 9503
rect 125241 9469 125275 9503
rect 127081 9469 127115 9503
rect 128645 9469 128679 9503
rect 131129 9469 131163 9503
rect 144837 9469 144871 9503
rect 152381 9469 152415 9503
rect 153485 9469 153519 9503
rect 155233 9469 155267 9503
rect 156337 9469 156371 9503
rect 163789 9469 163823 9503
rect 164893 9469 164927 9503
rect 166641 9469 166675 9503
rect 167745 9469 167779 9503
rect 169861 9469 169895 9503
rect 171425 9469 171459 9503
rect 172345 9469 172379 9503
rect 173725 9469 173759 9503
rect 175473 9469 175507 9503
rect 177037 9469 177071 9503
rect 178785 9469 178819 9503
rect 182833 9469 182867 9503
rect 184121 9469 184155 9503
rect 185685 9469 185719 9503
rect 188445 9469 188479 9503
rect 189457 9469 189491 9503
rect 191021 9469 191055 9503
rect 192677 9469 192711 9503
rect 194241 9469 194275 9503
rect 196725 9469 196759 9503
rect 68569 9401 68603 9435
rect 74181 9401 74215 9435
rect 86785 9401 86819 9435
rect 89637 9401 89671 9435
rect 102057 9401 102091 9435
rect 132417 9401 132451 9435
rect 136281 9401 136315 9435
rect 140973 9401 141007 9435
rect 162685 9401 162719 9435
rect 12633 9333 12667 9367
rect 27537 9333 27571 9367
rect 42717 9333 42751 9367
rect 46857 9333 46891 9367
rect 47869 9333 47903 9367
rect 59829 9333 59863 9367
rect 62681 9333 62715 9367
rect 64705 9333 64739 9367
rect 65717 9333 65751 9367
rect 70961 9333 70995 9367
rect 73077 9333 73111 9367
rect 75377 9333 75411 9367
rect 76389 9333 76423 9367
rect 78229 9333 78263 9367
rect 79701 9333 79735 9367
rect 82645 9333 82679 9367
rect 83933 9333 83967 9367
rect 84945 9333 84979 9367
rect 87797 9333 87831 9367
rect 96905 9333 96939 9367
rect 98193 9333 98227 9367
rect 99205 9333 99239 9367
rect 103897 9333 103931 9367
rect 108497 9333 108531 9367
rect 115305 9333 115339 9367
rect 116317 9333 116351 9367
rect 133429 9333 133463 9367
rect 135269 9333 135303 9367
rect 138121 9333 138155 9367
rect 139133 9333 139167 9367
rect 143825 9333 143859 9367
rect 146677 9333 146711 9367
rect 147689 9333 147723 9367
rect 149529 9333 149563 9367
rect 161673 9333 161707 9367
rect 179797 9333 179831 9367
rect 2973 9129 3007 9163
rect 7113 9129 7147 9163
rect 15301 9129 15335 9163
rect 62773 9129 62807 9163
rect 86785 9129 86819 9163
rect 105645 9129 105679 9163
rect 152105 9129 152139 9163
rect 160109 9129 160143 9163
rect 179613 9129 179647 9163
rect 197369 9129 197403 9163
rect 88257 9061 88291 9095
rect 5917 8993 5951 9027
rect 7021 8993 7055 9027
rect 11253 8993 11287 9027
rect 12357 8993 12391 9027
rect 17417 8993 17451 9027
rect 27905 8993 27939 9027
rect 29009 8993 29043 9027
rect 38853 8993 38887 9027
rect 40877 8993 40911 9027
rect 42441 8993 42475 9027
rect 44833 8993 44867 9027
rect 47317 8993 47351 9027
rect 56241 8993 56275 9027
rect 60473 8993 60507 9027
rect 60933 8993 60967 9027
rect 71421 8993 71455 9027
rect 72157 8993 72191 9027
rect 73721 8993 73755 9027
rect 75285 8993 75319 9027
rect 77033 8993 77067 9027
rect 77769 8993 77803 9027
rect 79517 8993 79551 9027
rect 80253 8993 80287 9027
rect 85957 8993 85991 9027
rect 91753 8993 91787 9027
rect 92213 8993 92247 9027
rect 96905 8993 96939 9027
rect 97917 8993 97951 9027
rect 98469 8993 98503 9027
rect 107945 8993 107979 9027
rect 108221 8993 108255 9027
rect 110981 8993 111015 9027
rect 111257 8993 111291 9027
rect 114477 8993 114511 9027
rect 119721 8993 119755 9027
rect 123033 8993 123067 9027
rect 124413 8993 124447 9027
rect 125977 8993 126011 9027
rect 128461 8993 128495 9027
rect 129565 8993 129599 9027
rect 134533 8993 134567 9027
rect 135637 8993 135671 9027
rect 136925 8993 136959 9027
rect 139869 8993 139903 9027
rect 143181 8993 143215 9027
rect 144377 8993 144411 9027
rect 145481 8993 145515 9027
rect 147873 8993 147907 9027
rect 154221 8993 154255 9027
rect 156705 8993 156739 9027
rect 164249 8993 164283 9027
rect 167469 8993 167503 9027
rect 169033 8993 169067 9027
rect 169953 8993 169987 9027
rect 171241 8993 171275 9027
rect 174921 8993 174955 9027
rect 182005 8993 182039 9027
rect 186237 8993 186271 9027
rect 190653 8993 190687 9027
rect 191941 8993 191975 9027
rect 193045 8993 193079 9027
rect 196449 8993 196483 9027
rect 197277 8993 197311 9027
rect 4629 8925 4663 8959
rect 5825 8925 5859 8959
rect 8033 8925 8067 8959
rect 12265 8925 12299 8959
rect 14197 8925 14231 8959
rect 16313 8925 16347 8959
rect 17325 8925 17359 8959
rect 21373 8925 21407 8959
rect 26893 8925 26927 8959
rect 29377 8925 29411 8959
rect 32137 8925 32171 8959
rect 33149 8925 33183 8959
rect 37749 8925 37783 8959
rect 39221 8925 39255 8959
rect 42349 8925 42383 8959
rect 43729 8925 43763 8959
rect 46121 8925 46155 8959
rect 47133 8925 47167 8959
rect 48973 8925 49007 8959
rect 55137 8925 55171 8959
rect 56149 8925 56183 8959
rect 59093 8925 59127 8959
rect 60565 8925 60599 8959
rect 61761 8925 61795 8959
rect 63785 8925 63819 8959
rect 65993 8925 66027 8959
rect 67005 8925 67039 8959
rect 68017 8925 68051 8959
rect 69305 8925 69339 8959
rect 70317 8925 70351 8959
rect 71789 8925 71823 8959
rect 75193 8925 75227 8959
rect 77401 8925 77435 8959
rect 81081 8925 81115 8959
rect 82645 8925 82679 8959
rect 84393 8925 84427 8959
rect 85865 8925 85899 8959
rect 89269 8925 89303 8959
rect 90373 8925 90407 8959
rect 91845 8925 91879 8959
rect 93869 8925 93903 8959
rect 95341 8925 95375 8959
rect 96813 8925 96847 8959
rect 98101 8925 98135 8959
rect 99481 8925 99515 8959
rect 100493 8925 100527 8959
rect 102057 8925 102091 8959
rect 103069 8925 103103 8959
rect 106657 8925 106691 8959
rect 109601 8925 109635 8959
rect 113005 8925 113039 8959
rect 114385 8925 114419 8959
rect 117145 8925 117179 8959
rect 118157 8925 118191 8959
rect 120549 8925 120583 8959
rect 121929 8925 121963 8959
rect 130853 8925 130887 8959
rect 131865 8925 131899 8959
rect 133153 8925 133187 8959
rect 138765 8925 138799 8959
rect 141157 8925 141191 8959
rect 142169 8925 142203 8959
rect 145849 8925 145883 8959
rect 146769 8925 146803 8959
rect 149989 8925 150023 8959
rect 151093 8925 151127 8959
rect 153117 8925 153151 8959
rect 154497 8925 154531 8959
rect 155601 8925 155635 8959
rect 157993 8925 158027 8959
rect 159097 8925 159131 8959
rect 161949 8925 161983 8959
rect 162961 8925 162995 8959
rect 165353 8925 165387 8959
rect 171425 8925 171459 8959
rect 172805 8925 172839 8959
rect 173817 8925 173851 8959
rect 176853 8925 176887 8959
rect 178049 8925 178083 8959
rect 180625 8925 180659 8959
rect 183661 8925 183695 8959
rect 184857 8925 184891 8959
rect 188169 8925 188203 8959
rect 189549 8925 189583 8959
rect 191021 8925 191055 8959
rect 192953 8925 192987 8959
rect 194885 8925 194919 8959
rect 196081 8925 196115 8959
rect 45017 8857 45051 8891
rect 119629 8857 119663 8891
rect 123401 8857 123435 8891
rect 125885 8857 125919 8891
rect 129749 8857 129783 8891
rect 136005 8857 136039 8891
rect 140237 8857 140271 8891
rect 148241 8857 148275 8891
rect 157073 8857 157107 8891
rect 164433 8857 164467 8891
rect 168941 8857 168975 8891
rect 175289 8857 175323 8891
rect 182097 8857 182131 8891
rect 186145 8857 186179 8891
rect 79609 8789 79643 8823
rect 107761 8789 107795 8823
rect 110797 8789 110831 8823
rect 87061 8585 87095 8619
rect 103253 8585 103287 8619
rect 105921 8585 105955 8619
rect 192125 8585 192159 8619
rect 196081 8585 196115 8619
rect 26433 8517 26467 8551
rect 30757 8517 30791 8551
rect 82185 8517 82219 8551
rect 100401 8517 100435 8551
rect 3341 8449 3375 8483
rect 5549 8449 5583 8483
rect 6837 8449 6871 8483
rect 7849 8449 7883 8483
rect 14381 8449 14415 8483
rect 15393 8449 15427 8483
rect 16773 8449 16807 8483
rect 20453 8449 20487 8483
rect 21465 8449 21499 8483
rect 29285 8449 29319 8483
rect 31953 8449 31987 8483
rect 33241 8449 33275 8483
rect 37749 8449 37783 8483
rect 39129 8449 39163 8483
rect 40969 8449 41003 8483
rect 42993 8449 43027 8483
rect 46121 8449 46155 8483
rect 47593 8449 47627 8483
rect 48605 8449 48639 8483
rect 55689 8449 55723 8483
rect 59553 8449 59587 8483
rect 60841 8449 60875 8483
rect 62957 8449 62991 8483
rect 66085 8449 66119 8483
rect 67097 8449 67131 8483
rect 76941 8449 76975 8483
rect 80713 8449 80747 8483
rect 83565 8449 83599 8483
rect 93685 8449 93719 8483
rect 95065 8449 95099 8483
rect 4353 8381 4387 8415
rect 5641 8381 5675 8415
rect 7941 8381 7975 8415
rect 15485 8381 15519 8415
rect 21557 8381 21591 8415
rect 24961 8381 24995 8415
rect 26065 8381 26099 8415
rect 30389 8381 30423 8415
rect 33057 8381 33091 8415
rect 36737 8381 36771 8415
rect 37841 8381 37875 8415
rect 41981 8381 42015 8415
rect 43545 8381 43579 8415
rect 48697 8381 48731 8415
rect 54677 8381 54711 8415
rect 55781 8381 55815 8415
rect 60657 8381 60691 8415
rect 67189 8381 67223 8415
rect 70961 8381 70995 8415
rect 71329 8381 71363 8415
rect 71513 8381 71547 8415
rect 72525 8381 72559 8415
rect 72893 8381 72927 8415
rect 73261 8381 73295 8415
rect 74457 8381 74491 8415
rect 74825 8381 74859 8415
rect 75193 8381 75227 8415
rect 76849 8381 76883 8415
rect 77217 8381 77251 8415
rect 82277 8381 82311 8415
rect 85681 8381 85715 8415
rect 85773 8381 85807 8415
rect 86141 8381 86175 8415
rect 87245 8381 87279 8415
rect 87705 8381 87739 8415
rect 88533 8381 88567 8415
rect 88901 8381 88935 8415
rect 89269 8381 89303 8415
rect 91109 8381 91143 8415
rect 92305 8381 92339 8415
rect 93777 8381 93811 8415
rect 94973 8381 95007 8415
rect 95433 8381 95467 8415
rect 96629 8381 96663 8415
rect 96997 8381 97031 8415
rect 97365 8381 97399 8415
rect 99113 8381 99147 8415
rect 100677 8381 100711 8415
rect 104817 8517 104851 8551
rect 116133 8517 116167 8551
rect 129289 8517 129323 8551
rect 146125 8517 146159 8551
rect 155325 8517 155359 8551
rect 159649 8517 159683 8551
rect 162961 8517 162995 8551
rect 172161 8517 172195 8551
rect 176761 8517 176795 8551
rect 179153 8517 179187 8551
rect 185409 8517 185443 8551
rect 187893 8517 187927 8551
rect 190285 8517 190319 8551
rect 103345 8449 103379 8483
rect 109044 8449 109078 8483
rect 110061 8449 110095 8483
rect 114661 8449 114695 8483
rect 121285 8449 121319 8483
rect 125149 8449 125183 8483
rect 126621 8449 126655 8483
rect 127817 8449 127851 8483
rect 131037 8449 131071 8483
rect 132417 8449 132451 8483
rect 133429 8449 133463 8483
rect 134901 8449 134935 8483
rect 136557 8449 136591 8483
rect 137937 8449 137971 8483
rect 138949 8449 138983 8483
rect 140421 8449 140455 8483
rect 143549 8449 143583 8483
rect 144653 8449 144687 8483
rect 147229 8449 147263 8483
rect 148701 8449 148735 8483
rect 149621 8449 149655 8483
rect 150633 8449 150667 8483
rect 151645 8449 151679 8483
rect 152841 8449 152875 8483
rect 156245 8449 156279 8483
rect 161489 8449 161523 8483
rect 167285 8449 167319 8483
rect 168481 8449 168515 8483
rect 169677 8449 169711 8483
rect 170689 8449 170723 8483
rect 174093 8449 174127 8483
rect 182833 8449 182867 8483
rect 183937 8449 183971 8483
rect 186421 8449 186455 8483
rect 193597 8449 193631 8483
rect 194977 8449 195011 8483
rect 104817 8381 104851 8415
rect 106105 8381 106139 8415
rect 106565 8381 106599 8415
rect 110153 8381 110187 8415
rect 111717 8381 111751 8415
rect 111809 8381 111843 8415
rect 111993 8381 112027 8415
rect 116225 8381 116259 8415
rect 119077 8381 119111 8415
rect 126713 8381 126747 8415
rect 129381 8381 129415 8415
rect 132141 8381 132175 8415
rect 134533 8381 134567 8415
rect 137661 8381 137695 8415
rect 140053 8381 140087 8415
rect 142537 8381 142571 8415
rect 146217 8381 146251 8415
rect 148333 8381 148367 8415
rect 153853 8381 153887 8415
rect 155417 8381 155451 8415
rect 157257 8381 157291 8415
rect 158361 8381 158395 8415
rect 159465 8381 159499 8415
rect 162593 8381 162627 8415
rect 165813 8381 165847 8415
rect 167377 8381 167411 8415
rect 171793 8381 171827 8415
rect 173081 8381 173115 8415
rect 175289 8381 175323 8415
rect 176393 8381 176427 8415
rect 177681 8381 177715 8415
rect 179061 8381 179095 8415
rect 181453 8381 181487 8415
rect 182925 8381 182959 8415
rect 185501 8381 185535 8415
rect 187985 8381 188019 8415
rect 188813 8381 188847 8415
rect 190377 8381 190411 8415
rect 192033 8381 192067 8415
rect 194701 8381 194735 8415
rect 195989 8381 196023 8415
rect 12449 8313 12483 8347
rect 49985 8313 50019 8347
rect 53665 8313 53699 8347
rect 69029 8313 69063 8347
rect 78597 8313 78631 8347
rect 103253 8313 103287 8347
rect 107853 8313 107887 8347
rect 117421 8313 117455 8347
rect 120273 8313 120307 8347
rect 122297 8313 122331 8347
rect 123585 8313 123619 8347
rect 11345 8245 11379 8279
rect 27353 8245 27387 8279
rect 34897 8245 34931 8279
rect 44373 8245 44407 8279
rect 58541 8245 58575 8279
rect 63969 8245 64003 8279
rect 64981 8245 65015 8279
rect 102241 8245 102275 8279
rect 113465 8245 113499 8279
rect 141525 8245 141559 8279
rect 164525 8245 164559 8279
rect 7389 8041 7423 8075
rect 23857 8041 23891 8075
rect 37749 8041 37783 8075
rect 42257 8041 42291 8075
rect 54861 8041 54895 8075
rect 55873 8041 55907 8075
rect 100493 8041 100527 8075
rect 163329 8041 163363 8075
rect 171333 8041 171367 8075
rect 184397 8041 184431 8075
rect 197369 8041 197403 8075
rect 48973 7973 49007 8007
rect 135545 7973 135579 8007
rect 6101 7905 6135 7939
rect 10701 7905 10735 7939
rect 11805 7905 11839 7939
rect 18061 7905 18095 7939
rect 26893 7905 26927 7939
rect 27997 7905 28031 7939
rect 32137 7905 32171 7939
rect 33241 7905 33275 7939
rect 34529 7905 34563 7939
rect 35633 7905 35667 7939
rect 43913 7905 43947 7939
rect 45017 7905 45051 7939
rect 47409 7905 47443 7939
rect 58541 7905 58575 7939
rect 59277 7905 59311 7939
rect 60197 7905 60231 7939
rect 61301 7905 61335 7939
rect 62865 7905 62899 7939
rect 63141 7905 63175 7939
rect 64429 7905 64463 7939
rect 64705 7905 64739 7939
rect 67833 7905 67867 7939
rect 68109 7905 68143 7939
rect 71421 7905 71455 7939
rect 72157 7905 72191 7939
rect 73445 7905 73479 7939
rect 73721 7905 73755 7939
rect 75285 7905 75319 7939
rect 75745 7905 75779 7939
rect 78229 7905 78263 7939
rect 78781 7905 78815 7939
rect 80529 7905 80563 7939
rect 80989 7905 81023 7939
rect 82829 7905 82863 7939
rect 83013 7905 83047 7939
rect 83197 7905 83231 7939
rect 84945 7905 84979 7939
rect 85681 7905 85715 7939
rect 86509 7905 86543 7939
rect 87245 7905 87279 7939
rect 88257 7905 88291 7939
rect 88993 7905 89027 7939
rect 90925 7905 90959 7939
rect 91385 7905 91419 7939
rect 92489 7905 92523 7939
rect 92949 7905 92983 7939
rect 94145 7905 94179 7939
rect 94605 7905 94639 7939
rect 95525 7905 95559 7939
rect 95801 7905 95835 7939
rect 96169 7905 96203 7939
rect 96997 7905 97031 7939
rect 98561 7905 98595 7939
rect 102425 7905 102459 7939
rect 103989 7905 104023 7939
rect 105369 7905 105403 7939
rect 105829 7905 105863 7939
rect 107577 7905 107611 7939
rect 107945 7905 107979 7939
rect 109233 7905 109267 7939
rect 109509 7905 109543 7939
rect 111257 7905 111291 7939
rect 112821 7905 112855 7939
rect 115213 7905 115247 7939
rect 118709 7905 118743 7939
rect 120273 7905 120307 7939
rect 123309 7905 123343 7939
rect 124873 7905 124907 7939
rect 127541 7905 127575 7939
rect 129105 7905 129139 7939
rect 130393 7905 130427 7939
rect 131497 7905 131531 7939
rect 134257 7905 134291 7939
rect 137569 7905 137603 7939
rect 139869 7905 139903 7939
rect 144377 7905 144411 7939
rect 146953 7905 146987 7939
rect 152105 7905 152139 7939
rect 154221 7905 154255 7939
rect 155601 7905 155635 7939
rect 156705 7905 156739 7939
rect 158637 7905 158671 7939
rect 159925 7905 159959 7939
rect 161305 7905 161339 7939
rect 164341 7905 164375 7939
rect 165905 7905 165939 7939
rect 169309 7905 169343 7939
rect 170137 7905 170171 7939
rect 172437 7905 172471 7939
rect 173541 7905 173575 7939
rect 174921 7905 174955 7939
rect 176485 7905 176519 7939
rect 178049 7905 178083 7939
rect 179613 7905 179647 7939
rect 182465 7905 182499 7939
rect 187249 7905 187283 7939
rect 188077 7905 188111 7939
rect 190653 7905 190687 7939
rect 191665 7905 191699 7939
rect 192769 7905 192803 7939
rect 194885 7905 194919 7939
rect 195989 7905 196023 7939
rect 197277 7905 197311 7939
rect 2973 7837 3007 7871
rect 4997 7837 5031 7871
rect 6009 7837 6043 7871
rect 8401 7837 8435 7871
rect 9689 7837 9723 7871
rect 11713 7837 11747 7871
rect 13093 7837 13127 7871
rect 14197 7837 14231 7871
rect 15577 7837 15611 7871
rect 16957 7837 16991 7871
rect 17969 7837 18003 7871
rect 19441 7837 19475 7871
rect 21741 7837 21775 7871
rect 22753 7837 22787 7871
rect 24869 7837 24903 7871
rect 27905 7837 27939 7871
rect 29561 7837 29595 7871
rect 30573 7837 30607 7871
rect 33149 7837 33183 7871
rect 35541 7837 35575 7871
rect 46305 7837 46339 7871
rect 47317 7837 47351 7871
rect 49985 7837 50019 7871
rect 51733 7837 51767 7871
rect 52745 7837 52779 7871
rect 61209 7837 61243 7871
rect 62957 7837 62991 7871
rect 64521 7837 64555 7871
rect 65809 7837 65843 7871
rect 67925 7837 67959 7871
rect 69121 7837 69155 7871
rect 70133 7837 70167 7871
rect 71789 7837 71823 7871
rect 73537 7837 73571 7871
rect 75377 7837 75411 7871
rect 77033 7837 77067 7871
rect 78413 7837 78447 7871
rect 80621 7837 80655 7871
rect 85313 7837 85347 7871
rect 88625 7837 88659 7871
rect 91017 7837 91051 7871
rect 92581 7837 92615 7871
rect 98377 7837 98411 7871
rect 99481 7837 99515 7871
rect 105461 7837 105495 7871
rect 107761 7837 107795 7871
rect 113649 7837 113683 7871
rect 116317 7837 116351 7871
rect 117697 7837 117731 7871
rect 122021 7837 122055 7871
rect 125701 7837 125735 7871
rect 128553 7837 128587 7871
rect 133153 7837 133187 7871
rect 136557 7837 136591 7871
rect 138765 7837 138799 7871
rect 141157 7837 141191 7871
rect 142629 7837 142663 7871
rect 145849 7837 145883 7871
rect 147321 7837 147355 7871
rect 148241 7837 148275 7871
rect 150081 7837 150115 7871
rect 151093 7837 151127 7871
rect 153117 7837 153151 7871
rect 157073 7837 157107 7871
rect 162317 7837 162351 7871
rect 165813 7837 165847 7871
rect 167745 7837 167779 7871
rect 179521 7837 179555 7871
rect 181177 7837 181211 7871
rect 182557 7837 182591 7871
rect 185685 7837 185719 7871
rect 188169 7837 188203 7871
rect 189273 7837 189307 7871
rect 192861 7837 192895 7871
rect 196081 7837 196115 7871
rect 45201 7769 45235 7803
rect 103897 7769 103931 7803
rect 112729 7769 112763 7803
rect 115121 7769 115155 7803
rect 120181 7769 120215 7803
rect 124597 7769 124631 7803
rect 131865 7769 131899 7803
rect 134625 7769 134659 7803
rect 140237 7769 140271 7803
rect 154589 7769 154623 7803
rect 160109 7769 160143 7803
rect 169217 7769 169251 7803
rect 173909 7769 173943 7803
rect 176209 7769 176243 7803
rect 187157 7769 187191 7803
rect 190561 7769 190595 7803
rect 58633 7701 58667 7735
rect 86601 7701 86635 7735
rect 93961 7701 93995 7735
rect 109049 7701 109083 7735
rect 101965 7497 101999 7531
rect 5825 7429 5859 7463
rect 8769 7429 8803 7463
rect 21925 7429 21959 7463
rect 47409 7429 47443 7463
rect 55413 7429 55447 7463
rect 59737 7429 59771 7463
rect 64613 7429 64647 7463
rect 70225 7429 70259 7463
rect 81357 7429 81391 7463
rect 94605 7429 94639 7463
rect 98469 7429 98503 7463
rect 3341 7361 3375 7395
rect 4353 7361 4387 7395
rect 7297 7361 7331 7395
rect 9965 7361 9999 7395
rect 11253 7361 11287 7395
rect 12449 7361 12483 7395
rect 13461 7361 13495 7395
rect 14841 7361 14875 7395
rect 15853 7361 15887 7395
rect 19073 7361 19107 7395
rect 20453 7361 20487 7395
rect 24869 7361 24903 7395
rect 25881 7361 25915 7395
rect 29469 7361 29503 7395
rect 30481 7361 30515 7395
rect 31861 7361 31895 7395
rect 32873 7361 32907 7395
rect 37841 7361 37875 7395
rect 41889 7361 41923 7395
rect 43913 7361 43947 7395
rect 49249 7361 49283 7395
rect 50261 7361 50295 7395
rect 51733 7361 51767 7395
rect 52745 7361 52779 7395
rect 54125 7361 54159 7395
rect 89729 7361 89763 7395
rect 96997 7361 97031 7395
rect 99757 7361 99791 7395
rect 100953 7361 100987 7395
rect 5917 7293 5951 7327
rect 8861 7293 8895 7327
rect 11069 7293 11103 7327
rect 13553 7293 13587 7327
rect 15945 7293 15979 7327
rect 18061 7293 18095 7327
rect 19165 7293 19199 7327
rect 22017 7293 22051 7327
rect 25973 7293 26007 7327
rect 30573 7293 30607 7327
rect 32965 7293 32999 7327
rect 36829 7293 36863 7327
rect 37933 7293 37967 7327
rect 42901 7293 42935 7327
rect 44465 7293 44499 7327
rect 46121 7293 46155 7327
rect 47225 7293 47259 7327
rect 50353 7293 50387 7327
rect 52837 7293 52871 7327
rect 55597 7293 55631 7327
rect 58357 7293 58391 7327
rect 58449 7293 58483 7327
rect 58817 7293 58851 7327
rect 59921 7293 59955 7327
rect 60197 7293 60231 7327
rect 61393 7293 61427 7327
rect 61577 7293 61611 7327
rect 61945 7293 61979 7327
rect 63141 7293 63175 7327
rect 63325 7293 63359 7327
rect 63509 7293 63543 7327
rect 64797 7293 64831 7327
rect 65073 7293 65107 7327
rect 68845 7293 68879 7327
rect 68937 7293 68971 7327
rect 69121 7293 69155 7327
rect 70317 7293 70351 7327
rect 70685 7293 70719 7327
rect 72801 7293 72835 7327
rect 72893 7293 72927 7327
rect 73261 7293 73295 7327
rect 74733 7293 74767 7327
rect 74917 7293 74951 7327
rect 75285 7293 75319 7327
rect 77861 7293 77895 7327
rect 77953 7293 77987 7327
rect 78321 7293 78355 7327
rect 81541 7293 81575 7327
rect 81817 7293 81851 7327
rect 82829 7293 82863 7327
rect 83197 7293 83231 7327
rect 83565 7293 83599 7327
rect 85589 7293 85623 7327
rect 85773 7293 85807 7327
rect 86141 7293 86175 7327
rect 87153 7293 87187 7327
rect 87337 7293 87371 7327
rect 87705 7293 87739 7327
rect 89637 7293 89671 7327
rect 90005 7293 90039 7327
rect 91293 7293 91327 7327
rect 91385 7293 91419 7327
rect 91753 7293 91787 7327
rect 92765 7293 92799 7327
rect 92949 7293 92983 7327
rect 93317 7293 93351 7327
rect 94789 7293 94823 7327
rect 95157 7293 95191 7327
rect 98561 7293 98595 7327
rect 99389 7293 99423 7327
rect 100125 7293 100159 7327
rect 157533 7497 157567 7531
rect 102885 7429 102919 7463
rect 107945 7429 107979 7463
rect 130117 7429 130151 7463
rect 137385 7429 137419 7463
rect 140513 7429 140547 7463
rect 109693 7361 109727 7395
rect 111165 7361 111199 7395
rect 112085 7361 112119 7395
rect 113741 7361 113775 7395
rect 115213 7361 115247 7395
rect 116593 7361 116627 7395
rect 118065 7361 118099 7395
rect 122113 7361 122147 7395
rect 127725 7361 127759 7395
rect 102793 7293 102827 7327
rect 103529 7293 103563 7327
rect 104357 7293 104391 7327
rect 104725 7293 104759 7327
rect 105093 7293 105127 7327
rect 105921 7293 105955 7327
rect 106289 7293 106323 7327
rect 106657 7293 106691 7327
rect 108129 7293 108163 7327
rect 108589 7293 108623 7327
rect 111257 7293 111291 7327
rect 115305 7293 115339 7327
rect 118157 7293 118191 7327
rect 119537 7293 119571 7327
rect 120641 7293 120675 7327
rect 121745 7293 121779 7327
rect 126253 7293 126287 7327
rect 127817 7293 127851 7327
rect 66085 7225 66119 7259
rect 79793 7225 79827 7259
rect 101965 7225 101999 7259
rect 132785 7361 132819 7395
rect 142261 7361 142295 7395
rect 143457 7361 143491 7395
rect 145941 7361 145975 7395
rect 148977 7361 149011 7395
rect 151737 7361 151771 7395
rect 152933 7361 152967 7395
rect 131313 7293 131347 7327
rect 132877 7293 132911 7327
rect 135913 7293 135947 7327
rect 137017 7293 137051 7327
rect 139041 7293 139075 7327
rect 140605 7293 140639 7327
rect 143365 7293 143399 7327
rect 147689 7293 147723 7327
rect 148885 7293 148919 7327
rect 150265 7293 150299 7327
rect 151369 7293 151403 7327
rect 130117 7225 130151 7259
rect 134717 7225 134751 7259
rect 23673 7157 23707 7191
rect 27261 7157 27295 7191
rect 67097 7157 67131 7191
rect 76113 7157 76147 7191
rect 123585 7157 123619 7191
rect 125241 7157 125275 7191
rect 128645 7157 128679 7191
rect 130301 7157 130335 7191
rect 133705 7157 133739 7191
rect 144653 7157 144687 7191
rect 17693 6953 17727 6987
rect 18705 6953 18739 6987
rect 99481 6953 99515 6987
rect 139777 6953 139811 6987
rect 110429 6885 110463 6919
rect 2973 6817 3007 6851
rect 3065 6817 3099 6851
rect 6285 6817 6319 6851
rect 8677 6817 8711 6851
rect 10609 6817 10643 6851
rect 11713 6817 11747 6851
rect 13001 6817 13035 6851
rect 15301 6817 15335 6851
rect 16589 6817 16623 6851
rect 21281 6817 21315 6851
rect 22385 6817 22419 6851
rect 23673 6817 23707 6851
rect 24961 6817 24995 6851
rect 26525 6817 26559 6851
rect 27721 6817 27755 6851
rect 33333 6817 33367 6851
rect 38117 6817 38151 6851
rect 42257 6817 42291 6851
rect 45569 6817 45603 6851
rect 46397 6817 46431 6851
rect 47593 6817 47627 6851
rect 48973 6817 49007 6851
rect 50077 6817 50111 6851
rect 51825 6817 51859 6851
rect 52929 6817 52963 6851
rect 57253 6817 57287 6851
rect 58817 6817 58851 6851
rect 59093 6817 59127 6851
rect 60473 6817 60507 6851
rect 60749 6817 60783 6851
rect 62497 6817 62531 6851
rect 62957 6817 62991 6851
rect 64061 6817 64095 6851
rect 64337 6817 64371 6851
rect 66177 6817 66211 6851
rect 66545 6817 66579 6851
rect 67557 6817 67591 6851
rect 68109 6817 68143 6851
rect 69121 6817 69155 6851
rect 69673 6817 69707 6851
rect 71421 6817 71455 6851
rect 71973 6817 72007 6851
rect 73261 6817 73295 6851
rect 73537 6817 73571 6851
rect 75561 6817 75595 6851
rect 75929 6817 75963 6851
rect 77585 6817 77619 6851
rect 77861 6817 77895 6851
rect 79885 6817 79919 6851
rect 81173 6817 81207 6851
rect 81633 6817 81667 6851
rect 82645 6817 82679 6851
rect 83381 6817 83415 6851
rect 85405 6817 85439 6851
rect 85681 6817 85715 6851
rect 88257 6817 88291 6851
rect 90373 6817 90407 6851
rect 90833 6817 90867 6851
rect 91937 6817 91971 6851
rect 92397 6817 92431 6851
rect 94789 6817 94823 6851
rect 95157 6817 95191 6851
rect 96445 6817 96479 6851
rect 96905 6817 96939 6851
rect 98009 6817 98043 6851
rect 98469 6817 98503 6851
rect 103989 6817 104023 6851
rect 106381 6817 106415 6851
rect 109233 6817 109267 6851
rect 4721 6749 4755 6783
rect 6193 6749 6227 6783
rect 7113 6749 7147 6783
rect 8585 6749 8619 6783
rect 12081 6749 12115 6783
rect 14013 6749 14047 6783
rect 16773 6749 16807 6783
rect 22293 6749 22327 6783
rect 24685 6749 24719 6783
rect 27537 6749 27571 6783
rect 28917 6749 28951 6783
rect 31033 6749 31067 6783
rect 32137 6749 32171 6783
rect 34529 6749 34563 6783
rect 36645 6749 36679 6783
rect 44005 6749 44039 6783
rect 45477 6749 45511 6783
rect 47409 6749 47443 6783
rect 49985 6749 50019 6783
rect 52837 6749 52871 6783
rect 54585 6749 54619 6783
rect 56149 6749 56183 6783
rect 69489 6749 69523 6783
rect 73353 6749 73387 6783
rect 78873 6749 78907 6783
rect 81265 6749 81299 6783
rect 83013 6749 83047 6783
rect 86693 6749 86727 6783
rect 96537 6749 96571 6783
rect 100769 6749 100803 6783
rect 102425 6749 102459 6783
rect 103897 6749 103931 6783
rect 105277 6749 105311 6783
rect 107669 6749 107703 6783
rect 108865 6749 108899 6783
rect 33425 6681 33459 6715
rect 57437 6681 57471 6715
rect 106749 6681 106783 6715
rect 110429 6681 110463 6715
rect 110521 6817 110555 6851
rect 110981 6817 111015 6851
rect 111257 6817 111291 6851
rect 115121 6817 115155 6851
rect 116317 6817 116351 6851
rect 117881 6817 117915 6851
rect 120181 6817 120215 6851
rect 122021 6817 122055 6851
rect 123585 6817 123619 6851
rect 124597 6817 124631 6851
rect 126161 6817 126195 6851
rect 129289 6817 129323 6851
rect 131497 6817 131531 6851
rect 134165 6817 134199 6851
rect 135729 6817 135763 6851
rect 138765 6817 138799 6851
rect 141341 6817 141375 6851
rect 142445 6817 142479 6851
rect 144377 6817 144411 6851
rect 146861 6817 146895 6851
rect 147965 6817 147999 6851
rect 150725 6817 150759 6851
rect 151737 6817 151771 6851
rect 153025 6817 153059 6851
rect 112453 6749 112487 6783
rect 113557 6749 113591 6783
rect 115029 6749 115063 6783
rect 117789 6749 117823 6783
rect 118709 6749 118743 6783
rect 123493 6749 123527 6783
rect 126069 6749 126103 6783
rect 127909 6749 127943 6783
rect 129381 6749 129415 6783
rect 130301 6749 130335 6783
rect 131773 6749 131807 6783
rect 133153 6749 133187 6783
rect 135637 6749 135671 6783
rect 136557 6749 136591 6783
rect 137569 6749 137603 6783
rect 145389 6749 145423 6783
rect 153117 6749 153151 6783
rect 161765 7361 161799 7395
rect 162041 7361 162075 7395
rect 182005 7361 182039 7395
rect 181729 7293 181763 7327
rect 110521 6681 110555 6715
rect 120181 6681 120215 6715
rect 142813 6681 142847 6715
rect 148333 6681 148367 6715
rect 157165 6681 157199 6715
rect 58633 6613 58667 6647
rect 60289 6613 60323 6647
rect 62313 6613 62347 6647
rect 63877 6613 63911 6647
rect 66085 6613 66119 6647
rect 67649 6613 67683 6647
rect 71513 6613 71547 6647
rect 75377 6613 75411 6647
rect 77401 6613 77435 6647
rect 85221 6613 85255 6647
rect 90189 6613 90223 6647
rect 91753 6613 91787 6647
rect 94605 6613 94639 6647
rect 97825 6613 97859 6647
rect 110797 6613 110831 6647
rect 70225 6409 70259 6443
rect 107669 6409 107703 6443
rect 13737 6341 13771 6375
rect 17049 6341 17083 6375
rect 36737 6341 36771 6375
rect 63693 6341 63727 6375
rect 74917 6341 74951 6375
rect 78229 6341 78263 6375
rect 79885 6341 79919 6375
rect 83013 6341 83047 6375
rect 88809 6341 88843 6375
rect 91201 6341 91235 6375
rect 3341 6273 3375 6307
rect 5825 6273 5859 6307
rect 8217 6273 8251 6307
rect 15577 6273 15611 6307
rect 19073 6273 19107 6307
rect 21833 6273 21867 6307
rect 23673 6273 23707 6307
rect 25053 6273 25087 6307
rect 27813 6273 27847 6307
rect 29653 6273 29687 6307
rect 30665 6273 30699 6307
rect 33057 6273 33091 6307
rect 37841 6273 37875 6307
rect 38853 6273 38887 6307
rect 42625 6273 42659 6307
rect 44833 6273 44867 6307
rect 47317 6273 47351 6307
rect 49525 6273 49559 6307
rect 53021 6273 53055 6307
rect 54033 6273 54067 6307
rect 57345 6273 57379 6307
rect 60197 6273 60231 6307
rect 66177 6273 66211 6307
rect 67189 6273 67223 6307
rect 68937 6273 68971 6307
rect 76757 6273 76791 6307
rect 100033 6273 100067 6307
rect 102609 6273 102643 6307
rect 105277 6273 105311 6307
rect 106289 6273 106323 6307
rect 111073 6341 111107 6375
rect 116317 6341 116351 6375
rect 118801 6341 118835 6375
rect 126161 6341 126195 6375
rect 128645 6341 128679 6375
rect 139961 6341 139995 6375
rect 117789 6273 117823 6307
rect 4353 6205 4387 6239
rect 5917 6205 5951 6239
rect 6837 6205 6871 6239
rect 7941 6205 7975 6239
rect 11345 6205 11379 6239
rect 12449 6205 12483 6239
rect 13553 6205 13587 6239
rect 16681 6205 16715 6239
rect 18061 6205 18095 6239
rect 19441 6205 19475 6239
rect 20821 6205 20855 6239
rect 22017 6205 22051 6239
rect 24869 6205 24903 6239
rect 26801 6205 26835 6239
rect 27905 6205 27939 6239
rect 31217 6205 31251 6239
rect 32045 6205 32079 6239
rect 33609 6205 33643 6239
rect 35449 6205 35483 6239
rect 36553 6205 36587 6239
rect 39405 6205 39439 6239
rect 43637 6205 43671 6239
rect 44741 6205 44775 6239
rect 46121 6205 46155 6239
rect 47225 6205 47259 6239
rect 48513 6205 48547 6239
rect 49709 6205 49743 6239
rect 54125 6205 54159 6239
rect 59185 6205 59219 6239
rect 60289 6205 60323 6239
rect 63877 6205 63911 6239
rect 64337 6205 64371 6239
rect 65165 6205 65199 6239
rect 68845 6205 68879 6239
rect 69121 6205 69155 6239
rect 70409 6205 70443 6239
rect 70685 6205 70719 6239
rect 71789 6205 71823 6239
rect 72065 6205 72099 6239
rect 72249 6205 72283 6239
rect 74733 6205 74767 6239
rect 74825 6205 74859 6239
rect 75377 6205 75411 6239
rect 76665 6205 76699 6239
rect 77125 6205 77159 6239
rect 78413 6205 78447 6239
rect 78873 6205 78907 6239
rect 80069 6205 80103 6239
rect 80345 6205 80379 6239
rect 81449 6205 81483 6239
rect 81725 6205 81759 6239
rect 81909 6205 81943 6239
rect 82921 6205 82955 6239
rect 83473 6205 83507 6239
rect 85405 6205 85439 6239
rect 85773 6205 85807 6239
rect 86141 6205 86175 6239
rect 87153 6205 87187 6239
rect 87521 6205 87555 6239
rect 87889 6205 87923 6239
rect 88993 6205 89027 6239
rect 89269 6205 89303 6239
rect 91385 6205 91419 6239
rect 91661 6205 91695 6239
rect 92949 6205 92983 6239
rect 93317 6205 93351 6239
rect 93685 6205 93719 6239
rect 94973 6205 95007 6239
rect 95157 6205 95191 6239
rect 95525 6205 95559 6239
rect 97089 6205 97123 6239
rect 97273 6205 97307 6239
rect 97641 6205 97675 6239
rect 98653 6205 98687 6239
rect 98837 6205 98871 6239
rect 99205 6205 99239 6239
rect 102517 6205 102551 6239
rect 102977 6205 103011 6239
rect 103897 6205 103931 6239
rect 105369 6205 105403 6239
rect 107669 6205 107703 6239
rect 108037 6205 108071 6239
rect 108221 6205 108255 6239
rect 108405 6205 108439 6239
rect 109601 6205 109635 6239
rect 109785 6205 109819 6239
rect 109969 6205 110003 6239
rect 111257 6205 111291 6239
rect 111717 6205 111751 6239
rect 113833 6205 113867 6239
rect 114845 6205 114879 6239
rect 116409 6205 116443 6239
rect 61577 6137 61611 6171
rect 101045 6137 101079 6171
rect 9229 6069 9263 6103
rect 10241 6069 10275 6103
rect 51733 6069 51767 6103
rect 55413 6069 55447 6103
rect 74733 6069 74767 6103
rect 119077 6273 119111 6307
rect 120549 6273 120583 6307
rect 121469 6273 121503 6307
rect 122941 6273 122975 6307
rect 127173 6273 127207 6307
rect 131405 6273 131439 6307
rect 132785 6273 132819 6307
rect 136097 6273 136131 6307
rect 137569 6273 137603 6307
rect 142537 6273 142571 6307
rect 145389 6273 145423 6307
rect 147137 6273 147171 6307
rect 150633 6273 150667 6307
rect 151645 6273 151679 6307
rect 153301 6273 153335 6307
rect 120641 6205 120675 6239
rect 122849 6205 122883 6239
rect 124689 6205 124723 6239
rect 125793 6205 125827 6239
rect 128737 6205 128771 6239
rect 132969 6205 133003 6239
rect 137201 6205 137235 6239
rect 138489 6205 138523 6239
rect 139593 6205 139627 6239
rect 141525 6205 141559 6239
rect 143917 6205 143951 6239
rect 145113 6205 145147 6239
rect 134809 6137 134843 6171
rect 118801 6069 118835 6103
rect 130301 6069 130335 6103
rect 133797 6069 133831 6103
rect 1961 5865 1995 5899
rect 8309 5865 8343 5899
rect 27629 5865 27663 5899
rect 32413 5865 32447 5899
rect 36093 5865 36127 5899
rect 44005 5865 44039 5899
rect 47409 5865 47443 5899
rect 85221 5865 85255 5899
rect 100493 5865 100527 5899
rect 101873 5865 101907 5899
rect 105093 5865 105127 5899
rect 126529 5865 126563 5899
rect 141157 5865 141191 5899
rect 142169 5865 142203 5899
rect 143273 5865 143307 5899
rect 145389 5865 145423 5899
rect 7297 5797 7331 5831
rect 6469 5729 6503 5763
rect 9689 5729 9723 5763
rect 10793 5729 10827 5763
rect 13461 5729 13495 5763
rect 15301 5729 15335 5763
rect 16405 5729 16439 5763
rect 19993 5729 20027 5763
rect 22385 5729 22419 5763
rect 25053 5729 25087 5763
rect 28641 5729 28675 5763
rect 29745 5729 29779 5763
rect 34529 5729 34563 5763
rect 39129 5729 39163 5763
rect 46581 5729 46615 5763
rect 48973 5729 49007 5763
rect 50537 5729 50571 5763
rect 51641 5729 51675 5763
rect 54585 5729 54619 5763
rect 55689 5729 55723 5763
rect 59277 5729 59311 5763
rect 61945 5729 61979 5763
rect 63049 5729 63083 5763
rect 63325 5729 63359 5763
rect 68845 5729 68879 5763
rect 72617 5729 72651 5763
rect 73813 5729 73847 5763
rect 74365 5729 74399 5763
rect 75377 5729 75411 5763
rect 76113 5729 76147 5763
rect 79149 5729 79183 5763
rect 81081 5729 81115 5763
rect 82829 5729 82863 5763
rect 83381 5729 83415 5763
rect 89637 5729 89671 5763
rect 91293 5729 91327 5763
rect 92029 5729 92063 5763
rect 95801 5729 95835 5763
rect 98469 5729 98503 5763
rect 103713 5729 103747 5763
rect 104081 5729 104115 5763
rect 107761 5729 107795 5763
rect 108773 5729 108807 5763
rect 109325 5729 109359 5763
rect 112269 5729 112303 5763
rect 114661 5729 114695 5763
rect 119905 5729 119939 5763
rect 123125 5729 123159 5763
rect 124689 5729 124723 5763
rect 126437 5729 126471 5763
rect 128829 5729 128863 5763
rect 131773 5729 131807 5763
rect 133153 5729 133187 5763
rect 134717 5729 134751 5763
rect 135545 5729 135579 5763
rect 137109 5729 137143 5763
rect 140329 5729 140363 5763
rect 144377 5729 144411 5763
rect 153485 5729 153519 5763
rect 2973 5661 3007 5695
rect 4905 5661 4939 5695
rect 6377 5661 6411 5695
rect 10701 5661 10735 5695
rect 12081 5661 12115 5695
rect 13553 5661 13587 5695
rect 16497 5661 16531 5695
rect 18429 5661 18463 5695
rect 19901 5661 19935 5695
rect 21281 5661 21315 5695
rect 22477 5661 22511 5695
rect 23673 5661 23707 5695
rect 26525 5661 26559 5695
rect 29653 5661 29687 5695
rect 31033 5661 31067 5695
rect 33425 5661 33459 5695
rect 37749 5661 37783 5695
rect 38761 5661 38795 5695
rect 40141 5661 40175 5695
rect 41981 5661 42015 5695
rect 45017 5661 45051 5695
rect 51549 5661 51583 5695
rect 52929 5661 52963 5695
rect 55597 5661 55631 5695
rect 57713 5661 57747 5695
rect 60381 5661 60415 5695
rect 61853 5661 61887 5695
rect 64337 5661 64371 5695
rect 66453 5661 66487 5695
rect 67465 5661 67499 5695
rect 68753 5661 68787 5695
rect 70225 5661 70259 5695
rect 71421 5661 71455 5695
rect 77585 5661 77619 5695
rect 79977 5661 80011 5695
rect 81449 5661 81483 5695
rect 84209 5661 84243 5695
rect 86785 5661 86819 5695
rect 88257 5661 88291 5695
rect 94237 5661 94271 5695
rect 95709 5661 95743 5695
rect 96905 5661 96939 5695
rect 98377 5661 98411 5695
rect 99481 5661 99515 5695
rect 106197 5661 106231 5695
rect 107669 5661 107703 5695
rect 110705 5661 110739 5695
rect 113097 5661 113131 5695
rect 114569 5661 114603 5695
rect 116317 5661 116351 5695
rect 117329 5661 117363 5695
rect 118341 5661 118375 5695
rect 120825 5661 120859 5695
rect 122113 5661 122147 5695
rect 127633 5661 127667 5695
rect 130669 5661 130703 5695
rect 138765 5661 138799 5695
rect 151921 5661 151955 5695
rect 24961 5593 24995 5627
rect 34713 5593 34747 5627
rect 46489 5593 46523 5627
rect 59185 5593 59219 5627
rect 72893 5593 72927 5627
rect 79057 5593 79091 5627
rect 82737 5593 82771 5627
rect 89729 5593 89763 5627
rect 112177 5593 112211 5627
rect 119813 5593 119847 5627
rect 124597 5593 124631 5627
rect 128921 5593 128955 5627
rect 131957 5593 131991 5627
rect 134625 5593 134659 5627
rect 137017 5593 137051 5627
rect 140237 5593 140271 5627
rect 153209 5593 153243 5627
rect 62865 5525 62899 5559
rect 73905 5525 73939 5559
rect 75469 5525 75503 5559
rect 91385 5525 91419 5559
rect 103529 5525 103563 5559
rect 108681 5525 108715 5559
rect 96445 5321 96479 5355
rect 5825 5253 5859 5287
rect 8125 5253 8159 5287
rect 37657 5253 37691 5287
rect 41981 5253 42015 5287
rect 45109 5253 45143 5287
rect 56149 5253 56183 5287
rect 57989 5253 58023 5287
rect 63049 5253 63083 5287
rect 67005 5253 67039 5287
rect 81449 5253 81483 5287
rect 90005 5253 90039 5287
rect 6837 5185 6871 5219
rect 9229 5185 9263 5219
rect 13645 5185 13679 5219
rect 15853 5185 15887 5219
rect 20269 5185 20303 5219
rect 21649 5185 21683 5219
rect 24685 5185 24719 5219
rect 30389 5185 30423 5219
rect 31769 5185 31803 5219
rect 32781 5185 32815 5219
rect 34897 5185 34931 5219
rect 40509 5185 40543 5219
rect 47133 5185 47167 5219
rect 49249 5185 49283 5219
rect 52285 5185 52319 5219
rect 53297 5185 53331 5219
rect 60473 5185 60507 5219
rect 64521 5185 64555 5219
rect 69305 5185 69339 5219
rect 76113 5185 76147 5219
rect 86877 5185 86911 5219
rect 94789 5185 94823 5219
rect 99573 5253 99607 5287
rect 101137 5253 101171 5287
rect 117421 5253 117455 5287
rect 126161 5253 126195 5287
rect 128737 5253 128771 5287
rect 137385 5253 137419 5287
rect 139777 5253 139811 5287
rect 3341 5117 3375 5151
rect 4353 5117 4387 5151
rect 5917 5117 5951 5151
rect 7941 5117 7975 5151
rect 12449 5117 12483 5151
rect 13829 5117 13863 5151
rect 14841 5117 14875 5151
rect 15945 5117 15979 5151
rect 19257 5117 19291 5151
rect 20729 5117 20763 5151
rect 23673 5117 23707 5151
rect 24777 5117 24811 5151
rect 29377 5117 29411 5151
rect 30481 5117 30515 5151
rect 32965 5117 32999 5151
rect 36185 5117 36219 5151
rect 37749 5117 37783 5151
rect 42073 5117 42107 5151
rect 43637 5117 43671 5151
rect 45201 5117 45235 5151
rect 46121 5117 46155 5151
rect 47225 5117 47259 5151
rect 53573 5117 53607 5151
rect 54861 5117 54895 5151
rect 55965 5117 55999 5151
rect 57989 5117 58023 5151
rect 58449 5117 58483 5151
rect 59461 5117 59495 5151
rect 60657 5117 60691 5151
rect 63233 5117 63267 5151
rect 63509 5117 63543 5151
rect 66913 5117 66947 5151
rect 67557 5117 67591 5151
rect 69029 5117 69063 5151
rect 69673 5117 69707 5151
rect 70501 5117 70535 5151
rect 70869 5117 70903 5151
rect 71053 5117 71087 5151
rect 72065 5117 72099 5151
rect 72433 5117 72467 5151
rect 72617 5117 72651 5151
rect 74181 5117 74215 5151
rect 74549 5117 74583 5151
rect 74733 5117 74767 5151
rect 77125 5117 77159 5151
rect 78229 5117 78263 5151
rect 79793 5117 79827 5151
rect 80161 5117 80195 5151
rect 80529 5117 80563 5151
rect 81633 5117 81667 5151
rect 82093 5117 82127 5151
rect 84301 5117 84335 5151
rect 85405 5117 85439 5151
rect 86785 5117 86819 5151
rect 88533 5117 88567 5151
rect 90097 5117 90131 5151
rect 91661 5117 91695 5151
rect 91753 5117 91787 5151
rect 93317 5117 93351 5151
rect 94881 5117 94915 5151
rect 96445 5117 96479 5151
rect 96629 5117 96663 5151
rect 96721 5117 96755 5151
rect 98193 5117 98227 5151
rect 61853 5049 61887 5083
rect 99665 5185 99699 5219
rect 105461 5185 105495 5219
rect 106381 5185 106415 5219
rect 112361 5185 112395 5219
rect 114937 5185 114971 5219
rect 115949 5185 115983 5219
rect 121745 5185 121779 5219
rect 131129 5185 131163 5219
rect 132417 5185 132451 5219
rect 133521 5185 133555 5219
rect 135913 5185 135947 5219
rect 143181 5185 143215 5219
rect 144377 5185 144411 5219
rect 153301 5185 153335 5219
rect 101229 5117 101263 5151
rect 102977 5117 103011 5151
rect 103989 5117 104023 5151
rect 105093 5117 105127 5151
rect 108129 5117 108163 5151
rect 108221 5117 108255 5151
rect 108589 5117 108623 5151
rect 110429 5117 110463 5151
rect 110613 5117 110647 5151
rect 110981 5117 111015 5151
rect 113465 5117 113499 5151
rect 115029 5117 115063 5151
rect 117513 5117 117547 5151
rect 119261 5117 119295 5151
rect 120273 5117 120307 5151
rect 121837 5117 121871 5151
rect 123577 5117 123611 5151
rect 124689 5117 124723 5151
rect 126253 5117 126287 5151
rect 127265 5117 127299 5151
rect 128829 5117 128863 5151
rect 132233 5117 132267 5151
rect 137477 5117 137511 5151
rect 138305 5117 138339 5151
rect 139869 5117 139903 5151
rect 144561 5117 144595 5151
rect 2329 4981 2363 5015
rect 10885 4981 10919 5015
rect 50629 4981 50663 5015
rect 65901 4981 65935 5015
rect 78413 4981 78447 5015
rect 82921 4981 82955 5015
rect 99573 4981 99607 5015
rect 123677 4981 123711 5015
rect 134533 4981 134567 5015
rect 141525 4981 141559 5015
rect 13369 4777 13403 4811
rect 15301 4777 15335 4811
rect 16773 4777 16807 4811
rect 19349 4777 19383 4811
rect 20913 4777 20947 4811
rect 21925 4777 21959 4811
rect 36093 4777 36127 4811
rect 37749 4777 37783 4811
rect 43453 4777 43487 4811
rect 47501 4777 47535 4811
rect 57069 4777 57103 4811
rect 62589 4777 62623 4811
rect 63601 4777 63635 4811
rect 66913 4777 66947 4811
rect 82645 4777 82679 4811
rect 87153 4777 87187 4811
rect 88717 4777 88751 4811
rect 111441 4777 111475 4811
rect 130853 4777 130887 4811
rect 131865 4777 131899 4811
rect 138765 4777 138799 4811
rect 106657 4709 106691 4743
rect 5733 4641 5767 4675
rect 7021 4641 7055 4675
rect 8309 4641 8343 4675
rect 10977 4641 11011 4675
rect 12541 4641 12575 4675
rect 24225 4641 24259 4675
rect 29837 4641 29871 4675
rect 34253 4641 34287 4675
rect 42349 4641 42383 4675
rect 43361 4641 43395 4675
rect 46673 4641 46707 4675
rect 50537 4641 50571 4675
rect 51733 4641 51767 4675
rect 53297 4641 53331 4675
rect 56241 4641 56275 4675
rect 61301 4641 61335 4675
rect 70501 4641 70535 4675
rect 72985 4641 73019 4675
rect 74549 4641 74583 4675
rect 77493 4641 77527 4675
rect 81081 4641 81115 4675
rect 83933 4641 83967 4675
rect 84393 4641 84427 4675
rect 85589 4641 85623 4675
rect 86233 4641 86267 4675
rect 87061 4641 87095 4675
rect 88901 4641 88935 4675
rect 92029 4641 92063 4675
rect 93961 4641 93995 4675
rect 97365 4641 97399 4675
rect 101045 4641 101079 4675
rect 104081 4641 104115 4675
rect 105369 4641 105403 4675
rect 105645 4641 105679 4675
rect 2973 4573 3007 4607
rect 4629 4573 4663 4607
rect 6101 4573 6135 4607
rect 8493 4573 8527 4607
rect 9689 4573 9723 4607
rect 12449 4573 12483 4607
rect 23121 4573 23155 4607
rect 24133 4573 24167 4607
rect 26985 4573 27019 4607
rect 28273 4573 28307 4607
rect 29745 4573 29779 4607
rect 30757 4573 30791 4607
rect 32689 4573 32723 4607
rect 33701 4573 33735 4607
rect 35081 4573 35115 4607
rect 40785 4573 40819 4607
rect 42073 4573 42107 4607
rect 45109 4573 45143 4607
rect 46581 4573 46615 4607
rect 48973 4573 49007 4607
rect 50445 4573 50479 4607
rect 53205 4573 53239 4607
rect 54677 4573 54711 4607
rect 58081 4573 58115 4607
rect 59093 4573 59127 4607
rect 60197 4573 60231 4607
rect 61209 4573 61243 4607
rect 67925 4573 67959 4607
rect 68937 4573 68971 4607
rect 70317 4573 70351 4607
rect 71421 4573 71455 4607
rect 72893 4573 72927 4607
rect 77033 4573 77067 4607
rect 79517 4573 79551 4607
rect 80989 4573 81023 4607
rect 119905 4709 119939 4743
rect 109325 4641 109359 4675
rect 113557 4641 113591 4675
rect 118709 4641 118743 4675
rect 90465 4573 90499 4607
rect 91937 4573 91971 4607
rect 93869 4573 93903 4607
rect 95801 4573 95835 4607
rect 98377 4573 98411 4607
rect 99481 4573 99515 4607
rect 100953 4573 100987 4607
rect 102517 4573 102551 4607
rect 103897 4573 103931 4607
rect 106657 4573 106691 4607
rect 106749 4573 106783 4607
rect 107761 4573 107795 4607
rect 112453 4573 112487 4607
rect 114845 4573 114879 4607
rect 117145 4573 117179 4607
rect 118525 4573 118559 4607
rect 56149 4505 56183 4539
rect 87061 4505 87095 4539
rect 97273 4505 97307 4539
rect 109233 4505 109267 4539
rect 113741 4505 113775 4539
rect 144193 4709 144227 4743
rect 119997 4641 120031 4675
rect 120089 4641 120123 4675
rect 123861 4641 123895 4675
rect 125057 4641 125091 4675
rect 126161 4641 126195 4675
rect 129933 4641 129967 4675
rect 130761 4641 130795 4675
rect 131773 4641 131807 4675
rect 133913 4641 133947 4675
rect 134993 4641 135027 4675
rect 136097 4641 136131 4675
rect 141617 4641 141651 4675
rect 122665 4573 122699 4607
rect 124137 4573 124171 4607
rect 128369 4573 128403 4607
rect 129841 4573 129875 4607
rect 137385 4573 137419 4607
rect 140053 4573 140087 4607
rect 142445 4573 142479 4607
rect 144193 4573 144227 4607
rect 126529 4505 126563 4539
rect 136465 4505 136499 4539
rect 141525 4505 141559 4539
rect 74733 4437 74767 4471
rect 85589 4437 85623 4471
rect 105185 4437 105219 4471
rect 119905 4437 119939 4471
rect 133981 4437 134015 4471
rect 123585 4233 123619 4267
rect 125057 4233 125091 4267
rect 136005 4233 136039 4267
rect 27997 4165 28031 4199
rect 32597 4165 32631 4199
rect 43729 4165 43763 4199
rect 53205 4165 53239 4199
rect 121929 4165 121963 4199
rect 124505 4165 124539 4199
rect 128461 4165 128495 4199
rect 131957 4165 131991 4199
rect 5365 4097 5399 4131
rect 8769 4097 8803 4131
rect 9689 4097 9723 4131
rect 10885 4097 10919 4131
rect 12449 4097 12483 4131
rect 21005 4097 21039 4131
rect 22569 4097 22603 4131
rect 25145 4097 25179 4131
rect 26525 4097 26559 4131
rect 29653 4097 29687 4131
rect 31125 4097 31159 4131
rect 33517 4097 33551 4131
rect 40509 4097 40543 4131
rect 42257 4097 42291 4131
rect 46489 4097 46523 4131
rect 47409 4097 47443 4131
rect 48605 4097 48639 4131
rect 59277 4097 59311 4131
rect 60657 4097 60691 4131
rect 71697 4097 71731 4131
rect 72709 4097 72743 4131
rect 75929 4097 75963 4131
rect 79793 4097 79827 4131
rect 80989 4097 81023 4131
rect 82001 4097 82035 4131
rect 85405 4097 85439 4131
rect 91017 4097 91051 4131
rect 94973 4097 95007 4131
rect 99021 4097 99055 4131
rect 102241 4097 102275 4131
rect 105553 4097 105587 4131
rect 107853 4097 107887 4131
rect 109417 4097 109451 4131
rect 111993 4097 112027 4131
rect 116041 4097 116075 4131
rect 117973 4097 118007 4131
rect 127449 4097 127483 4131
rect 132877 4097 132911 4131
rect 134257 4097 134291 4131
rect 139317 4097 139351 4131
rect 140421 4097 140455 4131
rect 141525 4097 141559 4131
rect 3249 4029 3283 4063
rect 4261 4029 4295 4063
rect 5273 4029 5307 4063
rect 7297 4029 7331 4063
rect 8861 4029 8895 4063
rect 11161 4029 11195 4063
rect 19533 4029 19567 4063
rect 21097 4029 21131 4063
rect 23673 4029 23707 4063
rect 24777 4029 24811 4063
rect 28089 4029 28123 4063
rect 32689 4029 32723 4063
rect 43361 4029 43395 4063
rect 46397 4029 46431 4063
rect 50629 4029 50663 4063
rect 51733 4029 51767 4063
rect 52837 4029 52871 4063
rect 54125 4029 54159 4063
rect 55137 4029 55171 4063
rect 55229 4029 55263 4063
rect 56149 4029 56183 4063
rect 58265 4029 58299 4063
rect 60473 4029 60507 4063
rect 63417 4029 63451 4063
rect 67465 4029 67499 4063
rect 68661 4029 68695 4063
rect 70133 4029 70167 4063
rect 70501 4029 70535 4063
rect 70869 4029 70903 4063
rect 74273 4029 74307 4063
rect 76021 4029 76055 4063
rect 78597 4029 78631 4063
rect 78873 4029 78907 4063
rect 83565 4029 83599 4063
rect 87337 4029 87371 4063
rect 87429 4029 87463 4063
rect 88901 4029 88935 4063
rect 88993 4029 89027 4063
rect 92489 4029 92523 4063
rect 96997 4029 97031 4063
rect 99113 4029 99147 4063
rect 100769 4029 100803 4063
rect 103345 4029 103379 4063
rect 104357 4029 104391 4063
rect 105829 4029 105863 4063
rect 106749 4029 106783 4063
rect 107945 4029 107979 4063
rect 110429 4029 110463 4063
rect 113465 4029 113499 4063
rect 114477 4029 114511 4063
rect 114569 4029 114603 4063
rect 116133 4029 116167 4063
rect 116961 4029 116995 4063
rect 119445 4029 119479 4063
rect 120457 4029 120491 4063
rect 121929 4029 121963 4063
rect 123493 4029 123527 4063
rect 124505 4029 124539 4063
rect 124965 4029 124999 4063
rect 125977 4029 126011 4063
rect 127173 4029 127207 4063
rect 128369 4029 128403 4063
rect 130393 4029 130427 4063
rect 130485 4029 130519 4063
rect 132049 4029 132083 4063
rect 134441 4029 134475 4063
rect 135913 4029 135947 4063
rect 136925 4029 136959 4063
rect 138029 4029 138063 4063
rect 139225 4029 139259 4063
rect 4353 3961 4387 3995
rect 13461 3961 13495 3995
rect 56241 3961 56275 3995
rect 58449 3961 58483 3995
rect 61669 3961 61703 3995
rect 68569 3961 68603 3995
rect 74181 3961 74215 3995
rect 92397 3961 92431 3995
rect 93961 3961 93995 3995
rect 96905 3961 96939 3995
rect 100585 3961 100619 3995
rect 142537 3961 142571 3995
rect 3341 3893 3375 3927
rect 44741 3893 44775 3927
rect 54217 3893 54251 3927
rect 63601 3893 63635 3927
rect 83933 3893 83967 3927
rect 113557 3893 113591 3927
rect 114477 3893 114511 3927
rect 117053 3893 117087 3927
rect 130393 3893 130427 3927
rect 7941 3689 7975 3723
rect 9689 3689 9723 3723
rect 18889 3689 18923 3723
rect 19809 3689 19843 3723
rect 22845 3689 22879 3723
rect 23857 3689 23891 3723
rect 24961 3689 24995 3723
rect 28365 3689 28399 3723
rect 37841 3689 37875 3723
rect 43453 3689 43487 3723
rect 50905 3689 50939 3723
rect 53021 3689 53055 3723
rect 55597 3689 55631 3723
rect 57161 3689 57195 3723
rect 59093 3689 59127 3723
rect 60197 3689 60231 3723
rect 68845 3689 68879 3723
rect 69857 3689 69891 3723
rect 73629 3689 73663 3723
rect 77033 3689 77067 3723
rect 83197 3689 83231 3723
rect 95433 3689 95467 3723
rect 101045 3689 101079 3723
rect 103069 3689 103103 3723
rect 113833 3689 113867 3723
rect 115213 3689 115247 3723
rect 117145 3689 117179 3723
rect 119353 3689 119387 3723
rect 122205 3689 122239 3723
rect 128553 3689 128587 3723
rect 133245 3689 133279 3723
rect 140789 3689 140823 3723
rect 142261 3689 142295 3723
rect 148977 3689 149011 3723
rect 4629 3621 4663 3655
rect 27261 3621 27295 3655
rect 41429 3621 41463 3655
rect 52009 3621 52043 3655
rect 106749 3621 106783 3655
rect 111717 3621 111751 3655
rect 121929 3621 121963 3655
rect 4537 3553 4571 3587
rect 5549 3553 5583 3587
rect 6561 3553 6595 3587
rect 7849 3553 7883 3587
rect 11253 3553 11287 3587
rect 12817 3553 12851 3587
rect 18797 3553 18831 3587
rect 24869 3553 24903 3587
rect 27169 3553 27203 3587
rect 32505 3553 32539 3587
rect 34069 3553 34103 3587
rect 37749 3553 37783 3587
rect 41337 3553 41371 3587
rect 43361 3553 43395 3587
rect 44649 3553 44683 3587
rect 46213 3553 46247 3587
rect 51917 3553 51951 3587
rect 52929 3553 52963 3587
rect 55505 3553 55539 3587
rect 61577 3553 61611 3587
rect 66545 3553 66579 3587
rect 72709 3553 72743 3587
rect 75469 3553 75503 3587
rect 79333 3553 79367 3587
rect 80345 3553 80379 3587
rect 84301 3553 84335 3587
rect 85865 3553 85899 3587
rect 89085 3553 89119 3587
rect 91569 3553 91603 3587
rect 93961 3553 93995 3587
rect 96445 3553 96479 3587
rect 97733 3553 97767 3587
rect 99573 3553 99607 3587
rect 102057 3553 102091 3587
rect 105829 3553 105863 3587
rect 107301 3553 107335 3587
rect 108957 3553 108991 3587
rect 110705 3553 110739 3587
rect 112721 3553 112755 3587
rect 113741 3553 113775 3587
rect 117053 3553 117087 3587
rect 118065 3553 118099 3587
rect 119261 3553 119295 3587
rect 120273 3553 120307 3587
rect 6653 3485 6687 3519
rect 12725 3485 12759 3519
rect 33977 3485 34011 3519
rect 45661 3485 45695 3519
rect 61485 3485 61519 3519
rect 66637 3485 66671 3519
rect 75377 3485 75411 3519
rect 78689 3485 78723 3519
rect 80989 3485 81023 3519
rect 88993 3485 89027 3519
rect 91477 3485 91511 3519
rect 99481 3485 99515 3519
rect 105185 3485 105219 3519
rect 108313 3485 108347 3519
rect 110797 3485 110831 3519
rect 112821 3485 112855 3519
rect 138581 3621 138615 3655
rect 139777 3621 139811 3655
rect 122113 3553 122147 3587
rect 123493 3553 123527 3587
rect 125057 3553 125091 3587
rect 125885 3553 125919 3587
rect 125977 3553 126011 3587
rect 126069 3553 126103 3587
rect 128461 3553 128495 3587
rect 129841 3553 129875 3587
rect 131129 3553 131163 3587
rect 133153 3553 133187 3587
rect 134165 3553 134199 3587
rect 135177 3553 135211 3587
rect 136373 3553 136407 3587
rect 137569 3553 137603 3587
rect 124965 3485 124999 3519
rect 136649 3485 136683 3519
rect 142169 3553 142203 3587
rect 144377 3553 144411 3587
rect 148885 3553 148919 3587
rect 138765 3485 138799 3519
rect 131129 3417 131163 3451
rect 138581 3417 138615 3451
rect 5641 3349 5675 3383
rect 72525 3349 72559 3383
rect 84485 3349 84519 3383
rect 86049 3349 86083 3383
rect 94329 3349 94363 3383
rect 98009 3349 98043 3383
rect 118157 3349 118191 3383
rect 120365 3349 120399 3383
rect 121929 3349 121963 3383
rect 134257 3349 134291 3383
rect 137477 3349 137511 3383
rect 137661 3349 137695 3383
rect 144469 3349 144503 3383
rect 144745 3349 144779 3383
rect 156981 3349 157015 3383
rect 4629 3145 4663 3179
rect 7941 3145 7975 3179
rect 8953 3145 8987 3179
rect 11437 3145 11471 3179
rect 12541 3145 12575 3179
rect 13553 3145 13587 3179
rect 14933 3145 14967 3179
rect 19993 3145 20027 3179
rect 21097 3145 21131 3179
rect 27077 3145 27111 3179
rect 29377 3145 29411 3179
rect 32321 3145 32355 3179
rect 33333 3145 33367 3179
rect 41245 3145 41279 3179
rect 42809 3145 42843 3179
rect 43821 3145 43855 3179
rect 46213 3145 46247 3179
rect 48605 3145 48639 3179
rect 50721 3145 50755 3179
rect 53573 3145 53607 3179
rect 54585 3145 54619 3179
rect 57897 3145 57931 3179
rect 104725 3145 104759 3179
rect 106197 3145 106231 3179
rect 111073 3145 111107 3179
rect 116501 3145 116535 3179
rect 117789 3145 117823 3179
rect 128737 3145 128771 3179
rect 128921 3145 128955 3179
rect 131313 3145 131347 3179
rect 134901 3145 134935 3179
rect 138489 3145 138523 3179
rect 121653 3077 121687 3111
rect 127909 3077 127943 3111
rect 133889 3077 133923 3111
rect 145205 3077 145239 3111
rect 151461 3077 151495 3111
rect 4445 3009 4479 3043
rect 24501 3009 24535 3043
rect 44741 3009 44775 3043
rect 52653 3009 52687 3043
rect 62957 3009 62991 3043
rect 74181 3009 74215 3043
rect 78689 3009 78723 3043
rect 81357 3009 81391 3043
rect 87153 3009 87187 3043
rect 89729 3009 89763 3043
rect 93685 3009 93719 3043
rect 112085 3009 112119 3043
rect 113833 3009 113867 3043
rect 120641 3009 120675 3043
rect 123585 3009 123619 3043
rect 126437 3009 126471 3043
rect 137201 3009 137235 3043
rect 4537 2941 4571 2975
rect 5549 2941 5583 2975
rect 6837 2941 6871 2975
rect 7849 2941 7883 2975
rect 8861 2941 8895 2975
rect 11345 2941 11379 2975
rect 12449 2941 12483 2975
rect 13461 2941 13495 2975
rect 14841 2941 14875 2975
rect 19901 2941 19935 2975
rect 21005 2941 21039 2975
rect 24409 2941 24443 2975
rect 25421 2941 25455 2975
rect 26985 2941 27019 2975
rect 29285 2941 29319 2975
rect 32229 2941 32263 2975
rect 33241 2941 33275 2975
rect 41153 2941 41187 2975
rect 42717 2941 42751 2975
rect 43729 2941 43763 2975
rect 46121 2941 46155 2975
rect 48513 2941 48547 2975
rect 50629 2941 50663 2975
rect 52377 2941 52411 2975
rect 53481 2941 53515 2975
rect 54493 2941 54527 2975
rect 57805 2941 57839 2975
rect 60381 2941 60415 2975
rect 63049 2941 63083 2975
rect 64889 2941 64923 2975
rect 67005 2941 67039 2975
rect 69213 2941 69247 2975
rect 70869 2941 70903 2975
rect 72709 2941 72743 2975
rect 76205 2941 76239 2975
rect 77769 2941 77803 2975
rect 80437 2941 80471 2975
rect 83381 2941 83415 2975
rect 85773 2941 85807 2975
rect 88257 2941 88291 2975
rect 91477 2941 91511 2975
rect 93593 2941 93627 2975
rect 94605 2941 94639 2975
rect 98837 2941 98871 2975
rect 100585 2941 100619 2975
rect 100677 2941 100711 2975
rect 103161 2941 103195 2975
rect 104633 2941 104667 2975
rect 106197 2941 106231 2975
rect 108497 2941 108531 2975
rect 109785 2941 109819 2975
rect 110981 2941 111015 2975
rect 111993 2941 112027 2975
rect 113465 2941 113499 2975
rect 115121 2941 115155 2975
rect 116409 2941 116443 2975
rect 117721 2941 117755 2975
rect 119561 2941 119595 2975
rect 120549 2941 120583 2975
rect 121561 2941 121595 2975
rect 123493 2941 123527 2975
rect 125425 2941 125459 2975
rect 125517 2941 125551 2975
rect 127541 2941 127575 2975
rect 128829 2941 128863 2975
rect 131221 2941 131255 2975
rect 132417 2941 132451 2975
rect 133981 2941 134015 2975
rect 134809 2941 134843 2975
rect 135913 2941 135947 2975
rect 136005 2941 136039 2975
rect 137377 2941 137411 2975
rect 137477 2941 137511 2975
rect 138397 2941 138431 2975
rect 145021 2941 145055 2975
rect 145113 2941 145147 2975
rect 151369 2941 151403 2975
rect 157257 3145 157291 3179
rect 6929 2873 6963 2907
rect 25513 2873 25547 2907
rect 60289 2873 60323 2907
rect 64797 2873 64831 2907
rect 66361 2873 66395 2907
rect 68569 2873 68603 2907
rect 70501 2873 70535 2907
rect 72065 2873 72099 2907
rect 75561 2873 75595 2907
rect 77125 2873 77159 2907
rect 80529 2873 80563 2907
rect 83289 2873 83323 2907
rect 85405 2873 85439 2907
rect 88901 2873 88935 2907
rect 91753 2873 91787 2907
rect 95249 2873 95283 2907
rect 98929 2873 98963 2907
rect 102517 2873 102551 2907
rect 107853 2873 107887 2907
rect 109417 2873 109451 2907
rect 113557 2873 113591 2907
rect 156981 2873 157015 2907
rect 157073 3009 157107 3043
rect 157441 2941 157475 2975
rect 157625 2941 157659 2975
rect 157073 2873 157107 2907
rect 157349 2873 157383 2907
rect 161305 2941 161339 2975
rect 162593 2941 162627 2975
rect 162961 2941 162995 2975
rect 164525 2873 164559 2907
rect 4445 2805 4479 2839
rect 5641 2805 5675 2839
rect 96629 2805 96663 2839
rect 115213 2805 115247 2839
rect 119629 2805 119663 2839
rect 139409 2805 139443 2839
rect 140421 2805 140455 2839
rect 141525 2805 141559 2839
rect 156889 2805 156923 2839
rect 157533 2805 157567 2839
rect 161305 2805 161339 2839
rect 164801 2805 164835 2839
rect 6561 2601 6595 2635
rect 7573 2601 7607 2635
rect 8585 2601 8619 2635
rect 11621 2601 11655 2635
rect 13921 2601 13955 2635
rect 15393 2601 15427 2635
rect 17233 2601 17267 2635
rect 21005 2601 21039 2635
rect 22017 2601 22051 2635
rect 23949 2601 23983 2635
rect 25145 2601 25179 2635
rect 26617 2601 26651 2635
rect 33333 2601 33367 2635
rect 35909 2601 35943 2635
rect 42349 2601 42383 2635
rect 44741 2601 44775 2635
rect 45753 2601 45787 2635
rect 46765 2601 46799 2635
rect 47777 2601 47811 2635
rect 50445 2601 50479 2635
rect 51825 2601 51859 2635
rect 52837 2601 52871 2635
rect 54769 2601 54803 2635
rect 55781 2601 55815 2635
rect 75469 2601 75503 2635
rect 83013 2601 83047 2635
rect 88257 2601 88291 2635
rect 92581 2601 92615 2635
rect 103069 2601 103103 2635
rect 114201 2601 114235 2635
rect 117237 2601 117271 2635
rect 118249 2601 118283 2635
rect 122021 2601 122055 2635
rect 123769 2601 123803 2635
rect 125793 2601 125827 2635
rect 128645 2601 128679 2635
rect 131957 2601 131991 2635
rect 138857 2601 138891 2635
rect 139869 2601 139903 2635
rect 144653 2601 144687 2635
rect 164801 2601 164835 2635
rect 169309 2601 169343 2635
rect 171241 2601 171275 2635
rect 175933 2601 175967 2635
rect 192677 2601 192711 2635
rect 193873 2601 193907 2635
rect 194977 2601 195011 2635
rect 195989 2601 196023 2635
rect 197001 2601 197035 2635
rect 37933 2533 37967 2567
rect 43453 2533 43487 2567
rect 95249 2533 95283 2567
rect 96077 2533 96111 2567
rect 97825 2533 97859 2567
rect 115213 2533 115247 2567
rect 124781 2533 124815 2567
rect 189365 2533 189399 2567
rect 5457 2465 5491 2499
rect 6469 2465 6503 2499
rect 7481 2465 7515 2499
rect 8493 2465 8527 2499
rect 11529 2465 11563 2499
rect 13829 2465 13863 2499
rect 15301 2465 15335 2499
rect 17133 2465 17167 2499
rect 20913 2465 20947 2499
rect 21925 2465 21959 2499
rect 23857 2465 23891 2499
rect 25053 2465 25087 2499
rect 26525 2465 26559 2499
rect 33241 2465 33275 2499
rect 35817 2465 35851 2499
rect 37841 2465 37875 2499
rect 42257 2465 42291 2499
rect 43361 2465 43395 2499
rect 44649 2465 44683 2499
rect 45661 2465 45695 2499
rect 46673 2465 46707 2499
rect 47685 2465 47719 2499
rect 50353 2465 50387 2499
rect 51733 2465 51767 2499
rect 52745 2465 52779 2499
rect 54677 2465 54711 2499
rect 55689 2465 55723 2499
rect 57805 2465 57839 2499
rect 60657 2465 60691 2499
rect 63417 2465 63451 2499
rect 67097 2465 67131 2499
rect 68661 2465 68695 2499
rect 70317 2465 70351 2499
rect 72709 2465 72743 2499
rect 74457 2465 74491 2499
rect 77309 2465 77343 2499
rect 78781 2465 78815 2499
rect 80713 2465 80747 2499
rect 84117 2465 84151 2499
rect 86233 2465 86267 2499
rect 89545 2465 89579 2499
rect 91109 2465 91143 2499
rect 94881 2465 94915 2499
rect 97273 2465 97307 2499
rect 99573 2465 99607 2499
rect 101689 2465 101723 2499
rect 103253 2465 103287 2499
rect 105185 2465 105219 2499
rect 106565 2465 106599 2499
rect 109601 2465 109635 2499
rect 110797 2465 110831 2499
rect 112269 2465 112303 2499
rect 114109 2465 114143 2499
rect 115121 2465 115155 2499
rect 117145 2465 117179 2499
rect 118157 2465 118191 2499
rect 119169 2465 119203 2499
rect 120181 2465 120215 2499
rect 120273 2465 120307 2499
rect 121929 2465 121963 2499
rect 123677 2465 123711 2499
rect 124597 2465 124631 2499
rect 124689 2465 124723 2499
rect 125609 2465 125643 2499
rect 125701 2465 125735 2499
rect 127541 2465 127575 2499
rect 128553 2465 128587 2499
rect 129565 2465 129599 2499
rect 130853 2465 130887 2499
rect 131865 2465 131899 2499
rect 133153 2465 133187 2499
rect 135913 2465 135947 2499
rect 137661 2465 137695 2499
rect 138789 2465 138823 2499
rect 139777 2465 139811 2499
rect 144561 2465 144595 2499
rect 157073 2465 157107 2499
rect 161205 2465 161239 2499
rect 163145 2465 163179 2499
rect 164709 2465 164743 2499
rect 167653 2465 167687 2499
rect 169217 2465 169251 2499
rect 171149 2465 171183 2499
rect 174001 2465 174035 2499
rect 174829 2465 174863 2499
rect 174921 2465 174955 2499
rect 175841 2465 175875 2499
rect 176945 2465 176979 2499
rect 178785 2465 178819 2499
rect 180349 2465 180383 2499
rect 182741 2465 182775 2499
rect 183661 2465 183695 2499
rect 185225 2465 185259 2499
rect 187617 2465 187651 2499
rect 189273 2465 189307 2499
rect 190561 2465 190595 2499
rect 190653 2465 190687 2499
rect 191573 2465 191607 2499
rect 192585 2465 192619 2499
rect 193781 2465 193815 2499
rect 194885 2465 194919 2499
rect 195897 2465 195931 2499
rect 196909 2465 196943 2499
rect 57161 2397 57195 2431
rect 66453 2397 66487 2431
rect 68017 2397 68051 2431
rect 69765 2397 69799 2431
rect 72065 2397 72099 2431
rect 73905 2397 73939 2431
rect 77125 2397 77159 2431
rect 78689 2397 78723 2431
rect 80253 2397 80287 2431
rect 84025 2397 84059 2431
rect 86877 2397 86911 2431
rect 89453 2397 89487 2431
rect 91753 2397 91787 2431
rect 99481 2397 99515 2431
rect 101781 2397 101815 2431
rect 107209 2397 107243 2431
rect 112361 2397 112395 2431
rect 129657 2397 129691 2431
rect 133245 2397 133279 2431
rect 134533 2397 134567 2431
rect 158085 2397 158119 2431
rect 159097 2397 159131 2431
rect 160109 2397 160143 2431
rect 165721 2397 165755 2431
rect 172437 2397 172471 2431
rect 173909 2397 173943 2431
rect 181172 2397 181206 2431
rect 186053 2397 186087 2431
rect 187433 2397 187467 2431
rect 191665 2397 191699 2431
rect 5549 2329 5583 2363
rect 105277 2329 105311 2363
rect 119261 2329 119295 2363
rect 127633 2329 127667 2363
rect 130945 2329 130979 2363
rect 135821 2329 135855 2363
rect 180257 2329 180291 2363
rect 182649 2329 182683 2363
rect 185133 2329 185167 2363
rect 60841 2261 60875 2295
rect 63233 2261 63267 2295
rect 109233 2261 109267 2295
rect 111165 2261 111199 2295
rect 120365 2261 120399 2295
rect 129473 2261 129507 2295
rect 137753 2261 137787 2295
rect 161305 2261 161339 2295
rect 163237 2261 163271 2295
rect 177037 2261 177071 2295
rect 5365 2057 5399 2091
rect 6929 2057 6963 2091
rect 7941 2057 7975 2091
rect 8953 2057 8987 2091
rect 9965 2057 9999 2091
rect 11437 2057 11471 2091
rect 12817 2057 12851 2091
rect 13829 2057 13863 2091
rect 16313 2057 16347 2091
rect 18153 2057 18187 2091
rect 20545 2057 20579 2091
rect 21649 2057 21683 2091
rect 23765 2057 23799 2091
rect 26709 2057 26743 2091
rect 30297 2057 30331 2091
rect 32321 2057 32355 2091
rect 33333 2057 33367 2091
rect 34989 2057 35023 2091
rect 37841 2057 37875 2091
rect 39405 2057 39439 2091
rect 41153 2057 41187 2091
rect 42349 2057 42383 2091
rect 43453 2057 43487 2091
rect 44465 2057 44499 2091
rect 46305 2057 46339 2091
rect 47317 2057 47351 2091
rect 48329 2057 48363 2091
rect 50721 2057 50755 2091
rect 57437 2057 57471 2091
rect 64981 2057 65015 2091
rect 100217 2057 100251 2091
rect 115213 2057 115247 2091
rect 116225 2057 116259 2091
rect 117421 2057 117455 2091
rect 120273 2057 120307 2091
rect 123585 2057 123619 2091
rect 124781 2057 124815 2091
rect 126713 2057 126747 2091
rect 129105 2057 129139 2091
rect 132877 2057 132911 2091
rect 133889 2057 133923 2091
rect 137477 2057 137511 2091
rect 138489 2057 138523 2091
rect 139501 2057 139535 2091
rect 140513 2057 140547 2091
rect 145021 2057 145055 2091
rect 146125 2057 146159 2091
rect 147229 2057 147263 2091
rect 148241 2057 148275 2091
rect 153209 2057 153243 2091
rect 160845 2057 160879 2091
rect 168573 2057 168607 2091
rect 173909 2057 173943 2091
rect 175289 2057 175323 2091
rect 179521 2057 179555 2091
rect 182005 2057 182039 2091
rect 183753 2057 183787 2091
rect 185409 2057 185443 2091
rect 192953 2057 192987 2091
rect 22661 1989 22695 2023
rect 31309 1989 31343 2023
rect 36369 1989 36403 2023
rect 101229 1989 101263 2023
rect 122573 1989 122607 2023
rect 125885 1989 125919 2023
rect 144009 1989 144043 2023
rect 165721 1989 165755 2023
rect 186513 1989 186547 2023
rect 187985 1989 188019 2023
rect 195805 1989 195839 2023
rect 55689 1921 55723 1955
rect 59553 1921 59587 1955
rect 63693 1921 63727 1955
rect 74181 1921 74215 1955
rect 95525 1921 95559 1955
rect 99205 1921 99239 1955
rect 105369 1921 105403 1955
rect 108589 1921 108623 1955
rect 113557 1921 113591 1955
rect 117237 1921 117271 1955
rect 155877 1921 155911 1955
rect 158729 1921 158763 1955
rect 159741 1921 159775 1955
rect 163789 1921 163823 1955
rect 164709 1921 164743 1955
rect 167469 1921 167503 1955
rect 171425 1921 171459 1955
rect 172897 1921 172931 1955
rect 177221 1921 177255 1955
rect 180993 1921 181027 1955
rect 194701 1921 194735 1955
rect 5273 1853 5307 1887
rect 6837 1853 6871 1887
rect 7849 1853 7883 1887
rect 8861 1853 8895 1887
rect 9873 1853 9907 1887
rect 11345 1853 11379 1887
rect 12725 1853 12759 1887
rect 13737 1853 13771 1887
rect 16221 1853 16255 1887
rect 18061 1853 18095 1887
rect 20453 1853 20487 1887
rect 21557 1853 21591 1887
rect 22569 1853 22603 1887
rect 23673 1853 23707 1887
rect 25605 1853 25639 1887
rect 26625 1853 26659 1887
rect 30205 1853 30239 1887
rect 31217 1853 31251 1887
rect 32237 1853 32271 1887
rect 33241 1853 33275 1887
rect 34897 1853 34931 1887
rect 36277 1853 36311 1887
rect 37749 1853 37783 1887
rect 39313 1853 39347 1887
rect 41061 1853 41095 1887
rect 42257 1853 42291 1887
rect 43361 1853 43395 1887
rect 44373 1853 44407 1887
rect 46213 1853 46247 1887
rect 47225 1853 47259 1887
rect 48237 1853 48271 1887
rect 50629 1853 50663 1887
rect 52377 1853 52411 1887
rect 52469 1853 52503 1887
rect 53757 1853 53791 1887
rect 54033 1853 54067 1887
rect 55137 1853 55171 1887
rect 57345 1853 57379 1887
rect 59277 1853 59311 1887
rect 61025 1853 61059 1887
rect 63417 1853 63451 1887
rect 65165 1853 65199 1887
rect 66269 1853 66303 1887
rect 68937 1853 68971 1887
rect 70593 1853 70627 1887
rect 72433 1853 72467 1887
rect 74273 1853 74307 1887
rect 76665 1853 76699 1887
rect 78229 1853 78263 1887
rect 80161 1853 80195 1887
rect 82001 1853 82035 1887
rect 83565 1853 83599 1887
rect 85865 1853 85899 1887
rect 87797 1853 87831 1887
rect 88809 1853 88843 1887
rect 91385 1853 91419 1887
rect 92857 1853 92891 1887
rect 95433 1853 95467 1887
rect 96721 1853 96755 1887
rect 98561 1853 98595 1887
rect 100125 1853 100159 1887
rect 101137 1853 101171 1887
rect 102793 1853 102827 1887
rect 105277 1853 105311 1887
rect 106841 1853 106875 1887
rect 108497 1853 108531 1887
rect 110337 1853 110371 1887
rect 111993 1853 112027 1887
rect 112085 1853 112119 1887
rect 113465 1853 113499 1887
rect 115121 1853 115155 1887
rect 116133 1853 116167 1887
rect 117329 1853 117363 1887
rect 119077 1853 119111 1887
rect 120181 1853 120215 1887
rect 121193 1853 121227 1887
rect 122481 1853 122515 1887
rect 123493 1853 123527 1887
rect 124689 1853 124723 1887
rect 125701 1853 125735 1887
rect 125793 1853 125827 1887
rect 126805 1853 126839 1887
rect 126897 1853 126931 1887
rect 128001 1853 128035 1887
rect 129013 1853 129047 1887
rect 130301 1853 130335 1887
rect 131313 1853 131347 1887
rect 132785 1853 132819 1887
rect 133797 1853 133831 1887
rect 134809 1853 134843 1887
rect 135913 1853 135947 1887
rect 137385 1853 137419 1887
rect 138397 1853 138431 1887
rect 139409 1853 139443 1887
rect 140421 1853 140455 1887
rect 143917 1853 143951 1887
rect 144929 1853 144963 1887
rect 146033 1853 146067 1887
rect 147137 1853 147171 1887
rect 148149 1853 148183 1887
rect 152473 1853 152507 1887
rect 153117 1853 153151 1887
rect 155785 1853 155819 1887
rect 157257 1853 157291 1887
rect 160753 1853 160787 1887
rect 161765 1853 161799 1887
rect 161857 1853 161891 1887
rect 162777 1853 162811 1887
rect 162869 1853 162903 1887
rect 25697 1785 25731 1819
rect 61117 1785 61151 1819
rect 66085 1785 66119 1819
rect 68569 1785 68603 1819
rect 70501 1785 70535 1819
rect 72065 1785 72099 1819
rect 76757 1785 76791 1819
rect 89453 1785 89487 1819
rect 91753 1785 91787 1819
rect 93317 1785 93351 1819
rect 97365 1785 97399 1819
rect 102977 1785 103011 1819
rect 106933 1785 106967 1819
rect 109785 1785 109819 1819
rect 119169 1785 119203 1819
rect 120089 1785 120123 1819
rect 131405 1785 131439 1819
rect 164617 1853 164651 1887
rect 165629 1853 165663 1887
rect 168481 1853 168515 1887
rect 169585 1853 169619 1887
rect 172989 1853 173023 1887
rect 173817 1853 173851 1887
rect 175197 1853 175231 1887
rect 177129 1853 177163 1887
rect 178417 1853 178451 1887
rect 179429 1853 179463 1887
rect 180901 1853 180935 1887
rect 181913 1853 181947 1887
rect 183661 1853 183695 1887
rect 185317 1853 185351 1887
rect 186421 1853 186455 1887
rect 187893 1853 187927 1887
rect 189549 1853 189583 1887
rect 190561 1853 190595 1887
rect 190653 1853 190687 1887
rect 192861 1853 192895 1887
rect 193873 1853 193907 1887
rect 195713 1853 195747 1887
rect 178509 1785 178543 1819
rect 78045 1717 78079 1751
rect 80069 1717 80103 1751
rect 81633 1717 81667 1751
rect 83381 1717 83415 1751
rect 85681 1717 85715 1751
rect 87429 1717 87463 1751
rect 121285 1717 121319 1751
rect 125057 1717 125091 1751
rect 128093 1717 128127 1751
rect 130393 1717 130427 1751
rect 134901 1717 134935 1751
rect 136005 1717 136039 1751
rect 152473 1717 152507 1751
rect 157349 1717 157383 1751
rect 163789 1717 163823 1751
rect 169677 1717 169711 1751
rect 189641 1717 189675 1751
rect 5365 1513 5399 1547
rect 7021 1513 7055 1547
rect 8033 1513 8067 1547
rect 15853 1513 15887 1547
rect 16865 1513 16899 1547
rect 20177 1513 20211 1547
rect 22477 1513 22511 1547
rect 24225 1513 24259 1547
rect 25237 1513 25271 1547
rect 28549 1513 28583 1547
rect 32965 1513 32999 1547
rect 33977 1513 34011 1547
rect 35541 1513 35575 1547
rect 39129 1513 39163 1547
rect 42993 1513 43027 1547
rect 44465 1513 44499 1547
rect 45477 1513 45511 1547
rect 49801 1513 49835 1547
rect 50813 1513 50847 1547
rect 52653 1513 52687 1547
rect 54125 1513 54159 1547
rect 59553 1513 59587 1547
rect 74089 1513 74123 1547
rect 79977 1513 80011 1547
rect 81817 1513 81851 1547
rect 82829 1513 82863 1547
rect 85589 1513 85623 1547
rect 91201 1513 91235 1547
rect 94053 1513 94087 1547
rect 96997 1513 97031 1547
rect 105737 1513 105771 1547
rect 109693 1513 109727 1547
rect 116409 1513 116443 1547
rect 118249 1513 118283 1547
rect 121469 1513 121503 1547
rect 122849 1513 122883 1547
rect 141249 1513 141283 1547
rect 146769 1513 146803 1547
rect 150357 1513 150391 1547
rect 152473 1513 152507 1547
rect 154221 1513 154255 1547
rect 161029 1513 161063 1547
rect 168389 1513 168423 1547
rect 169861 1513 169895 1547
rect 178233 1513 178267 1547
rect 179245 1513 179279 1547
rect 182373 1513 182407 1547
rect 184673 1513 184707 1547
rect 187341 1513 187375 1547
rect 188353 1513 188387 1547
rect 189549 1513 189583 1547
rect 191297 1513 191331 1547
rect 69673 1445 69707 1479
rect 78965 1445 78999 1479
rect 95341 1445 95375 1479
rect 102149 1445 102183 1479
rect 107485 1445 107519 1479
rect 114293 1445 114327 1479
rect 123953 1445 123987 1479
rect 124965 1445 124999 1479
rect 127541 1445 127575 1479
rect 128553 1445 128587 1479
rect 135361 1445 135395 1479
rect 136373 1445 136407 1479
rect 145113 1445 145147 1479
rect 159833 1445 159867 1479
rect 164525 1445 164559 1479
rect 165537 1445 165571 1479
rect 171333 1445 171367 1479
rect 173449 1445 173483 1479
rect 193137 1445 193171 1479
rect 5273 1377 5307 1411
rect 6929 1377 6963 1411
rect 7941 1377 7975 1411
rect 15761 1377 15795 1411
rect 16765 1377 16799 1411
rect 20085 1377 20119 1411
rect 21373 1377 21407 1411
rect 21465 1377 21499 1411
rect 22385 1377 22419 1411
rect 24133 1377 24167 1411
rect 25145 1377 25179 1411
rect 28457 1377 28491 1411
rect 32873 1377 32907 1411
rect 33885 1377 33919 1411
rect 35449 1377 35483 1411
rect 39037 1377 39071 1411
rect 42901 1377 42935 1411
rect 44373 1377 44407 1411
rect 45385 1377 45419 1411
rect 49709 1377 49743 1411
rect 50721 1377 50755 1411
rect 52561 1377 52595 1411
rect 54033 1377 54067 1411
rect 56885 1377 56919 1411
rect 59737 1377 59771 1411
rect 61117 1377 61151 1411
rect 61485 1377 61519 1411
rect 69765 1377 69799 1411
rect 72617 1377 72651 1411
rect 75469 1377 75503 1411
rect 76113 1377 76147 1411
rect 77125 1377 77159 1411
rect 78873 1377 78907 1411
rect 84485 1377 84519 1411
rect 84669 1377 84703 1411
rect 87429 1377 87463 1411
rect 88533 1377 88567 1411
rect 90189 1377 90223 1411
rect 90373 1377 90407 1411
rect 92489 1377 92523 1411
rect 93133 1377 93167 1411
rect 95433 1377 95467 1411
rect 96905 1377 96939 1411
rect 99113 1377 99147 1411
rect 102057 1377 102091 1411
rect 104633 1377 104667 1411
rect 105645 1377 105679 1411
rect 106841 1377 106875 1411
rect 108497 1377 108531 1411
rect 109601 1377 109635 1411
rect 110613 1377 110647 1411
rect 110705 1377 110739 1411
rect 112453 1377 112487 1411
rect 114201 1377 114235 1411
rect 115305 1377 115339 1411
rect 116317 1377 116351 1411
rect 118157 1377 118191 1411
rect 119169 1377 119203 1411
rect 121377 1377 121411 1411
rect 122757 1377 122791 1411
rect 123861 1377 123895 1411
rect 124873 1377 124907 1411
rect 127449 1377 127483 1411
rect 128461 1377 128495 1411
rect 129565 1377 129599 1411
rect 130577 1377 130611 1411
rect 130669 1377 130703 1411
rect 132417 1377 132451 1411
rect 132509 1377 132543 1411
rect 133429 1377 133463 1411
rect 133521 1377 133555 1411
rect 135269 1377 135303 1411
rect 136281 1377 136315 1411
rect 138949 1377 138983 1411
rect 139041 1377 139075 1411
rect 141157 1377 141191 1411
rect 144009 1377 144043 1411
rect 144101 1377 144135 1411
rect 145021 1377 145055 1411
rect 146677 1377 146711 1411
rect 150265 1377 150299 1411
rect 152381 1377 152415 1411
rect 154129 1377 154163 1411
rect 155225 1377 155259 1411
rect 159005 1377 159039 1411
rect 160937 1377 160971 1411
rect 162685 1377 162719 1411
rect 162777 1377 162811 1411
rect 169769 1377 169803 1411
rect 171241 1377 171275 1411
rect 172345 1377 172379 1411
rect 172437 1377 172471 1411
rect 173357 1377 173391 1411
rect 175197 1377 175231 1411
rect 176209 1377 176243 1411
rect 178141 1377 178175 1411
rect 179153 1377 179187 1411
rect 181269 1377 181303 1411
rect 182281 1377 182315 1411
rect 184581 1377 184615 1411
rect 187249 1377 187283 1411
rect 188261 1377 188295 1411
rect 189457 1377 189491 1411
rect 191213 1377 191247 1411
rect 193321 1377 193355 1411
rect 194057 1377 194091 1411
rect 195161 1377 195195 1411
rect 195989 1377 196023 1411
rect 56241 1309 56275 1343
rect 72525 1309 72559 1343
rect 86785 1309 86819 1343
rect 104725 1309 104759 1343
rect 108589 1309 108623 1343
rect 112545 1309 112579 1343
rect 140973 1309 141007 1343
rect 155325 1309 155359 1343
rect 167377 1309 167411 1343
rect 193137 1309 193171 1343
rect 115397 1241 115431 1275
rect 129657 1241 129691 1275
rect 133337 1241 133371 1275
rect 175289 1241 175323 1275
rect 176301 1241 176335 1275
rect 99205 1173 99239 1207
rect 119261 1173 119295 1207
rect 140973 1173 141007 1207
rect 181361 1173 181395 1207
rect 137569 969 137603 1003
rect 144929 969 144963 1003
rect 145021 969 145055 1003
rect 165997 969 166031 1003
rect 133245 901 133279 935
rect 129841 765 129875 799
rect 135085 697 135119 731
rect 135269 697 135303 731
rect 133245 629 133279 663
rect 129841 561 129875 595
rect 143733 901 143767 935
rect 141893 833 141927 867
rect 140789 561 140823 595
rect 140789 357 140823 391
rect 149805 901 149839 935
rect 145021 765 145055 799
rect 146033 765 146067 799
rect 149805 697 149839 731
rect 161949 901 161983 935
rect 143733 561 143767 595
rect 141893 357 141927 391
rect 161857 425 161891 459
rect 137569 289 137603 323
rect 161857 289 161891 323
rect 182189 901 182223 935
rect 182189 765 182223 799
rect 165997 697 166031 731
rect 161949 289 161983 323
rect 166825 493 166859 527
rect 166825 221 166859 255
<< metal1 >>
rect 94317 10591 94375 10597
rect 94317 10557 94329 10591
rect 94363 10588 94375 10591
rect 147306 10588 147312 10600
rect 94363 10560 147312 10588
rect 94363 10557 94375 10560
rect 94317 10551 94375 10557
rect 147306 10548 147312 10560
rect 147364 10548 147370 10600
rect 124398 10480 124404 10532
rect 124456 10520 124462 10532
rect 133598 10520 133604 10532
rect 124456 10492 133604 10520
rect 124456 10480 124462 10492
rect 133598 10480 133604 10492
rect 133656 10480 133662 10532
rect 82170 10412 82176 10464
rect 82228 10452 82234 10464
rect 132954 10452 132960 10464
rect 82228 10424 132960 10452
rect 82228 10412 82234 10424
rect 132954 10412 132960 10424
rect 133012 10412 133018 10464
rect 119798 10344 119804 10396
rect 119856 10384 119862 10396
rect 128906 10384 128912 10396
rect 119856 10356 128912 10384
rect 119856 10344 119862 10356
rect 128906 10344 128912 10356
rect 128964 10344 128970 10396
rect 97810 10276 97816 10328
rect 97868 10316 97874 10328
rect 145558 10316 145564 10328
rect 97868 10288 145564 10316
rect 97868 10276 97874 10288
rect 145558 10276 145564 10288
rect 145616 10276 145622 10328
rect 119706 10208 119712 10260
rect 119764 10248 119770 10260
rect 128538 10248 128544 10260
rect 119764 10220 128544 10248
rect 119764 10208 119770 10220
rect 128538 10208 128544 10220
rect 128596 10208 128602 10260
rect 130378 10208 130384 10260
rect 130436 10248 130442 10260
rect 140958 10248 140964 10260
rect 130436 10220 140964 10248
rect 130436 10208 130442 10220
rect 140958 10208 140964 10220
rect 141016 10208 141022 10260
rect 145834 10208 145840 10260
rect 145892 10248 145898 10260
rect 169570 10248 169576 10260
rect 145892 10220 169576 10248
rect 145892 10208 145898 10220
rect 169570 10208 169576 10220
rect 169628 10208 169634 10260
rect 75178 10140 75184 10192
rect 75236 10180 75242 10192
rect 142982 10180 142988 10192
rect 75236 10152 142988 10180
rect 75236 10140 75242 10152
rect 142982 10140 142988 10152
rect 143040 10140 143046 10192
rect 143537 10183 143595 10189
rect 143537 10149 143549 10183
rect 143583 10180 143595 10183
rect 153105 10183 153163 10189
rect 153105 10180 153117 10183
rect 143583 10152 153117 10180
rect 143583 10149 143595 10152
rect 143537 10143 143595 10149
rect 153105 10149 153117 10152
rect 153151 10149 153163 10183
rect 153105 10143 153163 10149
rect 153197 10183 153255 10189
rect 153197 10149 153209 10183
rect 153243 10180 153255 10183
rect 157981 10183 158039 10189
rect 157981 10180 157993 10183
rect 153243 10152 157993 10180
rect 153243 10149 153255 10152
rect 153197 10143 153255 10149
rect 157981 10149 157993 10152
rect 158027 10149 158039 10183
rect 157981 10143 158039 10149
rect 159082 10140 159088 10192
rect 159140 10180 159146 10192
rect 169938 10180 169944 10192
rect 159140 10152 169944 10180
rect 159140 10140 159146 10152
rect 169938 10140 169944 10152
rect 169996 10140 170002 10192
rect 171318 10140 171324 10192
rect 171376 10180 171382 10192
rect 185670 10180 185676 10192
rect 171376 10152 185676 10180
rect 171376 10140 171382 10152
rect 185670 10140 185676 10152
rect 185728 10140 185734 10192
rect 95694 10072 95700 10124
rect 95752 10112 95758 10124
rect 121270 10112 121276 10124
rect 95752 10084 121276 10112
rect 95752 10072 95758 10084
rect 121270 10072 121276 10084
rect 121328 10072 121334 10124
rect 128998 10072 129004 10124
rect 129056 10112 129062 10124
rect 144362 10112 144368 10124
rect 129056 10084 144368 10112
rect 129056 10072 129062 10084
rect 144362 10072 144368 10084
rect 144420 10072 144426 10124
rect 149698 10072 149704 10124
rect 149756 10112 149762 10124
rect 195146 10112 195152 10124
rect 149756 10084 195152 10112
rect 149756 10072 149762 10084
rect 195146 10072 195152 10084
rect 195204 10072 195210 10124
rect 97534 10004 97540 10056
rect 97592 10044 97598 10056
rect 105630 10044 105636 10056
rect 97592 10016 105636 10044
rect 97592 10004 97598 10016
rect 105630 10004 105636 10016
rect 105688 10004 105694 10056
rect 106090 10004 106096 10056
rect 106148 10044 106154 10056
rect 121178 10044 121184 10056
rect 106148 10016 121184 10044
rect 106148 10004 106154 10016
rect 121178 10004 121184 10016
rect 121236 10004 121242 10056
rect 125134 10004 125140 10056
rect 125192 10044 125198 10056
rect 136910 10044 136916 10056
rect 125192 10016 136916 10044
rect 125192 10004 125198 10016
rect 136910 10004 136916 10016
rect 136968 10004 136974 10056
rect 141786 10044 141792 10056
rect 137020 10016 141792 10044
rect 104434 9936 104440 9988
rect 104492 9976 104498 9988
rect 131758 9976 131764 9988
rect 104492 9948 131764 9976
rect 104492 9936 104498 9948
rect 131758 9936 131764 9948
rect 131816 9936 131822 9988
rect 135438 9936 135444 9988
rect 135496 9976 135502 9988
rect 137020 9976 137048 10016
rect 141786 10004 141792 10016
rect 141844 10004 141850 10056
rect 151262 10004 151268 10056
rect 151320 10044 151326 10056
rect 181254 10044 181260 10056
rect 151320 10016 181260 10044
rect 151320 10004 151326 10016
rect 181254 10004 181260 10016
rect 181312 10004 181318 10056
rect 182082 10004 182088 10056
rect 182140 10044 182146 10056
rect 187050 10044 187056 10056
rect 182140 10016 187056 10044
rect 182140 10004 182146 10016
rect 187050 10004 187056 10016
rect 187108 10004 187114 10056
rect 135496 9948 137048 9976
rect 135496 9936 135502 9948
rect 140406 9936 140412 9988
rect 140464 9976 140470 9988
rect 143353 9979 143411 9985
rect 143353 9976 143365 9979
rect 140464 9948 143365 9976
rect 140464 9936 140470 9948
rect 143353 9945 143365 9948
rect 143399 9945 143411 9979
rect 143353 9939 143411 9945
rect 143445 9979 143503 9985
rect 143445 9945 143457 9979
rect 143491 9976 143503 9979
rect 143537 9979 143595 9985
rect 143537 9976 143549 9979
rect 143491 9948 143549 9976
rect 143491 9945 143503 9948
rect 143445 9939 143503 9945
rect 143537 9945 143549 9948
rect 143583 9945 143595 9979
rect 143537 9939 143595 9945
rect 153197 9979 153255 9985
rect 153197 9945 153209 9979
rect 153243 9945 153255 9979
rect 153197 9939 153255 9945
rect 77846 9868 77852 9920
rect 77904 9908 77910 9920
rect 86034 9908 86040 9920
rect 77904 9880 86040 9908
rect 77904 9868 77910 9880
rect 86034 9868 86040 9880
rect 86092 9868 86098 9920
rect 94314 9908 94320 9920
rect 94275 9880 94320 9908
rect 94314 9868 94320 9880
rect 94372 9868 94378 9920
rect 96062 9868 96068 9920
rect 96120 9908 96126 9920
rect 99926 9908 99932 9920
rect 96120 9880 99932 9908
rect 96120 9868 96126 9880
rect 99926 9868 99932 9880
rect 99984 9868 99990 9920
rect 107930 9868 107936 9920
rect 107988 9908 107994 9920
rect 140774 9908 140780 9920
rect 107988 9880 140780 9908
rect 107988 9868 107994 9880
rect 140774 9868 140780 9880
rect 140832 9868 140838 9920
rect 153105 9911 153163 9917
rect 153105 9877 153117 9911
rect 153151 9908 153163 9911
rect 153212 9908 153240 9939
rect 156046 9936 156052 9988
rect 156104 9976 156110 9988
rect 159174 9976 159180 9988
rect 156104 9948 159180 9976
rect 156104 9936 156110 9948
rect 159174 9936 159180 9948
rect 159232 9936 159238 9988
rect 165246 9936 165252 9988
rect 165304 9976 165310 9988
rect 177022 9976 177028 9988
rect 165304 9948 177028 9976
rect 165304 9936 165310 9948
rect 177022 9936 177028 9948
rect 177080 9936 177086 9988
rect 181530 9976 181536 9988
rect 179432 9948 181536 9976
rect 153151 9880 153240 9908
rect 157981 9911 158039 9917
rect 153151 9877 153163 9880
rect 153105 9871 153163 9877
rect 157981 9877 157993 9911
rect 158027 9908 158039 9911
rect 166166 9908 166172 9920
rect 158027 9880 166172 9908
rect 158027 9877 158039 9880
rect 157981 9871 158039 9877
rect 166166 9868 166172 9880
rect 166224 9868 166230 9920
rect 166258 9868 166264 9920
rect 166316 9908 166322 9920
rect 179432 9908 179460 9948
rect 181530 9936 181536 9948
rect 181588 9936 181594 9988
rect 182726 9936 182732 9988
rect 182784 9976 182790 9988
rect 198826 9976 198832 9988
rect 182784 9948 198832 9976
rect 182784 9936 182790 9948
rect 198826 9936 198832 9948
rect 198884 9936 198890 9988
rect 166316 9880 179460 9908
rect 166316 9868 166322 9880
rect 179506 9868 179512 9920
rect 179564 9908 179570 9920
rect 183186 9908 183192 9920
rect 179564 9880 183192 9908
rect 179564 9868 179570 9880
rect 183186 9868 183192 9880
rect 183244 9868 183250 9920
rect 191098 9868 191104 9920
rect 191156 9908 191162 9920
rect 197998 9908 198004 9920
rect 191156 9880 198004 9908
rect 191156 9868 191162 9880
rect 197998 9868 198004 9880
rect 198056 9868 198062 9920
rect 1104 9818 198812 9840
rect 1104 9766 4078 9818
rect 4130 9766 44078 9818
rect 44130 9766 84078 9818
rect 84130 9766 124078 9818
rect 124130 9766 164078 9818
rect 164130 9766 198812 9818
rect 1104 9744 198812 9766
rect 1026 9664 1032 9716
rect 1084 9704 1090 9716
rect 3053 9707 3111 9713
rect 3053 9704 3065 9707
rect 1084 9676 3065 9704
rect 1084 9664 1090 9676
rect 3053 9673 3065 9676
rect 3099 9673 3111 9707
rect 3053 9667 3111 9673
rect 85850 9664 85856 9716
rect 85908 9704 85914 9716
rect 134794 9704 134800 9716
rect 85908 9676 134800 9704
rect 85908 9664 85914 9676
rect 134794 9664 134800 9676
rect 134852 9664 134858 9716
rect 136174 9664 136180 9716
rect 136232 9704 136238 9716
rect 139118 9704 139124 9716
rect 136232 9676 139124 9704
rect 136232 9664 136238 9676
rect 139118 9664 139124 9676
rect 139176 9664 139182 9716
rect 152090 9664 152096 9716
rect 152148 9704 152154 9716
rect 152148 9676 181484 9704
rect 152148 9664 152154 9676
rect 73154 9636 73160 9648
rect 69860 9608 73160 9636
rect 198 9528 204 9580
rect 256 9568 262 9580
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 256 9540 5457 9568
rect 256 9528 262 9540
rect 5445 9537 5457 9540
rect 5491 9537 5503 9571
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 5445 9531 5503 9537
rect 5644 9540 7941 9568
rect 1486 9460 1492 9512
rect 1544 9500 1550 9512
rect 2961 9503 3019 9509
rect 2961 9500 2973 9503
rect 1544 9472 2973 9500
rect 1544 9460 1550 9472
rect 2961 9469 2973 9472
rect 3007 9469 3019 9503
rect 2961 9463 3019 9469
rect 2976 9432 3004 9463
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 3384 9472 4445 9500
rect 3384 9460 3390 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 5534 9500 5540 9512
rect 5495 9472 5540 9500
rect 4433 9463 4491 9469
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 5644 9432 5672 9540
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 11330 9528 11336 9580
rect 11388 9568 11394 9580
rect 16485 9571 16543 9577
rect 16485 9568 16497 9571
rect 11388 9540 16497 9568
rect 11388 9528 11394 9540
rect 16485 9537 16497 9540
rect 16531 9537 16543 9571
rect 16485 9531 16543 9537
rect 43714 9528 43720 9580
rect 43772 9568 43778 9580
rect 69860 9577 69888 9608
rect 73154 9596 73160 9608
rect 73212 9596 73218 9648
rect 75362 9596 75368 9648
rect 75420 9636 75426 9648
rect 83826 9636 83832 9648
rect 75420 9608 83832 9636
rect 75420 9596 75426 9608
rect 83826 9596 83832 9608
rect 83884 9596 83890 9648
rect 85942 9596 85948 9648
rect 86000 9636 86006 9648
rect 110322 9636 110328 9648
rect 86000 9608 110328 9636
rect 86000 9596 86006 9608
rect 110322 9596 110328 9608
rect 110380 9596 110386 9648
rect 111702 9596 111708 9648
rect 111760 9636 111766 9648
rect 111760 9608 133184 9636
rect 111760 9596 111766 9608
rect 45005 9571 45063 9577
rect 45005 9568 45017 9571
rect 43772 9540 45017 9568
rect 43772 9528 43778 9540
rect 45005 9537 45017 9540
rect 45051 9537 45063 9571
rect 45005 9531 45063 9537
rect 69845 9571 69903 9577
rect 69845 9537 69857 9571
rect 69891 9537 69903 9571
rect 69845 9531 69903 9537
rect 81437 9571 81495 9577
rect 81437 9537 81449 9571
rect 81483 9568 81495 9571
rect 86126 9568 86132 9580
rect 81483 9540 86132 9568
rect 81483 9537 81495 9540
rect 81437 9531 81495 9537
rect 86126 9528 86132 9540
rect 86184 9528 86190 9580
rect 94314 9568 94320 9580
rect 94275 9540 94320 9568
rect 94314 9528 94320 9540
rect 94372 9528 94378 9580
rect 101033 9571 101091 9577
rect 101033 9568 101045 9571
rect 95620 9540 101045 9568
rect 6914 9500 6920 9512
rect 6875 9472 6920 9500
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7156 9472 8033 9500
rect 7156 9460 7162 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15344 9472 15485 9500
rect 15344 9460 15350 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 17034 9500 17040 9512
rect 16995 9472 17040 9500
rect 15473 9463 15531 9469
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 40954 9460 40960 9512
rect 41012 9500 41018 9512
rect 43993 9503 44051 9509
rect 43993 9500 44005 9503
rect 41012 9472 44005 9500
rect 41012 9460 41018 9472
rect 43993 9469 44005 9472
rect 44039 9469 44051 9503
rect 43993 9463 44051 9469
rect 45097 9503 45155 9509
rect 45097 9469 45109 9503
rect 45143 9469 45155 9503
rect 61286 9500 61292 9512
rect 61247 9472 61292 9500
rect 45097 9463 45155 9469
rect 2976 9404 5672 9432
rect 43622 9392 43628 9444
rect 43680 9432 43686 9444
rect 45112 9432 45140 9463
rect 61286 9460 61292 9472
rect 61344 9460 61350 9512
rect 61470 9500 61476 9512
rect 61431 9472 61476 9500
rect 61470 9460 61476 9472
rect 61528 9460 61534 9512
rect 61562 9460 61568 9512
rect 61620 9500 61626 9512
rect 61657 9503 61715 9509
rect 61657 9500 61669 9503
rect 61620 9472 61669 9500
rect 61620 9460 61626 9472
rect 61657 9469 61669 9472
rect 61703 9469 61715 9503
rect 61657 9463 61715 9469
rect 67545 9503 67603 9509
rect 67545 9469 67557 9503
rect 67591 9500 67603 9503
rect 71406 9500 71412 9512
rect 67591 9472 71412 9500
rect 67591 9469 67603 9472
rect 67545 9463 67603 9469
rect 71406 9460 71412 9472
rect 71464 9460 71470 9512
rect 81345 9503 81403 9509
rect 81345 9469 81357 9503
rect 81391 9469 81403 9503
rect 81345 9463 81403 9469
rect 81805 9503 81863 9509
rect 81805 9469 81817 9503
rect 81851 9500 81863 9503
rect 89438 9500 89444 9512
rect 81851 9472 89444 9500
rect 81851 9469 81863 9472
rect 81805 9463 81863 9469
rect 43680 9404 45140 9432
rect 68557 9435 68615 9441
rect 43680 9392 43686 9404
rect 68557 9401 68569 9435
rect 68603 9432 68615 9435
rect 71590 9432 71596 9444
rect 68603 9404 71596 9432
rect 68603 9401 68615 9404
rect 68557 9395 68615 9401
rect 71590 9392 71596 9404
rect 71648 9392 71654 9444
rect 73430 9392 73436 9444
rect 73488 9432 73494 9444
rect 74169 9435 74227 9441
rect 74169 9432 74181 9435
rect 73488 9404 74181 9432
rect 73488 9392 73494 9404
rect 74169 9401 74181 9404
rect 74215 9401 74227 9435
rect 81360 9432 81388 9463
rect 89438 9460 89444 9472
rect 89496 9460 89502 9512
rect 91281 9503 91339 9509
rect 91281 9469 91293 9503
rect 91327 9500 91339 9503
rect 92845 9503 92903 9509
rect 92845 9500 92857 9503
rect 91327 9472 92857 9500
rect 91327 9469 91339 9472
rect 91281 9463 91339 9469
rect 92845 9469 92857 9472
rect 92891 9469 92903 9503
rect 92845 9463 92903 9469
rect 94409 9503 94467 9509
rect 94409 9469 94421 9503
rect 94455 9500 94467 9503
rect 95418 9500 95424 9512
rect 94455 9472 95424 9500
rect 94455 9469 94467 9472
rect 94409 9463 94467 9469
rect 95418 9460 95424 9472
rect 95476 9460 95482 9512
rect 95620 9509 95648 9540
rect 101033 9537 101045 9540
rect 101079 9537 101091 9571
rect 101033 9531 101091 9537
rect 108206 9528 108212 9580
rect 108264 9568 108270 9580
rect 111242 9568 111248 9580
rect 108264 9540 111248 9568
rect 108264 9528 108270 9540
rect 111242 9528 111248 9540
rect 111300 9528 111306 9580
rect 111429 9571 111487 9577
rect 111429 9537 111441 9571
rect 111475 9568 111487 9571
rect 113910 9568 113916 9580
rect 111475 9540 113680 9568
rect 113871 9540 113916 9568
rect 111475 9537 111487 9540
rect 111429 9531 111487 9537
rect 95605 9503 95663 9509
rect 95605 9469 95617 9503
rect 95651 9469 95663 9503
rect 95605 9463 95663 9469
rect 95697 9503 95755 9509
rect 95697 9469 95709 9503
rect 95743 9469 95755 9503
rect 96062 9500 96068 9512
rect 96023 9472 96068 9500
rect 95697 9463 95755 9469
rect 86773 9435 86831 9441
rect 86773 9432 86785 9435
rect 81360 9404 86785 9432
rect 74169 9395 74227 9401
rect 86773 9401 86785 9404
rect 86819 9401 86831 9435
rect 86773 9395 86831 9401
rect 87230 9392 87236 9444
rect 87288 9432 87294 9444
rect 89625 9435 89683 9441
rect 89625 9432 89637 9435
rect 87288 9404 89637 9432
rect 87288 9392 87294 9404
rect 89625 9401 89637 9404
rect 89671 9401 89683 9435
rect 95712 9432 95740 9463
rect 96062 9460 96068 9472
rect 96120 9460 96126 9512
rect 97994 9460 98000 9512
rect 98052 9500 98058 9512
rect 98638 9500 98644 9512
rect 98052 9472 98644 9500
rect 98052 9460 98058 9472
rect 98638 9460 98644 9472
rect 98696 9460 98702 9512
rect 99374 9460 99380 9512
rect 99432 9500 99438 9512
rect 104897 9503 104955 9509
rect 104897 9500 104909 9503
rect 99432 9472 104909 9500
rect 99432 9460 99438 9472
rect 104897 9469 104909 9472
rect 104943 9469 104955 9503
rect 104897 9463 104955 9469
rect 107473 9503 107531 9509
rect 107473 9469 107485 9503
rect 107519 9500 107531 9503
rect 109957 9503 110015 9509
rect 109957 9500 109969 9503
rect 107519 9472 109969 9500
rect 107519 9469 107531 9472
rect 107473 9463 107531 9469
rect 109957 9469 109969 9472
rect 110003 9469 110015 9503
rect 111518 9500 111524 9512
rect 111479 9472 111524 9500
rect 109957 9463 110015 9469
rect 111518 9460 111524 9472
rect 111576 9460 111582 9512
rect 112441 9503 112499 9509
rect 112441 9469 112453 9503
rect 112487 9469 112499 9503
rect 112441 9463 112499 9469
rect 95970 9432 95976 9444
rect 95712 9404 95976 9432
rect 89625 9395 89683 9401
rect 95970 9392 95976 9404
rect 96028 9392 96034 9444
rect 97902 9392 97908 9444
rect 97960 9432 97966 9444
rect 102045 9435 102103 9441
rect 102045 9432 102057 9435
rect 97960 9404 102057 9432
rect 97960 9392 97966 9404
rect 102045 9401 102057 9404
rect 102091 9401 102103 9435
rect 102045 9395 102103 9401
rect 105630 9392 105636 9444
rect 105688 9432 105694 9444
rect 112456 9432 112484 9463
rect 105688 9404 112484 9432
rect 113652 9432 113680 9540
rect 113910 9528 113916 9540
rect 113968 9528 113974 9580
rect 119430 9568 119436 9580
rect 114020 9540 119436 9568
rect 114020 9509 114048 9540
rect 119430 9528 119436 9540
rect 119488 9528 119494 9580
rect 119614 9568 119620 9580
rect 119575 9540 119620 9568
rect 119614 9528 119620 9540
rect 119672 9528 119678 9580
rect 120997 9571 121055 9577
rect 120997 9537 121009 9571
rect 121043 9568 121055 9571
rect 124674 9568 124680 9580
rect 121043 9540 124680 9568
rect 121043 9537 121055 9540
rect 120997 9531 121055 9537
rect 124674 9528 124680 9540
rect 124732 9528 124738 9580
rect 125502 9568 125508 9580
rect 125463 9540 125508 9568
rect 125502 9528 125508 9540
rect 125560 9528 125566 9580
rect 128541 9571 128599 9577
rect 128541 9537 128553 9571
rect 128587 9568 128599 9571
rect 129274 9568 129280 9580
rect 128587 9540 129280 9568
rect 128587 9537 128599 9540
rect 128541 9531 128599 9537
rect 129274 9528 129280 9540
rect 129332 9528 129338 9580
rect 129553 9571 129611 9577
rect 129553 9537 129565 9571
rect 129599 9568 129611 9571
rect 130378 9568 130384 9580
rect 129599 9540 130384 9568
rect 129599 9537 129611 9540
rect 129553 9531 129611 9537
rect 130378 9528 130384 9540
rect 130436 9528 130442 9580
rect 130562 9568 130568 9580
rect 130523 9540 130568 9568
rect 130562 9528 130568 9540
rect 130620 9528 130626 9580
rect 114005 9503 114063 9509
rect 114005 9469 114017 9503
rect 114051 9469 114063 9503
rect 114005 9463 114063 9469
rect 115198 9460 115204 9512
rect 115256 9500 115262 9512
rect 118145 9503 118203 9509
rect 118145 9500 118157 9503
rect 115256 9472 118157 9500
rect 115256 9460 115262 9472
rect 118145 9469 118157 9472
rect 118191 9469 118203 9503
rect 118145 9463 118203 9469
rect 119709 9503 119767 9509
rect 119709 9469 119721 9503
rect 119755 9500 119767 9503
rect 119798 9500 119804 9512
rect 119755 9472 119804 9500
rect 119755 9469 119767 9472
rect 119709 9463 119767 9469
rect 119798 9460 119804 9472
rect 119856 9460 119862 9512
rect 122745 9503 122803 9509
rect 122745 9469 122757 9503
rect 122791 9500 122803 9503
rect 124125 9503 124183 9509
rect 124125 9500 124137 9503
rect 122791 9472 124137 9500
rect 122791 9469 122803 9472
rect 122745 9463 122803 9469
rect 124125 9469 124137 9472
rect 124171 9469 124183 9503
rect 124125 9463 124183 9469
rect 124490 9460 124496 9512
rect 124548 9500 124554 9512
rect 125229 9503 125287 9509
rect 125229 9500 125241 9503
rect 124548 9472 125241 9500
rect 124548 9460 124554 9472
rect 125229 9469 125241 9472
rect 125275 9469 125287 9503
rect 125229 9463 125287 9469
rect 127069 9503 127127 9509
rect 127069 9469 127081 9503
rect 127115 9469 127127 9503
rect 127069 9463 127127 9469
rect 128633 9503 128691 9509
rect 128633 9469 128645 9503
rect 128679 9500 128691 9503
rect 129458 9500 129464 9512
rect 128679 9472 129464 9500
rect 128679 9469 128691 9472
rect 128633 9463 128691 9469
rect 127084 9432 127112 9463
rect 129458 9460 129464 9472
rect 129516 9460 129522 9512
rect 131117 9503 131175 9509
rect 131117 9469 131129 9503
rect 131163 9500 131175 9503
rect 132310 9500 132316 9512
rect 131163 9472 132316 9500
rect 131163 9469 131175 9472
rect 131117 9463 131175 9469
rect 132310 9460 132316 9472
rect 132368 9460 132374 9512
rect 133156 9500 133184 9608
rect 136266 9596 136272 9648
rect 136324 9636 136330 9648
rect 142614 9636 142620 9648
rect 136324 9608 142620 9636
rect 136324 9596 136330 9608
rect 142614 9596 142620 9608
rect 142672 9596 142678 9648
rect 156690 9636 156696 9648
rect 156651 9608 156696 9636
rect 156690 9596 156696 9608
rect 156748 9596 156754 9648
rect 158070 9596 158076 9648
rect 158128 9636 158134 9648
rect 164142 9636 164148 9648
rect 158128 9608 164148 9636
rect 158128 9596 158134 9608
rect 164142 9596 164148 9608
rect 164200 9596 164206 9648
rect 165246 9636 165252 9648
rect 165207 9608 165252 9636
rect 165246 9596 165252 9608
rect 165304 9596 165310 9648
rect 165338 9596 165344 9648
rect 165396 9636 165402 9648
rect 168374 9636 168380 9648
rect 165396 9608 168380 9636
rect 165396 9596 165402 9608
rect 168374 9596 168380 9608
rect 168432 9596 168438 9648
rect 171318 9636 171324 9648
rect 171279 9608 171324 9636
rect 171318 9596 171324 9608
rect 171376 9596 171382 9648
rect 179230 9636 179236 9648
rect 176672 9608 179236 9636
rect 134518 9528 134524 9580
rect 134576 9568 134582 9580
rect 141973 9571 142031 9577
rect 141973 9568 141985 9571
rect 134576 9540 141985 9568
rect 134576 9528 134582 9540
rect 141973 9537 141985 9540
rect 142019 9537 142031 9571
rect 151262 9568 151268 9580
rect 151223 9540 151268 9568
rect 141973 9531 142031 9537
rect 151262 9528 151268 9540
rect 151320 9528 151326 9580
rect 153838 9568 153844 9580
rect 153799 9540 153844 9568
rect 153838 9528 153844 9540
rect 153896 9528 153902 9580
rect 158809 9571 158867 9577
rect 158809 9537 158821 9571
rect 158855 9568 158867 9571
rect 159082 9568 159088 9580
rect 158855 9540 159088 9568
rect 158855 9537 158867 9540
rect 158809 9531 158867 9537
rect 159082 9528 159088 9540
rect 159140 9528 159146 9580
rect 159821 9571 159879 9577
rect 159821 9537 159833 9571
rect 159867 9568 159879 9571
rect 159867 9540 165016 9568
rect 159867 9537 159879 9540
rect 159821 9531 159879 9537
rect 144825 9503 144883 9509
rect 144825 9500 144837 9503
rect 133156 9472 144837 9500
rect 144825 9469 144837 9472
rect 144871 9469 144883 9503
rect 144825 9463 144883 9469
rect 150618 9460 150624 9512
rect 150676 9500 150682 9512
rect 152369 9503 152427 9509
rect 152369 9500 152381 9503
rect 150676 9472 152381 9500
rect 150676 9460 150682 9472
rect 152369 9469 152381 9472
rect 152415 9469 152427 9503
rect 153470 9500 153476 9512
rect 153431 9472 153476 9500
rect 152369 9463 152427 9469
rect 153470 9460 153476 9472
rect 153528 9460 153534 9512
rect 155221 9503 155279 9509
rect 155221 9469 155233 9503
rect 155267 9469 155279 9503
rect 156322 9500 156328 9512
rect 156283 9472 156328 9500
rect 155221 9463 155279 9469
rect 132405 9435 132463 9441
rect 132405 9432 132417 9435
rect 113652 9404 116716 9432
rect 127084 9404 132417 9432
rect 105688 9392 105694 9404
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 12621 9367 12679 9373
rect 12621 9364 12633 9367
rect 11296 9336 12633 9364
rect 11296 9324 11302 9336
rect 12621 9333 12633 9336
rect 12667 9333 12679 9367
rect 12621 9327 12679 9333
rect 27525 9367 27583 9373
rect 27525 9333 27537 9367
rect 27571 9364 27583 9367
rect 27890 9364 27896 9376
rect 27571 9336 27896 9364
rect 27571 9333 27583 9336
rect 27525 9327 27583 9333
rect 27890 9324 27896 9336
rect 27948 9324 27954 9376
rect 40862 9324 40868 9376
rect 40920 9364 40926 9376
rect 42705 9367 42763 9373
rect 42705 9364 42717 9367
rect 40920 9336 42717 9364
rect 40920 9324 40926 9336
rect 42705 9333 42717 9336
rect 42751 9333 42763 9367
rect 42705 9327 42763 9333
rect 46106 9324 46112 9376
rect 46164 9364 46170 9376
rect 46845 9367 46903 9373
rect 46845 9364 46857 9367
rect 46164 9336 46857 9364
rect 46164 9324 46170 9336
rect 46845 9333 46857 9336
rect 46891 9333 46903 9367
rect 46845 9327 46903 9333
rect 46934 9324 46940 9376
rect 46992 9364 46998 9376
rect 47857 9367 47915 9373
rect 47857 9364 47869 9367
rect 46992 9336 47869 9364
rect 46992 9324 46998 9336
rect 47857 9333 47869 9336
rect 47903 9333 47915 9367
rect 47857 9327 47915 9333
rect 59354 9324 59360 9376
rect 59412 9364 59418 9376
rect 59817 9367 59875 9373
rect 59817 9364 59829 9367
rect 59412 9336 59829 9364
rect 59412 9324 59418 9336
rect 59817 9333 59829 9336
rect 59863 9333 59875 9367
rect 62666 9364 62672 9376
rect 62627 9336 62672 9364
rect 59817 9327 59875 9333
rect 62666 9324 62672 9336
rect 62724 9324 62730 9376
rect 64690 9364 64696 9376
rect 64651 9336 64696 9364
rect 64690 9324 64696 9336
rect 64748 9324 64754 9376
rect 65702 9364 65708 9376
rect 65663 9336 65708 9364
rect 65702 9324 65708 9336
rect 65760 9324 65766 9376
rect 70486 9324 70492 9376
rect 70544 9364 70550 9376
rect 70949 9367 71007 9373
rect 70949 9364 70961 9367
rect 70544 9336 70961 9364
rect 70544 9324 70550 9336
rect 70949 9333 70961 9336
rect 70995 9333 71007 9367
rect 70949 9327 71007 9333
rect 73065 9367 73123 9373
rect 73065 9333 73077 9367
rect 73111 9364 73123 9367
rect 73706 9364 73712 9376
rect 73111 9336 73712 9364
rect 73111 9333 73123 9336
rect 73065 9327 73123 9333
rect 73706 9324 73712 9336
rect 73764 9324 73770 9376
rect 73982 9324 73988 9376
rect 74040 9364 74046 9376
rect 75365 9367 75423 9373
rect 75365 9364 75377 9367
rect 74040 9336 75377 9364
rect 74040 9324 74046 9336
rect 75365 9333 75377 9336
rect 75411 9333 75423 9367
rect 76374 9364 76380 9376
rect 76335 9336 76380 9364
rect 75365 9327 75423 9333
rect 76374 9324 76380 9336
rect 76432 9324 76438 9376
rect 78214 9364 78220 9376
rect 78175 9336 78220 9364
rect 78214 9324 78220 9336
rect 78272 9324 78278 9376
rect 79689 9367 79747 9373
rect 79689 9333 79701 9367
rect 79735 9364 79747 9367
rect 80698 9364 80704 9376
rect 79735 9336 80704 9364
rect 79735 9333 79747 9336
rect 79689 9327 79747 9333
rect 80698 9324 80704 9336
rect 80756 9324 80762 9376
rect 82630 9364 82636 9376
rect 82591 9336 82636 9364
rect 82630 9324 82636 9336
rect 82688 9324 82694 9376
rect 82722 9324 82728 9376
rect 82780 9364 82786 9376
rect 83921 9367 83979 9373
rect 83921 9364 83933 9367
rect 82780 9336 83933 9364
rect 82780 9324 82786 9336
rect 83921 9333 83933 9336
rect 83967 9333 83979 9367
rect 83921 9327 83979 9333
rect 84933 9367 84991 9373
rect 84933 9333 84945 9367
rect 84979 9364 84991 9367
rect 85574 9364 85580 9376
rect 84979 9336 85580 9364
rect 84979 9333 84991 9336
rect 84933 9327 84991 9333
rect 85574 9324 85580 9336
rect 85632 9324 85638 9376
rect 85666 9324 85672 9376
rect 85724 9364 85730 9376
rect 87785 9367 87843 9373
rect 87785 9364 87797 9367
rect 85724 9336 87797 9364
rect 85724 9324 85730 9336
rect 87785 9333 87797 9336
rect 87831 9333 87843 9367
rect 96890 9364 96896 9376
rect 96851 9336 96896 9364
rect 87785 9327 87843 9333
rect 96890 9324 96896 9336
rect 96948 9324 96954 9376
rect 96982 9324 96988 9376
rect 97040 9364 97046 9376
rect 98181 9367 98239 9373
rect 98181 9364 98193 9367
rect 97040 9336 98193 9364
rect 97040 9324 97046 9336
rect 98181 9333 98193 9336
rect 98227 9333 98239 9367
rect 99190 9364 99196 9376
rect 99151 9336 99196 9364
rect 98181 9327 98239 9333
rect 99190 9324 99196 9336
rect 99248 9324 99254 9376
rect 99558 9324 99564 9376
rect 99616 9364 99622 9376
rect 103885 9367 103943 9373
rect 103885 9364 103897 9367
rect 99616 9336 103897 9364
rect 99616 9324 99622 9336
rect 103885 9333 103897 9336
rect 103931 9333 103943 9367
rect 103885 9327 103943 9333
rect 108485 9367 108543 9373
rect 108485 9333 108497 9367
rect 108531 9364 108543 9367
rect 110414 9364 110420 9376
rect 108531 9336 110420 9364
rect 108531 9333 108543 9336
rect 108485 9327 108543 9333
rect 110414 9324 110420 9336
rect 110472 9324 110478 9376
rect 114646 9324 114652 9376
rect 114704 9364 114710 9376
rect 115293 9367 115351 9373
rect 115293 9364 115305 9367
rect 114704 9336 115305 9364
rect 114704 9324 114710 9336
rect 115293 9333 115305 9336
rect 115339 9333 115351 9367
rect 115293 9327 115351 9333
rect 116305 9367 116363 9373
rect 116305 9333 116317 9367
rect 116351 9364 116363 9367
rect 116578 9364 116584 9376
rect 116351 9336 116584 9364
rect 116351 9333 116363 9336
rect 116305 9327 116363 9333
rect 116578 9324 116584 9336
rect 116636 9324 116642 9376
rect 116688 9364 116716 9404
rect 132405 9401 132417 9404
rect 132451 9401 132463 9435
rect 136269 9435 136327 9441
rect 136269 9432 136281 9435
rect 132405 9395 132463 9401
rect 132512 9404 136281 9432
rect 128354 9364 128360 9376
rect 116688 9336 128360 9364
rect 128354 9324 128360 9336
rect 128412 9324 128418 9376
rect 128446 9324 128452 9376
rect 128504 9364 128510 9376
rect 132512 9364 132540 9404
rect 136269 9401 136281 9404
rect 136315 9401 136327 9435
rect 136269 9395 136327 9401
rect 136358 9392 136364 9444
rect 136416 9432 136422 9444
rect 140958 9432 140964 9444
rect 136416 9404 140820 9432
rect 140919 9404 140964 9432
rect 136416 9392 136422 9404
rect 133414 9364 133420 9376
rect 128504 9336 132540 9364
rect 133375 9336 133420 9364
rect 128504 9324 128510 9336
rect 133414 9324 133420 9336
rect 133472 9324 133478 9376
rect 133598 9324 133604 9376
rect 133656 9364 133662 9376
rect 135257 9367 135315 9373
rect 135257 9364 135269 9367
rect 133656 9336 135269 9364
rect 133656 9324 133662 9336
rect 135257 9333 135269 9336
rect 135303 9333 135315 9367
rect 135257 9327 135315 9333
rect 135714 9324 135720 9376
rect 135772 9364 135778 9376
rect 138109 9367 138167 9373
rect 138109 9364 138121 9367
rect 135772 9336 138121 9364
rect 135772 9324 135778 9336
rect 138109 9333 138121 9336
rect 138155 9333 138167 9367
rect 139118 9364 139124 9376
rect 139079 9336 139124 9364
rect 138109 9327 138167 9333
rect 139118 9324 139124 9336
rect 139176 9324 139182 9376
rect 140792 9364 140820 9404
rect 140958 9392 140964 9404
rect 141016 9392 141022 9444
rect 146110 9432 146116 9444
rect 141068 9404 146116 9432
rect 141068 9364 141096 9404
rect 146110 9392 146116 9404
rect 146168 9392 146174 9444
rect 151630 9392 151636 9444
rect 151688 9432 151694 9444
rect 155236 9432 155264 9463
rect 156322 9460 156328 9472
rect 156380 9460 156386 9512
rect 160094 9460 160100 9512
rect 160152 9500 160158 9512
rect 163777 9503 163835 9509
rect 163777 9500 163789 9503
rect 160152 9472 163789 9500
rect 160152 9460 160158 9472
rect 163777 9469 163789 9472
rect 163823 9469 163835 9503
rect 164878 9500 164884 9512
rect 164839 9472 164884 9500
rect 163777 9463 163835 9469
rect 164878 9460 164884 9472
rect 164936 9460 164942 9512
rect 164988 9500 165016 9540
rect 165062 9528 165068 9580
rect 165120 9568 165126 9580
rect 166258 9568 166264 9580
rect 165120 9540 166264 9568
rect 165120 9528 165126 9540
rect 166258 9528 166264 9540
rect 166316 9528 166322 9580
rect 168101 9571 168159 9577
rect 168101 9537 168113 9571
rect 168147 9568 168159 9571
rect 172146 9568 172152 9580
rect 168147 9540 172152 9568
rect 168147 9537 168159 9540
rect 168101 9531 168159 9537
rect 172146 9528 172152 9540
rect 172204 9528 172210 9580
rect 173805 9571 173863 9577
rect 173805 9537 173817 9571
rect 173851 9568 173863 9571
rect 173851 9540 176608 9568
rect 173851 9537 173863 9540
rect 173805 9531 173863 9537
rect 166629 9503 166687 9509
rect 166629 9500 166641 9503
rect 164988 9472 166641 9500
rect 166629 9469 166641 9472
rect 166675 9469 166687 9503
rect 167730 9500 167736 9512
rect 167691 9472 167736 9500
rect 166629 9463 166687 9469
rect 167730 9460 167736 9472
rect 167788 9460 167794 9512
rect 169754 9460 169760 9512
rect 169812 9500 169818 9512
rect 169849 9503 169907 9509
rect 169849 9500 169861 9503
rect 169812 9472 169861 9500
rect 169812 9460 169818 9472
rect 169849 9469 169861 9472
rect 169895 9469 169907 9503
rect 171410 9500 171416 9512
rect 171371 9472 171416 9500
rect 169849 9463 169907 9469
rect 171410 9460 171416 9472
rect 171468 9460 171474 9512
rect 172330 9500 172336 9512
rect 172291 9472 172336 9500
rect 172330 9460 172336 9472
rect 172388 9460 172394 9512
rect 173710 9500 173716 9512
rect 173671 9472 173716 9500
rect 173710 9460 173716 9472
rect 173768 9460 173774 9512
rect 175458 9500 175464 9512
rect 175419 9472 175464 9500
rect 175458 9460 175464 9472
rect 175516 9460 175522 9512
rect 176580 9500 176608 9540
rect 176672 9500 176700 9608
rect 179230 9596 179236 9608
rect 179288 9596 179294 9648
rect 176933 9571 176991 9577
rect 176933 9537 176945 9571
rect 176979 9537 176991 9571
rect 181254 9568 181260 9580
rect 181215 9540 181260 9568
rect 176933 9531 176991 9537
rect 176580 9472 176700 9500
rect 151688 9404 155264 9432
rect 151688 9392 151694 9404
rect 155586 9392 155592 9444
rect 155644 9432 155650 9444
rect 157426 9432 157432 9444
rect 155644 9404 157432 9432
rect 155644 9392 155650 9404
rect 157426 9392 157432 9404
rect 157484 9392 157490 9444
rect 162210 9432 162216 9444
rect 157536 9404 162216 9432
rect 140792 9336 141096 9364
rect 142062 9324 142068 9376
rect 142120 9364 142126 9376
rect 143813 9367 143871 9373
rect 143813 9364 143825 9367
rect 142120 9336 143825 9364
rect 142120 9324 142126 9336
rect 143813 9333 143825 9336
rect 143859 9333 143871 9367
rect 143813 9327 143871 9333
rect 144914 9324 144920 9376
rect 144972 9364 144978 9376
rect 146665 9367 146723 9373
rect 146665 9364 146677 9367
rect 144972 9336 146677 9364
rect 144972 9324 144978 9336
rect 146665 9333 146677 9336
rect 146711 9333 146723 9367
rect 146665 9327 146723 9333
rect 147674 9324 147680 9376
rect 147732 9364 147738 9376
rect 147732 9336 147777 9364
rect 147732 9324 147738 9336
rect 148410 9324 148416 9376
rect 148468 9364 148474 9376
rect 149517 9367 149575 9373
rect 149517 9364 149529 9367
rect 148468 9336 149529 9364
rect 148468 9324 148474 9336
rect 149517 9333 149529 9336
rect 149563 9333 149575 9367
rect 149517 9327 149575 9333
rect 155494 9324 155500 9376
rect 155552 9364 155558 9376
rect 156598 9364 156604 9376
rect 155552 9336 156604 9364
rect 155552 9324 155558 9336
rect 156598 9324 156604 9336
rect 156656 9324 156662 9376
rect 157334 9324 157340 9376
rect 157392 9364 157398 9376
rect 157536 9364 157564 9404
rect 162210 9392 162216 9404
rect 162268 9392 162274 9444
rect 162673 9435 162731 9441
rect 162673 9401 162685 9435
rect 162719 9432 162731 9435
rect 175918 9432 175924 9444
rect 162719 9404 175924 9432
rect 162719 9401 162731 9404
rect 162673 9395 162731 9401
rect 175918 9392 175924 9404
rect 175976 9392 175982 9444
rect 176948 9432 176976 9531
rect 181254 9528 181260 9540
rect 181312 9528 181318 9580
rect 181456 9568 181484 9676
rect 181530 9664 181536 9716
rect 181588 9704 181594 9716
rect 183922 9704 183928 9716
rect 181588 9676 183928 9704
rect 181588 9664 181594 9676
rect 183922 9664 183928 9676
rect 183980 9664 183986 9716
rect 187418 9664 187424 9716
rect 187476 9704 187482 9716
rect 191926 9704 191932 9716
rect 187476 9676 191932 9704
rect 187476 9664 187482 9676
rect 191926 9664 191932 9676
rect 191984 9664 191990 9716
rect 181622 9596 181628 9648
rect 181680 9636 181686 9648
rect 182542 9636 182548 9648
rect 181680 9608 182548 9636
rect 181680 9596 181686 9608
rect 182542 9596 182548 9608
rect 182600 9596 182606 9648
rect 182726 9636 182732 9648
rect 182687 9608 182732 9636
rect 182726 9596 182732 9608
rect 182784 9596 182790 9648
rect 185581 9639 185639 9645
rect 185581 9605 185593 9639
rect 185627 9636 185639 9639
rect 191098 9636 191104 9648
rect 185627 9608 191104 9636
rect 185627 9605 185639 9608
rect 185581 9599 185639 9605
rect 191098 9596 191104 9608
rect 191156 9596 191162 9648
rect 194137 9639 194195 9645
rect 194137 9605 194149 9639
rect 194183 9636 194195 9639
rect 196250 9636 196256 9648
rect 194183 9608 196256 9636
rect 194183 9605 194195 9608
rect 194137 9599 194195 9605
rect 196250 9596 196256 9608
rect 196308 9596 196314 9648
rect 196621 9639 196679 9645
rect 196621 9605 196633 9639
rect 196667 9636 196679 9639
rect 199746 9636 199752 9648
rect 196667 9608 199752 9636
rect 196667 9605 196679 9608
rect 196621 9599 196679 9605
rect 199746 9596 199752 9608
rect 199804 9596 199810 9648
rect 186869 9571 186927 9577
rect 186869 9568 186881 9571
rect 181456 9540 186881 9568
rect 186869 9537 186881 9540
rect 186915 9537 186927 9571
rect 186869 9531 186927 9537
rect 188341 9571 188399 9577
rect 188341 9537 188353 9571
rect 188387 9568 188399 9571
rect 190178 9568 190184 9580
rect 188387 9540 190184 9568
rect 188387 9537 188399 9540
rect 188341 9531 188399 9537
rect 190178 9528 190184 9540
rect 190236 9528 190242 9580
rect 190917 9571 190975 9577
rect 190917 9537 190929 9571
rect 190963 9568 190975 9571
rect 194502 9568 194508 9580
rect 190963 9540 194508 9568
rect 190963 9537 190975 9540
rect 190917 9531 190975 9537
rect 194502 9528 194508 9540
rect 194560 9528 194566 9580
rect 195146 9568 195152 9580
rect 195107 9540 195152 9568
rect 195146 9528 195152 9540
rect 195204 9528 195210 9580
rect 177025 9503 177083 9509
rect 177025 9469 177037 9503
rect 177071 9500 177083 9503
rect 177850 9500 177856 9512
rect 177071 9472 177856 9500
rect 177071 9469 177083 9472
rect 177025 9463 177083 9469
rect 177850 9460 177856 9472
rect 177908 9460 177914 9512
rect 178773 9503 178831 9509
rect 178773 9469 178785 9503
rect 178819 9500 178831 9503
rect 182634 9500 182640 9512
rect 178819 9472 182640 9500
rect 178819 9469 178831 9472
rect 178773 9463 178831 9469
rect 182634 9460 182640 9472
rect 182692 9460 182698 9512
rect 182818 9500 182824 9512
rect 182779 9472 182824 9500
rect 182818 9460 182824 9472
rect 182876 9460 182882 9512
rect 183738 9460 183744 9512
rect 183796 9500 183802 9512
rect 184109 9503 184167 9509
rect 184109 9500 184121 9503
rect 183796 9472 184121 9500
rect 183796 9460 183802 9472
rect 184109 9469 184121 9472
rect 184155 9469 184167 9503
rect 184109 9463 184167 9469
rect 185673 9503 185731 9509
rect 185673 9469 185685 9503
rect 185719 9469 185731 9503
rect 185673 9463 185731 9469
rect 188433 9503 188491 9509
rect 188433 9469 188445 9503
rect 188479 9500 188491 9503
rect 188982 9500 188988 9512
rect 188479 9472 188988 9500
rect 188479 9469 188491 9472
rect 188433 9463 188491 9469
rect 184014 9432 184020 9444
rect 176948 9404 184020 9432
rect 184014 9392 184020 9404
rect 184072 9392 184078 9444
rect 185688 9432 185716 9463
rect 188982 9460 188988 9472
rect 189040 9460 189046 9512
rect 189442 9500 189448 9512
rect 189403 9472 189448 9500
rect 189442 9460 189448 9472
rect 189500 9460 189506 9512
rect 191009 9503 191067 9509
rect 191009 9469 191021 9503
rect 191055 9500 191067 9503
rect 192662 9500 192668 9512
rect 191055 9472 192524 9500
rect 192623 9472 192668 9500
rect 191055 9469 191067 9472
rect 191009 9463 191067 9469
rect 191190 9432 191196 9444
rect 185688 9404 191196 9432
rect 191190 9392 191196 9404
rect 191248 9392 191254 9444
rect 192496 9432 192524 9472
rect 192662 9460 192668 9472
rect 192720 9460 192726 9512
rect 194226 9500 194232 9512
rect 194187 9472 194232 9500
rect 194226 9460 194232 9472
rect 194284 9460 194290 9512
rect 196713 9503 196771 9509
rect 196713 9469 196725 9503
rect 196759 9500 196771 9503
rect 197354 9500 197360 9512
rect 196759 9472 197360 9500
rect 196759 9469 196771 9472
rect 196713 9463 196771 9469
rect 197354 9460 197360 9472
rect 197412 9460 197418 9512
rect 195054 9432 195060 9444
rect 192496 9404 195060 9432
rect 195054 9392 195060 9404
rect 195112 9392 195118 9444
rect 157392 9336 157564 9364
rect 161661 9367 161719 9373
rect 157392 9324 157398 9336
rect 161661 9333 161673 9367
rect 161707 9364 161719 9367
rect 164326 9364 164332 9376
rect 161707 9336 164332 9364
rect 161707 9333 161719 9336
rect 161661 9327 161719 9333
rect 164326 9324 164332 9336
rect 164384 9324 164390 9376
rect 169110 9324 169116 9376
rect 169168 9364 169174 9376
rect 174906 9364 174912 9376
rect 169168 9336 174912 9364
rect 169168 9324 169174 9336
rect 174906 9324 174912 9336
rect 174964 9324 174970 9376
rect 179785 9367 179843 9373
rect 179785 9333 179797 9367
rect 179831 9364 179843 9367
rect 191926 9364 191932 9376
rect 179831 9336 191932 9364
rect 179831 9333 179843 9336
rect 179785 9327 179843 9333
rect 191926 9324 191932 9336
rect 191984 9324 191990 9376
rect 1104 9274 198812 9296
rect 1104 9222 24078 9274
rect 24130 9222 64078 9274
rect 64130 9222 104078 9274
rect 104130 9222 144078 9274
rect 144130 9222 184078 9274
rect 184130 9222 198812 9274
rect 1104 9200 198812 9222
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 6914 9160 6920 9172
rect 3007 9132 6920 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7098 9160 7104 9172
rect 7059 9132 7104 9160
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 61286 9120 61292 9172
rect 61344 9160 61350 9172
rect 62761 9163 62819 9169
rect 62761 9160 62773 9163
rect 61344 9132 62773 9160
rect 61344 9120 61350 9132
rect 62761 9129 62773 9132
rect 62807 9129 62819 9163
rect 62761 9123 62819 9129
rect 64690 9120 64696 9172
rect 64748 9160 64754 9172
rect 74442 9160 74448 9172
rect 64748 9132 74448 9160
rect 64748 9120 64754 9132
rect 74442 9120 74448 9132
rect 74500 9120 74506 9172
rect 86773 9163 86831 9169
rect 86773 9160 86785 9163
rect 79520 9132 86785 9160
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 4120 9064 7052 9092
rect 4120 9052 4126 9064
rect 5902 9024 5908 9036
rect 5863 8996 5908 9024
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 7024 9033 7052 9064
rect 27062 9052 27068 9104
rect 27120 9092 27126 9104
rect 27120 9064 29040 9092
rect 27120 9052 27126 9064
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 8993 7067 9027
rect 11238 9024 11244 9036
rect 11199 8996 11244 9024
rect 7009 8987 7067 8993
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 12345 9027 12403 9033
rect 12345 9024 12357 9027
rect 11664 8996 12357 9024
rect 11664 8984 11670 8996
rect 12345 8993 12357 8996
rect 12391 8993 12403 9027
rect 12345 8987 12403 8993
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 15252 8996 17417 9024
rect 15252 8984 15258 8996
rect 17405 8993 17417 8996
rect 17451 8993 17463 9027
rect 27890 9024 27896 9036
rect 27851 8996 27896 9024
rect 17405 8987 17463 8993
rect 27890 8984 27896 8996
rect 27948 8984 27954 9036
rect 29012 9033 29040 9064
rect 41322 9052 41328 9104
rect 41380 9092 41386 9104
rect 41380 9064 43576 9092
rect 41380 9052 41386 9064
rect 28997 9027 29055 9033
rect 28997 8993 29009 9027
rect 29043 8993 29055 9027
rect 28997 8987 29055 8993
rect 38286 8984 38292 9036
rect 38344 9024 38350 9036
rect 38841 9027 38899 9033
rect 38841 9024 38853 9027
rect 38344 8996 38853 9024
rect 38344 8984 38350 8996
rect 38841 8993 38853 8996
rect 38887 8993 38899 9027
rect 40862 9024 40868 9036
rect 40823 8996 40868 9024
rect 38841 8987 38899 8993
rect 40862 8984 40868 8996
rect 40920 8984 40926 9036
rect 42429 9027 42487 9033
rect 42429 8993 42441 9027
rect 42475 9024 42487 9027
rect 43438 9024 43444 9036
rect 42475 8996 43444 9024
rect 42475 8993 42487 8996
rect 42429 8987 42487 8993
rect 43438 8984 43444 8996
rect 43496 8984 43502 9036
rect 43548 9024 43576 9064
rect 43806 9052 43812 9104
rect 43864 9092 43870 9104
rect 77202 9092 77208 9104
rect 43864 9064 47348 9092
rect 43864 9052 43870 9064
rect 47320 9033 47348 9064
rect 72160 9064 77208 9092
rect 44821 9027 44879 9033
rect 44821 9024 44833 9027
rect 43548 8996 44833 9024
rect 44821 8993 44833 8996
rect 44867 8993 44879 9027
rect 47305 9027 47363 9033
rect 44821 8987 44879 8993
rect 46032 8996 47164 9024
rect 4614 8956 4620 8968
rect 4575 8928 4620 8956
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 5810 8956 5816 8968
rect 5771 8928 5816 8956
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 6880 8928 8033 8956
rect 6880 8916 6886 8928
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 8021 8919 8079 8925
rect 9692 8928 12265 8956
rect 4522 8848 4528 8900
rect 4580 8888 4586 8900
rect 9692 8888 9720 8928
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8956 14243 8959
rect 14366 8956 14372 8968
rect 14231 8928 14372 8956
rect 14231 8925 14243 8928
rect 14185 8919 14243 8925
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 16758 8956 16764 8968
rect 16347 8928 16764 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 17328 8888 17356 8919
rect 20438 8916 20444 8968
rect 20496 8956 20502 8968
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 20496 8928 21373 8956
rect 20496 8916 20502 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 26881 8959 26939 8965
rect 26881 8925 26893 8959
rect 26927 8956 26939 8959
rect 29270 8956 29276 8968
rect 26927 8928 29276 8956
rect 26927 8925 26939 8928
rect 26881 8919 26939 8925
rect 29270 8916 29276 8928
rect 29328 8916 29334 8968
rect 29365 8959 29423 8965
rect 29365 8925 29377 8959
rect 29411 8956 29423 8959
rect 31110 8956 31116 8968
rect 29411 8928 31116 8956
rect 29411 8925 29423 8928
rect 29365 8919 29423 8925
rect 31110 8916 31116 8928
rect 31168 8916 31174 8968
rect 32122 8956 32128 8968
rect 32083 8928 32128 8956
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 32214 8916 32220 8968
rect 32272 8956 32278 8968
rect 33137 8959 33195 8965
rect 33137 8956 33149 8959
rect 32272 8928 33149 8956
rect 32272 8916 32278 8928
rect 33137 8925 33149 8928
rect 33183 8925 33195 8959
rect 33137 8919 33195 8925
rect 37737 8959 37795 8965
rect 37737 8925 37749 8959
rect 37783 8956 37795 8959
rect 39114 8956 39120 8968
rect 37783 8928 39120 8956
rect 37783 8925 37795 8928
rect 37737 8919 37795 8925
rect 39114 8916 39120 8928
rect 39172 8916 39178 8968
rect 39209 8959 39267 8965
rect 39209 8925 39221 8959
rect 39255 8956 39267 8959
rect 39390 8956 39396 8968
rect 39255 8928 39396 8956
rect 39255 8925 39267 8928
rect 39209 8919 39267 8925
rect 39390 8916 39396 8928
rect 39448 8916 39454 8968
rect 42337 8959 42395 8965
rect 42337 8925 42349 8959
rect 42383 8956 42395 8959
rect 42702 8956 42708 8968
rect 42383 8928 42708 8956
rect 42383 8925 42395 8928
rect 42337 8919 42395 8925
rect 42702 8916 42708 8928
rect 42760 8916 42766 8968
rect 43714 8956 43720 8968
rect 43675 8928 43720 8956
rect 43714 8916 43720 8928
rect 43772 8916 43778 8968
rect 44174 8916 44180 8968
rect 44232 8956 44238 8968
rect 46032 8956 46060 8996
rect 44232 8928 46060 8956
rect 46109 8959 46167 8965
rect 44232 8916 44238 8928
rect 46109 8925 46121 8959
rect 46155 8956 46167 8959
rect 46934 8956 46940 8968
rect 46155 8928 46940 8956
rect 46155 8925 46167 8928
rect 46109 8919 46167 8925
rect 46934 8916 46940 8928
rect 46992 8916 46998 8968
rect 47136 8965 47164 8996
rect 47305 8993 47317 9027
rect 47351 8993 47363 9027
rect 47305 8987 47363 8993
rect 49050 8984 49056 9036
rect 49108 9024 49114 9036
rect 56229 9027 56287 9033
rect 49108 8996 56180 9024
rect 49108 8984 49114 8996
rect 47121 8959 47179 8965
rect 47121 8925 47133 8959
rect 47167 8925 47179 8959
rect 47121 8919 47179 8925
rect 47578 8916 47584 8968
rect 47636 8956 47642 8968
rect 48961 8959 49019 8965
rect 48961 8956 48973 8959
rect 47636 8928 48973 8956
rect 47636 8916 47642 8928
rect 48961 8925 48973 8928
rect 49007 8925 49019 8959
rect 48961 8919 49019 8925
rect 55125 8959 55183 8965
rect 55125 8925 55137 8959
rect 55171 8956 55183 8959
rect 55858 8956 55864 8968
rect 55171 8928 55864 8956
rect 55171 8925 55183 8928
rect 55125 8919 55183 8925
rect 55858 8916 55864 8928
rect 55916 8916 55922 8968
rect 56152 8965 56180 8996
rect 56229 8993 56241 9027
rect 56275 8993 56287 9027
rect 60458 9024 60464 9036
rect 60419 8996 60464 9024
rect 56229 8987 56287 8993
rect 56137 8959 56195 8965
rect 56137 8925 56149 8959
rect 56183 8925 56195 8959
rect 56137 8919 56195 8925
rect 4580 8860 9720 8888
rect 12268 8860 17356 8888
rect 4580 8848 4586 8860
rect 12268 8832 12296 8860
rect 40218 8848 40224 8900
rect 40276 8888 40282 8900
rect 45005 8891 45063 8897
rect 45005 8888 45017 8891
rect 40276 8860 45017 8888
rect 40276 8848 40282 8860
rect 45005 8857 45017 8860
rect 45051 8857 45063 8891
rect 45005 8851 45063 8857
rect 53098 8848 53104 8900
rect 53156 8888 53162 8900
rect 56244 8888 56272 8987
rect 60458 8984 60464 8996
rect 60516 8984 60522 9036
rect 60921 9027 60979 9033
rect 60921 8993 60933 9027
rect 60967 9024 60979 9027
rect 61194 9024 61200 9036
rect 60967 8996 61200 9024
rect 60967 8993 60979 8996
rect 60921 8987 60979 8993
rect 61194 8984 61200 8996
rect 61252 8984 61258 9036
rect 65702 8984 65708 9036
rect 65760 9024 65766 9036
rect 72160 9033 72188 9064
rect 77202 9052 77208 9064
rect 77260 9052 77266 9104
rect 71409 9027 71467 9033
rect 71409 9024 71421 9027
rect 65760 8996 71421 9024
rect 65760 8984 65766 8996
rect 71409 8993 71421 8996
rect 71455 8993 71467 9027
rect 71409 8987 71467 8993
rect 72145 9027 72203 9033
rect 72145 8993 72157 9027
rect 72191 8993 72203 9027
rect 73706 9024 73712 9036
rect 73667 8996 73712 9024
rect 72145 8987 72203 8993
rect 73706 8984 73712 8996
rect 73764 8984 73770 9036
rect 75270 9024 75276 9036
rect 75231 8996 75276 9024
rect 75270 8984 75276 8996
rect 75328 8984 75334 9036
rect 75454 8984 75460 9036
rect 75512 9024 75518 9036
rect 77021 9027 77079 9033
rect 77021 9024 77033 9027
rect 75512 8996 77033 9024
rect 75512 8984 75518 8996
rect 77021 8993 77033 8996
rect 77067 8993 77079 9027
rect 77021 8987 77079 8993
rect 77757 9027 77815 9033
rect 77757 8993 77769 9027
rect 77803 9024 77815 9027
rect 77846 9024 77852 9036
rect 77803 8996 77852 9024
rect 77803 8993 77815 8996
rect 77757 8987 77815 8993
rect 77846 8984 77852 8996
rect 77904 8984 77910 9036
rect 79520 9033 79548 9132
rect 86773 9129 86785 9132
rect 86819 9129 86831 9163
rect 86773 9123 86831 9129
rect 86954 9120 86960 9172
rect 87012 9160 87018 9172
rect 99282 9160 99288 9172
rect 87012 9132 99288 9160
rect 87012 9120 87018 9132
rect 99282 9120 99288 9132
rect 99340 9120 99346 9172
rect 105630 9160 105636 9172
rect 105591 9132 105636 9160
rect 105630 9120 105636 9132
rect 105688 9120 105694 9172
rect 105722 9120 105728 9172
rect 105780 9160 105786 9172
rect 110782 9160 110788 9172
rect 105780 9132 110788 9160
rect 105780 9120 105786 9132
rect 110782 9120 110788 9132
rect 110840 9120 110846 9172
rect 142062 9160 142068 9172
rect 110984 9132 142068 9160
rect 85482 9052 85488 9104
rect 85540 9092 85546 9104
rect 88245 9095 88303 9101
rect 88245 9092 88257 9095
rect 85540 9064 88257 9092
rect 85540 9052 85546 9064
rect 88245 9061 88257 9064
rect 88291 9061 88303 9095
rect 99190 9092 99196 9104
rect 88245 9055 88303 9061
rect 91756 9064 99196 9092
rect 79505 9027 79563 9033
rect 79505 8993 79517 9027
rect 79551 8993 79563 9027
rect 79505 8987 79563 8993
rect 80241 9027 80299 9033
rect 80241 8993 80253 9027
rect 80287 9024 80299 9027
rect 85942 9024 85948 9036
rect 80287 8996 82952 9024
rect 85903 8996 85948 9024
rect 80287 8993 80299 8996
rect 80241 8987 80299 8993
rect 59081 8959 59139 8965
rect 59081 8925 59093 8959
rect 59127 8956 59139 8959
rect 59538 8956 59544 8968
rect 59127 8928 59544 8956
rect 59127 8925 59139 8928
rect 59081 8919 59139 8925
rect 59538 8916 59544 8928
rect 59596 8916 59602 8968
rect 60550 8956 60556 8968
rect 60511 8928 60556 8956
rect 60550 8916 60556 8928
rect 60608 8916 60614 8968
rect 61102 8916 61108 8968
rect 61160 8956 61166 8968
rect 61749 8959 61807 8965
rect 61749 8956 61761 8959
rect 61160 8928 61761 8956
rect 61160 8916 61166 8928
rect 61749 8925 61761 8928
rect 61795 8925 61807 8959
rect 61749 8919 61807 8925
rect 62574 8916 62580 8968
rect 62632 8956 62638 8968
rect 63773 8959 63831 8965
rect 63773 8956 63785 8959
rect 62632 8928 63785 8956
rect 62632 8916 62638 8928
rect 63773 8925 63785 8928
rect 63819 8925 63831 8959
rect 63773 8919 63831 8925
rect 65981 8959 66039 8965
rect 65981 8925 65993 8959
rect 66027 8925 66039 8959
rect 65981 8919 66039 8925
rect 53156 8860 56272 8888
rect 65996 8888 66024 8919
rect 66070 8916 66076 8968
rect 66128 8956 66134 8968
rect 66993 8959 67051 8965
rect 66993 8956 67005 8959
rect 66128 8928 67005 8956
rect 66128 8916 66134 8928
rect 66993 8925 67005 8928
rect 67039 8925 67051 8959
rect 66993 8919 67051 8925
rect 67818 8916 67824 8968
rect 67876 8956 67882 8968
rect 68005 8959 68063 8965
rect 68005 8956 68017 8959
rect 67876 8928 68017 8956
rect 67876 8916 67882 8928
rect 68005 8925 68017 8928
rect 68051 8925 68063 8959
rect 68005 8919 68063 8925
rect 69293 8959 69351 8965
rect 69293 8925 69305 8959
rect 69339 8956 69351 8959
rect 69934 8956 69940 8968
rect 69339 8928 69940 8956
rect 69339 8925 69351 8928
rect 69293 8919 69351 8925
rect 69934 8916 69940 8928
rect 69992 8916 69998 8968
rect 70302 8956 70308 8968
rect 70263 8928 70308 8956
rect 70302 8916 70308 8928
rect 70360 8916 70366 8968
rect 71777 8959 71835 8965
rect 71777 8925 71789 8959
rect 71823 8956 71835 8959
rect 72234 8956 72240 8968
rect 71823 8928 72240 8956
rect 71823 8925 71835 8928
rect 71777 8919 71835 8925
rect 72234 8916 72240 8928
rect 72292 8916 72298 8968
rect 75178 8956 75184 8968
rect 75139 8928 75184 8956
rect 75178 8916 75184 8928
rect 75236 8916 75242 8968
rect 77386 8956 77392 8968
rect 77347 8928 77392 8956
rect 77386 8916 77392 8928
rect 77444 8916 77450 8968
rect 81069 8959 81127 8965
rect 81069 8956 81081 8959
rect 79704 8928 81081 8956
rect 70946 8888 70952 8900
rect 65996 8860 70952 8888
rect 53156 8848 53162 8860
rect 70946 8848 70952 8860
rect 71004 8848 71010 8900
rect 76834 8848 76840 8900
rect 76892 8888 76898 8900
rect 79704 8888 79732 8928
rect 81069 8925 81081 8928
rect 81115 8925 81127 8959
rect 81069 8919 81127 8925
rect 81526 8916 81532 8968
rect 81584 8956 81590 8968
rect 82633 8959 82691 8965
rect 82633 8956 82645 8959
rect 81584 8928 82645 8956
rect 81584 8916 81590 8928
rect 82633 8925 82645 8928
rect 82679 8925 82691 8959
rect 82633 8919 82691 8925
rect 76892 8860 79732 8888
rect 76892 8848 76898 8860
rect 12250 8780 12256 8832
rect 12308 8780 12314 8832
rect 79597 8823 79655 8829
rect 79597 8789 79609 8823
rect 79643 8820 79655 8823
rect 82814 8820 82820 8832
rect 79643 8792 82820 8820
rect 79643 8789 79655 8792
rect 79597 8783 79655 8789
rect 82814 8780 82820 8792
rect 82872 8780 82878 8832
rect 82924 8820 82952 8996
rect 85942 8984 85948 8996
rect 86000 8984 86006 9036
rect 91756 9033 91784 9064
rect 99190 9052 99196 9064
rect 99248 9052 99254 9104
rect 106918 9052 106924 9104
rect 106976 9092 106982 9104
rect 106976 9064 108252 9092
rect 106976 9052 106982 9064
rect 91741 9027 91799 9033
rect 91741 8993 91753 9027
rect 91787 8993 91799 9027
rect 91741 8987 91799 8993
rect 92201 9027 92259 9033
rect 92201 8993 92213 9027
rect 92247 9024 92259 9027
rect 95142 9024 95148 9036
rect 92247 8996 95148 9024
rect 92247 8993 92259 8996
rect 92201 8987 92259 8993
rect 95142 8984 95148 8996
rect 95200 8984 95206 9036
rect 96893 9027 96951 9033
rect 96893 8993 96905 9027
rect 96939 9024 96951 9027
rect 97074 9024 97080 9036
rect 96939 8996 97080 9024
rect 96939 8993 96951 8996
rect 96893 8987 96951 8993
rect 97074 8984 97080 8996
rect 97132 8984 97138 9036
rect 97902 9024 97908 9036
rect 97863 8996 97908 9024
rect 97902 8984 97908 8996
rect 97960 8984 97966 9036
rect 98457 9027 98515 9033
rect 98457 8993 98469 9027
rect 98503 9024 98515 9027
rect 100846 9024 100852 9036
rect 98503 8996 100852 9024
rect 98503 8993 98515 8996
rect 98457 8987 98515 8993
rect 100846 8984 100852 8996
rect 100904 8984 100910 9036
rect 107930 9024 107936 9036
rect 107891 8996 107936 9024
rect 107930 8984 107936 8996
rect 107988 8984 107994 9036
rect 108224 9033 108252 9064
rect 110984 9033 111012 9132
rect 142062 9120 142068 9132
rect 142120 9120 142126 9172
rect 148318 9160 148324 9172
rect 142264 9132 148324 9160
rect 142264 9092 142292 9132
rect 148318 9120 148324 9132
rect 148376 9120 148382 9172
rect 152090 9160 152096 9172
rect 152051 9132 152096 9160
rect 152090 9120 152096 9132
rect 152148 9120 152154 9172
rect 155770 9120 155776 9172
rect 155828 9160 155834 9172
rect 158806 9160 158812 9172
rect 155828 9132 158812 9160
rect 155828 9120 155834 9132
rect 158806 9120 158812 9132
rect 158864 9120 158870 9172
rect 160094 9160 160100 9172
rect 160055 9132 160100 9160
rect 160094 9120 160100 9132
rect 160152 9120 160158 9172
rect 160278 9120 160284 9172
rect 160336 9160 160342 9172
rect 166626 9160 166632 9172
rect 160336 9132 166632 9160
rect 160336 9120 160342 9132
rect 166626 9120 166632 9132
rect 166684 9120 166690 9172
rect 179506 9160 179512 9172
rect 171428 9132 179512 9160
rect 147674 9092 147680 9104
rect 114388 9064 142292 9092
rect 144380 9064 147680 9092
rect 108209 9027 108267 9033
rect 108209 8993 108221 9027
rect 108255 8993 108267 9027
rect 108209 8987 108267 8993
rect 110969 9027 111027 9033
rect 110969 8993 110981 9027
rect 111015 8993 111027 9027
rect 111242 9024 111248 9036
rect 111203 8996 111248 9024
rect 110969 8987 111027 8993
rect 111242 8984 111248 8996
rect 111300 8984 111306 9036
rect 83550 8916 83556 8968
rect 83608 8956 83614 8968
rect 84381 8959 84439 8965
rect 84381 8956 84393 8959
rect 83608 8928 84393 8956
rect 83608 8916 83614 8928
rect 84381 8925 84393 8928
rect 84427 8925 84439 8959
rect 85850 8956 85856 8968
rect 85811 8928 85856 8956
rect 84381 8919 84439 8925
rect 85850 8916 85856 8928
rect 85908 8916 85914 8968
rect 89254 8956 89260 8968
rect 89215 8928 89260 8956
rect 89254 8916 89260 8928
rect 89312 8916 89318 8968
rect 90358 8956 90364 8968
rect 90319 8928 90364 8956
rect 90358 8916 90364 8928
rect 90416 8916 90422 8968
rect 91830 8956 91836 8968
rect 91791 8928 91836 8956
rect 91830 8916 91836 8928
rect 91888 8916 91894 8968
rect 93857 8959 93915 8965
rect 93857 8925 93869 8959
rect 93903 8956 93915 8959
rect 95329 8959 95387 8965
rect 95329 8956 95341 8959
rect 93903 8928 95341 8956
rect 93903 8925 93915 8928
rect 93857 8919 93915 8925
rect 95329 8925 95341 8928
rect 95375 8925 95387 8959
rect 95329 8919 95387 8925
rect 95418 8916 95424 8968
rect 95476 8956 95482 8968
rect 96801 8959 96859 8965
rect 95476 8928 96752 8956
rect 95476 8916 95482 8928
rect 96724 8888 96752 8928
rect 96801 8925 96813 8959
rect 96847 8956 96859 8959
rect 97810 8956 97816 8968
rect 96847 8928 97816 8956
rect 96847 8925 96859 8928
rect 96801 8919 96859 8925
rect 97810 8916 97816 8928
rect 97868 8916 97874 8968
rect 98086 8956 98092 8968
rect 98047 8928 98092 8956
rect 98086 8916 98092 8928
rect 98144 8916 98150 8968
rect 99098 8916 99104 8968
rect 99156 8956 99162 8968
rect 99469 8959 99527 8965
rect 99469 8956 99481 8959
rect 99156 8928 99481 8956
rect 99156 8916 99162 8928
rect 99469 8925 99481 8928
rect 99515 8925 99527 8959
rect 99469 8919 99527 8925
rect 99926 8916 99932 8968
rect 99984 8956 99990 8968
rect 100481 8959 100539 8965
rect 100481 8956 100493 8959
rect 99984 8928 100493 8956
rect 99984 8916 99990 8928
rect 100481 8925 100493 8928
rect 100527 8925 100539 8959
rect 102042 8956 102048 8968
rect 102003 8928 102048 8956
rect 100481 8919 100539 8925
rect 102042 8916 102048 8928
rect 102100 8916 102106 8968
rect 103054 8956 103060 8968
rect 103015 8928 103060 8956
rect 103054 8916 103060 8928
rect 103112 8916 103118 8968
rect 106645 8959 106703 8965
rect 106645 8925 106657 8959
rect 106691 8956 106703 8959
rect 109218 8956 109224 8968
rect 106691 8928 109224 8956
rect 106691 8925 106703 8928
rect 106645 8919 106703 8925
rect 109218 8916 109224 8928
rect 109276 8916 109282 8968
rect 114388 8965 114416 9064
rect 114465 9027 114523 9033
rect 114465 8993 114477 9027
rect 114511 9024 114523 9027
rect 119706 9024 119712 9036
rect 114511 8996 118280 9024
rect 119667 8996 119712 9024
rect 114511 8993 114523 8996
rect 114465 8987 114523 8993
rect 109589 8959 109647 8965
rect 109589 8925 109601 8959
rect 109635 8956 109647 8959
rect 112993 8959 113051 8965
rect 112993 8956 113005 8959
rect 109635 8928 113005 8956
rect 109635 8925 109647 8928
rect 109589 8919 109647 8925
rect 112993 8925 113005 8928
rect 113039 8925 113051 8959
rect 112993 8919 113051 8925
rect 114373 8959 114431 8965
rect 114373 8925 114385 8959
rect 114419 8925 114431 8959
rect 114373 8919 114431 8925
rect 117133 8959 117191 8965
rect 117133 8925 117145 8959
rect 117179 8956 117191 8959
rect 118145 8959 118203 8965
rect 118145 8956 118157 8959
rect 117179 8928 118157 8956
rect 117179 8925 117191 8928
rect 117133 8919 117191 8925
rect 118145 8925 118157 8928
rect 118191 8925 118203 8959
rect 118252 8956 118280 8996
rect 119706 8984 119712 8996
rect 119764 8984 119770 9036
rect 122190 8984 122196 9036
rect 122248 9024 122254 9036
rect 123021 9027 123079 9033
rect 123021 9024 123033 9027
rect 122248 8996 123033 9024
rect 122248 8984 122254 8996
rect 123021 8993 123033 8996
rect 123067 8993 123079 9027
rect 124398 9024 124404 9036
rect 124359 8996 124404 9024
rect 123021 8987 123079 8993
rect 124398 8984 124404 8996
rect 124456 8984 124462 9036
rect 125965 9027 126023 9033
rect 125965 8993 125977 9027
rect 126011 9024 126023 9027
rect 128078 9024 128084 9036
rect 126011 8996 128084 9024
rect 126011 8993 126023 8996
rect 125965 8987 126023 8993
rect 128078 8984 128084 8996
rect 128136 8984 128142 9036
rect 128446 9024 128452 9036
rect 128407 8996 128452 9024
rect 128446 8984 128452 8996
rect 128504 8984 128510 9036
rect 129550 9024 129556 9036
rect 129511 8996 129556 9024
rect 129550 8984 129556 8996
rect 129608 8984 129614 9036
rect 130378 8984 130384 9036
rect 130436 9024 130442 9036
rect 134518 9024 134524 9036
rect 130436 8996 134380 9024
rect 134479 8996 134524 9024
rect 130436 8984 130442 8996
rect 120350 8956 120356 8968
rect 118252 8928 120356 8956
rect 118145 8919 118203 8925
rect 120350 8916 120356 8928
rect 120408 8916 120414 8968
rect 120537 8959 120595 8965
rect 120537 8925 120549 8959
rect 120583 8956 120595 8959
rect 121917 8959 121975 8965
rect 121917 8956 121929 8959
rect 120583 8928 121929 8956
rect 120583 8925 120595 8928
rect 120537 8919 120595 8925
rect 121917 8925 121929 8928
rect 121963 8925 121975 8959
rect 130470 8956 130476 8968
rect 121917 8919 121975 8925
rect 125612 8928 130476 8956
rect 117222 8888 117228 8900
rect 96724 8860 117228 8888
rect 117222 8848 117228 8860
rect 117280 8848 117286 8900
rect 119617 8891 119675 8897
rect 119617 8857 119629 8891
rect 119663 8888 119675 8891
rect 119706 8888 119712 8900
rect 119663 8860 119712 8888
rect 119663 8857 119675 8860
rect 119617 8851 119675 8857
rect 119706 8848 119712 8860
rect 119764 8848 119770 8900
rect 123389 8891 123447 8897
rect 123389 8857 123401 8891
rect 123435 8888 123447 8891
rect 125612 8888 125640 8928
rect 130470 8916 130476 8928
rect 130528 8916 130534 8968
rect 130838 8956 130844 8968
rect 130799 8928 130844 8956
rect 130838 8916 130844 8928
rect 130896 8916 130902 8968
rect 131853 8959 131911 8965
rect 131853 8925 131865 8959
rect 131899 8925 131911 8959
rect 131853 8919 131911 8925
rect 133141 8959 133199 8965
rect 133141 8925 133153 8959
rect 133187 8956 133199 8959
rect 133322 8956 133328 8968
rect 133187 8928 133328 8956
rect 133187 8925 133199 8928
rect 133141 8919 133199 8925
rect 125870 8888 125876 8900
rect 123435 8860 125640 8888
rect 125831 8860 125876 8888
rect 123435 8857 123447 8860
rect 123389 8851 123447 8857
rect 125870 8848 125876 8860
rect 125928 8848 125934 8900
rect 129366 8848 129372 8900
rect 129424 8888 129430 8900
rect 129737 8891 129795 8897
rect 129737 8888 129749 8891
rect 129424 8860 129749 8888
rect 129424 8848 129430 8860
rect 129737 8857 129749 8860
rect 129783 8857 129795 8891
rect 129737 8851 129795 8857
rect 88610 8820 88616 8832
rect 82924 8792 88616 8820
rect 88610 8780 88616 8792
rect 88668 8780 88674 8832
rect 97442 8780 97448 8832
rect 97500 8820 97506 8832
rect 102594 8820 102600 8832
rect 97500 8792 102600 8820
rect 97500 8780 97506 8792
rect 102594 8780 102600 8792
rect 102652 8780 102658 8832
rect 107286 8780 107292 8832
rect 107344 8820 107350 8832
rect 107749 8823 107807 8829
rect 107749 8820 107761 8823
rect 107344 8792 107761 8820
rect 107344 8780 107350 8792
rect 107749 8789 107761 8792
rect 107795 8789 107807 8823
rect 107749 8783 107807 8789
rect 110785 8823 110843 8829
rect 110785 8789 110797 8823
rect 110831 8820 110843 8823
rect 111150 8820 111156 8832
rect 110831 8792 111156 8820
rect 110831 8789 110843 8792
rect 110785 8783 110843 8789
rect 111150 8780 111156 8792
rect 111208 8780 111214 8832
rect 118418 8780 118424 8832
rect 118476 8820 118482 8832
rect 125226 8820 125232 8832
rect 118476 8792 125232 8820
rect 118476 8780 118482 8792
rect 125226 8780 125232 8792
rect 125284 8780 125290 8832
rect 127802 8780 127808 8832
rect 127860 8820 127866 8832
rect 131868 8820 131896 8919
rect 133322 8916 133328 8928
rect 133380 8916 133386 8968
rect 134352 8956 134380 8996
rect 134518 8984 134524 8996
rect 134576 8984 134582 9036
rect 135070 8984 135076 9036
rect 135128 9024 135134 9036
rect 135625 9027 135683 9033
rect 135625 9024 135637 9027
rect 135128 8996 135637 9024
rect 135128 8984 135134 8996
rect 135625 8993 135637 8996
rect 135671 8993 135683 9027
rect 136910 9024 136916 9036
rect 136871 8996 136916 9024
rect 135625 8987 135683 8993
rect 136910 8984 136916 8996
rect 136968 8984 136974 9036
rect 138382 8984 138388 9036
rect 138440 9024 138446 9036
rect 144380 9033 144408 9064
rect 147674 9052 147680 9064
rect 147732 9052 147738 9104
rect 150710 9052 150716 9104
rect 150768 9092 150774 9104
rect 162118 9092 162124 9104
rect 150768 9064 162124 9092
rect 150768 9052 150774 9064
rect 162118 9052 162124 9064
rect 162176 9052 162182 9104
rect 165614 9092 165620 9104
rect 164252 9064 165620 9092
rect 139857 9027 139915 9033
rect 139857 9024 139869 9027
rect 138440 8996 139869 9024
rect 138440 8984 138446 8996
rect 139857 8993 139869 8996
rect 139903 8993 139915 9027
rect 143169 9027 143227 9033
rect 143169 9024 143181 9027
rect 139857 8987 139915 8993
rect 140976 8996 143181 9024
rect 137830 8956 137836 8968
rect 134352 8928 137836 8956
rect 137830 8916 137836 8928
rect 137888 8916 137894 8968
rect 138753 8959 138811 8965
rect 138753 8925 138765 8959
rect 138799 8956 138811 8959
rect 140976 8956 141004 8996
rect 143169 8993 143181 8996
rect 143215 8993 143227 9027
rect 143169 8987 143227 8993
rect 144365 9027 144423 9033
rect 144365 8993 144377 9027
rect 144411 8993 144423 9027
rect 145466 9024 145472 9036
rect 145427 8996 145472 9024
rect 144365 8987 144423 8993
rect 145466 8984 145472 8996
rect 145524 8984 145530 9036
rect 147861 9027 147919 9033
rect 147861 9024 147873 9027
rect 145576 8996 147873 9024
rect 141142 8956 141148 8968
rect 138799 8928 141004 8956
rect 141103 8928 141148 8956
rect 138799 8925 138811 8928
rect 138753 8919 138811 8925
rect 141142 8916 141148 8928
rect 141200 8916 141206 8968
rect 142154 8956 142160 8968
rect 142115 8928 142160 8956
rect 142154 8916 142160 8928
rect 142212 8916 142218 8968
rect 144730 8916 144736 8968
rect 144788 8956 144794 8968
rect 145576 8956 145604 8996
rect 147861 8993 147873 8996
rect 147907 8993 147919 9027
rect 147861 8987 147919 8993
rect 150434 8984 150440 9036
rect 150492 9024 150498 9036
rect 154209 9027 154267 9033
rect 154209 9024 154221 9027
rect 150492 8996 154221 9024
rect 150492 8984 150498 8996
rect 154209 8993 154221 8996
rect 154255 8993 154267 9027
rect 156690 9024 156696 9036
rect 156651 8996 156696 9024
rect 154209 8987 154267 8993
rect 156690 8984 156696 8996
rect 156748 8984 156754 9036
rect 156874 8984 156880 9036
rect 156932 9024 156938 9036
rect 160186 9024 160192 9036
rect 156932 8996 160192 9024
rect 156932 8984 156938 8996
rect 160186 8984 160192 8996
rect 160244 8984 160250 9036
rect 164252 9033 164280 9064
rect 165614 9052 165620 9064
rect 165672 9052 165678 9104
rect 166442 9052 166448 9104
rect 166500 9092 166506 9104
rect 170950 9092 170956 9104
rect 166500 9064 170956 9092
rect 166500 9052 166506 9064
rect 170950 9052 170956 9064
rect 171008 9052 171014 9104
rect 164237 9027 164295 9033
rect 164237 8993 164249 9027
rect 164283 8993 164295 9027
rect 164237 8987 164295 8993
rect 164326 8984 164332 9036
rect 164384 9024 164390 9036
rect 167457 9027 167515 9033
rect 167457 9024 167469 9027
rect 164384 8996 167469 9024
rect 164384 8984 164390 8996
rect 167457 8993 167469 8996
rect 167503 8993 167515 9027
rect 169018 9024 169024 9036
rect 168979 8996 169024 9024
rect 167457 8987 167515 8993
rect 169018 8984 169024 8996
rect 169076 8984 169082 9036
rect 169938 9024 169944 9036
rect 169899 8996 169944 9024
rect 169938 8984 169944 8996
rect 169996 8984 170002 9036
rect 171226 9024 171232 9036
rect 171187 8996 171232 9024
rect 171226 8984 171232 8996
rect 171284 8984 171290 9036
rect 145834 8956 145840 8968
rect 144788 8928 145604 8956
rect 145795 8928 145840 8956
rect 144788 8916 144794 8928
rect 145834 8916 145840 8928
rect 145892 8916 145898 8968
rect 146757 8959 146815 8965
rect 146757 8925 146769 8959
rect 146803 8956 146815 8959
rect 149977 8959 150035 8965
rect 149977 8956 149989 8959
rect 146803 8928 149989 8956
rect 146803 8925 146815 8928
rect 146757 8919 146815 8925
rect 149977 8925 149989 8928
rect 150023 8925 150035 8959
rect 151078 8956 151084 8968
rect 151039 8928 151084 8956
rect 149977 8919 150035 8925
rect 151078 8916 151084 8928
rect 151136 8916 151142 8968
rect 152826 8916 152832 8968
rect 152884 8956 152890 8968
rect 153105 8959 153163 8965
rect 153105 8956 153117 8959
rect 152884 8928 153117 8956
rect 152884 8916 152890 8928
rect 153105 8925 153117 8928
rect 153151 8925 153163 8959
rect 154482 8956 154488 8968
rect 154443 8928 154488 8956
rect 153105 8919 153163 8925
rect 154482 8916 154488 8928
rect 154540 8916 154546 8968
rect 155589 8959 155647 8965
rect 155589 8925 155601 8959
rect 155635 8956 155647 8959
rect 156230 8956 156236 8968
rect 155635 8928 156236 8956
rect 155635 8925 155647 8928
rect 155589 8919 155647 8925
rect 156230 8916 156236 8928
rect 156288 8916 156294 8968
rect 157978 8956 157984 8968
rect 157939 8928 157984 8956
rect 157978 8916 157984 8928
rect 158036 8916 158042 8968
rect 159085 8959 159143 8965
rect 159085 8925 159097 8959
rect 159131 8956 159143 8959
rect 160002 8956 160008 8968
rect 159131 8928 160008 8956
rect 159131 8925 159143 8928
rect 159085 8919 159143 8925
rect 160002 8916 160008 8928
rect 160060 8916 160066 8968
rect 161934 8956 161940 8968
rect 161895 8928 161940 8956
rect 161934 8916 161940 8928
rect 161992 8916 161998 8968
rect 162949 8959 163007 8965
rect 162949 8925 162961 8959
rect 162995 8956 163007 8959
rect 165341 8959 165399 8965
rect 165341 8956 165353 8959
rect 162995 8928 165353 8956
rect 162995 8925 163007 8928
rect 162949 8919 163007 8925
rect 165341 8925 165353 8928
rect 165387 8925 165399 8959
rect 169202 8956 169208 8968
rect 165341 8919 165399 8925
rect 165448 8928 169208 8956
rect 135993 8891 136051 8897
rect 135993 8857 136005 8891
rect 136039 8888 136051 8891
rect 140222 8888 140228 8900
rect 136039 8860 140084 8888
rect 140183 8860 140228 8888
rect 136039 8857 136051 8860
rect 135993 8851 136051 8857
rect 127860 8792 131896 8820
rect 127860 8780 127866 8792
rect 132218 8780 132224 8832
rect 132276 8820 132282 8832
rect 139118 8820 139124 8832
rect 132276 8792 139124 8820
rect 132276 8780 132282 8792
rect 139118 8780 139124 8792
rect 139176 8780 139182 8832
rect 140056 8820 140084 8860
rect 140222 8848 140228 8860
rect 140280 8848 140286 8900
rect 148226 8888 148232 8900
rect 148187 8860 148232 8888
rect 148226 8848 148232 8860
rect 148284 8848 148290 8900
rect 157061 8891 157119 8897
rect 157061 8857 157073 8891
rect 157107 8888 157119 8891
rect 164418 8888 164424 8900
rect 157107 8860 162164 8888
rect 164379 8860 164424 8888
rect 157107 8857 157119 8860
rect 157061 8851 157119 8857
rect 141234 8820 141240 8832
rect 140056 8792 141240 8820
rect 141234 8780 141240 8792
rect 141292 8780 141298 8832
rect 157150 8780 157156 8832
rect 157208 8820 157214 8832
rect 160462 8820 160468 8832
rect 157208 8792 160468 8820
rect 157208 8780 157214 8792
rect 160462 8780 160468 8792
rect 160520 8780 160526 8832
rect 162136 8820 162164 8860
rect 164418 8848 164424 8860
rect 164476 8848 164482 8900
rect 164786 8848 164792 8900
rect 164844 8888 164850 8900
rect 165448 8888 165476 8928
rect 169202 8916 169208 8928
rect 169260 8916 169266 8968
rect 171428 8965 171456 9132
rect 179506 9120 179512 9132
rect 179564 9120 179570 9172
rect 179601 9163 179659 9169
rect 179601 9129 179613 9163
rect 179647 9160 179659 9163
rect 184474 9160 184480 9172
rect 179647 9132 184480 9160
rect 179647 9129 179659 9132
rect 179601 9123 179659 9129
rect 184474 9120 184480 9132
rect 184532 9120 184538 9172
rect 192110 9160 192116 9172
rect 187804 9132 192116 9160
rect 171502 9052 171508 9104
rect 171560 9092 171566 9104
rect 187804 9092 187832 9132
rect 192110 9120 192116 9132
rect 192168 9120 192174 9172
rect 197354 9160 197360 9172
rect 197315 9132 197360 9160
rect 197354 9120 197360 9132
rect 197412 9120 197418 9172
rect 171560 9064 187832 9092
rect 171560 9052 171566 9064
rect 187878 9052 187884 9104
rect 187936 9092 187942 9104
rect 198458 9092 198464 9104
rect 187936 9064 198464 9092
rect 187936 9052 187942 9064
rect 198458 9052 198464 9064
rect 198516 9052 198522 9104
rect 174906 9024 174912 9036
rect 174867 8996 174912 9024
rect 174906 8984 174912 8996
rect 174964 8984 174970 9036
rect 181622 9024 181628 9036
rect 179708 8996 181628 9024
rect 171413 8959 171471 8965
rect 171413 8925 171425 8959
rect 171459 8925 171471 8959
rect 171413 8919 171471 8925
rect 172793 8959 172851 8965
rect 172793 8925 172805 8959
rect 172839 8956 172851 8959
rect 173710 8956 173716 8968
rect 172839 8928 173716 8956
rect 172839 8925 172851 8928
rect 172793 8919 172851 8925
rect 173710 8916 173716 8928
rect 173768 8916 173774 8968
rect 173805 8959 173863 8965
rect 173805 8925 173817 8959
rect 173851 8956 173863 8959
rect 176841 8959 176899 8965
rect 176841 8956 176853 8959
rect 173851 8928 176853 8956
rect 173851 8925 173863 8928
rect 173805 8919 173863 8925
rect 176841 8925 176853 8928
rect 176887 8925 176899 8959
rect 178034 8956 178040 8968
rect 177995 8928 178040 8956
rect 176841 8919 176899 8925
rect 178034 8916 178040 8928
rect 178092 8916 178098 8968
rect 164844 8860 165476 8888
rect 168929 8891 168987 8897
rect 164844 8848 164850 8860
rect 168929 8857 168941 8891
rect 168975 8888 168987 8891
rect 172514 8888 172520 8900
rect 168975 8860 172520 8888
rect 168975 8857 168987 8860
rect 168929 8851 168987 8857
rect 172514 8848 172520 8860
rect 172572 8848 172578 8900
rect 175277 8891 175335 8897
rect 175277 8857 175289 8891
rect 175323 8888 175335 8891
rect 179708 8888 179736 8996
rect 181622 8984 181628 8996
rect 181680 8984 181686 9036
rect 181990 9024 181996 9036
rect 181951 8996 181996 9024
rect 181990 8984 181996 8996
rect 182048 8984 182054 9036
rect 182634 8984 182640 9036
rect 182692 9024 182698 9036
rect 184566 9024 184572 9036
rect 182692 8996 184572 9024
rect 182692 8984 182698 8996
rect 184566 8984 184572 8996
rect 184624 8984 184630 9036
rect 186222 9024 186228 9036
rect 186183 8996 186228 9024
rect 186222 8984 186228 8996
rect 186280 8984 186286 9036
rect 189350 8984 189356 9036
rect 189408 9024 189414 9036
rect 190641 9027 190699 9033
rect 190641 9024 190653 9027
rect 189408 8996 190653 9024
rect 189408 8984 189414 8996
rect 190641 8993 190653 8996
rect 190687 8993 190699 9027
rect 191926 9024 191932 9036
rect 191887 8996 191932 9024
rect 190641 8987 190699 8993
rect 191926 8984 191932 8996
rect 191984 8984 191990 9036
rect 193033 9027 193091 9033
rect 193033 8993 193045 9027
rect 193079 8993 193091 9027
rect 196434 9024 196440 9036
rect 196395 8996 196440 9024
rect 193033 8987 193091 8993
rect 180613 8959 180671 8965
rect 180613 8925 180625 8959
rect 180659 8956 180671 8959
rect 183649 8959 183707 8965
rect 183649 8956 183661 8959
rect 180659 8928 183661 8956
rect 180659 8925 180671 8928
rect 180613 8919 180671 8925
rect 183649 8925 183661 8928
rect 183695 8925 183707 8959
rect 184842 8956 184848 8968
rect 184803 8928 184848 8956
rect 183649 8919 183707 8925
rect 184842 8916 184848 8928
rect 184900 8916 184906 8968
rect 184934 8916 184940 8968
rect 184992 8956 184998 8968
rect 187510 8956 187516 8968
rect 184992 8928 187516 8956
rect 184992 8916 184998 8928
rect 187510 8916 187516 8928
rect 187568 8916 187574 8968
rect 188157 8959 188215 8965
rect 188157 8925 188169 8959
rect 188203 8956 188215 8959
rect 189537 8959 189595 8965
rect 189537 8956 189549 8959
rect 188203 8928 189549 8956
rect 188203 8925 188215 8928
rect 188157 8919 188215 8925
rect 189537 8925 189549 8928
rect 189583 8925 189595 8959
rect 189537 8919 189595 8925
rect 191009 8959 191067 8965
rect 191009 8925 191021 8959
rect 191055 8956 191067 8959
rect 191466 8956 191472 8968
rect 191055 8928 191472 8956
rect 191055 8925 191067 8928
rect 191009 8919 191067 8925
rect 191466 8916 191472 8928
rect 191524 8916 191530 8968
rect 192294 8916 192300 8968
rect 192352 8956 192358 8968
rect 192941 8959 192999 8965
rect 192941 8956 192953 8959
rect 192352 8928 192953 8956
rect 192352 8916 192358 8928
rect 192941 8925 192953 8928
rect 192987 8925 192999 8959
rect 192941 8919 192999 8925
rect 182082 8888 182088 8900
rect 175323 8860 179736 8888
rect 182043 8860 182088 8888
rect 175323 8857 175335 8860
rect 175277 8851 175335 8857
rect 182082 8848 182088 8860
rect 182140 8848 182146 8900
rect 183554 8888 183560 8900
rect 182192 8860 183560 8888
rect 173158 8820 173164 8832
rect 162136 8792 173164 8820
rect 173158 8780 173164 8792
rect 173216 8780 173222 8832
rect 174262 8780 174268 8832
rect 174320 8820 174326 8832
rect 176746 8820 176752 8832
rect 174320 8792 176752 8820
rect 174320 8780 174326 8792
rect 176746 8780 176752 8792
rect 176804 8780 176810 8832
rect 176838 8780 176844 8832
rect 176896 8820 176902 8832
rect 182192 8820 182220 8860
rect 183554 8848 183560 8860
rect 183612 8848 183618 8900
rect 186133 8891 186191 8897
rect 186133 8857 186145 8891
rect 186179 8888 186191 8891
rect 189718 8888 189724 8900
rect 186179 8860 189724 8888
rect 186179 8857 186191 8860
rect 186133 8851 186191 8857
rect 189718 8848 189724 8860
rect 189776 8848 189782 8900
rect 190730 8848 190736 8900
rect 190788 8888 190794 8900
rect 193048 8888 193076 8987
rect 196434 8984 196440 8996
rect 196492 8984 196498 9036
rect 197262 9024 197268 9036
rect 197223 8996 197268 9024
rect 197262 8984 197268 8996
rect 197320 8984 197326 9036
rect 194870 8956 194876 8968
rect 194831 8928 194876 8956
rect 194870 8916 194876 8928
rect 194928 8916 194934 8968
rect 195330 8916 195336 8968
rect 195388 8956 195394 8968
rect 196069 8959 196127 8965
rect 196069 8956 196081 8959
rect 195388 8928 196081 8956
rect 195388 8916 195394 8928
rect 196069 8925 196081 8928
rect 196115 8925 196127 8959
rect 196069 8919 196127 8925
rect 190788 8860 193076 8888
rect 190788 8848 190794 8860
rect 176896 8792 182220 8820
rect 176896 8780 176902 8792
rect 182818 8780 182824 8832
rect 182876 8820 182882 8832
rect 197354 8820 197360 8832
rect 182876 8792 197360 8820
rect 182876 8780 182882 8792
rect 197354 8780 197360 8792
rect 197412 8780 197418 8832
rect 1104 8730 198812 8752
rect 1104 8678 4078 8730
rect 4130 8678 44078 8730
rect 44130 8678 84078 8730
rect 84130 8678 124078 8730
rect 124130 8678 164078 8730
rect 164130 8678 198812 8730
rect 1104 8656 198812 8678
rect 48498 8576 48504 8628
rect 48556 8616 48562 8628
rect 48556 8588 52224 8616
rect 48556 8576 48562 8588
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 11572 8520 15424 8548
rect 11572 8508 11578 8520
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5040 8452 5549 8480
rect 5040 8440 5046 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 6822 8480 6828 8492
rect 6783 8452 6828 8480
rect 5537 8443 5595 8449
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 7834 8480 7840 8492
rect 7795 8452 7840 8480
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 14366 8480 14372 8492
rect 14327 8452 14372 8480
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 15396 8489 15424 8520
rect 19794 8508 19800 8560
rect 19852 8548 19858 8560
rect 26421 8551 26479 8557
rect 19852 8520 21496 8548
rect 19852 8508 19858 8520
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 16758 8480 16764 8492
rect 16719 8452 16764 8480
rect 15381 8443 15439 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 20438 8480 20444 8492
rect 20399 8452 20444 8480
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 21468 8489 21496 8520
rect 26421 8517 26433 8551
rect 26467 8548 26479 8551
rect 28074 8548 28080 8560
rect 26467 8520 28080 8548
rect 26467 8517 26479 8520
rect 26421 8511 26479 8517
rect 28074 8508 28080 8520
rect 28132 8508 28138 8560
rect 30745 8551 30803 8557
rect 30745 8517 30757 8551
rect 30791 8548 30803 8551
rect 31570 8548 31576 8560
rect 30791 8520 31576 8548
rect 30791 8517 30803 8520
rect 30745 8511 30803 8517
rect 31570 8508 31576 8520
rect 31628 8508 31634 8560
rect 46382 8508 46388 8560
rect 46440 8548 46446 8560
rect 46440 8520 48636 8548
rect 46440 8508 46446 8520
rect 21453 8483 21511 8489
rect 21453 8449 21465 8483
rect 21499 8449 21511 8483
rect 29270 8480 29276 8492
rect 29231 8452 29276 8480
rect 21453 8443 21511 8449
rect 29270 8440 29276 8452
rect 29328 8440 29334 8492
rect 31941 8483 31999 8489
rect 31941 8449 31953 8483
rect 31987 8480 31999 8483
rect 32214 8480 32220 8492
rect 31987 8452 32220 8480
rect 31987 8449 31999 8452
rect 31941 8443 31999 8449
rect 32214 8440 32220 8452
rect 32272 8440 32278 8492
rect 33226 8480 33232 8492
rect 33187 8452 33232 8480
rect 33226 8440 33232 8452
rect 33284 8440 33290 8492
rect 34146 8440 34152 8492
rect 34204 8480 34210 8492
rect 37737 8483 37795 8489
rect 37737 8480 37749 8483
rect 34204 8452 37749 8480
rect 34204 8440 34210 8452
rect 37737 8449 37749 8452
rect 37783 8449 37795 8483
rect 39114 8480 39120 8492
rect 39075 8452 39120 8480
rect 37737 8443 37795 8449
rect 39114 8440 39120 8452
rect 39172 8440 39178 8492
rect 40954 8480 40960 8492
rect 40915 8452 40960 8480
rect 40954 8440 40960 8452
rect 41012 8440 41018 8492
rect 41414 8440 41420 8492
rect 41472 8480 41478 8492
rect 42981 8483 43039 8489
rect 42981 8480 42993 8483
rect 41472 8452 42993 8480
rect 41472 8440 41478 8452
rect 42981 8449 42993 8452
rect 43027 8449 43039 8483
rect 42981 8443 43039 8449
rect 43714 8440 43720 8492
rect 43772 8480 43778 8492
rect 46109 8483 46167 8489
rect 46109 8480 46121 8483
rect 43772 8452 46121 8480
rect 43772 8440 43778 8452
rect 46109 8449 46121 8452
rect 46155 8449 46167 8483
rect 47578 8480 47584 8492
rect 47539 8452 47584 8480
rect 46109 8443 46167 8449
rect 47578 8440 47584 8452
rect 47636 8440 47642 8492
rect 48608 8489 48636 8520
rect 48593 8483 48651 8489
rect 48593 8449 48605 8483
rect 48639 8449 48651 8483
rect 52196 8480 52224 8588
rect 77386 8576 77392 8628
rect 77444 8616 77450 8628
rect 82262 8616 82268 8628
rect 77444 8588 82268 8616
rect 77444 8576 77450 8588
rect 82262 8576 82268 8588
rect 82320 8576 82326 8628
rect 82814 8576 82820 8628
rect 82872 8616 82878 8628
rect 83918 8616 83924 8628
rect 82872 8588 83924 8616
rect 82872 8576 82878 8588
rect 83918 8576 83924 8588
rect 83976 8576 83982 8628
rect 87049 8619 87107 8625
rect 87049 8585 87061 8619
rect 87095 8616 87107 8619
rect 91094 8616 91100 8628
rect 87095 8588 91100 8616
rect 87095 8585 87107 8588
rect 87049 8579 87107 8585
rect 91094 8576 91100 8588
rect 91152 8576 91158 8628
rect 96706 8576 96712 8628
rect 96764 8616 96770 8628
rect 99558 8616 99564 8628
rect 96764 8588 99564 8616
rect 96764 8576 96770 8588
rect 99558 8576 99564 8588
rect 99616 8576 99622 8628
rect 103241 8619 103299 8625
rect 103241 8616 103253 8619
rect 100404 8588 103253 8616
rect 60458 8508 60464 8560
rect 60516 8548 60522 8560
rect 75822 8548 75828 8560
rect 60516 8520 62988 8548
rect 60516 8508 60522 8520
rect 55677 8483 55735 8489
rect 55677 8480 55689 8483
rect 52196 8452 55689 8480
rect 48593 8443 48651 8449
rect 55677 8449 55689 8452
rect 55723 8449 55735 8483
rect 59538 8480 59544 8492
rect 59499 8452 59544 8480
rect 55677 8443 55735 8449
rect 59538 8440 59544 8452
rect 59596 8440 59602 8492
rect 60826 8480 60832 8492
rect 60787 8452 60832 8480
rect 60826 8440 60832 8452
rect 60884 8440 60890 8492
rect 62960 8489 62988 8520
rect 71792 8520 75828 8548
rect 62945 8483 63003 8489
rect 62945 8449 62957 8483
rect 62991 8449 63003 8483
rect 66070 8480 66076 8492
rect 66031 8452 66076 8480
rect 62945 8443 63003 8449
rect 66070 8440 66076 8452
rect 66128 8440 66134 8492
rect 67082 8480 67088 8492
rect 67043 8452 67088 8480
rect 67082 8440 67088 8452
rect 67140 8440 67146 8492
rect 71792 8480 71820 8520
rect 75822 8508 75828 8520
rect 75880 8508 75886 8560
rect 80238 8548 80244 8560
rect 76944 8520 80244 8548
rect 75086 8480 75092 8492
rect 71516 8452 71820 8480
rect 73264 8452 75092 8480
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8381 4399 8415
rect 5626 8412 5632 8424
rect 5587 8384 5632 8412
rect 4341 8375 4399 8381
rect 4356 8344 4384 8375
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 5776 8384 7941 8412
rect 5776 8372 5782 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 11422 8372 11428 8424
rect 11480 8412 11486 8424
rect 15473 8415 15531 8421
rect 15473 8412 15485 8415
rect 11480 8384 15485 8412
rect 11480 8372 11486 8384
rect 15473 8381 15485 8384
rect 15519 8381 15531 8415
rect 15473 8375 15531 8381
rect 18966 8372 18972 8424
rect 19024 8412 19030 8424
rect 21545 8415 21603 8421
rect 21545 8412 21557 8415
rect 19024 8384 21557 8412
rect 19024 8372 19030 8384
rect 21545 8381 21557 8384
rect 21591 8381 21603 8415
rect 24946 8412 24952 8424
rect 24907 8384 24952 8412
rect 21545 8375 21603 8381
rect 24946 8372 24952 8384
rect 25004 8372 25010 8424
rect 26050 8412 26056 8424
rect 26011 8384 26056 8412
rect 26050 8372 26056 8384
rect 26108 8372 26114 8424
rect 29086 8372 29092 8424
rect 29144 8412 29150 8424
rect 30377 8415 30435 8421
rect 30377 8412 30389 8415
rect 29144 8384 30389 8412
rect 29144 8372 29150 8384
rect 30377 8381 30389 8384
rect 30423 8381 30435 8415
rect 33042 8412 33048 8424
rect 33003 8384 33048 8412
rect 30377 8375 30435 8381
rect 33042 8372 33048 8384
rect 33100 8372 33106 8424
rect 36725 8415 36783 8421
rect 36725 8381 36737 8415
rect 36771 8412 36783 8415
rect 37550 8412 37556 8424
rect 36771 8384 37556 8412
rect 36771 8381 36783 8384
rect 36725 8375 36783 8381
rect 37550 8372 37556 8384
rect 37608 8372 37614 8424
rect 37829 8415 37887 8421
rect 37829 8381 37841 8415
rect 37875 8381 37887 8415
rect 41966 8412 41972 8424
rect 41927 8384 41972 8412
rect 37829 8375 37887 8381
rect 7374 8344 7380 8356
rect 4356 8316 7380 8344
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 11514 8304 11520 8356
rect 11572 8344 11578 8356
rect 12437 8347 12495 8353
rect 12437 8344 12449 8347
rect 11572 8316 12449 8344
rect 11572 8304 11578 8316
rect 12437 8313 12449 8316
rect 12483 8313 12495 8347
rect 12437 8307 12495 8313
rect 35986 8304 35992 8356
rect 36044 8344 36050 8356
rect 37844 8344 37872 8375
rect 41966 8372 41972 8384
rect 42024 8372 42030 8424
rect 43530 8412 43536 8424
rect 43491 8384 43536 8412
rect 43530 8372 43536 8384
rect 43588 8372 43594 8424
rect 46474 8372 46480 8424
rect 46532 8412 46538 8424
rect 48685 8415 48743 8421
rect 48685 8412 48697 8415
rect 46532 8384 48697 8412
rect 46532 8372 46538 8384
rect 48685 8381 48697 8384
rect 48731 8381 48743 8415
rect 48685 8375 48743 8381
rect 52086 8372 52092 8424
rect 52144 8412 52150 8424
rect 54662 8412 54668 8424
rect 52144 8384 54248 8412
rect 54623 8384 54668 8412
rect 52144 8372 52150 8384
rect 36044 8316 37872 8344
rect 36044 8304 36050 8316
rect 48958 8304 48964 8356
rect 49016 8344 49022 8356
rect 49973 8347 50031 8353
rect 49973 8344 49985 8347
rect 49016 8316 49985 8344
rect 49016 8304 49022 8316
rect 49973 8313 49985 8316
rect 50019 8313 50031 8347
rect 49973 8307 50031 8313
rect 53653 8347 53711 8353
rect 53653 8313 53665 8347
rect 53699 8344 53711 8347
rect 54110 8344 54116 8356
rect 53699 8316 54116 8344
rect 53699 8313 53711 8316
rect 53653 8307 53711 8313
rect 54110 8304 54116 8316
rect 54168 8304 54174 8356
rect 54220 8344 54248 8384
rect 54662 8372 54668 8384
rect 54720 8372 54726 8424
rect 55769 8415 55827 8421
rect 55769 8381 55781 8415
rect 55815 8381 55827 8415
rect 55769 8375 55827 8381
rect 55784 8344 55812 8375
rect 59630 8372 59636 8424
rect 59688 8412 59694 8424
rect 60645 8415 60703 8421
rect 60645 8412 60657 8415
rect 59688 8384 60657 8412
rect 59688 8372 59694 8384
rect 60645 8381 60657 8384
rect 60691 8381 60703 8415
rect 60645 8375 60703 8381
rect 63678 8372 63684 8424
rect 63736 8412 63742 8424
rect 67177 8415 67235 8421
rect 67177 8412 67189 8415
rect 63736 8384 67189 8412
rect 63736 8372 63742 8384
rect 67177 8381 67189 8384
rect 67223 8381 67235 8415
rect 70946 8412 70952 8424
rect 70907 8384 70952 8412
rect 67177 8375 67235 8381
rect 70946 8372 70952 8384
rect 71004 8372 71010 8424
rect 71314 8412 71320 8424
rect 71275 8384 71320 8412
rect 71314 8372 71320 8384
rect 71372 8372 71378 8424
rect 71516 8421 71544 8452
rect 71501 8415 71559 8421
rect 71501 8381 71513 8415
rect 71547 8381 71559 8415
rect 71501 8375 71559 8381
rect 71590 8372 71596 8424
rect 71648 8412 71654 8424
rect 72513 8415 72571 8421
rect 72513 8412 72525 8415
rect 71648 8384 72525 8412
rect 71648 8372 71654 8384
rect 72513 8381 72525 8384
rect 72559 8381 72571 8415
rect 72513 8375 72571 8381
rect 72881 8415 72939 8421
rect 72881 8381 72893 8415
rect 72927 8412 72939 8415
rect 73062 8412 73068 8424
rect 72927 8384 73068 8412
rect 72927 8381 72939 8384
rect 72881 8375 72939 8381
rect 73062 8372 73068 8384
rect 73120 8372 73126 8424
rect 73264 8421 73292 8452
rect 75086 8440 75092 8452
rect 75144 8440 75150 8492
rect 76944 8489 76972 8520
rect 80238 8508 80244 8520
rect 80296 8508 80302 8560
rect 82170 8548 82176 8560
rect 82131 8520 82176 8548
rect 82170 8508 82176 8520
rect 82228 8508 82234 8560
rect 92382 8548 92388 8560
rect 87708 8520 92388 8548
rect 76929 8483 76987 8489
rect 76929 8449 76941 8483
rect 76975 8449 76987 8483
rect 80698 8480 80704 8492
rect 80659 8452 80704 8480
rect 76929 8443 76987 8449
rect 80698 8440 80704 8452
rect 80756 8440 80762 8492
rect 82906 8480 82912 8492
rect 82096 8452 82912 8480
rect 73249 8415 73307 8421
rect 73249 8381 73261 8415
rect 73295 8381 73307 8415
rect 74442 8412 74448 8424
rect 74403 8384 74448 8412
rect 73249 8375 73307 8381
rect 74442 8372 74448 8384
rect 74500 8372 74506 8424
rect 74813 8415 74871 8421
rect 74813 8381 74825 8415
rect 74859 8381 74871 8415
rect 74813 8375 74871 8381
rect 75181 8415 75239 8421
rect 75181 8381 75193 8415
rect 75227 8412 75239 8415
rect 75362 8412 75368 8424
rect 75227 8384 75368 8412
rect 75227 8381 75239 8384
rect 75181 8375 75239 8381
rect 69014 8344 69020 8356
rect 54220 8316 55812 8344
rect 68975 8316 69020 8344
rect 69014 8304 69020 8316
rect 69072 8304 69078 8356
rect 74828 8344 74856 8375
rect 75362 8372 75368 8384
rect 75420 8372 75426 8424
rect 76834 8412 76840 8424
rect 76795 8384 76840 8412
rect 76834 8372 76840 8384
rect 76892 8372 76898 8424
rect 77205 8415 77263 8421
rect 77205 8381 77217 8415
rect 77251 8412 77263 8415
rect 82096 8412 82124 8452
rect 82906 8440 82912 8452
rect 82964 8440 82970 8492
rect 83550 8480 83556 8492
rect 83511 8452 83556 8480
rect 83550 8440 83556 8452
rect 83608 8440 83614 8492
rect 86954 8480 86960 8492
rect 85500 8452 86960 8480
rect 77251 8384 82124 8412
rect 82265 8415 82323 8421
rect 77251 8381 77263 8384
rect 77205 8375 77263 8381
rect 82265 8381 82277 8415
rect 82311 8412 82323 8415
rect 85500 8412 85528 8452
rect 86954 8440 86960 8452
rect 87012 8440 87018 8492
rect 85666 8412 85672 8424
rect 82311 8384 85528 8412
rect 85627 8384 85672 8412
rect 82311 8381 82323 8384
rect 82265 8375 82323 8381
rect 85666 8372 85672 8384
rect 85724 8372 85730 8424
rect 85761 8415 85819 8421
rect 85761 8381 85773 8415
rect 85807 8412 85819 8415
rect 85942 8412 85948 8424
rect 85807 8384 85948 8412
rect 85807 8381 85819 8384
rect 85761 8375 85819 8381
rect 85942 8372 85948 8384
rect 86000 8372 86006 8424
rect 86129 8415 86187 8421
rect 86129 8381 86141 8415
rect 86175 8381 86187 8415
rect 87230 8412 87236 8424
rect 87191 8384 87236 8412
rect 86129 8375 86187 8381
rect 74828 8316 78352 8344
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11333 8279 11391 8285
rect 11333 8276 11345 8279
rect 11204 8248 11345 8276
rect 11204 8236 11210 8248
rect 11333 8245 11345 8248
rect 11379 8245 11391 8279
rect 27338 8276 27344 8288
rect 27299 8248 27344 8276
rect 11333 8239 11391 8245
rect 27338 8236 27344 8248
rect 27396 8236 27402 8288
rect 34882 8276 34888 8288
rect 34843 8248 34888 8276
rect 34882 8236 34888 8248
rect 34940 8236 34946 8288
rect 44358 8276 44364 8288
rect 44319 8248 44364 8276
rect 44358 8236 44364 8248
rect 44416 8236 44422 8288
rect 58526 8276 58532 8288
rect 58487 8248 58532 8276
rect 58526 8236 58532 8248
rect 58584 8236 58590 8288
rect 63954 8276 63960 8288
rect 63915 8248 63960 8276
rect 63954 8236 63960 8248
rect 64012 8236 64018 8288
rect 64966 8276 64972 8288
rect 64927 8248 64972 8276
rect 64966 8236 64972 8248
rect 65024 8236 65030 8288
rect 78324 8276 78352 8316
rect 78398 8304 78404 8356
rect 78456 8344 78462 8356
rect 78585 8347 78643 8353
rect 78585 8344 78597 8347
rect 78456 8316 78597 8344
rect 78456 8304 78462 8316
rect 78585 8313 78597 8316
rect 78631 8313 78643 8347
rect 84378 8344 84384 8356
rect 78585 8307 78643 8313
rect 78692 8316 84384 8344
rect 78692 8276 78720 8316
rect 84378 8304 84384 8316
rect 84436 8304 84442 8356
rect 86144 8344 86172 8375
rect 87230 8372 87236 8384
rect 87288 8372 87294 8424
rect 87708 8421 87736 8520
rect 92382 8508 92388 8520
rect 92440 8508 92446 8560
rect 98546 8548 98552 8560
rect 95068 8520 98552 8548
rect 93394 8480 93400 8492
rect 89272 8452 93400 8480
rect 87693 8415 87751 8421
rect 87693 8381 87705 8415
rect 87739 8381 87751 8415
rect 87693 8375 87751 8381
rect 88334 8372 88340 8424
rect 88392 8412 88398 8424
rect 88521 8415 88579 8421
rect 88521 8412 88533 8415
rect 88392 8384 88533 8412
rect 88392 8372 88398 8384
rect 88521 8381 88533 8384
rect 88567 8381 88579 8415
rect 88886 8412 88892 8424
rect 88847 8384 88892 8412
rect 88521 8375 88579 8381
rect 88886 8372 88892 8384
rect 88944 8372 88950 8424
rect 89272 8421 89300 8452
rect 93394 8440 93400 8452
rect 93452 8440 93458 8492
rect 93670 8480 93676 8492
rect 93631 8452 93676 8480
rect 93670 8440 93676 8452
rect 93728 8440 93734 8492
rect 95068 8489 95096 8520
rect 98546 8508 98552 8520
rect 98604 8508 98610 8560
rect 100404 8557 100432 8588
rect 103241 8585 103253 8588
rect 103287 8585 103299 8619
rect 103241 8579 103299 8585
rect 103514 8576 103520 8628
rect 103572 8616 103578 8628
rect 105909 8619 105967 8625
rect 105909 8616 105921 8619
rect 103572 8588 105921 8616
rect 103572 8576 103578 8588
rect 105909 8585 105921 8588
rect 105955 8585 105967 8619
rect 105909 8579 105967 8585
rect 108850 8576 108856 8628
rect 108908 8616 108914 8628
rect 136358 8616 136364 8628
rect 108908 8588 129228 8616
rect 108908 8576 108914 8588
rect 100389 8551 100447 8557
rect 100389 8517 100401 8551
rect 100435 8517 100447 8551
rect 100389 8511 100447 8517
rect 104805 8551 104863 8557
rect 104805 8517 104817 8551
rect 104851 8548 104863 8551
rect 105262 8548 105268 8560
rect 104851 8520 105268 8548
rect 104851 8517 104863 8520
rect 104805 8511 104863 8517
rect 105262 8508 105268 8520
rect 105320 8508 105326 8560
rect 109126 8508 109132 8560
rect 109184 8548 109190 8560
rect 116121 8551 116179 8557
rect 109184 8520 112024 8548
rect 109184 8508 109190 8520
rect 95053 8483 95111 8489
rect 95053 8449 95065 8483
rect 95099 8449 95111 8483
rect 97258 8480 97264 8492
rect 95053 8443 95111 8449
rect 95436 8452 97264 8480
rect 89257 8415 89315 8421
rect 89257 8381 89269 8415
rect 89303 8381 89315 8415
rect 89257 8375 89315 8381
rect 91097 8415 91155 8421
rect 91097 8381 91109 8415
rect 91143 8412 91155 8415
rect 92293 8415 92351 8421
rect 92293 8412 92305 8415
rect 91143 8384 92305 8412
rect 91143 8381 91155 8384
rect 91097 8375 91155 8381
rect 92293 8381 92305 8384
rect 92339 8381 92351 8415
rect 93762 8412 93768 8424
rect 93723 8384 93768 8412
rect 92293 8375 92351 8381
rect 93762 8372 93768 8384
rect 93820 8372 93826 8424
rect 95436 8421 95464 8452
rect 97258 8440 97264 8452
rect 97316 8440 97322 8492
rect 102042 8440 102048 8492
rect 102100 8480 102106 8492
rect 103333 8483 103391 8489
rect 103333 8480 103345 8483
rect 102100 8452 103345 8480
rect 102100 8440 102106 8452
rect 103333 8449 103345 8452
rect 103379 8449 103391 8483
rect 108758 8480 108764 8492
rect 103333 8443 103391 8449
rect 106476 8452 108764 8480
rect 94961 8415 95019 8421
rect 94961 8381 94973 8415
rect 95007 8381 95019 8415
rect 94961 8375 95019 8381
rect 95421 8415 95479 8421
rect 95421 8381 95433 8415
rect 95467 8381 95479 8415
rect 96614 8412 96620 8424
rect 96575 8384 96620 8412
rect 95421 8375 95479 8381
rect 90818 8344 90824 8356
rect 86144 8316 90824 8344
rect 90818 8304 90824 8316
rect 90876 8304 90882 8356
rect 94976 8344 95004 8375
rect 96614 8372 96620 8384
rect 96672 8372 96678 8424
rect 96985 8415 97043 8421
rect 96985 8381 96997 8415
rect 97031 8412 97043 8415
rect 97074 8412 97080 8424
rect 97031 8384 97080 8412
rect 97031 8381 97043 8384
rect 96985 8375 97043 8381
rect 97074 8372 97080 8384
rect 97132 8372 97138 8424
rect 97353 8415 97411 8421
rect 97353 8381 97365 8415
rect 97399 8412 97411 8415
rect 97534 8412 97540 8424
rect 97399 8384 97540 8412
rect 97399 8381 97411 8384
rect 97353 8375 97411 8381
rect 97534 8372 97540 8384
rect 97592 8372 97598 8424
rect 99098 8412 99104 8424
rect 99059 8384 99104 8412
rect 99098 8372 99104 8384
rect 99156 8372 99162 8424
rect 100665 8415 100723 8421
rect 100665 8381 100677 8415
rect 100711 8412 100723 8415
rect 104526 8412 104532 8424
rect 100711 8384 104532 8412
rect 100711 8381 100723 8384
rect 100665 8375 100723 8381
rect 104526 8372 104532 8384
rect 104584 8372 104590 8424
rect 104805 8415 104863 8421
rect 104805 8381 104817 8415
rect 104851 8412 104863 8415
rect 105722 8412 105728 8424
rect 104851 8384 105728 8412
rect 104851 8381 104863 8384
rect 104805 8375 104863 8381
rect 105722 8372 105728 8384
rect 105780 8372 105786 8424
rect 106090 8412 106096 8424
rect 106051 8384 106096 8412
rect 106090 8372 106096 8384
rect 106148 8372 106154 8424
rect 97994 8344 98000 8356
rect 94976 8316 98000 8344
rect 97994 8304 98000 8316
rect 98052 8304 98058 8356
rect 99466 8344 99472 8356
rect 99208 8316 99472 8344
rect 78324 8248 78720 8276
rect 80974 8236 80980 8288
rect 81032 8276 81038 8288
rect 84654 8276 84660 8288
rect 81032 8248 84660 8276
rect 81032 8236 81038 8248
rect 84654 8236 84660 8248
rect 84712 8236 84718 8288
rect 85666 8236 85672 8288
rect 85724 8276 85730 8288
rect 90266 8276 90272 8288
rect 85724 8248 90272 8276
rect 85724 8236 85730 8248
rect 90266 8236 90272 8248
rect 90324 8236 90330 8288
rect 91370 8236 91376 8288
rect 91428 8276 91434 8288
rect 99208 8276 99236 8316
rect 99466 8304 99472 8316
rect 99524 8304 99530 8356
rect 103241 8347 103299 8353
rect 102060 8316 102364 8344
rect 91428 8248 99236 8276
rect 91428 8236 91434 8248
rect 99282 8236 99288 8288
rect 99340 8276 99346 8288
rect 102060 8276 102088 8316
rect 102226 8276 102232 8288
rect 99340 8248 102088 8276
rect 102187 8248 102232 8276
rect 99340 8236 99346 8248
rect 102226 8236 102232 8248
rect 102284 8236 102290 8288
rect 102336 8276 102364 8316
rect 103241 8313 103253 8347
rect 103287 8344 103299 8347
rect 106476 8344 106504 8452
rect 108758 8440 108764 8452
rect 108816 8440 108822 8492
rect 109032 8483 109090 8489
rect 109032 8449 109044 8483
rect 109078 8480 109090 8483
rect 109218 8480 109224 8492
rect 109078 8452 109224 8480
rect 109078 8449 109090 8452
rect 109032 8443 109090 8449
rect 109218 8440 109224 8452
rect 109276 8440 109282 8492
rect 109954 8440 109960 8492
rect 110012 8480 110018 8492
rect 110049 8483 110107 8489
rect 110049 8480 110061 8483
rect 110012 8452 110061 8480
rect 110012 8440 110018 8452
rect 110049 8449 110061 8452
rect 110095 8449 110107 8483
rect 110049 8443 110107 8449
rect 106553 8415 106611 8421
rect 106553 8381 106565 8415
rect 106599 8412 106611 8415
rect 110138 8412 110144 8424
rect 106599 8384 109816 8412
rect 110099 8384 110144 8412
rect 106599 8381 106611 8384
rect 106553 8375 106611 8381
rect 103287 8316 106504 8344
rect 107841 8347 107899 8353
rect 103287 8313 103299 8316
rect 103241 8307 103299 8313
rect 107841 8313 107853 8347
rect 107887 8344 107899 8347
rect 109678 8344 109684 8356
rect 107887 8316 109684 8344
rect 107887 8313 107899 8316
rect 107841 8307 107899 8313
rect 109678 8304 109684 8316
rect 109736 8304 109742 8356
rect 109788 8344 109816 8384
rect 110138 8372 110144 8384
rect 110196 8372 110202 8424
rect 111702 8412 111708 8424
rect 111663 8384 111708 8412
rect 111702 8372 111708 8384
rect 111760 8372 111766 8424
rect 111797 8415 111855 8421
rect 111797 8381 111809 8415
rect 111843 8412 111855 8415
rect 111886 8412 111892 8424
rect 111843 8384 111892 8412
rect 111843 8381 111855 8384
rect 111797 8375 111855 8381
rect 111886 8372 111892 8384
rect 111944 8372 111950 8424
rect 111996 8421 112024 8520
rect 116121 8517 116133 8551
rect 116167 8548 116179 8551
rect 128998 8548 129004 8560
rect 116167 8520 129004 8548
rect 116167 8517 116179 8520
rect 116121 8511 116179 8517
rect 128998 8508 129004 8520
rect 129056 8508 129062 8560
rect 114646 8480 114652 8492
rect 114607 8452 114652 8480
rect 114646 8440 114652 8452
rect 114704 8440 114710 8492
rect 121086 8480 121092 8492
rect 116228 8452 121092 8480
rect 116228 8421 116256 8452
rect 121086 8440 121092 8452
rect 121144 8440 121150 8492
rect 121273 8483 121331 8489
rect 121273 8449 121285 8483
rect 121319 8480 121331 8483
rect 124582 8480 124588 8492
rect 121319 8452 124588 8480
rect 121319 8449 121331 8452
rect 121273 8443 121331 8449
rect 124582 8440 124588 8452
rect 124640 8440 124646 8492
rect 125134 8480 125140 8492
rect 125095 8452 125140 8480
rect 125134 8440 125140 8452
rect 125192 8440 125198 8492
rect 126606 8480 126612 8492
rect 126567 8452 126612 8480
rect 126606 8440 126612 8452
rect 126664 8440 126670 8492
rect 127802 8480 127808 8492
rect 127763 8452 127808 8480
rect 127802 8440 127808 8452
rect 127860 8440 127866 8492
rect 129200 8480 129228 8588
rect 129292 8588 136364 8616
rect 129292 8557 129320 8588
rect 136358 8576 136364 8588
rect 136416 8576 136422 8628
rect 138198 8576 138204 8628
rect 138256 8616 138262 8628
rect 144822 8616 144828 8628
rect 138256 8588 144828 8616
rect 138256 8576 138262 8588
rect 144822 8576 144828 8588
rect 144880 8576 144886 8628
rect 151078 8576 151084 8628
rect 151136 8616 151142 8628
rect 159818 8616 159824 8628
rect 151136 8588 159824 8616
rect 151136 8576 151142 8588
rect 159818 8576 159824 8588
rect 159876 8576 159882 8628
rect 159910 8576 159916 8628
rect 159968 8616 159974 8628
rect 164326 8616 164332 8628
rect 159968 8588 164332 8616
rect 159968 8576 159974 8588
rect 164326 8576 164332 8588
rect 164384 8576 164390 8628
rect 164418 8576 164424 8628
rect 164476 8616 164482 8628
rect 175734 8616 175740 8628
rect 164476 8588 175740 8616
rect 164476 8576 164482 8588
rect 175734 8576 175740 8588
rect 175792 8576 175798 8628
rect 176194 8576 176200 8628
rect 176252 8616 176258 8628
rect 178954 8616 178960 8628
rect 176252 8588 178960 8616
rect 176252 8576 176258 8588
rect 178954 8576 178960 8588
rect 179012 8576 179018 8628
rect 184658 8616 184664 8628
rect 179064 8588 184664 8616
rect 129277 8551 129335 8557
rect 129277 8517 129289 8551
rect 129323 8517 129335 8551
rect 131298 8548 131304 8560
rect 129277 8511 129335 8517
rect 129384 8520 131304 8548
rect 129384 8480 129412 8520
rect 131298 8508 131304 8520
rect 131356 8508 131362 8560
rect 135714 8548 135720 8560
rect 133432 8520 135720 8548
rect 129200 8452 129412 8480
rect 131025 8483 131083 8489
rect 131025 8449 131037 8483
rect 131071 8480 131083 8483
rect 132218 8480 132224 8492
rect 131071 8452 132224 8480
rect 131071 8449 131083 8452
rect 131025 8443 131083 8449
rect 132218 8440 132224 8452
rect 132276 8440 132282 8492
rect 132402 8480 132408 8492
rect 132363 8452 132408 8480
rect 132402 8440 132408 8452
rect 132460 8440 132466 8492
rect 133432 8489 133460 8520
rect 135714 8508 135720 8520
rect 135772 8508 135778 8560
rect 142154 8548 142160 8560
rect 136560 8520 138888 8548
rect 133417 8483 133475 8489
rect 133417 8449 133429 8483
rect 133463 8449 133475 8483
rect 133417 8443 133475 8449
rect 134889 8483 134947 8489
rect 134889 8449 134901 8483
rect 134935 8480 134947 8483
rect 135162 8480 135168 8492
rect 134935 8452 135168 8480
rect 134935 8449 134947 8452
rect 134889 8443 134947 8449
rect 135162 8440 135168 8452
rect 135220 8440 135226 8492
rect 135530 8440 135536 8492
rect 135588 8480 135594 8492
rect 136082 8480 136088 8492
rect 135588 8452 136088 8480
rect 135588 8440 135594 8452
rect 136082 8440 136088 8452
rect 136140 8440 136146 8492
rect 136560 8489 136588 8520
rect 136545 8483 136603 8489
rect 136545 8449 136557 8483
rect 136591 8449 136603 8483
rect 137922 8480 137928 8492
rect 137883 8452 137928 8480
rect 136545 8443 136603 8449
rect 137922 8440 137928 8452
rect 137980 8440 137986 8492
rect 111981 8415 112039 8421
rect 111981 8381 111993 8415
rect 112027 8381 112039 8415
rect 111981 8375 112039 8381
rect 116213 8415 116271 8421
rect 116213 8381 116225 8415
rect 116259 8381 116271 8415
rect 116213 8375 116271 8381
rect 119065 8415 119123 8421
rect 119065 8381 119077 8415
rect 119111 8412 119123 8415
rect 121454 8412 121460 8424
rect 119111 8384 121460 8412
rect 119111 8381 119123 8384
rect 119065 8375 119123 8381
rect 121454 8372 121460 8384
rect 121512 8372 121518 8424
rect 126698 8412 126704 8424
rect 126659 8384 126704 8412
rect 126698 8372 126704 8384
rect 126756 8372 126762 8424
rect 129369 8415 129427 8421
rect 129369 8381 129381 8415
rect 129415 8412 129427 8415
rect 129642 8412 129648 8424
rect 129415 8384 129648 8412
rect 129415 8381 129427 8384
rect 129369 8375 129427 8381
rect 129642 8372 129648 8384
rect 129700 8372 129706 8424
rect 132126 8412 132132 8424
rect 132087 8384 132132 8412
rect 132126 8372 132132 8384
rect 132184 8372 132190 8424
rect 132954 8372 132960 8424
rect 133012 8412 133018 8424
rect 134521 8415 134579 8421
rect 134521 8412 134533 8415
rect 133012 8384 134533 8412
rect 133012 8372 133018 8384
rect 134521 8381 134533 8384
rect 134567 8381 134579 8415
rect 134521 8375 134579 8381
rect 135990 8372 135996 8424
rect 136048 8412 136054 8424
rect 137649 8415 137707 8421
rect 137649 8412 137661 8415
rect 136048 8384 137661 8412
rect 136048 8372 136054 8384
rect 137649 8381 137661 8384
rect 137695 8381 137707 8415
rect 138860 8412 138888 8520
rect 138952 8520 142160 8548
rect 138952 8489 138980 8520
rect 142154 8508 142160 8520
rect 142212 8508 142218 8560
rect 146110 8548 146116 8560
rect 146071 8520 146116 8548
rect 146110 8508 146116 8520
rect 146168 8508 146174 8560
rect 155313 8551 155371 8557
rect 155313 8517 155325 8551
rect 155359 8548 155371 8551
rect 159542 8548 159548 8560
rect 155359 8520 159548 8548
rect 155359 8517 155371 8520
rect 155313 8511 155371 8517
rect 159542 8508 159548 8520
rect 159600 8508 159606 8560
rect 159637 8551 159695 8557
rect 159637 8517 159649 8551
rect 159683 8548 159695 8551
rect 162949 8551 163007 8557
rect 159683 8520 162900 8548
rect 159683 8517 159695 8520
rect 159637 8511 159695 8517
rect 138937 8483 138995 8489
rect 138937 8449 138949 8483
rect 138983 8449 138995 8483
rect 140406 8480 140412 8492
rect 138937 8443 138995 8449
rect 139044 8452 140176 8480
rect 140367 8452 140412 8480
rect 139044 8412 139072 8452
rect 138860 8384 139072 8412
rect 137649 8375 137707 8381
rect 139118 8372 139124 8424
rect 139176 8412 139182 8424
rect 140041 8415 140099 8421
rect 140041 8412 140053 8415
rect 139176 8384 140053 8412
rect 139176 8372 139182 8384
rect 140041 8381 140053 8384
rect 140087 8381 140099 8415
rect 140148 8412 140176 8452
rect 140406 8440 140412 8452
rect 140464 8440 140470 8492
rect 140774 8440 140780 8492
rect 140832 8480 140838 8492
rect 143537 8483 143595 8489
rect 143537 8480 143549 8483
rect 140832 8452 143549 8480
rect 140832 8440 140838 8452
rect 143537 8449 143549 8452
rect 143583 8449 143595 8483
rect 143537 8443 143595 8449
rect 144641 8483 144699 8489
rect 144641 8449 144653 8483
rect 144687 8480 144699 8483
rect 144914 8480 144920 8492
rect 144687 8452 144920 8480
rect 144687 8449 144699 8452
rect 144641 8443 144699 8449
rect 144914 8440 144920 8452
rect 144972 8440 144978 8492
rect 147217 8483 147275 8489
rect 147217 8449 147229 8483
rect 147263 8480 147275 8483
rect 148410 8480 148416 8492
rect 147263 8452 148416 8480
rect 147263 8449 147275 8452
rect 147217 8443 147275 8449
rect 148410 8440 148416 8452
rect 148468 8440 148474 8492
rect 148686 8480 148692 8492
rect 148647 8452 148692 8480
rect 148686 8440 148692 8452
rect 148744 8440 148750 8492
rect 149609 8483 149667 8489
rect 149609 8449 149621 8483
rect 149655 8480 149667 8483
rect 149698 8480 149704 8492
rect 149655 8452 149704 8480
rect 149655 8449 149667 8452
rect 149609 8443 149667 8449
rect 149698 8440 149704 8452
rect 149756 8440 149762 8492
rect 150621 8483 150679 8489
rect 150621 8449 150633 8483
rect 150667 8480 150679 8483
rect 150710 8480 150716 8492
rect 150667 8452 150716 8480
rect 150667 8449 150679 8452
rect 150621 8443 150679 8449
rect 150710 8440 150716 8452
rect 150768 8440 150774 8492
rect 151630 8480 151636 8492
rect 151591 8452 151636 8480
rect 151630 8440 151636 8452
rect 151688 8440 151694 8492
rect 152826 8480 152832 8492
rect 152787 8452 152832 8480
rect 152826 8440 152832 8452
rect 152884 8440 152890 8492
rect 156230 8480 156236 8492
rect 156191 8452 156236 8480
rect 156230 8440 156236 8452
rect 156288 8440 156294 8492
rect 159910 8480 159916 8492
rect 156340 8452 159916 8480
rect 142525 8415 142583 8421
rect 142525 8412 142537 8415
rect 140148 8384 142537 8412
rect 140041 8375 140099 8381
rect 142525 8381 142537 8384
rect 142571 8381 142583 8415
rect 146202 8412 146208 8424
rect 146163 8384 146208 8412
rect 142525 8375 142583 8381
rect 146202 8372 146208 8384
rect 146260 8372 146266 8424
rect 148321 8415 148379 8421
rect 148321 8381 148333 8415
rect 148367 8381 148379 8415
rect 153838 8412 153844 8424
rect 153799 8384 153844 8412
rect 148321 8375 148379 8381
rect 112162 8344 112168 8356
rect 109788 8316 112168 8344
rect 112162 8304 112168 8316
rect 112220 8304 112226 8356
rect 117409 8347 117467 8353
rect 117409 8313 117421 8347
rect 117455 8344 117467 8347
rect 118694 8344 118700 8356
rect 117455 8316 118700 8344
rect 117455 8313 117467 8316
rect 117409 8307 117467 8313
rect 118694 8304 118700 8316
rect 118752 8304 118758 8356
rect 120258 8344 120264 8356
rect 120219 8316 120264 8344
rect 120258 8304 120264 8316
rect 120316 8304 120322 8356
rect 122285 8347 122343 8353
rect 122285 8313 122297 8347
rect 122331 8344 122343 8347
rect 123294 8344 123300 8356
rect 122331 8316 123300 8344
rect 122331 8313 122343 8316
rect 122285 8307 122343 8313
rect 123294 8304 123300 8316
rect 123352 8304 123358 8356
rect 123573 8347 123631 8353
rect 123573 8313 123585 8347
rect 123619 8344 123631 8347
rect 126146 8344 126152 8356
rect 123619 8316 126152 8344
rect 123619 8313 123631 8316
rect 123573 8307 123631 8313
rect 126146 8304 126152 8316
rect 126204 8304 126210 8356
rect 127894 8304 127900 8356
rect 127952 8344 127958 8356
rect 130838 8344 130844 8356
rect 127952 8316 130844 8344
rect 127952 8304 127958 8316
rect 130838 8304 130844 8316
rect 130896 8304 130902 8356
rect 140700 8316 141648 8344
rect 112806 8276 112812 8288
rect 102336 8248 112812 8276
rect 112806 8236 112812 8248
rect 112864 8236 112870 8288
rect 113450 8276 113456 8288
rect 113411 8248 113456 8276
rect 113450 8236 113456 8248
rect 113508 8236 113514 8288
rect 119982 8236 119988 8288
rect 120040 8276 120046 8288
rect 133782 8276 133788 8288
rect 120040 8248 133788 8276
rect 120040 8236 120046 8248
rect 133782 8236 133788 8248
rect 133840 8236 133846 8288
rect 133874 8236 133880 8288
rect 133932 8276 133938 8288
rect 140700 8276 140728 8316
rect 133932 8248 140728 8276
rect 133932 8236 133938 8248
rect 140774 8236 140780 8288
rect 140832 8276 140838 8288
rect 141513 8279 141571 8285
rect 141513 8276 141525 8279
rect 140832 8248 141525 8276
rect 140832 8236 140838 8248
rect 141513 8245 141525 8248
rect 141559 8245 141571 8279
rect 141620 8276 141648 8316
rect 142448 8316 142660 8344
rect 142448 8276 142476 8316
rect 141620 8248 142476 8276
rect 142632 8276 142660 8316
rect 143460 8316 143672 8344
rect 143460 8276 143488 8316
rect 142632 8248 143488 8276
rect 143644 8276 143672 8316
rect 145558 8304 145564 8356
rect 145616 8344 145622 8356
rect 148336 8344 148364 8375
rect 153838 8372 153844 8384
rect 153896 8372 153902 8424
rect 155402 8412 155408 8424
rect 155363 8384 155408 8412
rect 155402 8372 155408 8384
rect 155460 8372 155466 8424
rect 156138 8372 156144 8424
rect 156196 8412 156202 8424
rect 156340 8412 156368 8452
rect 159910 8440 159916 8452
rect 159968 8440 159974 8492
rect 160002 8440 160008 8492
rect 160060 8480 160066 8492
rect 161477 8483 161535 8489
rect 161477 8480 161489 8483
rect 160060 8452 161489 8480
rect 160060 8440 160066 8452
rect 161477 8449 161489 8452
rect 161523 8449 161535 8483
rect 162872 8480 162900 8520
rect 162949 8517 162961 8551
rect 162995 8548 163007 8551
rect 170030 8548 170036 8560
rect 162995 8520 170036 8548
rect 162995 8517 163007 8520
rect 162949 8511 163007 8517
rect 170030 8508 170036 8520
rect 170088 8508 170094 8560
rect 171502 8548 171508 8560
rect 170600 8520 171508 8548
rect 165338 8480 165344 8492
rect 162872 8452 165344 8480
rect 161477 8443 161535 8449
rect 165338 8440 165344 8452
rect 165396 8440 165402 8492
rect 166810 8440 166816 8492
rect 166868 8480 166874 8492
rect 167273 8483 167331 8489
rect 166868 8452 167132 8480
rect 166868 8440 166874 8452
rect 156196 8384 156368 8412
rect 157245 8415 157303 8421
rect 156196 8372 156202 8384
rect 157245 8381 157257 8415
rect 157291 8412 157303 8415
rect 158349 8415 158407 8421
rect 158349 8412 158361 8415
rect 157291 8384 158361 8412
rect 157291 8381 157303 8384
rect 157245 8375 157303 8381
rect 158349 8381 158361 8384
rect 158395 8381 158407 8415
rect 158349 8375 158407 8381
rect 159453 8415 159511 8421
rect 159453 8381 159465 8415
rect 159499 8381 159511 8415
rect 162578 8412 162584 8424
rect 162539 8384 162584 8412
rect 159453 8375 159511 8381
rect 145616 8316 148364 8344
rect 149532 8316 149744 8344
rect 145616 8304 145622 8316
rect 149532 8276 149560 8316
rect 143644 8248 149560 8276
rect 149716 8276 149744 8316
rect 150544 8316 150756 8344
rect 150544 8276 150572 8316
rect 149716 8248 150572 8276
rect 150728 8276 150756 8316
rect 151556 8316 151768 8344
rect 151556 8276 151584 8316
rect 150728 8248 151584 8276
rect 151740 8276 151768 8316
rect 154022 8304 154028 8356
rect 154080 8344 154086 8356
rect 159468 8344 159496 8375
rect 162578 8372 162584 8384
rect 162636 8372 162642 8424
rect 164234 8372 164240 8424
rect 164292 8412 164298 8424
rect 165801 8415 165859 8421
rect 165801 8412 165813 8415
rect 164292 8384 165813 8412
rect 164292 8372 164298 8384
rect 165801 8381 165813 8384
rect 165847 8381 165859 8415
rect 167104 8412 167132 8452
rect 167273 8449 167285 8483
rect 167319 8449 167331 8483
rect 168466 8480 168472 8492
rect 168427 8452 168472 8480
rect 167273 8443 167331 8449
rect 167178 8412 167184 8424
rect 167104 8384 167184 8412
rect 165801 8375 165859 8381
rect 167178 8372 167184 8384
rect 167236 8372 167242 8424
rect 154080 8316 159496 8344
rect 154080 8304 154086 8316
rect 159542 8304 159548 8356
rect 159600 8344 159606 8356
rect 166534 8344 166540 8356
rect 159600 8316 166540 8344
rect 159600 8304 159606 8316
rect 166534 8304 166540 8316
rect 166592 8304 166598 8356
rect 167288 8344 167316 8443
rect 168466 8440 168472 8452
rect 168524 8440 168530 8492
rect 169665 8483 169723 8489
rect 169665 8449 169677 8483
rect 169711 8480 169723 8483
rect 170600 8480 170628 8520
rect 171502 8508 171508 8520
rect 171560 8508 171566 8560
rect 172149 8551 172207 8557
rect 172149 8517 172161 8551
rect 172195 8548 172207 8551
rect 176749 8551 176807 8557
rect 172195 8520 176700 8548
rect 172195 8517 172207 8520
rect 172149 8511 172207 8517
rect 169711 8452 170628 8480
rect 170677 8483 170735 8489
rect 169711 8449 169723 8452
rect 169665 8443 169723 8449
rect 170677 8449 170689 8483
rect 170723 8480 170735 8483
rect 174081 8483 174139 8489
rect 174081 8480 174093 8483
rect 170723 8452 174093 8480
rect 170723 8449 170735 8452
rect 170677 8443 170735 8449
rect 174081 8449 174093 8452
rect 174127 8449 174139 8483
rect 176672 8480 176700 8520
rect 176749 8517 176761 8551
rect 176795 8548 176807 8551
rect 176838 8548 176844 8560
rect 176795 8520 176844 8548
rect 176795 8517 176807 8520
rect 176749 8511 176807 8517
rect 176838 8508 176844 8520
rect 176896 8508 176902 8560
rect 176672 8452 177804 8480
rect 174081 8443 174139 8449
rect 167365 8415 167423 8421
rect 167365 8381 167377 8415
rect 167411 8412 167423 8415
rect 170766 8412 170772 8424
rect 167411 8384 170772 8412
rect 167411 8381 167423 8384
rect 167365 8375 167423 8381
rect 170766 8372 170772 8384
rect 170824 8372 170830 8424
rect 171778 8412 171784 8424
rect 171739 8384 171784 8412
rect 171778 8372 171784 8384
rect 171836 8372 171842 8424
rect 173069 8415 173127 8421
rect 173069 8381 173081 8415
rect 173115 8412 173127 8415
rect 175277 8415 175335 8421
rect 175277 8412 175289 8415
rect 173115 8384 175289 8412
rect 173115 8381 173127 8384
rect 173069 8375 173127 8381
rect 175277 8381 175289 8384
rect 175323 8381 175335 8415
rect 176378 8412 176384 8424
rect 176339 8384 176384 8412
rect 175277 8375 175335 8381
rect 176378 8372 176384 8384
rect 176436 8372 176442 8424
rect 176562 8372 176568 8424
rect 176620 8412 176626 8424
rect 177669 8415 177727 8421
rect 177669 8412 177681 8415
rect 176620 8384 177681 8412
rect 176620 8372 176626 8384
rect 177669 8381 177681 8384
rect 177715 8381 177727 8415
rect 177669 8375 177727 8381
rect 171042 8344 171048 8356
rect 167288 8316 171048 8344
rect 171042 8304 171048 8316
rect 171100 8304 171106 8356
rect 176470 8344 176476 8356
rect 173820 8316 176476 8344
rect 159634 8276 159640 8288
rect 151740 8248 159640 8276
rect 141513 8239 141571 8245
rect 159634 8236 159640 8248
rect 159692 8236 159698 8288
rect 160646 8236 160652 8288
rect 160704 8276 160710 8288
rect 163958 8276 163964 8288
rect 160704 8248 163964 8276
rect 160704 8236 160710 8248
rect 163958 8236 163964 8248
rect 164016 8236 164022 8288
rect 164510 8276 164516 8288
rect 164471 8248 164516 8276
rect 164510 8236 164516 8248
rect 164568 8236 164574 8288
rect 164602 8236 164608 8288
rect 164660 8276 164666 8288
rect 167086 8276 167092 8288
rect 164660 8248 167092 8276
rect 164660 8236 164666 8248
rect 167086 8236 167092 8248
rect 167144 8236 167150 8288
rect 171134 8236 171140 8288
rect 171192 8276 171198 8288
rect 173820 8276 173848 8316
rect 176470 8304 176476 8316
rect 176528 8304 176534 8356
rect 177776 8344 177804 8452
rect 179064 8421 179092 8588
rect 184658 8576 184664 8588
rect 184716 8576 184722 8628
rect 185412 8588 189120 8616
rect 179141 8551 179199 8557
rect 179141 8517 179153 8551
rect 179187 8548 179199 8551
rect 184934 8548 184940 8560
rect 179187 8520 184940 8548
rect 179187 8517 179199 8520
rect 179141 8511 179199 8517
rect 184934 8508 184940 8520
rect 184992 8508 184998 8560
rect 185412 8557 185440 8588
rect 185397 8551 185455 8557
rect 185397 8517 185409 8551
rect 185443 8517 185455 8551
rect 187878 8548 187884 8560
rect 187839 8520 187884 8548
rect 185397 8511 185455 8517
rect 187878 8508 187884 8520
rect 187936 8508 187942 8560
rect 182821 8483 182879 8489
rect 182821 8449 182833 8483
rect 182867 8449 182879 8483
rect 183830 8480 183836 8492
rect 182821 8443 182879 8449
rect 182928 8452 183836 8480
rect 179049 8415 179107 8421
rect 179049 8381 179061 8415
rect 179095 8381 179107 8415
rect 181438 8412 181444 8424
rect 181399 8384 181444 8412
rect 179049 8375 179107 8381
rect 181438 8372 181444 8384
rect 181496 8372 181502 8424
rect 180978 8344 180984 8356
rect 177776 8316 180984 8344
rect 180978 8304 180984 8316
rect 181036 8304 181042 8356
rect 182836 8344 182864 8443
rect 182928 8421 182956 8452
rect 183830 8440 183836 8452
rect 183888 8440 183894 8492
rect 183922 8440 183928 8492
rect 183980 8480 183986 8492
rect 183980 8452 184025 8480
rect 183980 8440 183986 8452
rect 184106 8440 184112 8492
rect 184164 8480 184170 8492
rect 184750 8480 184756 8492
rect 184164 8452 184756 8480
rect 184164 8440 184170 8452
rect 184750 8440 184756 8452
rect 184808 8440 184814 8492
rect 186409 8483 186467 8489
rect 186409 8480 186421 8483
rect 184860 8452 186421 8480
rect 182913 8415 182971 8421
rect 182913 8381 182925 8415
rect 182959 8381 182971 8415
rect 182913 8375 182971 8381
rect 183002 8372 183008 8424
rect 183060 8412 183066 8424
rect 184860 8412 184888 8452
rect 186409 8449 186421 8452
rect 186455 8449 186467 8483
rect 188430 8480 188436 8492
rect 186409 8443 186467 8449
rect 187436 8452 188436 8480
rect 185486 8412 185492 8424
rect 183060 8384 184888 8412
rect 185447 8384 185492 8412
rect 183060 8372 183066 8384
rect 185486 8372 185492 8384
rect 185544 8372 185550 8424
rect 187436 8344 187464 8452
rect 188430 8440 188436 8452
rect 188488 8440 188494 8492
rect 187973 8415 188031 8421
rect 187973 8381 187985 8415
rect 188019 8381 188031 8415
rect 187973 8375 188031 8381
rect 182836 8316 187464 8344
rect 187988 8344 188016 8375
rect 188062 8372 188068 8424
rect 188120 8412 188126 8424
rect 188801 8415 188859 8421
rect 188801 8412 188813 8415
rect 188120 8384 188813 8412
rect 188120 8372 188126 8384
rect 188801 8381 188813 8384
rect 188847 8381 188859 8415
rect 188801 8375 188859 8381
rect 188890 8344 188896 8356
rect 187988 8316 188896 8344
rect 188890 8304 188896 8316
rect 188948 8304 188954 8356
rect 189092 8344 189120 8588
rect 191190 8576 191196 8628
rect 191248 8616 191254 8628
rect 192113 8619 192171 8625
rect 192113 8616 192125 8619
rect 191248 8588 192125 8616
rect 191248 8576 191254 8588
rect 192113 8585 192125 8588
rect 192159 8585 192171 8619
rect 192113 8579 192171 8585
rect 194226 8576 194232 8628
rect 194284 8616 194290 8628
rect 196069 8619 196127 8625
rect 196069 8616 196081 8619
rect 194284 8588 196081 8616
rect 194284 8576 194290 8588
rect 196069 8585 196081 8588
rect 196115 8585 196127 8619
rect 196069 8579 196127 8585
rect 190273 8551 190331 8557
rect 190273 8517 190285 8551
rect 190319 8548 190331 8551
rect 191006 8548 191012 8560
rect 190319 8520 191012 8548
rect 190319 8517 190331 8520
rect 190273 8511 190331 8517
rect 191006 8508 191012 8520
rect 191064 8508 191070 8560
rect 196250 8548 196256 8560
rect 192036 8520 196256 8548
rect 190365 8415 190423 8421
rect 190365 8381 190377 8415
rect 190411 8412 190423 8415
rect 190638 8412 190644 8424
rect 190411 8384 190644 8412
rect 190411 8381 190423 8384
rect 190365 8375 190423 8381
rect 190638 8372 190644 8384
rect 190696 8372 190702 8424
rect 192036 8421 192064 8520
rect 196250 8508 196256 8520
rect 196308 8508 196314 8560
rect 192110 8440 192116 8492
rect 192168 8480 192174 8492
rect 193585 8483 193643 8489
rect 193585 8480 193597 8483
rect 192168 8452 193597 8480
rect 192168 8440 192174 8452
rect 193585 8449 193597 8452
rect 193631 8449 193643 8483
rect 194962 8480 194968 8492
rect 194923 8452 194968 8480
rect 193585 8443 193643 8449
rect 194962 8440 194968 8452
rect 195020 8440 195026 8492
rect 197538 8480 197544 8492
rect 195072 8452 197544 8480
rect 192021 8415 192079 8421
rect 192021 8381 192033 8415
rect 192067 8381 192079 8415
rect 192021 8375 192079 8381
rect 193858 8372 193864 8424
rect 193916 8412 193922 8424
rect 194689 8415 194747 8421
rect 194689 8412 194701 8415
rect 193916 8384 194701 8412
rect 193916 8372 193922 8384
rect 194689 8381 194701 8384
rect 194735 8381 194747 8415
rect 194689 8375 194747 8381
rect 195072 8344 195100 8452
rect 197538 8440 197544 8452
rect 197596 8440 197602 8492
rect 195977 8415 196035 8421
rect 195977 8381 195989 8415
rect 196023 8381 196035 8415
rect 195977 8375 196035 8381
rect 195992 8344 196020 8375
rect 189092 8316 195100 8344
rect 195164 8316 196020 8344
rect 171192 8248 173848 8276
rect 171192 8236 171198 8248
rect 173894 8236 173900 8288
rect 173952 8276 173958 8288
rect 177482 8276 177488 8288
rect 173952 8248 177488 8276
rect 173952 8236 173958 8248
rect 177482 8236 177488 8248
rect 177540 8236 177546 8288
rect 179506 8236 179512 8288
rect 179564 8276 179570 8288
rect 190546 8276 190552 8288
rect 179564 8248 190552 8276
rect 179564 8236 179570 8248
rect 190546 8236 190552 8248
rect 190604 8236 190610 8288
rect 194502 8236 194508 8288
rect 194560 8276 194566 8288
rect 195164 8276 195192 8316
rect 194560 8248 195192 8276
rect 194560 8236 194566 8248
rect 1104 8186 198812 8208
rect 1104 8134 24078 8186
rect 24130 8134 64078 8186
rect 64130 8134 104078 8186
rect 104130 8134 144078 8186
rect 144130 8134 184078 8186
rect 184130 8134 198812 8186
rect 1104 8112 198812 8134
rect 7374 8072 7380 8084
rect 7335 8044 7380 8072
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 23845 8075 23903 8081
rect 23845 8041 23857 8075
rect 23891 8072 23903 8075
rect 24946 8072 24952 8084
rect 23891 8044 24952 8072
rect 23891 8041 23903 8044
rect 23845 8035 23903 8041
rect 24946 8032 24952 8044
rect 25004 8032 25010 8084
rect 37550 8032 37556 8084
rect 37608 8072 37614 8084
rect 37737 8075 37795 8081
rect 37737 8072 37749 8075
rect 37608 8044 37749 8072
rect 37608 8032 37614 8044
rect 37737 8041 37749 8044
rect 37783 8041 37795 8075
rect 37737 8035 37795 8041
rect 41966 8032 41972 8084
rect 42024 8072 42030 8084
rect 42245 8075 42303 8081
rect 42245 8072 42257 8075
rect 42024 8044 42257 8072
rect 42024 8032 42030 8044
rect 42245 8041 42257 8044
rect 42291 8041 42303 8075
rect 42245 8035 42303 8041
rect 54662 8032 54668 8084
rect 54720 8072 54726 8084
rect 54849 8075 54907 8081
rect 54849 8072 54861 8075
rect 54720 8044 54861 8072
rect 54720 8032 54726 8044
rect 54849 8041 54861 8044
rect 54895 8041 54907 8075
rect 55858 8072 55864 8084
rect 55819 8044 55864 8072
rect 54849 8035 54907 8041
rect 55858 8032 55864 8044
rect 55916 8032 55922 8084
rect 75270 8032 75276 8084
rect 75328 8072 75334 8084
rect 81250 8072 81256 8084
rect 75328 8044 81256 8072
rect 75328 8032 75334 8044
rect 81250 8032 81256 8044
rect 81308 8032 81314 8084
rect 83090 8032 83096 8084
rect 83148 8072 83154 8084
rect 91646 8072 91652 8084
rect 83148 8044 86540 8072
rect 83148 8032 83154 8044
rect 29546 7964 29552 8016
rect 29604 8004 29610 8016
rect 29604 7976 32260 8004
rect 29604 7964 29610 7976
rect 6086 7936 6092 7948
rect 6047 7908 6092 7936
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7936 10747 7939
rect 11514 7936 11520 7948
rect 10735 7908 11520 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 11790 7936 11796 7948
rect 11751 7908 11796 7936
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 16850 7896 16856 7948
rect 16908 7936 16914 7948
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 16908 7908 18061 7936
rect 16908 7896 16914 7908
rect 18049 7905 18061 7908
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 26881 7939 26939 7945
rect 26881 7905 26893 7939
rect 26927 7936 26939 7939
rect 27338 7936 27344 7948
rect 26927 7908 27344 7936
rect 26927 7905 26939 7908
rect 26881 7899 26939 7905
rect 27338 7896 27344 7908
rect 27396 7896 27402 7948
rect 27985 7939 28043 7945
rect 27985 7905 27997 7939
rect 28031 7905 28043 7939
rect 32122 7936 32128 7948
rect 32083 7908 32128 7936
rect 27985 7899 28043 7905
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 4338 7868 4344 7880
rect 3007 7840 4344 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 3326 7760 3332 7812
rect 3384 7800 3390 7812
rect 5000 7800 5028 7831
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5408 7840 6009 7868
rect 5408 7828 5414 7840
rect 5997 7837 6009 7840
rect 6043 7837 6055 7871
rect 5997 7831 6055 7837
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 7524 7840 8401 7868
rect 7524 7828 7530 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 9674 7868 9680 7880
rect 9635 7840 9680 7868
rect 8389 7831 8447 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7837 11759 7871
rect 11701 7831 11759 7837
rect 3384 7772 5028 7800
rect 3384 7760 3390 7772
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 11716 7800 11744 7831
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 12492 7840 13093 7868
rect 12492 7828 12498 7840
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 14185 7871 14243 7877
rect 14185 7837 14197 7871
rect 14231 7868 14243 7871
rect 14826 7868 14832 7880
rect 14231 7840 14832 7868
rect 14231 7837 14243 7840
rect 14185 7831 14243 7837
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 15562 7868 15568 7880
rect 15523 7840 15568 7868
rect 15562 7828 15568 7840
rect 15620 7828 15626 7880
rect 16942 7868 16948 7880
rect 16903 7840 16948 7868
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7868 19487 7871
rect 20438 7868 20444 7880
rect 19475 7840 20444 7868
rect 19475 7837 19487 7840
rect 19429 7831 19487 7837
rect 7340 7772 11744 7800
rect 7340 7760 7346 7772
rect 15838 7760 15844 7812
rect 15896 7800 15902 7812
rect 17972 7800 18000 7831
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 21726 7868 21732 7880
rect 21687 7840 21732 7868
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7868 22799 7871
rect 23566 7868 23572 7880
rect 22787 7840 23572 7868
rect 22787 7837 22799 7840
rect 22741 7831 22799 7837
rect 23566 7828 23572 7840
rect 23624 7828 23630 7880
rect 24854 7868 24860 7880
rect 24815 7840 24860 7868
rect 24854 7828 24860 7840
rect 24912 7828 24918 7880
rect 25866 7828 25872 7880
rect 25924 7868 25930 7880
rect 27893 7871 27951 7877
rect 27893 7868 27905 7871
rect 25924 7840 27905 7868
rect 25924 7828 25930 7840
rect 27893 7837 27905 7840
rect 27939 7837 27951 7871
rect 27893 7831 27951 7837
rect 15896 7772 18000 7800
rect 15896 7760 15902 7772
rect 25130 7760 25136 7812
rect 25188 7800 25194 7812
rect 28000 7800 28028 7899
rect 32122 7896 32128 7908
rect 32180 7896 32186 7948
rect 32232 7936 32260 7976
rect 32582 7964 32588 8016
rect 32640 8004 32646 8016
rect 32640 7976 35664 8004
rect 32640 7964 32646 7976
rect 33229 7939 33287 7945
rect 33229 7936 33241 7939
rect 32232 7908 33241 7936
rect 33229 7905 33241 7908
rect 33275 7905 33287 7939
rect 33229 7899 33287 7905
rect 34517 7939 34575 7945
rect 34517 7905 34529 7939
rect 34563 7936 34575 7939
rect 34882 7936 34888 7948
rect 34563 7908 34888 7936
rect 34563 7905 34575 7908
rect 34517 7899 34575 7905
rect 34882 7896 34888 7908
rect 34940 7896 34946 7948
rect 35636 7945 35664 7976
rect 47302 7964 47308 8016
rect 47360 8004 47366 8016
rect 48961 8007 49019 8013
rect 48961 8004 48973 8007
rect 47360 7976 48973 8004
rect 47360 7964 47366 7976
rect 48961 7973 48973 7976
rect 49007 7973 49019 8007
rect 60734 8004 60740 8016
rect 48961 7967 49019 7973
rect 59280 7976 60740 8004
rect 35621 7939 35679 7945
rect 35621 7905 35633 7939
rect 35667 7905 35679 7939
rect 35621 7899 35679 7905
rect 43901 7939 43959 7945
rect 43901 7905 43913 7939
rect 43947 7936 43959 7939
rect 44358 7936 44364 7948
rect 43947 7908 44364 7936
rect 43947 7905 43959 7908
rect 43901 7899 43959 7905
rect 44358 7896 44364 7908
rect 44416 7896 44422 7948
rect 44450 7896 44456 7948
rect 44508 7936 44514 7948
rect 45005 7939 45063 7945
rect 45005 7936 45017 7939
rect 44508 7908 45017 7936
rect 44508 7896 44514 7908
rect 45005 7905 45017 7908
rect 45051 7905 45063 7939
rect 47394 7936 47400 7948
rect 47355 7908 47400 7936
rect 45005 7899 45063 7905
rect 47394 7896 47400 7908
rect 47452 7896 47458 7948
rect 58526 7936 58532 7948
rect 58487 7908 58532 7936
rect 58526 7896 58532 7908
rect 58584 7896 58590 7948
rect 59280 7945 59308 7976
rect 60734 7964 60740 7976
rect 60792 7964 60798 8016
rect 63954 8004 63960 8016
rect 62868 7976 63960 8004
rect 59265 7939 59323 7945
rect 59265 7905 59277 7939
rect 59311 7905 59323 7939
rect 59265 7899 59323 7905
rect 60185 7939 60243 7945
rect 60185 7905 60197 7939
rect 60231 7936 60243 7939
rect 61102 7936 61108 7948
rect 60231 7908 61108 7936
rect 60231 7905 60243 7908
rect 60185 7899 60243 7905
rect 61102 7896 61108 7908
rect 61160 7896 61166 7948
rect 61286 7936 61292 7948
rect 61247 7908 61292 7936
rect 61286 7896 61292 7908
rect 61344 7896 61350 7948
rect 62868 7945 62896 7976
rect 63954 7964 63960 7976
rect 64012 7964 64018 8016
rect 64966 8004 64972 8016
rect 64432 7976 64972 8004
rect 64432 7945 64460 7976
rect 64966 7964 64972 7976
rect 65024 7964 65030 8016
rect 67266 7964 67272 8016
rect 67324 8004 67330 8016
rect 67324 7976 68140 8004
rect 67324 7964 67330 7976
rect 62853 7939 62911 7945
rect 62853 7905 62865 7939
rect 62899 7905 62911 7939
rect 62853 7899 62911 7905
rect 63129 7939 63187 7945
rect 63129 7905 63141 7939
rect 63175 7905 63187 7939
rect 63129 7899 63187 7905
rect 64417 7939 64475 7945
rect 64417 7905 64429 7939
rect 64463 7905 64475 7939
rect 64417 7899 64475 7905
rect 64693 7939 64751 7945
rect 64693 7905 64705 7939
rect 64739 7905 64751 7939
rect 67818 7936 67824 7948
rect 67779 7908 67824 7936
rect 64693 7899 64751 7905
rect 29454 7828 29460 7880
rect 29512 7868 29518 7880
rect 29549 7871 29607 7877
rect 29549 7868 29561 7871
rect 29512 7840 29561 7868
rect 29512 7828 29518 7840
rect 29549 7837 29561 7840
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 30561 7871 30619 7877
rect 30561 7837 30573 7871
rect 30607 7868 30619 7871
rect 31846 7868 31852 7880
rect 30607 7840 31852 7868
rect 30607 7837 30619 7840
rect 30561 7831 30619 7837
rect 31846 7828 31852 7840
rect 31904 7828 31910 7880
rect 33137 7871 33195 7877
rect 33137 7837 33149 7871
rect 33183 7837 33195 7871
rect 33137 7831 33195 7837
rect 25188 7772 28028 7800
rect 25188 7760 25194 7772
rect 30282 7760 30288 7812
rect 30340 7800 30346 7812
rect 33152 7800 33180 7831
rect 34974 7828 34980 7880
rect 35032 7868 35038 7880
rect 35529 7871 35587 7877
rect 35529 7868 35541 7871
rect 35032 7840 35541 7868
rect 35032 7828 35038 7840
rect 35529 7837 35541 7840
rect 35575 7837 35587 7871
rect 35529 7831 35587 7837
rect 41874 7828 41880 7880
rect 41932 7868 41938 7880
rect 46293 7871 46351 7877
rect 46293 7868 46305 7871
rect 41932 7840 46305 7868
rect 41932 7828 41938 7840
rect 46293 7837 46305 7840
rect 46339 7837 46351 7871
rect 46293 7831 46351 7837
rect 47305 7871 47363 7877
rect 47305 7837 47317 7871
rect 47351 7837 47363 7871
rect 47305 7831 47363 7837
rect 30340 7772 33180 7800
rect 30340 7760 30346 7772
rect 38930 7760 38936 7812
rect 38988 7800 38994 7812
rect 45189 7803 45247 7809
rect 45189 7800 45201 7803
rect 38988 7772 45201 7800
rect 38988 7760 38994 7772
rect 45189 7769 45201 7772
rect 45235 7769 45247 7803
rect 45189 7763 45247 7769
rect 41506 7692 41512 7744
rect 41564 7732 41570 7744
rect 47320 7732 47348 7831
rect 49234 7828 49240 7880
rect 49292 7868 49298 7880
rect 49973 7871 50031 7877
rect 49973 7868 49985 7871
rect 49292 7840 49985 7868
rect 49292 7828 49298 7840
rect 49973 7837 49985 7840
rect 50019 7837 50031 7871
rect 51718 7868 51724 7880
rect 51679 7840 51724 7868
rect 49973 7831 50031 7837
rect 51718 7828 51724 7840
rect 51776 7828 51782 7880
rect 52546 7828 52552 7880
rect 52604 7868 52610 7880
rect 52733 7871 52791 7877
rect 52733 7868 52745 7871
rect 52604 7840 52745 7868
rect 52604 7828 52610 7840
rect 52733 7837 52745 7840
rect 52779 7837 52791 7871
rect 52733 7831 52791 7837
rect 61197 7871 61255 7877
rect 61197 7837 61209 7871
rect 61243 7837 61255 7871
rect 61197 7831 61255 7837
rect 62945 7871 63003 7877
rect 62945 7837 62957 7871
rect 62991 7868 63003 7871
rect 63034 7868 63040 7880
rect 62991 7840 63040 7868
rect 62991 7837 63003 7840
rect 62945 7831 63003 7837
rect 51166 7760 51172 7812
rect 51224 7800 51230 7812
rect 61212 7800 61240 7831
rect 63034 7828 63040 7840
rect 63092 7828 63098 7880
rect 51224 7772 61240 7800
rect 51224 7760 51230 7772
rect 62114 7760 62120 7812
rect 62172 7800 62178 7812
rect 63144 7800 63172 7899
rect 64506 7868 64512 7880
rect 64467 7840 64512 7868
rect 64506 7828 64512 7840
rect 64564 7828 64570 7880
rect 62172 7772 63172 7800
rect 62172 7760 62178 7772
rect 63494 7760 63500 7812
rect 63552 7800 63558 7812
rect 64708 7800 64736 7899
rect 67818 7896 67824 7908
rect 67876 7896 67882 7948
rect 68112 7945 68140 7976
rect 71774 7964 71780 8016
rect 71832 8004 71838 8016
rect 80330 8004 80336 8016
rect 71832 7976 73752 8004
rect 71832 7964 71838 7976
rect 68097 7939 68155 7945
rect 68097 7905 68109 7939
rect 68143 7905 68155 7939
rect 71406 7936 71412 7948
rect 71367 7908 71412 7936
rect 68097 7899 68155 7905
rect 71406 7896 71412 7908
rect 71464 7896 71470 7948
rect 72145 7939 72203 7945
rect 72145 7905 72157 7939
rect 72191 7905 72203 7939
rect 73430 7936 73436 7948
rect 73391 7908 73436 7936
rect 72145 7899 72203 7905
rect 64782 7828 64788 7880
rect 64840 7868 64846 7880
rect 65797 7871 65855 7877
rect 65797 7868 65809 7871
rect 64840 7840 65809 7868
rect 64840 7828 64846 7840
rect 65797 7837 65809 7840
rect 65843 7837 65855 7871
rect 67910 7868 67916 7880
rect 67871 7840 67916 7868
rect 65797 7831 65855 7837
rect 67910 7828 67916 7840
rect 67968 7828 67974 7880
rect 68830 7828 68836 7880
rect 68888 7868 68894 7880
rect 69109 7871 69167 7877
rect 69109 7868 69121 7871
rect 68888 7840 69121 7868
rect 68888 7828 68894 7840
rect 69109 7837 69121 7840
rect 69155 7837 69167 7871
rect 70118 7868 70124 7880
rect 70079 7840 70124 7868
rect 69109 7831 69167 7837
rect 70118 7828 70124 7840
rect 70176 7828 70182 7880
rect 71777 7871 71835 7877
rect 71777 7837 71789 7871
rect 71823 7868 71835 7871
rect 71958 7868 71964 7880
rect 71823 7840 71964 7868
rect 71823 7837 71835 7840
rect 71777 7831 71835 7837
rect 71958 7828 71964 7840
rect 72016 7828 72022 7880
rect 63552 7772 64736 7800
rect 72160 7800 72188 7899
rect 73430 7896 73436 7908
rect 73488 7896 73494 7948
rect 73724 7945 73752 7976
rect 78784 7976 80336 8004
rect 73709 7939 73767 7945
rect 73709 7905 73721 7939
rect 73755 7905 73767 7939
rect 75270 7936 75276 7948
rect 75231 7908 75276 7936
rect 73709 7899 73767 7905
rect 75270 7896 75276 7908
rect 75328 7896 75334 7948
rect 75733 7939 75791 7945
rect 75733 7905 75745 7939
rect 75779 7936 75791 7939
rect 78214 7936 78220 7948
rect 75779 7908 77892 7936
rect 78175 7908 78220 7936
rect 75779 7905 75791 7908
rect 75733 7899 75791 7905
rect 73522 7868 73528 7880
rect 73483 7840 73528 7868
rect 73522 7828 73528 7840
rect 73580 7828 73586 7880
rect 75365 7871 75423 7877
rect 75365 7837 75377 7871
rect 75411 7868 75423 7871
rect 75822 7868 75828 7880
rect 75411 7840 75828 7868
rect 75411 7837 75423 7840
rect 75365 7831 75423 7837
rect 75822 7828 75828 7840
rect 75880 7828 75886 7880
rect 77018 7868 77024 7880
rect 76979 7840 77024 7868
rect 77018 7828 77024 7840
rect 77076 7828 77082 7880
rect 75546 7800 75552 7812
rect 72160 7772 75552 7800
rect 63552 7760 63558 7772
rect 75546 7760 75552 7772
rect 75604 7760 75610 7812
rect 41564 7704 47348 7732
rect 41564 7692 41570 7704
rect 58250 7692 58256 7744
rect 58308 7732 58314 7744
rect 58621 7735 58679 7741
rect 58621 7732 58633 7735
rect 58308 7704 58633 7732
rect 58308 7692 58314 7704
rect 58621 7701 58633 7704
rect 58667 7701 58679 7735
rect 77864 7732 77892 7908
rect 78214 7896 78220 7908
rect 78272 7896 78278 7948
rect 78784 7945 78812 7976
rect 80330 7964 80336 7976
rect 80388 7964 80394 8016
rect 82722 8004 82728 8016
rect 80532 7976 82728 8004
rect 80532 7945 80560 7976
rect 82722 7964 82728 7976
rect 82780 7964 82786 8016
rect 85482 8004 85488 8016
rect 82832 7976 85488 8004
rect 78769 7939 78827 7945
rect 78769 7905 78781 7939
rect 78815 7905 78827 7939
rect 78769 7899 78827 7905
rect 80517 7939 80575 7945
rect 80517 7905 80529 7939
rect 80563 7905 80575 7939
rect 80974 7936 80980 7948
rect 80935 7908 80980 7936
rect 80517 7899 80575 7905
rect 80974 7896 80980 7908
rect 81032 7896 81038 7948
rect 82832 7945 82860 7976
rect 85482 7964 85488 7976
rect 85540 7964 85546 8016
rect 82817 7939 82875 7945
rect 82817 7905 82829 7939
rect 82863 7905 82875 7939
rect 82998 7936 83004 7948
rect 82959 7908 83004 7936
rect 82817 7899 82875 7905
rect 82998 7896 83004 7908
rect 83056 7896 83062 7948
rect 83185 7939 83243 7945
rect 83185 7936 83197 7939
rect 83108 7908 83197 7936
rect 78401 7871 78459 7877
rect 78401 7837 78413 7871
rect 78447 7868 78459 7871
rect 78490 7868 78496 7880
rect 78447 7840 78496 7868
rect 78447 7837 78459 7840
rect 78401 7831 78459 7837
rect 78490 7828 78496 7840
rect 78548 7828 78554 7880
rect 80606 7868 80612 7880
rect 80567 7840 80612 7868
rect 80606 7828 80612 7840
rect 80664 7828 80670 7880
rect 79502 7760 79508 7812
rect 79560 7800 79566 7812
rect 81894 7800 81900 7812
rect 79560 7772 81900 7800
rect 79560 7760 79566 7772
rect 81894 7760 81900 7772
rect 81952 7760 81958 7812
rect 83108 7800 83136 7908
rect 83185 7905 83197 7908
rect 83231 7905 83243 7939
rect 83185 7899 83243 7905
rect 83274 7896 83280 7948
rect 83332 7936 83338 7948
rect 84933 7939 84991 7945
rect 84933 7936 84945 7939
rect 83332 7908 84945 7936
rect 83332 7896 83338 7908
rect 84933 7905 84945 7908
rect 84979 7905 84991 7939
rect 85666 7936 85672 7948
rect 85627 7908 85672 7936
rect 84933 7899 84991 7905
rect 85666 7896 85672 7908
rect 85724 7896 85730 7948
rect 86512 7945 86540 8044
rect 87248 8044 91652 8072
rect 87248 7945 87276 8044
rect 91646 8032 91652 8044
rect 91704 8032 91710 8084
rect 94590 8032 94596 8084
rect 94648 8072 94654 8084
rect 97902 8072 97908 8084
rect 94648 8044 97908 8072
rect 94648 8032 94654 8044
rect 97902 8032 97908 8044
rect 97960 8032 97966 8084
rect 97994 8032 98000 8084
rect 98052 8072 98058 8084
rect 100481 8075 100539 8081
rect 100481 8072 100493 8075
rect 98052 8044 100493 8072
rect 98052 8032 98058 8044
rect 100481 8041 100493 8044
rect 100527 8041 100539 8075
rect 110966 8072 110972 8084
rect 100481 8035 100539 8041
rect 105832 8044 110972 8072
rect 99926 8004 99932 8016
rect 92492 7976 99932 8004
rect 86497 7939 86555 7945
rect 86497 7905 86509 7939
rect 86543 7905 86555 7939
rect 86497 7899 86555 7905
rect 87233 7939 87291 7945
rect 87233 7905 87245 7939
rect 87279 7905 87291 7939
rect 87233 7899 87291 7905
rect 88245 7939 88303 7945
rect 88245 7905 88257 7939
rect 88291 7905 88303 7939
rect 88245 7899 88303 7905
rect 88981 7939 89039 7945
rect 88981 7905 88993 7939
rect 89027 7936 89039 7939
rect 90910 7936 90916 7948
rect 89027 7908 89484 7936
rect 90871 7908 90916 7936
rect 89027 7905 89039 7908
rect 88981 7899 89039 7905
rect 85298 7868 85304 7880
rect 85259 7840 85304 7868
rect 85298 7828 85304 7840
rect 85356 7828 85362 7880
rect 86310 7828 86316 7880
rect 86368 7868 86374 7880
rect 88260 7868 88288 7899
rect 86368 7840 88288 7868
rect 88613 7871 88671 7877
rect 86368 7828 86374 7840
rect 88613 7837 88625 7871
rect 88659 7868 88671 7871
rect 89346 7868 89352 7880
rect 88659 7840 89352 7868
rect 88659 7837 88671 7840
rect 88613 7831 88671 7837
rect 89346 7828 89352 7840
rect 89404 7828 89410 7880
rect 86954 7800 86960 7812
rect 83108 7772 86960 7800
rect 86954 7760 86960 7772
rect 87012 7760 87018 7812
rect 88794 7800 88800 7812
rect 87708 7772 88800 7800
rect 85758 7732 85764 7744
rect 77864 7704 85764 7732
rect 58621 7695 58679 7701
rect 85758 7692 85764 7704
rect 85816 7692 85822 7744
rect 86589 7735 86647 7741
rect 86589 7701 86601 7735
rect 86635 7732 86647 7735
rect 87708 7732 87736 7772
rect 88794 7760 88800 7772
rect 88852 7760 88858 7812
rect 89456 7800 89484 7908
rect 90910 7896 90916 7908
rect 90968 7896 90974 7948
rect 91370 7936 91376 7948
rect 91331 7908 91376 7936
rect 91370 7896 91376 7908
rect 91428 7896 91434 7948
rect 92492 7945 92520 7976
rect 99926 7964 99932 7976
rect 99984 7964 99990 8016
rect 92477 7939 92535 7945
rect 92477 7905 92489 7939
rect 92523 7905 92535 7939
rect 92477 7899 92535 7905
rect 92937 7939 92995 7945
rect 92937 7905 92949 7939
rect 92983 7905 92995 7939
rect 92937 7899 92995 7905
rect 94133 7939 94191 7945
rect 94133 7905 94145 7939
rect 94179 7905 94191 7939
rect 94590 7936 94596 7948
rect 94551 7908 94596 7936
rect 94133 7899 94191 7905
rect 91002 7868 91008 7880
rect 90963 7840 91008 7868
rect 91002 7828 91008 7840
rect 91060 7828 91066 7880
rect 92566 7868 92572 7880
rect 92527 7840 92572 7868
rect 92566 7828 92572 7840
rect 92624 7828 92630 7880
rect 92842 7800 92848 7812
rect 89456 7772 92848 7800
rect 92842 7760 92848 7772
rect 92900 7760 92906 7812
rect 92952 7800 92980 7899
rect 94148 7868 94176 7899
rect 94590 7896 94596 7908
rect 94648 7896 94654 7948
rect 95510 7936 95516 7948
rect 95471 7908 95516 7936
rect 95510 7896 95516 7908
rect 95568 7896 95574 7948
rect 95789 7939 95847 7945
rect 95789 7905 95801 7939
rect 95835 7936 95847 7939
rect 96062 7936 96068 7948
rect 95835 7908 96068 7936
rect 95835 7905 95847 7908
rect 95789 7899 95847 7905
rect 96062 7896 96068 7908
rect 96120 7896 96126 7948
rect 96157 7939 96215 7945
rect 96157 7905 96169 7939
rect 96203 7905 96215 7939
rect 96982 7936 96988 7948
rect 96943 7908 96988 7936
rect 96157 7899 96215 7905
rect 96172 7868 96200 7899
rect 96982 7896 96988 7908
rect 97040 7896 97046 7948
rect 98454 7936 98460 7948
rect 97092 7908 98460 7936
rect 97092 7868 97120 7908
rect 98454 7896 98460 7908
rect 98512 7896 98518 7948
rect 98549 7939 98607 7945
rect 98549 7905 98561 7939
rect 98595 7936 98607 7939
rect 98595 7908 98776 7936
rect 98595 7905 98607 7908
rect 98549 7899 98607 7905
rect 98362 7868 98368 7880
rect 94148 7840 95740 7868
rect 96172 7840 97120 7868
rect 98323 7840 98368 7868
rect 95602 7800 95608 7812
rect 92952 7772 95608 7800
rect 95602 7760 95608 7772
rect 95660 7760 95666 7812
rect 86635 7704 87736 7732
rect 93949 7735 94007 7741
rect 86635 7701 86647 7704
rect 86589 7695 86647 7701
rect 93949 7701 93961 7735
rect 93995 7732 94007 7735
rect 94590 7732 94596 7744
rect 93995 7704 94596 7732
rect 93995 7701 94007 7704
rect 93949 7695 94007 7701
rect 94590 7692 94596 7704
rect 94648 7692 94654 7744
rect 95712 7732 95740 7840
rect 98362 7828 98368 7840
rect 98420 7828 98426 7880
rect 95786 7760 95792 7812
rect 95844 7800 95850 7812
rect 98638 7800 98644 7812
rect 95844 7772 98644 7800
rect 95844 7760 95850 7772
rect 98638 7760 98644 7772
rect 98696 7760 98702 7812
rect 98748 7800 98776 7908
rect 98822 7896 98828 7948
rect 98880 7936 98886 7948
rect 102134 7936 102140 7948
rect 98880 7908 102140 7936
rect 98880 7896 98886 7908
rect 102134 7896 102140 7908
rect 102192 7896 102198 7948
rect 102226 7896 102232 7948
rect 102284 7936 102290 7948
rect 102413 7939 102471 7945
rect 102413 7936 102425 7939
rect 102284 7908 102425 7936
rect 102284 7896 102290 7908
rect 102413 7905 102425 7908
rect 102459 7905 102471 7939
rect 102413 7899 102471 7905
rect 103977 7939 104035 7945
rect 103977 7905 103989 7939
rect 104023 7936 104035 7939
rect 104066 7936 104072 7948
rect 104023 7908 104072 7936
rect 104023 7905 104035 7908
rect 103977 7899 104035 7905
rect 104066 7896 104072 7908
rect 104124 7896 104130 7948
rect 105354 7936 105360 7948
rect 105315 7908 105360 7936
rect 105354 7896 105360 7908
rect 105412 7896 105418 7948
rect 105832 7945 105860 8044
rect 110966 8032 110972 8044
rect 111024 8032 111030 8084
rect 111058 8032 111064 8084
rect 111116 8072 111122 8084
rect 124766 8072 124772 8084
rect 111116 8044 124772 8072
rect 111116 8032 111122 8044
rect 124766 8032 124772 8044
rect 124824 8032 124830 8084
rect 141142 8072 141148 8084
rect 127544 8044 141148 8072
rect 107746 7964 107752 8016
rect 107804 8004 107810 8016
rect 122282 8004 122288 8016
rect 107804 7976 109540 8004
rect 107804 7964 107810 7976
rect 105817 7939 105875 7945
rect 105817 7905 105829 7939
rect 105863 7905 105875 7939
rect 107562 7936 107568 7948
rect 107523 7908 107568 7936
rect 105817 7899 105875 7905
rect 107562 7896 107568 7908
rect 107620 7896 107626 7948
rect 107654 7896 107660 7948
rect 107712 7936 107718 7948
rect 107933 7939 107991 7945
rect 107933 7936 107945 7939
rect 107712 7908 107945 7936
rect 107712 7896 107718 7908
rect 107933 7905 107945 7908
rect 107979 7905 107991 7939
rect 109218 7936 109224 7948
rect 109179 7908 109224 7936
rect 107933 7899 107991 7905
rect 109218 7896 109224 7908
rect 109276 7896 109282 7948
rect 109512 7945 109540 7976
rect 112824 7976 122288 8004
rect 109497 7939 109555 7945
rect 109497 7905 109509 7939
rect 109543 7905 109555 7939
rect 109497 7899 109555 7905
rect 110414 7896 110420 7948
rect 110472 7936 110478 7948
rect 112824 7945 112852 7976
rect 122282 7964 122288 7976
rect 122340 7964 122346 8016
rect 123202 7964 123208 8016
rect 123260 8004 123266 8016
rect 123260 7976 124996 8004
rect 123260 7964 123266 7976
rect 111245 7939 111303 7945
rect 111245 7936 111257 7939
rect 110472 7908 111257 7936
rect 110472 7896 110478 7908
rect 111245 7905 111257 7908
rect 111291 7905 111303 7939
rect 111245 7899 111303 7905
rect 112809 7939 112867 7945
rect 112809 7905 112821 7939
rect 112855 7905 112867 7939
rect 112809 7899 112867 7905
rect 115201 7939 115259 7945
rect 115201 7905 115213 7939
rect 115247 7936 115259 7939
rect 115842 7936 115848 7948
rect 115247 7908 115848 7936
rect 115247 7905 115259 7908
rect 115201 7899 115259 7905
rect 115842 7896 115848 7908
rect 115900 7896 115906 7948
rect 118694 7896 118700 7948
rect 118752 7936 118758 7948
rect 120261 7939 120319 7945
rect 118752 7908 118797 7936
rect 118752 7896 118758 7908
rect 120261 7905 120273 7939
rect 120307 7936 120319 7939
rect 123294 7936 123300 7948
rect 120307 7908 123156 7936
rect 123255 7908 123300 7936
rect 120307 7905 120319 7908
rect 120261 7899 120319 7905
rect 99466 7868 99472 7880
rect 99427 7840 99472 7868
rect 99466 7828 99472 7840
rect 99524 7828 99530 7880
rect 99558 7828 99564 7880
rect 99616 7868 99622 7880
rect 103422 7868 103428 7880
rect 99616 7840 103428 7868
rect 99616 7828 99622 7840
rect 103422 7828 103428 7840
rect 103480 7828 103486 7880
rect 105449 7871 105507 7877
rect 105449 7837 105461 7871
rect 105495 7868 105507 7871
rect 106734 7868 106740 7880
rect 105495 7840 106740 7868
rect 105495 7837 105507 7840
rect 105449 7831 105507 7837
rect 106734 7828 106740 7840
rect 106792 7828 106798 7880
rect 107746 7868 107752 7880
rect 107707 7840 107752 7868
rect 107746 7828 107752 7840
rect 107804 7828 107810 7880
rect 112070 7828 112076 7880
rect 112128 7868 112134 7880
rect 113637 7871 113695 7877
rect 113637 7868 113649 7871
rect 112128 7840 113649 7868
rect 112128 7828 112134 7840
rect 113637 7837 113649 7840
rect 113683 7837 113695 7871
rect 116302 7868 116308 7880
rect 116263 7840 116308 7868
rect 113637 7831 113695 7837
rect 116302 7828 116308 7840
rect 116360 7828 116366 7880
rect 117685 7871 117743 7877
rect 117685 7837 117697 7871
rect 117731 7868 117743 7871
rect 119062 7868 119068 7880
rect 117731 7840 119068 7868
rect 117731 7837 117743 7840
rect 117685 7831 117743 7837
rect 119062 7828 119068 7840
rect 119120 7828 119126 7880
rect 122009 7871 122067 7877
rect 122009 7837 122021 7871
rect 122055 7868 122067 7871
rect 122650 7868 122656 7880
rect 122055 7840 122656 7868
rect 122055 7837 122067 7840
rect 122009 7831 122067 7837
rect 122650 7828 122656 7840
rect 122708 7828 122714 7880
rect 103882 7800 103888 7812
rect 98748 7772 103744 7800
rect 103843 7772 103888 7800
rect 100938 7732 100944 7744
rect 95712 7704 100944 7732
rect 100938 7692 100944 7704
rect 100996 7692 101002 7744
rect 103716 7732 103744 7772
rect 103882 7760 103888 7772
rect 103940 7760 103946 7812
rect 106274 7760 106280 7812
rect 106332 7800 106338 7812
rect 112717 7803 112775 7809
rect 106332 7772 112576 7800
rect 106332 7760 106338 7772
rect 104802 7732 104808 7744
rect 103716 7704 104808 7732
rect 104802 7692 104808 7704
rect 104860 7692 104866 7744
rect 109034 7692 109040 7744
rect 109092 7732 109098 7744
rect 109092 7704 109137 7732
rect 109092 7692 109098 7704
rect 110782 7692 110788 7744
rect 110840 7732 110846 7744
rect 111978 7732 111984 7744
rect 110840 7704 111984 7732
rect 110840 7692 110846 7704
rect 111978 7692 111984 7704
rect 112036 7692 112042 7744
rect 112548 7732 112576 7772
rect 112717 7769 112729 7803
rect 112763 7800 112775 7803
rect 114186 7800 114192 7812
rect 112763 7772 114192 7800
rect 112763 7769 112775 7772
rect 112717 7763 112775 7769
rect 114186 7760 114192 7772
rect 114244 7760 114250 7812
rect 115109 7803 115167 7809
rect 115109 7769 115121 7803
rect 115155 7800 115167 7803
rect 119982 7800 119988 7812
rect 115155 7772 119988 7800
rect 115155 7769 115167 7772
rect 115109 7763 115167 7769
rect 119982 7760 119988 7772
rect 120040 7760 120046 7812
rect 120166 7800 120172 7812
rect 120127 7772 120172 7800
rect 120166 7760 120172 7772
rect 120224 7760 120230 7812
rect 118234 7732 118240 7744
rect 112548 7704 118240 7732
rect 118234 7692 118240 7704
rect 118292 7692 118298 7744
rect 123128 7732 123156 7908
rect 123294 7896 123300 7908
rect 123352 7896 123358 7948
rect 124858 7936 124864 7948
rect 124819 7908 124864 7936
rect 124858 7896 124864 7908
rect 124916 7896 124922 7948
rect 124398 7760 124404 7812
rect 124456 7800 124462 7812
rect 124585 7803 124643 7809
rect 124585 7800 124597 7803
rect 124456 7772 124597 7800
rect 124456 7760 124462 7772
rect 124585 7769 124597 7772
rect 124631 7769 124643 7803
rect 124968 7800 124996 7976
rect 127544 7945 127572 8044
rect 141142 8032 141148 8044
rect 141200 8032 141206 8084
rect 141234 8032 141240 8084
rect 141292 8072 141298 8084
rect 163317 8075 163375 8081
rect 141292 8044 162164 8072
rect 141292 8032 141298 8044
rect 135533 8007 135591 8013
rect 135533 8004 135545 8007
rect 130396 7976 135545 8004
rect 130396 7945 130424 7976
rect 135533 7973 135545 7976
rect 135579 7973 135591 8007
rect 135533 7967 135591 7973
rect 137830 7964 137836 8016
rect 137888 8004 137894 8016
rect 137888 7976 140636 8004
rect 137888 7964 137894 7976
rect 127529 7939 127587 7945
rect 127529 7905 127541 7939
rect 127575 7905 127587 7939
rect 127529 7899 127587 7905
rect 129093 7939 129151 7945
rect 129093 7905 129105 7939
rect 129139 7905 129151 7939
rect 129093 7899 129151 7905
rect 130381 7939 130439 7945
rect 130381 7905 130393 7939
rect 130427 7905 130439 7939
rect 130381 7899 130439 7905
rect 125686 7868 125692 7880
rect 125647 7840 125692 7868
rect 125686 7828 125692 7840
rect 125744 7828 125750 7880
rect 128354 7828 128360 7880
rect 128412 7868 128418 7880
rect 128541 7871 128599 7877
rect 128541 7868 128553 7871
rect 128412 7840 128553 7868
rect 128412 7828 128418 7840
rect 128541 7837 128553 7840
rect 128587 7837 128599 7871
rect 129108 7868 129136 7899
rect 131390 7896 131396 7948
rect 131448 7936 131454 7948
rect 131485 7939 131543 7945
rect 131485 7936 131497 7939
rect 131448 7908 131497 7936
rect 131448 7896 131454 7908
rect 131485 7905 131497 7908
rect 131531 7905 131543 7939
rect 131485 7899 131543 7905
rect 133230 7896 133236 7948
rect 133288 7936 133294 7948
rect 134245 7939 134303 7945
rect 134245 7936 134257 7939
rect 133288 7908 134257 7936
rect 133288 7896 133294 7908
rect 134245 7905 134257 7908
rect 134291 7905 134303 7939
rect 134245 7899 134303 7905
rect 134334 7896 134340 7948
rect 134392 7936 134398 7948
rect 137557 7939 137615 7945
rect 137557 7936 137569 7939
rect 134392 7908 137569 7936
rect 134392 7896 134398 7908
rect 137557 7905 137569 7908
rect 137603 7905 137615 7939
rect 137557 7899 137615 7905
rect 139486 7896 139492 7948
rect 139544 7936 139550 7948
rect 139857 7939 139915 7945
rect 139857 7936 139869 7939
rect 139544 7908 139869 7936
rect 139544 7896 139550 7908
rect 139857 7905 139869 7908
rect 139903 7905 139915 7939
rect 139857 7899 139915 7905
rect 139946 7896 139952 7948
rect 140004 7936 140010 7948
rect 140498 7936 140504 7948
rect 140004 7908 140504 7936
rect 140004 7896 140010 7908
rect 140498 7896 140504 7908
rect 140556 7896 140562 7948
rect 140608 7936 140636 7976
rect 141970 7964 141976 8016
rect 142028 8004 142034 8016
rect 147214 8004 147220 8016
rect 142028 7976 147220 8004
rect 142028 7964 142034 7976
rect 147214 7964 147220 7976
rect 147272 7964 147278 8016
rect 160646 8004 160652 8016
rect 147324 7976 160652 8004
rect 144365 7939 144423 7945
rect 144365 7936 144377 7939
rect 140608 7908 144377 7936
rect 144365 7905 144377 7908
rect 144411 7905 144423 7939
rect 144365 7899 144423 7905
rect 145006 7896 145012 7948
rect 145064 7936 145070 7948
rect 146941 7939 146999 7945
rect 146941 7936 146953 7939
rect 145064 7908 146953 7936
rect 145064 7896 145070 7908
rect 146941 7905 146953 7908
rect 146987 7905 146999 7939
rect 146941 7899 146999 7905
rect 130838 7868 130844 7880
rect 129108 7840 130844 7868
rect 128541 7831 128599 7837
rect 130838 7828 130844 7840
rect 130896 7828 130902 7880
rect 133141 7871 133199 7877
rect 130948 7840 131988 7868
rect 130948 7800 130976 7840
rect 124968 7772 130976 7800
rect 131853 7803 131911 7809
rect 124585 7763 124643 7769
rect 131853 7769 131865 7803
rect 131899 7769 131911 7803
rect 131960 7800 131988 7840
rect 133141 7837 133153 7871
rect 133187 7868 133199 7871
rect 136545 7871 136603 7877
rect 136545 7868 136557 7871
rect 133187 7840 136557 7868
rect 133187 7837 133199 7840
rect 133141 7831 133199 7837
rect 136545 7837 136557 7840
rect 136591 7837 136603 7871
rect 136545 7831 136603 7837
rect 138753 7871 138811 7877
rect 138753 7837 138765 7871
rect 138799 7868 138811 7871
rect 140774 7868 140780 7880
rect 138799 7840 140780 7868
rect 138799 7837 138811 7840
rect 138753 7831 138811 7837
rect 140774 7828 140780 7840
rect 140832 7828 140838 7880
rect 141142 7868 141148 7880
rect 141103 7840 141148 7868
rect 141142 7828 141148 7840
rect 141200 7828 141206 7880
rect 142246 7828 142252 7880
rect 142304 7868 142310 7880
rect 142617 7871 142675 7877
rect 142617 7868 142629 7871
rect 142304 7840 142629 7868
rect 142304 7828 142310 7840
rect 142617 7837 142629 7840
rect 142663 7837 142675 7871
rect 142617 7831 142675 7837
rect 145837 7871 145895 7877
rect 145837 7837 145849 7871
rect 145883 7868 145895 7871
rect 145926 7868 145932 7880
rect 145883 7840 145932 7868
rect 145883 7837 145895 7840
rect 145837 7831 145895 7837
rect 145926 7828 145932 7840
rect 145984 7828 145990 7880
rect 147324 7877 147352 7976
rect 160646 7964 160652 7976
rect 160704 7964 160710 8016
rect 162136 8004 162164 8044
rect 163317 8041 163329 8075
rect 163363 8072 163375 8075
rect 164234 8072 164240 8084
rect 163363 8044 164240 8072
rect 163363 8041 163375 8044
rect 163317 8035 163375 8041
rect 164234 8032 164240 8044
rect 164292 8032 164298 8084
rect 164326 8032 164332 8084
rect 164384 8072 164390 8084
rect 165062 8072 165068 8084
rect 164384 8044 165068 8072
rect 164384 8032 164390 8044
rect 165062 8032 165068 8044
rect 165120 8032 165126 8084
rect 167270 8032 167276 8084
rect 167328 8072 167334 8084
rect 171134 8072 171140 8084
rect 167328 8044 171140 8072
rect 167328 8032 167334 8044
rect 171134 8032 171140 8044
rect 171192 8032 171198 8084
rect 171321 8075 171379 8081
rect 171321 8041 171333 8075
rect 171367 8072 171379 8075
rect 172330 8072 172336 8084
rect 171367 8044 172336 8072
rect 171367 8041 171379 8044
rect 171321 8035 171379 8041
rect 172330 8032 172336 8044
rect 172388 8032 172394 8084
rect 172698 8032 172704 8084
rect 172756 8072 172762 8084
rect 181346 8072 181352 8084
rect 172756 8044 181352 8072
rect 172756 8032 172762 8044
rect 181346 8032 181352 8044
rect 181404 8032 181410 8084
rect 181530 8032 181536 8084
rect 181588 8072 181594 8084
rect 183738 8072 183744 8084
rect 181588 8044 183744 8072
rect 181588 8032 181594 8044
rect 183738 8032 183744 8044
rect 183796 8032 183802 8084
rect 184385 8075 184443 8081
rect 184385 8041 184397 8075
rect 184431 8072 184443 8075
rect 184842 8072 184848 8084
rect 184431 8044 184848 8072
rect 184431 8041 184443 8044
rect 184385 8035 184443 8041
rect 184842 8032 184848 8044
rect 184900 8032 184906 8084
rect 184934 8032 184940 8084
rect 184992 8072 184998 8084
rect 189442 8072 189448 8084
rect 184992 8044 189448 8072
rect 184992 8032 184998 8044
rect 189442 8032 189448 8044
rect 189500 8032 189506 8084
rect 190546 8032 190552 8084
rect 190604 8072 190610 8084
rect 195330 8072 195336 8084
rect 190604 8044 195336 8072
rect 190604 8032 190610 8044
rect 195330 8032 195336 8044
rect 195388 8032 195394 8084
rect 197354 8072 197360 8084
rect 197315 8044 197360 8072
rect 197354 8032 197360 8044
rect 197412 8032 197418 8084
rect 164602 8004 164608 8016
rect 162136 7976 164608 8004
rect 164602 7964 164608 7976
rect 164660 7964 164666 8016
rect 168466 7964 168472 8016
rect 168524 8004 168530 8016
rect 168524 7976 194916 8004
rect 168524 7964 168530 7976
rect 152093 7939 152151 7945
rect 152093 7905 152105 7939
rect 152139 7936 152151 7939
rect 154114 7936 154120 7948
rect 152139 7908 154120 7936
rect 152139 7905 152151 7908
rect 152093 7899 152151 7905
rect 154114 7896 154120 7908
rect 154172 7896 154178 7948
rect 154209 7939 154267 7945
rect 154209 7905 154221 7939
rect 154255 7905 154267 7939
rect 154209 7899 154267 7905
rect 147309 7871 147367 7877
rect 147309 7837 147321 7871
rect 147355 7837 147367 7871
rect 147309 7831 147367 7837
rect 147766 7828 147772 7880
rect 147824 7868 147830 7880
rect 148229 7871 148287 7877
rect 148229 7868 148241 7871
rect 147824 7840 148241 7868
rect 147824 7828 147830 7840
rect 148229 7837 148241 7840
rect 148275 7837 148287 7871
rect 150066 7868 150072 7880
rect 150027 7840 150072 7868
rect 148229 7831 148287 7837
rect 150066 7828 150072 7840
rect 150124 7828 150130 7880
rect 151078 7868 151084 7880
rect 151039 7840 151084 7868
rect 151078 7828 151084 7840
rect 151136 7828 151142 7880
rect 153010 7868 153016 7880
rect 151188 7840 153016 7868
rect 133506 7800 133512 7812
rect 131960 7772 133512 7800
rect 131853 7763 131911 7769
rect 129826 7732 129832 7744
rect 123128 7704 129832 7732
rect 129826 7692 129832 7704
rect 129884 7692 129890 7744
rect 131868 7732 131896 7763
rect 133506 7760 133512 7772
rect 133564 7760 133570 7812
rect 133598 7760 133604 7812
rect 133656 7800 133662 7812
rect 134426 7800 134432 7812
rect 133656 7772 134432 7800
rect 133656 7760 133662 7772
rect 134426 7760 134432 7772
rect 134484 7760 134490 7812
rect 134610 7800 134616 7812
rect 134571 7772 134616 7800
rect 134610 7760 134616 7772
rect 134668 7760 134674 7812
rect 134702 7760 134708 7812
rect 134760 7800 134766 7812
rect 139946 7800 139952 7812
rect 134760 7772 139952 7800
rect 134760 7760 134766 7772
rect 139946 7760 139952 7772
rect 140004 7760 140010 7812
rect 140222 7800 140228 7812
rect 140183 7772 140228 7800
rect 140222 7760 140228 7772
rect 140280 7760 140286 7812
rect 140314 7760 140320 7812
rect 140372 7800 140378 7812
rect 151188 7800 151216 7840
rect 153010 7828 153016 7840
rect 153068 7828 153074 7880
rect 153105 7871 153163 7877
rect 153105 7837 153117 7871
rect 153151 7868 153163 7871
rect 153286 7868 153292 7880
rect 153151 7840 153292 7868
rect 153151 7837 153163 7840
rect 153105 7831 153163 7837
rect 153286 7828 153292 7840
rect 153344 7828 153350 7880
rect 140372 7772 151216 7800
rect 140372 7760 140378 7772
rect 152458 7760 152464 7812
rect 152516 7800 152522 7812
rect 154224 7800 154252 7899
rect 154298 7896 154304 7948
rect 154356 7936 154362 7948
rect 155589 7939 155647 7945
rect 155589 7936 155601 7939
rect 154356 7908 155601 7936
rect 154356 7896 154362 7908
rect 155589 7905 155601 7908
rect 155635 7905 155647 7939
rect 155589 7899 155647 7905
rect 155862 7896 155868 7948
rect 155920 7936 155926 7948
rect 156693 7939 156751 7945
rect 156693 7936 156705 7939
rect 155920 7908 156705 7936
rect 155920 7896 155926 7908
rect 156693 7905 156705 7908
rect 156739 7905 156751 7939
rect 156693 7899 156751 7905
rect 156782 7896 156788 7948
rect 156840 7936 156846 7948
rect 156840 7908 157840 7936
rect 156840 7896 156846 7908
rect 156598 7868 156604 7880
rect 152516 7772 154252 7800
rect 154316 7840 156604 7868
rect 152516 7760 152522 7772
rect 154316 7732 154344 7840
rect 156598 7828 156604 7840
rect 156656 7828 156662 7880
rect 157061 7871 157119 7877
rect 157061 7837 157073 7871
rect 157107 7868 157119 7871
rect 157702 7868 157708 7880
rect 157107 7840 157708 7868
rect 157107 7837 157119 7840
rect 157061 7831 157119 7837
rect 157702 7828 157708 7840
rect 157760 7828 157766 7880
rect 157812 7868 157840 7908
rect 157978 7896 157984 7948
rect 158036 7936 158042 7948
rect 158625 7939 158683 7945
rect 158625 7936 158637 7939
rect 158036 7908 158637 7936
rect 158036 7896 158042 7908
rect 158625 7905 158637 7908
rect 158671 7905 158683 7939
rect 159910 7936 159916 7948
rect 159871 7908 159916 7936
rect 158625 7899 158683 7905
rect 159910 7896 159916 7908
rect 159968 7896 159974 7948
rect 161293 7939 161351 7945
rect 161293 7905 161305 7939
rect 161339 7936 161351 7939
rect 164234 7936 164240 7948
rect 161339 7908 164240 7936
rect 161339 7905 161351 7908
rect 161293 7899 161351 7905
rect 164234 7896 164240 7908
rect 164292 7896 164298 7948
rect 164329 7939 164387 7945
rect 164329 7905 164341 7939
rect 164375 7936 164387 7939
rect 164510 7936 164516 7948
rect 164375 7908 164516 7936
rect 164375 7905 164387 7908
rect 164329 7899 164387 7905
rect 164510 7896 164516 7908
rect 164568 7896 164574 7948
rect 165893 7939 165951 7945
rect 165893 7905 165905 7939
rect 165939 7936 165951 7939
rect 169297 7939 169355 7945
rect 165939 7908 167500 7936
rect 165939 7905 165951 7908
rect 165893 7899 165951 7905
rect 158346 7868 158352 7880
rect 157812 7840 158352 7868
rect 158346 7828 158352 7840
rect 158404 7828 158410 7880
rect 161198 7868 161204 7880
rect 160020 7840 161204 7868
rect 154577 7803 154635 7809
rect 154577 7769 154589 7803
rect 154623 7769 154635 7803
rect 154577 7763 154635 7769
rect 131868 7704 154344 7732
rect 154592 7732 154620 7763
rect 155954 7760 155960 7812
rect 156012 7800 156018 7812
rect 160020 7800 160048 7840
rect 161198 7828 161204 7840
rect 161256 7828 161262 7880
rect 162302 7868 162308 7880
rect 162263 7840 162308 7868
rect 162302 7828 162308 7840
rect 162360 7828 162366 7880
rect 165801 7871 165859 7877
rect 165801 7837 165813 7871
rect 165847 7868 165859 7871
rect 167270 7868 167276 7880
rect 165847 7840 167276 7868
rect 165847 7837 165859 7840
rect 165801 7831 165859 7837
rect 167270 7828 167276 7840
rect 167328 7828 167334 7880
rect 156012 7772 160048 7800
rect 160097 7803 160155 7809
rect 156012 7760 156018 7772
rect 160097 7769 160109 7803
rect 160143 7800 160155 7803
rect 166994 7800 167000 7812
rect 160143 7772 167000 7800
rect 160143 7769 160155 7772
rect 160097 7763 160155 7769
rect 166994 7760 167000 7772
rect 167052 7760 167058 7812
rect 167472 7800 167500 7908
rect 169297 7905 169309 7939
rect 169343 7905 169355 7939
rect 169297 7899 169355 7905
rect 170125 7939 170183 7945
rect 170125 7905 170137 7939
rect 170171 7936 170183 7939
rect 172425 7939 172483 7945
rect 172425 7936 172437 7939
rect 170171 7908 172437 7936
rect 170171 7905 170183 7908
rect 170125 7899 170183 7905
rect 172425 7905 172437 7908
rect 172471 7905 172483 7939
rect 173526 7936 173532 7948
rect 173487 7908 173532 7936
rect 172425 7899 172483 7905
rect 167730 7868 167736 7880
rect 167691 7840 167736 7868
rect 167730 7828 167736 7840
rect 167788 7828 167794 7880
rect 169312 7868 169340 7899
rect 173526 7896 173532 7908
rect 173584 7896 173590 7948
rect 173710 7896 173716 7948
rect 173768 7936 173774 7948
rect 174909 7939 174967 7945
rect 174909 7936 174921 7939
rect 173768 7908 174921 7936
rect 173768 7896 173774 7908
rect 174909 7905 174921 7908
rect 174955 7905 174967 7939
rect 176470 7936 176476 7948
rect 176431 7908 176476 7936
rect 174909 7899 174967 7905
rect 176470 7896 176476 7908
rect 176528 7896 176534 7948
rect 178034 7936 178040 7948
rect 177995 7908 178040 7936
rect 178034 7896 178040 7908
rect 178092 7896 178098 7948
rect 179601 7939 179659 7945
rect 179601 7905 179613 7939
rect 179647 7936 179659 7939
rect 182082 7936 182088 7948
rect 179647 7908 182088 7936
rect 179647 7905 179659 7908
rect 179601 7899 179659 7905
rect 182082 7896 182088 7908
rect 182140 7896 182146 7948
rect 182450 7936 182456 7948
rect 182411 7908 182456 7936
rect 182450 7896 182456 7908
rect 182508 7896 182514 7948
rect 183554 7896 183560 7948
rect 183612 7936 183618 7948
rect 187237 7939 187295 7945
rect 183612 7908 185900 7936
rect 183612 7896 183618 7908
rect 179506 7868 179512 7880
rect 169312 7840 178540 7868
rect 179467 7840 179512 7868
rect 169205 7803 169263 7809
rect 167472 7772 168512 7800
rect 166442 7732 166448 7744
rect 154592 7704 166448 7732
rect 166442 7692 166448 7704
rect 166500 7692 166506 7744
rect 168484 7732 168512 7772
rect 169205 7769 169217 7803
rect 169251 7800 169263 7803
rect 172698 7800 172704 7812
rect 169251 7772 172704 7800
rect 169251 7769 169263 7772
rect 169205 7763 169263 7769
rect 172698 7760 172704 7772
rect 172756 7760 172762 7812
rect 173894 7800 173900 7812
rect 173855 7772 173900 7800
rect 173894 7760 173900 7772
rect 173952 7760 173958 7812
rect 176194 7800 176200 7812
rect 176155 7772 176200 7800
rect 176194 7760 176200 7772
rect 176252 7760 176258 7812
rect 176378 7760 176384 7812
rect 176436 7800 176442 7812
rect 178402 7800 178408 7812
rect 176436 7772 178408 7800
rect 176436 7760 176442 7772
rect 178402 7760 178408 7772
rect 178460 7760 178466 7812
rect 178512 7800 178540 7840
rect 179506 7828 179512 7840
rect 179564 7828 179570 7880
rect 181162 7868 181168 7880
rect 181123 7840 181168 7868
rect 181162 7828 181168 7840
rect 181220 7828 181226 7880
rect 182542 7868 182548 7880
rect 182503 7840 182548 7868
rect 182542 7828 182548 7840
rect 182600 7828 182606 7880
rect 182818 7828 182824 7880
rect 182876 7868 182882 7880
rect 185673 7871 185731 7877
rect 185673 7868 185685 7871
rect 182876 7840 185685 7868
rect 182876 7828 182882 7840
rect 185673 7837 185685 7840
rect 185719 7837 185731 7871
rect 185872 7868 185900 7908
rect 187237 7905 187249 7939
rect 187283 7936 187295 7939
rect 187878 7936 187884 7948
rect 187283 7908 187884 7936
rect 187283 7905 187295 7908
rect 187237 7899 187295 7905
rect 187878 7896 187884 7908
rect 187936 7896 187942 7948
rect 188065 7939 188123 7945
rect 188065 7905 188077 7939
rect 188111 7936 188123 7939
rect 190546 7936 190552 7948
rect 188111 7908 190552 7936
rect 188111 7905 188123 7908
rect 188065 7899 188123 7905
rect 190546 7896 190552 7908
rect 190604 7896 190610 7948
rect 190641 7939 190699 7945
rect 190641 7905 190653 7939
rect 190687 7905 190699 7939
rect 191650 7936 191656 7948
rect 191611 7908 191656 7936
rect 190641 7899 190699 7905
rect 188157 7871 188215 7877
rect 188157 7868 188169 7871
rect 185872 7840 188169 7868
rect 185673 7831 185731 7837
rect 188157 7837 188169 7840
rect 188203 7837 188215 7871
rect 188157 7831 188215 7837
rect 189261 7871 189319 7877
rect 189261 7837 189273 7871
rect 189307 7837 189319 7871
rect 189261 7831 189319 7837
rect 183554 7800 183560 7812
rect 178512 7772 183560 7800
rect 183554 7760 183560 7772
rect 183612 7760 183618 7812
rect 184658 7760 184664 7812
rect 184716 7800 184722 7812
rect 184842 7800 184848 7812
rect 184716 7772 184848 7800
rect 184716 7760 184722 7772
rect 184842 7760 184848 7772
rect 184900 7760 184906 7812
rect 187145 7803 187203 7809
rect 187145 7769 187157 7803
rect 187191 7800 187203 7803
rect 189166 7800 189172 7812
rect 187191 7772 189172 7800
rect 187191 7769 187203 7772
rect 187145 7763 187203 7769
rect 189166 7760 189172 7772
rect 189224 7760 189230 7812
rect 170030 7732 170036 7744
rect 168484 7704 170036 7732
rect 170030 7692 170036 7704
rect 170088 7692 170094 7744
rect 171042 7692 171048 7744
rect 171100 7732 171106 7744
rect 176562 7732 176568 7744
rect 171100 7704 176568 7732
rect 171100 7692 171106 7704
rect 176562 7692 176568 7704
rect 176620 7692 176626 7744
rect 176654 7692 176660 7744
rect 176712 7732 176718 7744
rect 181806 7732 181812 7744
rect 176712 7704 181812 7732
rect 176712 7692 176718 7704
rect 181806 7692 181812 7704
rect 181864 7692 181870 7744
rect 182634 7692 182640 7744
rect 182692 7732 182698 7744
rect 189276 7732 189304 7831
rect 190549 7803 190607 7809
rect 190549 7769 190561 7803
rect 190595 7769 190607 7803
rect 190656 7800 190684 7899
rect 191650 7896 191656 7908
rect 191708 7896 191714 7948
rect 192754 7936 192760 7948
rect 192715 7908 192760 7936
rect 192754 7896 192760 7908
rect 192812 7896 192818 7948
rect 194888 7945 194916 7976
rect 194873 7939 194931 7945
rect 194873 7905 194885 7939
rect 194919 7905 194931 7939
rect 194873 7899 194931 7905
rect 194962 7896 194968 7948
rect 195020 7936 195026 7948
rect 195977 7939 196035 7945
rect 195977 7936 195989 7939
rect 195020 7908 195989 7936
rect 195020 7896 195026 7908
rect 195977 7905 195989 7908
rect 196023 7905 196035 7939
rect 195977 7899 196035 7905
rect 197078 7896 197084 7948
rect 197136 7936 197142 7948
rect 197265 7939 197323 7945
rect 197265 7936 197277 7939
rect 197136 7908 197277 7936
rect 197136 7896 197142 7908
rect 197265 7905 197277 7908
rect 197311 7905 197323 7939
rect 197265 7899 197323 7905
rect 192846 7868 192852 7880
rect 192807 7840 192852 7868
rect 192846 7828 192852 7840
rect 192904 7828 192910 7880
rect 195790 7828 195796 7880
rect 195848 7868 195854 7880
rect 196069 7871 196127 7877
rect 196069 7868 196081 7871
rect 195848 7840 196081 7868
rect 195848 7828 195854 7840
rect 196069 7837 196081 7840
rect 196115 7837 196127 7871
rect 196069 7831 196127 7837
rect 192938 7800 192944 7812
rect 190656 7772 192944 7800
rect 190549 7763 190607 7769
rect 182692 7704 189304 7732
rect 190564 7732 190592 7763
rect 192938 7760 192944 7772
rect 192996 7760 193002 7812
rect 199286 7732 199292 7744
rect 190564 7704 199292 7732
rect 182692 7692 182698 7704
rect 199286 7692 199292 7704
rect 199344 7692 199350 7744
rect 1104 7642 198812 7664
rect 1104 7590 4078 7642
rect 4130 7590 44078 7642
rect 44130 7590 84078 7642
rect 84130 7590 124078 7642
rect 124130 7590 164078 7642
rect 164130 7590 198812 7642
rect 1104 7568 198812 7590
rect 17586 7488 17592 7540
rect 17644 7528 17650 7540
rect 17644 7500 24992 7528
rect 17644 7488 17650 7500
rect 5813 7463 5871 7469
rect 5813 7429 5825 7463
rect 5859 7460 5871 7463
rect 7006 7460 7012 7472
rect 5859 7432 7012 7460
rect 5859 7429 5871 7432
rect 5813 7423 5871 7429
rect 7006 7420 7012 7432
rect 7064 7420 7070 7472
rect 8757 7463 8815 7469
rect 8757 7429 8769 7463
rect 8803 7460 8815 7463
rect 11054 7460 11060 7472
rect 8803 7432 11060 7460
rect 8803 7429 8815 7432
rect 8757 7423 8815 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 21913 7463 21971 7469
rect 21913 7429 21925 7463
rect 21959 7460 21971 7463
rect 22370 7460 22376 7472
rect 21959 7432 22376 7460
rect 21959 7429 21971 7432
rect 21913 7423 21971 7429
rect 22370 7420 22376 7432
rect 22428 7420 22434 7472
rect 3326 7392 3332 7404
rect 3287 7364 3332 7392
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 4338 7392 4344 7404
rect 4299 7364 4344 7392
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 7466 7392 7472 7404
rect 7331 7364 7472 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7392 10011 7395
rect 11146 7392 11152 7404
rect 9999 7364 11152 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7361 11299 7395
rect 11241 7355 11299 7361
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6362 7324 6368 7336
rect 5951 7296 6368 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 8846 7324 8852 7336
rect 8807 7296 8852 7324
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 11054 7324 11060 7336
rect 11015 7296 11060 7324
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 11256 7256 11284 7355
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 13446 7392 13452 7404
rect 12492 7364 12537 7392
rect 13407 7364 13452 7392
rect 12492 7352 12498 7364
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 14826 7392 14832 7404
rect 14787 7364 14832 7392
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 13044 7296 13553 7324
rect 13044 7284 13050 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 13541 7287 13599 7293
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 15856 7324 15884 7355
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 16724 7364 19073 7392
rect 16724 7352 16730 7364
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 20438 7392 20444 7404
rect 20399 7364 20444 7392
rect 19061 7355 19119 7361
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 24854 7392 24860 7404
rect 24815 7364 24860 7392
rect 24854 7352 24860 7364
rect 24912 7352 24918 7404
rect 24964 7392 24992 7500
rect 82998 7488 83004 7540
rect 83056 7528 83062 7540
rect 83826 7528 83832 7540
rect 83056 7500 83832 7528
rect 83056 7488 83062 7500
rect 83826 7488 83832 7500
rect 83884 7488 83890 7540
rect 87782 7528 87788 7540
rect 85408 7500 87788 7528
rect 25406 7420 25412 7472
rect 25464 7460 25470 7472
rect 25464 7432 32904 7460
rect 25464 7420 25470 7432
rect 25869 7395 25927 7401
rect 25869 7392 25881 7395
rect 24964 7364 25881 7392
rect 25869 7361 25881 7364
rect 25915 7361 25927 7395
rect 29454 7392 29460 7404
rect 29415 7364 29460 7392
rect 25869 7355 25927 7361
rect 29454 7352 29460 7364
rect 29512 7352 29518 7404
rect 30469 7395 30527 7401
rect 30469 7392 30481 7395
rect 29564 7364 30481 7392
rect 13780 7296 15884 7324
rect 15933 7327 15991 7333
rect 13780 7284 13786 7296
rect 15933 7293 15945 7327
rect 15979 7293 15991 7327
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 15933 7287 15991 7293
rect 6972 7228 11284 7256
rect 6972 7216 6978 7228
rect 14182 7216 14188 7268
rect 14240 7256 14246 7268
rect 15948 7256 15976 7287
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 19153 7327 19211 7333
rect 19153 7293 19165 7327
rect 19199 7293 19211 7327
rect 22002 7324 22008 7336
rect 21963 7296 22008 7324
rect 19153 7287 19211 7293
rect 14240 7228 15976 7256
rect 14240 7216 14246 7228
rect 17218 7216 17224 7268
rect 17276 7256 17282 7268
rect 19168 7256 19196 7287
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 25961 7327 26019 7333
rect 25961 7324 25973 7327
rect 22112 7296 25973 7324
rect 17276 7228 19196 7256
rect 17276 7216 17282 7228
rect 20530 7216 20536 7268
rect 20588 7256 20594 7268
rect 22112 7256 22140 7296
rect 25961 7293 25973 7296
rect 26007 7293 26019 7327
rect 25961 7287 26019 7293
rect 20588 7228 22140 7256
rect 20588 7216 20594 7228
rect 24210 7216 24216 7268
rect 24268 7256 24274 7268
rect 29564 7256 29592 7364
rect 30469 7361 30481 7364
rect 30515 7361 30527 7395
rect 31846 7392 31852 7404
rect 31807 7364 31852 7392
rect 30469 7355 30527 7361
rect 31846 7352 31852 7364
rect 31904 7352 31910 7404
rect 32876 7401 32904 7432
rect 41138 7420 41144 7472
rect 41196 7460 41202 7472
rect 47397 7463 47455 7469
rect 47397 7460 47409 7463
rect 41196 7432 47409 7460
rect 41196 7420 41202 7432
rect 47397 7429 47409 7432
rect 47443 7429 47455 7463
rect 47397 7423 47455 7429
rect 51534 7420 51540 7472
rect 51592 7460 51598 7472
rect 51592 7432 52776 7460
rect 51592 7420 51598 7432
rect 32861 7395 32919 7401
rect 32861 7361 32873 7395
rect 32907 7361 32919 7395
rect 32861 7355 32919 7361
rect 33318 7352 33324 7404
rect 33376 7392 33382 7404
rect 37829 7395 37887 7401
rect 37829 7392 37841 7395
rect 33376 7364 37841 7392
rect 33376 7352 33382 7364
rect 37829 7361 37841 7364
rect 37875 7361 37887 7395
rect 41874 7392 41880 7404
rect 41835 7364 41880 7392
rect 37829 7355 37887 7361
rect 41874 7352 41880 7364
rect 41932 7352 41938 7404
rect 43901 7395 43959 7401
rect 43901 7392 43913 7395
rect 41984 7364 43913 7392
rect 30558 7324 30564 7336
rect 30519 7296 30564 7324
rect 30558 7284 30564 7296
rect 30616 7284 30622 7336
rect 32953 7327 33011 7333
rect 32953 7293 32965 7327
rect 32999 7293 33011 7327
rect 32953 7287 33011 7293
rect 36817 7327 36875 7333
rect 36817 7293 36829 7327
rect 36863 7324 36875 7327
rect 37734 7324 37740 7336
rect 36863 7296 37740 7324
rect 36863 7293 36875 7296
rect 36817 7287 36875 7293
rect 24268 7228 29592 7256
rect 24268 7216 24274 7228
rect 23658 7188 23664 7200
rect 23619 7160 23664 7188
rect 23658 7148 23664 7160
rect 23716 7148 23722 7200
rect 27246 7188 27252 7200
rect 27207 7160 27252 7188
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 28534 7148 28540 7200
rect 28592 7188 28598 7200
rect 32968 7188 32996 7287
rect 37734 7284 37740 7296
rect 37792 7284 37798 7336
rect 37918 7324 37924 7336
rect 37879 7296 37924 7324
rect 37918 7284 37924 7296
rect 37976 7284 37982 7336
rect 39942 7284 39948 7336
rect 40000 7324 40006 7336
rect 41984 7324 42012 7364
rect 43901 7361 43913 7364
rect 43947 7361 43959 7395
rect 49234 7392 49240 7404
rect 49195 7364 49240 7392
rect 43901 7355 43959 7361
rect 49234 7352 49240 7364
rect 49292 7352 49298 7404
rect 49326 7352 49332 7404
rect 49384 7392 49390 7404
rect 50249 7395 50307 7401
rect 50249 7392 50261 7395
rect 49384 7364 50261 7392
rect 49384 7352 49390 7364
rect 50249 7361 50261 7364
rect 50295 7361 50307 7395
rect 51718 7392 51724 7404
rect 51679 7364 51724 7392
rect 50249 7355 50307 7361
rect 51718 7352 51724 7364
rect 51776 7352 51782 7404
rect 52748 7401 52776 7432
rect 55214 7420 55220 7472
rect 55272 7460 55278 7472
rect 55401 7463 55459 7469
rect 55401 7460 55413 7463
rect 55272 7432 55413 7460
rect 55272 7420 55278 7432
rect 55401 7429 55413 7432
rect 55447 7429 55459 7463
rect 55401 7423 55459 7429
rect 55674 7420 55680 7472
rect 55732 7460 55738 7472
rect 59725 7463 59783 7469
rect 59725 7460 59737 7463
rect 55732 7432 59737 7460
rect 55732 7420 55738 7432
rect 59725 7429 59737 7432
rect 59771 7429 59783 7463
rect 59725 7423 59783 7429
rect 63402 7420 63408 7472
rect 63460 7460 63466 7472
rect 64601 7463 64659 7469
rect 64601 7460 64613 7463
rect 63460 7432 64613 7460
rect 63460 7420 63466 7432
rect 64601 7429 64613 7432
rect 64647 7429 64659 7463
rect 64601 7423 64659 7429
rect 68462 7420 68468 7472
rect 68520 7460 68526 7472
rect 70213 7463 70271 7469
rect 70213 7460 70225 7463
rect 68520 7432 70225 7460
rect 68520 7420 68526 7432
rect 70213 7429 70225 7432
rect 70259 7429 70271 7463
rect 70213 7423 70271 7429
rect 80698 7420 80704 7472
rect 80756 7460 80762 7472
rect 81345 7463 81403 7469
rect 81345 7460 81357 7463
rect 80756 7432 81357 7460
rect 80756 7420 80762 7432
rect 81345 7429 81357 7432
rect 81391 7429 81403 7463
rect 81345 7423 81403 7429
rect 52733 7395 52791 7401
rect 52733 7361 52745 7395
rect 52779 7361 52791 7395
rect 54110 7392 54116 7404
rect 54071 7364 54116 7392
rect 52733 7355 52791 7361
rect 54110 7352 54116 7364
rect 54168 7352 54174 7404
rect 59354 7392 59360 7404
rect 58360 7364 59360 7392
rect 42886 7324 42892 7336
rect 40000 7296 42012 7324
rect 42847 7296 42892 7324
rect 40000 7284 40006 7296
rect 42886 7284 42892 7296
rect 42944 7284 42950 7336
rect 44453 7327 44511 7333
rect 44453 7293 44465 7327
rect 44499 7324 44511 7327
rect 45370 7324 45376 7336
rect 44499 7296 45376 7324
rect 44499 7293 44511 7296
rect 44453 7287 44511 7293
rect 45370 7284 45376 7296
rect 45428 7284 45434 7336
rect 46106 7324 46112 7336
rect 46067 7296 46112 7324
rect 46106 7284 46112 7296
rect 46164 7284 46170 7336
rect 47213 7327 47271 7333
rect 47213 7293 47225 7327
rect 47259 7293 47271 7327
rect 50338 7324 50344 7336
rect 50299 7296 50344 7324
rect 47213 7287 47271 7293
rect 43070 7216 43076 7268
rect 43128 7256 43134 7268
rect 47228 7256 47256 7287
rect 50338 7284 50344 7296
rect 50396 7284 50402 7336
rect 51810 7284 51816 7336
rect 51868 7324 51874 7336
rect 52825 7327 52883 7333
rect 52825 7324 52837 7327
rect 51868 7296 52837 7324
rect 51868 7284 51874 7296
rect 52825 7293 52837 7296
rect 52871 7293 52883 7327
rect 55582 7324 55588 7336
rect 55543 7296 55588 7324
rect 52825 7287 52883 7293
rect 55582 7284 55588 7296
rect 55640 7284 55646 7336
rect 58360 7333 58388 7364
rect 59354 7352 59360 7364
rect 59412 7352 59418 7404
rect 59446 7352 59452 7404
rect 59504 7392 59510 7404
rect 62666 7392 62672 7404
rect 59504 7364 60228 7392
rect 59504 7352 59510 7364
rect 58345 7327 58403 7333
rect 58345 7293 58357 7327
rect 58391 7293 58403 7327
rect 58345 7287 58403 7293
rect 58434 7284 58440 7336
rect 58492 7324 58498 7336
rect 60200 7333 60228 7364
rect 61396 7364 62672 7392
rect 61396 7333 61424 7364
rect 62666 7352 62672 7364
rect 62724 7352 62730 7404
rect 62942 7352 62948 7404
rect 63000 7392 63006 7404
rect 63000 7364 63540 7392
rect 63000 7352 63006 7364
rect 58805 7327 58863 7333
rect 58492 7296 58537 7324
rect 58492 7284 58498 7296
rect 58805 7293 58817 7327
rect 58851 7324 58863 7327
rect 59909 7327 59967 7333
rect 58851 7296 59492 7324
rect 58851 7293 58863 7296
rect 58805 7287 58863 7293
rect 43128 7228 47256 7256
rect 43128 7216 43134 7228
rect 28592 7160 32996 7188
rect 59464 7188 59492 7296
rect 59909 7293 59921 7327
rect 59955 7324 59967 7327
rect 60185 7327 60243 7333
rect 59955 7296 60136 7324
rect 59955 7293 59967 7296
rect 59909 7287 59967 7293
rect 60108 7256 60136 7296
rect 60185 7293 60197 7327
rect 60231 7293 60243 7327
rect 60185 7287 60243 7293
rect 61381 7327 61439 7333
rect 61381 7293 61393 7327
rect 61427 7293 61439 7327
rect 61562 7324 61568 7336
rect 61523 7296 61568 7324
rect 61381 7287 61439 7293
rect 61562 7284 61568 7296
rect 61620 7284 61626 7336
rect 61933 7327 61991 7333
rect 61933 7293 61945 7327
rect 61979 7324 61991 7327
rect 62482 7324 62488 7336
rect 61979 7296 62488 7324
rect 61979 7293 61991 7296
rect 61933 7287 61991 7293
rect 62482 7284 62488 7296
rect 62540 7284 62546 7336
rect 63129 7327 63187 7333
rect 63129 7293 63141 7327
rect 63175 7293 63187 7327
rect 63310 7324 63316 7336
rect 63271 7296 63316 7324
rect 63129 7287 63187 7293
rect 63144 7256 63172 7287
rect 63310 7284 63316 7296
rect 63368 7284 63374 7336
rect 63512 7333 63540 7364
rect 68554 7352 68560 7404
rect 68612 7392 68618 7404
rect 73982 7392 73988 7404
rect 68612 7364 70716 7392
rect 68612 7352 68618 7364
rect 63497 7327 63555 7333
rect 63497 7293 63509 7327
rect 63543 7293 63555 7327
rect 64782 7324 64788 7336
rect 64743 7296 64788 7324
rect 63497 7287 63555 7293
rect 64782 7284 64788 7296
rect 64840 7284 64846 7336
rect 65058 7324 65064 7336
rect 65019 7296 65064 7324
rect 65058 7284 65064 7296
rect 65116 7284 65122 7336
rect 68830 7324 68836 7336
rect 68791 7296 68836 7324
rect 68830 7284 68836 7296
rect 68888 7284 68894 7336
rect 68922 7284 68928 7336
rect 68980 7324 68986 7336
rect 69109 7327 69167 7333
rect 68980 7296 69025 7324
rect 68980 7284 68986 7296
rect 69109 7293 69121 7327
rect 69155 7293 69167 7327
rect 69109 7287 69167 7293
rect 70305 7327 70363 7333
rect 70305 7293 70317 7327
rect 70351 7324 70363 7327
rect 70486 7324 70492 7336
rect 70351 7296 70492 7324
rect 70351 7293 70363 7296
rect 70305 7287 70363 7293
rect 66073 7259 66131 7265
rect 66073 7256 66085 7259
rect 60108 7228 60412 7256
rect 63144 7228 66085 7256
rect 60274 7188 60280 7200
rect 59464 7160 60280 7188
rect 28592 7148 28598 7160
rect 60274 7148 60280 7160
rect 60332 7148 60338 7200
rect 60384 7188 60412 7228
rect 66073 7225 66085 7228
rect 66119 7225 66131 7259
rect 66073 7219 66131 7225
rect 66254 7216 66260 7268
rect 66312 7256 66318 7268
rect 69124 7256 69152 7287
rect 70486 7284 70492 7296
rect 70544 7284 70550 7336
rect 70688 7333 70716 7364
rect 72804 7364 73988 7392
rect 72804 7333 72832 7364
rect 73982 7352 73988 7364
rect 74040 7352 74046 7404
rect 76374 7392 76380 7404
rect 74736 7364 76380 7392
rect 70673 7327 70731 7333
rect 70673 7293 70685 7327
rect 70719 7293 70731 7327
rect 70673 7287 70731 7293
rect 72789 7327 72847 7333
rect 72789 7293 72801 7327
rect 72835 7293 72847 7327
rect 72789 7287 72847 7293
rect 72881 7327 72939 7333
rect 72881 7293 72893 7327
rect 72927 7324 72939 7327
rect 72970 7324 72976 7336
rect 72927 7296 72976 7324
rect 72927 7293 72939 7296
rect 72881 7287 72939 7293
rect 72970 7284 72976 7296
rect 73028 7284 73034 7336
rect 73249 7327 73307 7333
rect 73249 7293 73261 7327
rect 73295 7324 73307 7327
rect 74626 7324 74632 7336
rect 73295 7296 74632 7324
rect 73295 7293 73307 7296
rect 73249 7287 73307 7293
rect 74626 7284 74632 7296
rect 74684 7284 74690 7336
rect 74736 7333 74764 7364
rect 76374 7352 76380 7364
rect 76432 7352 76438 7404
rect 81158 7352 81164 7404
rect 81216 7392 81222 7404
rect 81216 7364 81848 7392
rect 81216 7352 81222 7364
rect 74721 7327 74779 7333
rect 74721 7293 74733 7327
rect 74767 7293 74779 7327
rect 74902 7324 74908 7336
rect 74863 7296 74908 7324
rect 74721 7287 74779 7293
rect 74902 7284 74908 7296
rect 74960 7284 74966 7336
rect 75273 7327 75331 7333
rect 75273 7293 75285 7327
rect 75319 7324 75331 7327
rect 76742 7324 76748 7336
rect 75319 7296 76748 7324
rect 75319 7293 75331 7296
rect 75273 7287 75331 7293
rect 76742 7284 76748 7296
rect 76800 7284 76806 7336
rect 77849 7327 77907 7333
rect 77849 7293 77861 7327
rect 77895 7293 77907 7327
rect 77849 7287 77907 7293
rect 66312 7228 69152 7256
rect 77864 7256 77892 7287
rect 77938 7284 77944 7336
rect 77996 7324 78002 7336
rect 78309 7327 78367 7333
rect 77996 7296 78041 7324
rect 77996 7284 78002 7296
rect 78309 7293 78321 7327
rect 78355 7324 78367 7327
rect 78582 7324 78588 7336
rect 78355 7296 78588 7324
rect 78355 7293 78367 7296
rect 78309 7287 78367 7293
rect 78582 7284 78588 7296
rect 78640 7284 78646 7336
rect 81526 7324 81532 7336
rect 81487 7296 81532 7324
rect 81526 7284 81532 7296
rect 81584 7284 81590 7336
rect 81820 7333 81848 7364
rect 81805 7327 81863 7333
rect 81805 7293 81817 7327
rect 81851 7293 81863 7327
rect 81805 7287 81863 7293
rect 82817 7327 82875 7333
rect 82817 7293 82829 7327
rect 82863 7293 82875 7327
rect 83182 7324 83188 7336
rect 83143 7296 83188 7324
rect 82817 7287 82875 7293
rect 79781 7259 79839 7265
rect 79781 7256 79793 7259
rect 77864 7228 79793 7256
rect 66312 7216 66318 7228
rect 79781 7225 79793 7228
rect 79827 7225 79839 7259
rect 79781 7219 79839 7225
rect 81342 7216 81348 7268
rect 81400 7256 81406 7268
rect 82832 7256 82860 7287
rect 83182 7284 83188 7296
rect 83240 7284 83246 7336
rect 83553 7327 83611 7333
rect 83553 7293 83565 7327
rect 83599 7324 83611 7327
rect 85408 7324 85436 7500
rect 87782 7488 87788 7500
rect 87840 7488 87846 7540
rect 99466 7528 99472 7540
rect 89640 7500 99472 7528
rect 87322 7460 87328 7472
rect 86144 7432 87328 7460
rect 85574 7324 85580 7336
rect 83599 7296 85436 7324
rect 85535 7296 85580 7324
rect 83599 7293 83611 7296
rect 83553 7287 83611 7293
rect 85574 7284 85580 7296
rect 85632 7284 85638 7336
rect 85761 7327 85819 7333
rect 85761 7293 85773 7327
rect 85807 7324 85819 7327
rect 85850 7324 85856 7336
rect 85807 7296 85856 7324
rect 85807 7293 85819 7296
rect 85761 7287 85819 7293
rect 85850 7284 85856 7296
rect 85908 7284 85914 7336
rect 86144 7333 86172 7432
rect 87322 7420 87328 7432
rect 87380 7420 87386 7472
rect 89254 7392 89260 7404
rect 87156 7364 89260 7392
rect 87156 7333 87184 7364
rect 89254 7352 89260 7364
rect 89312 7352 89318 7404
rect 86129 7327 86187 7333
rect 86129 7293 86141 7327
rect 86175 7293 86187 7327
rect 86129 7287 86187 7293
rect 87141 7327 87199 7333
rect 87141 7293 87153 7327
rect 87187 7293 87199 7327
rect 87322 7324 87328 7336
rect 87283 7296 87328 7324
rect 87141 7287 87199 7293
rect 87322 7284 87328 7296
rect 87380 7284 87386 7336
rect 89640 7333 89668 7500
rect 99466 7488 99472 7500
rect 99524 7488 99530 7540
rect 101953 7531 102011 7537
rect 101953 7497 101965 7531
rect 101999 7528 102011 7531
rect 112162 7528 112168 7540
rect 101999 7500 112168 7528
rect 101999 7497 102011 7500
rect 101953 7491 102011 7497
rect 112162 7488 112168 7500
rect 112220 7488 112226 7540
rect 123202 7528 123208 7540
rect 115216 7500 123208 7528
rect 94498 7420 94504 7472
rect 94556 7460 94562 7472
rect 94593 7463 94651 7469
rect 94593 7460 94605 7463
rect 94556 7432 94605 7460
rect 94556 7420 94562 7432
rect 94593 7429 94605 7432
rect 94639 7429 94651 7463
rect 98270 7460 98276 7472
rect 94593 7423 94651 7429
rect 94792 7432 98276 7460
rect 89717 7395 89775 7401
rect 89717 7361 89729 7395
rect 89763 7392 89775 7395
rect 90082 7392 90088 7404
rect 89763 7364 90088 7392
rect 89763 7361 89775 7364
rect 89717 7355 89775 7361
rect 90082 7352 90088 7364
rect 90140 7352 90146 7404
rect 94222 7392 94228 7404
rect 90928 7364 94228 7392
rect 87693 7327 87751 7333
rect 87693 7293 87705 7327
rect 87739 7293 87751 7327
rect 87693 7287 87751 7293
rect 89625 7327 89683 7333
rect 89625 7293 89637 7327
rect 89671 7293 89683 7327
rect 89625 7287 89683 7293
rect 89993 7327 90051 7333
rect 89993 7293 90005 7327
rect 90039 7324 90051 7327
rect 90928 7324 90956 7364
rect 94222 7352 94228 7364
rect 94280 7352 94286 7404
rect 90039 7296 90956 7324
rect 91281 7327 91339 7333
rect 90039 7293 90051 7296
rect 89993 7287 90051 7293
rect 91281 7293 91293 7327
rect 91327 7293 91339 7327
rect 91281 7287 91339 7293
rect 91373 7327 91431 7333
rect 91373 7293 91385 7327
rect 91419 7324 91431 7327
rect 91462 7324 91468 7336
rect 91419 7296 91468 7324
rect 91419 7293 91431 7296
rect 91373 7287 91431 7293
rect 81400 7228 82860 7256
rect 87708 7256 87736 7287
rect 91186 7256 91192 7268
rect 87708 7228 91192 7256
rect 81400 7216 81406 7228
rect 91186 7216 91192 7228
rect 91244 7216 91250 7268
rect 64690 7188 64696 7200
rect 60384 7160 64696 7188
rect 64690 7148 64696 7160
rect 64748 7148 64754 7200
rect 66346 7148 66352 7200
rect 66404 7188 66410 7200
rect 67085 7191 67143 7197
rect 67085 7188 67097 7191
rect 66404 7160 67097 7188
rect 66404 7148 66410 7160
rect 67085 7157 67097 7160
rect 67131 7157 67143 7191
rect 67085 7151 67143 7157
rect 74534 7148 74540 7200
rect 74592 7188 74598 7200
rect 76101 7191 76159 7197
rect 76101 7188 76113 7191
rect 74592 7160 76113 7188
rect 74592 7148 74598 7160
rect 76101 7157 76113 7160
rect 76147 7157 76159 7191
rect 91296 7188 91324 7287
rect 91462 7284 91468 7296
rect 91520 7284 91526 7336
rect 91738 7324 91744 7336
rect 91699 7296 91744 7324
rect 91738 7284 91744 7296
rect 91796 7284 91802 7336
rect 92753 7327 92811 7333
rect 92753 7293 92765 7327
rect 92799 7293 92811 7327
rect 92753 7287 92811 7293
rect 92768 7256 92796 7287
rect 92842 7284 92848 7336
rect 92900 7324 92906 7336
rect 92937 7327 92995 7333
rect 92937 7324 92949 7327
rect 92900 7296 92949 7324
rect 92900 7284 92906 7296
rect 92937 7293 92949 7296
rect 92983 7293 92995 7327
rect 93302 7324 93308 7336
rect 93263 7296 93308 7324
rect 92937 7287 92995 7293
rect 93302 7284 93308 7296
rect 93360 7284 93366 7336
rect 94792 7333 94820 7432
rect 98270 7420 98276 7432
rect 98328 7420 98334 7472
rect 98454 7460 98460 7472
rect 98415 7432 98460 7460
rect 98454 7420 98460 7432
rect 98512 7420 98518 7472
rect 102778 7420 102784 7472
rect 102836 7460 102842 7472
rect 102873 7463 102931 7469
rect 102873 7460 102885 7463
rect 102836 7432 102885 7460
rect 102836 7420 102842 7432
rect 102873 7429 102885 7432
rect 102919 7429 102931 7463
rect 105998 7460 106004 7472
rect 102873 7423 102931 7429
rect 103532 7432 106004 7460
rect 96890 7352 96896 7404
rect 96948 7392 96954 7404
rect 96985 7395 97043 7401
rect 96985 7392 96997 7395
rect 96948 7364 96997 7392
rect 96948 7352 96954 7364
rect 96985 7361 96997 7364
rect 97031 7361 97043 7395
rect 99650 7392 99656 7404
rect 96985 7355 97043 7361
rect 98288 7364 99656 7392
rect 94777 7327 94835 7333
rect 94777 7293 94789 7327
rect 94823 7293 94835 7327
rect 94777 7287 94835 7293
rect 95145 7327 95203 7333
rect 95145 7293 95157 7327
rect 95191 7324 95203 7327
rect 95786 7324 95792 7336
rect 95191 7296 95792 7324
rect 95191 7293 95203 7296
rect 95145 7287 95203 7293
rect 95786 7284 95792 7296
rect 95844 7284 95850 7336
rect 96154 7284 96160 7336
rect 96212 7324 96218 7336
rect 98178 7324 98184 7336
rect 96212 7296 98184 7324
rect 96212 7284 96218 7296
rect 98178 7284 98184 7296
rect 98236 7284 98242 7336
rect 98288 7256 98316 7364
rect 99650 7352 99656 7364
rect 99708 7352 99714 7404
rect 99745 7395 99803 7401
rect 99745 7361 99757 7395
rect 99791 7392 99803 7395
rect 100754 7392 100760 7404
rect 99791 7364 100760 7392
rect 99791 7361 99803 7364
rect 99745 7355 99803 7361
rect 100754 7352 100760 7364
rect 100812 7352 100818 7404
rect 100938 7392 100944 7404
rect 100899 7364 100944 7392
rect 100938 7352 100944 7364
rect 100996 7352 101002 7404
rect 98549 7327 98607 7333
rect 98549 7293 98561 7327
rect 98595 7293 98607 7327
rect 99374 7324 99380 7336
rect 99335 7296 99380 7324
rect 98549 7287 98607 7293
rect 92768 7228 98316 7256
rect 98564 7256 98592 7287
rect 99374 7284 99380 7296
rect 99432 7284 99438 7336
rect 100113 7327 100171 7333
rect 100113 7293 100125 7327
rect 100159 7324 100171 7327
rect 100386 7324 100392 7336
rect 100159 7296 100392 7324
rect 100159 7293 100171 7296
rect 100113 7287 100171 7293
rect 100386 7284 100392 7296
rect 100444 7284 100450 7336
rect 101490 7284 101496 7336
rect 101548 7324 101554 7336
rect 103532 7333 103560 7432
rect 105998 7420 106004 7432
rect 106056 7420 106062 7472
rect 107838 7420 107844 7472
rect 107896 7460 107902 7472
rect 107933 7463 107991 7469
rect 107933 7460 107945 7463
rect 107896 7432 107945 7460
rect 107896 7420 107902 7432
rect 107933 7429 107945 7432
rect 107979 7429 107991 7463
rect 107933 7423 107991 7429
rect 108022 7420 108028 7472
rect 108080 7460 108086 7472
rect 111058 7460 111064 7472
rect 108080 7432 111064 7460
rect 108080 7420 108086 7432
rect 111058 7420 111064 7432
rect 111116 7420 111122 7472
rect 104066 7352 104072 7404
rect 104124 7392 104130 7404
rect 109402 7392 109408 7404
rect 104124 7364 109408 7392
rect 104124 7352 104130 7364
rect 109402 7352 109408 7364
rect 109460 7352 109466 7404
rect 109678 7392 109684 7404
rect 109639 7364 109684 7392
rect 109678 7352 109684 7364
rect 109736 7352 109742 7404
rect 111153 7395 111211 7401
rect 111153 7361 111165 7395
rect 111199 7361 111211 7395
rect 112070 7392 112076 7404
rect 112031 7364 112076 7392
rect 111153 7355 111211 7361
rect 102781 7327 102839 7333
rect 102781 7324 102793 7327
rect 101548 7296 102793 7324
rect 101548 7284 101554 7296
rect 102781 7293 102793 7296
rect 102827 7293 102839 7327
rect 102781 7287 102839 7293
rect 103517 7327 103575 7333
rect 103517 7293 103529 7327
rect 103563 7293 103575 7327
rect 103517 7287 103575 7293
rect 103606 7284 103612 7336
rect 103664 7324 103670 7336
rect 104345 7327 104403 7333
rect 104345 7324 104357 7327
rect 103664 7296 104357 7324
rect 103664 7284 103670 7296
rect 104345 7293 104357 7296
rect 104391 7293 104403 7327
rect 104345 7287 104403 7293
rect 104713 7327 104771 7333
rect 104713 7293 104725 7327
rect 104759 7293 104771 7327
rect 104713 7287 104771 7293
rect 105081 7327 105139 7333
rect 105081 7293 105093 7327
rect 105127 7293 105139 7327
rect 105906 7324 105912 7336
rect 105867 7296 105912 7324
rect 105081 7287 105139 7293
rect 101953 7259 102011 7265
rect 101953 7256 101965 7259
rect 98564 7228 101965 7256
rect 101953 7225 101965 7228
rect 101999 7225 102011 7259
rect 101953 7219 102011 7225
rect 99466 7188 99472 7200
rect 91296 7160 99472 7188
rect 76101 7151 76159 7157
rect 99466 7148 99472 7160
rect 99524 7148 99530 7200
rect 102226 7148 102232 7200
rect 102284 7188 102290 7200
rect 104728 7188 104756 7287
rect 105096 7256 105124 7287
rect 105906 7284 105912 7296
rect 105964 7284 105970 7336
rect 106277 7327 106335 7333
rect 106277 7293 106289 7327
rect 106323 7324 106335 7327
rect 106366 7324 106372 7336
rect 106323 7296 106372 7324
rect 106323 7293 106335 7296
rect 106277 7287 106335 7293
rect 106366 7284 106372 7296
rect 106424 7284 106430 7336
rect 106645 7327 106703 7333
rect 106645 7293 106657 7327
rect 106691 7293 106703 7327
rect 108114 7324 108120 7336
rect 108075 7296 108120 7324
rect 106645 7287 106703 7293
rect 106458 7256 106464 7268
rect 105096 7228 106464 7256
rect 106458 7216 106464 7228
rect 106516 7216 106522 7268
rect 106660 7256 106688 7287
rect 108114 7284 108120 7296
rect 108172 7284 108178 7336
rect 108577 7327 108635 7333
rect 108577 7293 108589 7327
rect 108623 7324 108635 7327
rect 109862 7324 109868 7336
rect 108623 7296 109868 7324
rect 108623 7293 108635 7296
rect 108577 7287 108635 7293
rect 109862 7284 109868 7296
rect 109920 7284 109926 7336
rect 110506 7256 110512 7268
rect 106660 7228 110512 7256
rect 110506 7216 110512 7228
rect 110564 7216 110570 7268
rect 111168 7256 111196 7355
rect 112070 7352 112076 7364
rect 112128 7352 112134 7404
rect 113450 7352 113456 7404
rect 113508 7392 113514 7404
rect 113729 7395 113787 7401
rect 113729 7392 113741 7395
rect 113508 7364 113741 7392
rect 113508 7352 113514 7364
rect 113729 7361 113741 7364
rect 113775 7361 113787 7395
rect 113729 7355 113787 7361
rect 113910 7352 113916 7404
rect 113968 7392 113974 7404
rect 114370 7392 114376 7404
rect 113968 7364 114376 7392
rect 113968 7352 113974 7364
rect 114370 7352 114376 7364
rect 114428 7352 114434 7404
rect 115216 7401 115244 7500
rect 123202 7488 123208 7500
rect 123260 7488 123266 7540
rect 132586 7528 132592 7540
rect 123312 7500 132592 7528
rect 123312 7460 123340 7500
rect 132586 7488 132592 7500
rect 132644 7488 132650 7540
rect 133966 7488 133972 7540
rect 134024 7528 134030 7540
rect 134024 7500 142476 7528
rect 134024 7488 134030 7500
rect 117884 7432 123340 7460
rect 115201 7395 115259 7401
rect 115201 7361 115213 7395
rect 115247 7361 115259 7395
rect 116578 7392 116584 7404
rect 116539 7364 116584 7392
rect 115201 7355 115259 7361
rect 116578 7352 116584 7364
rect 116636 7352 116642 7404
rect 111245 7327 111303 7333
rect 111245 7293 111257 7327
rect 111291 7324 111303 7327
rect 111702 7324 111708 7336
rect 111291 7296 111708 7324
rect 111291 7293 111303 7296
rect 111245 7287 111303 7293
rect 111702 7284 111708 7296
rect 111760 7284 111766 7336
rect 115290 7324 115296 7336
rect 115251 7296 115296 7324
rect 115290 7284 115296 7296
rect 115348 7284 115354 7336
rect 117884 7256 117912 7432
rect 124766 7420 124772 7472
rect 124824 7460 124830 7472
rect 126054 7460 126060 7472
rect 124824 7432 126060 7460
rect 124824 7420 124830 7432
rect 126054 7420 126060 7432
rect 126112 7420 126118 7472
rect 130105 7463 130163 7469
rect 130105 7460 130117 7463
rect 127544 7432 130117 7460
rect 118050 7392 118056 7404
rect 118011 7364 118056 7392
rect 118050 7352 118056 7364
rect 118108 7352 118114 7404
rect 122101 7395 122159 7401
rect 122101 7361 122113 7395
rect 122147 7392 122159 7395
rect 127544 7392 127572 7432
rect 130105 7429 130117 7432
rect 130151 7429 130163 7463
rect 134702 7460 134708 7472
rect 130105 7423 130163 7429
rect 130212 7432 134708 7460
rect 127710 7392 127716 7404
rect 122147 7364 127572 7392
rect 127671 7364 127716 7392
rect 122147 7361 122159 7364
rect 122101 7355 122159 7361
rect 127710 7352 127716 7364
rect 127768 7352 127774 7404
rect 118145 7327 118203 7333
rect 118145 7293 118157 7327
rect 118191 7293 118203 7327
rect 118145 7287 118203 7293
rect 119525 7327 119583 7333
rect 119525 7293 119537 7327
rect 119571 7324 119583 7327
rect 120629 7327 120687 7333
rect 120629 7324 120641 7327
rect 119571 7296 120641 7324
rect 119571 7293 119583 7296
rect 119525 7287 119583 7293
rect 120629 7293 120641 7296
rect 120675 7293 120687 7327
rect 120629 7287 120687 7293
rect 111168 7228 117912 7256
rect 118160 7256 118188 7287
rect 121546 7284 121552 7336
rect 121604 7324 121610 7336
rect 121733 7327 121791 7333
rect 121733 7324 121745 7327
rect 121604 7296 121745 7324
rect 121604 7284 121610 7296
rect 121733 7293 121745 7296
rect 121779 7293 121791 7327
rect 121733 7287 121791 7293
rect 126146 7284 126152 7336
rect 126204 7324 126210 7336
rect 126241 7327 126299 7333
rect 126241 7324 126253 7327
rect 126204 7296 126253 7324
rect 126204 7284 126210 7296
rect 126241 7293 126253 7296
rect 126287 7293 126299 7327
rect 127802 7324 127808 7336
rect 127763 7296 127808 7324
rect 126241 7287 126299 7293
rect 127802 7284 127808 7296
rect 127860 7284 127866 7336
rect 130212 7324 130240 7432
rect 134702 7420 134708 7432
rect 134760 7420 134766 7472
rect 134812 7432 135024 7460
rect 132773 7395 132831 7401
rect 132773 7361 132785 7395
rect 132819 7392 132831 7395
rect 134812 7392 134840 7432
rect 132819 7364 134840 7392
rect 132819 7361 132831 7364
rect 132773 7355 132831 7361
rect 130028 7296 130240 7324
rect 131301 7327 131359 7333
rect 120994 7256 121000 7268
rect 118160 7228 121000 7256
rect 120994 7216 121000 7228
rect 121052 7216 121058 7268
rect 124214 7216 124220 7268
rect 124272 7256 124278 7268
rect 130028 7256 130056 7296
rect 131301 7293 131313 7327
rect 131347 7293 131359 7327
rect 131301 7287 131359 7293
rect 132865 7327 132923 7333
rect 132865 7293 132877 7327
rect 132911 7324 132923 7327
rect 133046 7324 133052 7336
rect 132911 7296 133052 7324
rect 132911 7293 132923 7296
rect 132865 7287 132923 7293
rect 124272 7228 130056 7256
rect 130105 7259 130163 7265
rect 124272 7216 124278 7228
rect 130105 7225 130117 7259
rect 130151 7256 130163 7259
rect 131316 7256 131344 7287
rect 133046 7284 133052 7296
rect 133104 7284 133110 7336
rect 133138 7284 133144 7336
rect 133196 7324 133202 7336
rect 134610 7324 134616 7336
rect 133196 7296 134616 7324
rect 133196 7284 133202 7296
rect 134610 7284 134616 7296
rect 134668 7284 134674 7336
rect 134996 7324 135024 7432
rect 135162 7420 135168 7472
rect 135220 7460 135226 7472
rect 137186 7460 137192 7472
rect 135220 7432 137192 7460
rect 135220 7420 135226 7432
rect 137186 7420 137192 7432
rect 137244 7420 137250 7472
rect 137370 7460 137376 7472
rect 137331 7432 137376 7460
rect 137370 7420 137376 7432
rect 137428 7420 137434 7472
rect 137462 7420 137468 7472
rect 137520 7460 137526 7472
rect 140314 7460 140320 7472
rect 137520 7432 140320 7460
rect 137520 7420 137526 7432
rect 140314 7420 140320 7432
rect 140372 7420 140378 7472
rect 140498 7460 140504 7472
rect 140459 7432 140504 7460
rect 140498 7420 140504 7432
rect 140556 7420 140562 7472
rect 142448 7460 142476 7500
rect 142522 7488 142528 7540
rect 142580 7528 142586 7540
rect 156782 7528 156788 7540
rect 142580 7500 156788 7528
rect 142580 7488 142586 7500
rect 156782 7488 156788 7500
rect 156840 7488 156846 7540
rect 157521 7531 157579 7537
rect 157521 7497 157533 7531
rect 157567 7528 157579 7531
rect 157567 7500 157840 7528
rect 157567 7497 157579 7500
rect 157521 7491 157579 7497
rect 140608 7432 142384 7460
rect 142448 7432 150020 7460
rect 136726 7352 136732 7404
rect 136784 7392 136790 7404
rect 140608 7392 140636 7432
rect 142246 7392 142252 7404
rect 136784 7364 140636 7392
rect 142207 7364 142252 7392
rect 136784 7352 136790 7364
rect 142246 7352 142252 7364
rect 142304 7352 142310 7404
rect 142356 7392 142384 7432
rect 142522 7392 142528 7404
rect 142356 7364 142528 7392
rect 142522 7352 142528 7364
rect 142580 7352 142586 7404
rect 143442 7392 143448 7404
rect 143403 7364 143448 7392
rect 143442 7352 143448 7364
rect 143500 7352 143506 7404
rect 145926 7392 145932 7404
rect 145887 7364 145932 7392
rect 145926 7352 145932 7364
rect 145984 7352 145990 7404
rect 148962 7392 148968 7404
rect 148923 7364 148968 7392
rect 148962 7352 148968 7364
rect 149020 7352 149026 7404
rect 149992 7392 150020 7432
rect 150066 7420 150072 7472
rect 150124 7460 150130 7472
rect 150124 7432 153976 7460
rect 150124 7420 150130 7432
rect 151722 7392 151728 7404
rect 149992 7364 151492 7392
rect 151683 7364 151728 7392
rect 135806 7324 135812 7336
rect 134996 7296 135812 7324
rect 135806 7284 135812 7296
rect 135864 7284 135870 7336
rect 135901 7327 135959 7333
rect 135901 7293 135913 7327
rect 135947 7293 135959 7327
rect 137002 7324 137008 7336
rect 136963 7296 137008 7324
rect 135901 7287 135959 7293
rect 133874 7256 133880 7268
rect 130151 7228 130424 7256
rect 131316 7228 133880 7256
rect 130151 7225 130163 7228
rect 130105 7219 130163 7225
rect 102284 7160 104756 7188
rect 102284 7148 102290 7160
rect 104802 7148 104808 7200
rect 104860 7188 104866 7200
rect 109310 7188 109316 7200
rect 104860 7160 109316 7188
rect 104860 7148 104866 7160
rect 109310 7148 109316 7160
rect 109368 7148 109374 7200
rect 109402 7148 109408 7200
rect 109460 7188 109466 7200
rect 111334 7188 111340 7200
rect 109460 7160 111340 7188
rect 109460 7148 109466 7160
rect 111334 7148 111340 7160
rect 111392 7148 111398 7200
rect 120074 7148 120080 7200
rect 120132 7188 120138 7200
rect 120810 7188 120816 7200
rect 120132 7160 120816 7188
rect 120132 7148 120138 7160
rect 120810 7148 120816 7160
rect 120868 7148 120874 7200
rect 123573 7191 123631 7197
rect 123573 7157 123585 7191
rect 123619 7188 123631 7191
rect 125042 7188 125048 7200
rect 123619 7160 125048 7188
rect 123619 7157 123631 7160
rect 123573 7151 123631 7157
rect 125042 7148 125048 7160
rect 125100 7148 125106 7200
rect 125226 7188 125232 7200
rect 125187 7160 125232 7188
rect 125226 7148 125232 7160
rect 125284 7148 125290 7200
rect 126146 7148 126152 7200
rect 126204 7188 126210 7200
rect 127434 7188 127440 7200
rect 126204 7160 127440 7188
rect 126204 7148 126210 7160
rect 127434 7148 127440 7160
rect 127492 7148 127498 7200
rect 128630 7188 128636 7200
rect 128591 7160 128636 7188
rect 128630 7148 128636 7160
rect 128688 7148 128694 7200
rect 130286 7188 130292 7200
rect 130247 7160 130292 7188
rect 130286 7148 130292 7160
rect 130344 7148 130350 7200
rect 130396 7188 130424 7228
rect 133874 7216 133880 7228
rect 133932 7216 133938 7268
rect 134705 7259 134763 7265
rect 134705 7225 134717 7259
rect 134751 7256 134763 7259
rect 135346 7256 135352 7268
rect 134751 7228 135352 7256
rect 134751 7225 134763 7228
rect 134705 7219 134763 7225
rect 135346 7216 135352 7228
rect 135404 7216 135410 7268
rect 135916 7256 135944 7287
rect 137002 7284 137008 7296
rect 137060 7284 137066 7336
rect 137094 7284 137100 7336
rect 137152 7324 137158 7336
rect 138750 7324 138756 7336
rect 137152 7296 138756 7324
rect 137152 7284 137158 7296
rect 138750 7284 138756 7296
rect 138808 7284 138814 7336
rect 139029 7327 139087 7333
rect 139029 7293 139041 7327
rect 139075 7324 139087 7327
rect 140498 7324 140504 7336
rect 139075 7296 140504 7324
rect 139075 7293 139087 7296
rect 139029 7287 139087 7293
rect 140498 7284 140504 7296
rect 140556 7284 140562 7336
rect 140593 7327 140651 7333
rect 140593 7293 140605 7327
rect 140639 7324 140651 7327
rect 141970 7324 141976 7336
rect 140639 7296 141976 7324
rect 140639 7293 140651 7296
rect 140593 7287 140651 7293
rect 141970 7284 141976 7296
rect 142028 7284 142034 7336
rect 143353 7327 143411 7333
rect 143353 7324 143365 7327
rect 142448 7296 143365 7324
rect 139762 7256 139768 7268
rect 135916 7228 139768 7256
rect 139762 7216 139768 7228
rect 139820 7216 139826 7268
rect 141234 7216 141240 7268
rect 141292 7256 141298 7268
rect 142448 7256 142476 7296
rect 143353 7293 143365 7296
rect 143399 7293 143411 7327
rect 143353 7287 143411 7293
rect 147674 7284 147680 7336
rect 147732 7324 147738 7336
rect 148870 7324 148876 7336
rect 147732 7296 147777 7324
rect 148831 7296 148876 7324
rect 147732 7284 147738 7296
rect 148870 7284 148876 7296
rect 148928 7284 148934 7336
rect 150253 7327 150311 7333
rect 150253 7293 150265 7327
rect 150299 7324 150311 7327
rect 150710 7324 150716 7336
rect 150299 7296 150716 7324
rect 150299 7293 150311 7296
rect 150253 7287 150311 7293
rect 150710 7284 150716 7296
rect 150768 7284 150774 7336
rect 151357 7327 151415 7333
rect 151357 7293 151369 7327
rect 151403 7293 151415 7327
rect 151464 7324 151492 7364
rect 151722 7352 151728 7364
rect 151780 7352 151786 7404
rect 152921 7395 152979 7401
rect 152921 7361 152933 7395
rect 152967 7392 152979 7395
rect 153838 7392 153844 7404
rect 152967 7364 153844 7392
rect 152967 7361 152979 7364
rect 152921 7355 152979 7361
rect 153838 7352 153844 7364
rect 153896 7352 153902 7404
rect 153948 7392 153976 7432
rect 157334 7420 157340 7472
rect 157392 7460 157398 7472
rect 157702 7460 157708 7472
rect 157392 7432 157708 7460
rect 157392 7420 157398 7432
rect 157702 7420 157708 7432
rect 157760 7420 157766 7472
rect 157812 7460 157840 7500
rect 158898 7488 158904 7540
rect 158956 7528 158962 7540
rect 158956 7500 181300 7528
rect 158956 7488 158962 7500
rect 160278 7460 160284 7472
rect 157812 7432 160284 7460
rect 160278 7420 160284 7432
rect 160336 7420 160342 7472
rect 162302 7420 162308 7472
rect 162360 7460 162366 7472
rect 180886 7460 180892 7472
rect 162360 7432 180892 7460
rect 162360 7420 162366 7432
rect 180886 7420 180892 7432
rect 180944 7420 180950 7472
rect 181272 7460 181300 7500
rect 181346 7488 181352 7540
rect 181404 7528 181410 7540
rect 187970 7528 187976 7540
rect 181404 7500 187976 7528
rect 181404 7488 181410 7500
rect 187970 7488 187976 7500
rect 188028 7488 188034 7540
rect 188356 7500 188936 7528
rect 184934 7460 184940 7472
rect 181272 7432 184940 7460
rect 184934 7420 184940 7432
rect 184992 7420 184998 7472
rect 161753 7395 161811 7401
rect 161753 7392 161765 7395
rect 153948 7364 161765 7392
rect 161753 7361 161765 7364
rect 161799 7361 161811 7395
rect 161753 7355 161811 7361
rect 161842 7352 161848 7404
rect 161900 7352 161906 7404
rect 161934 7352 161940 7404
rect 161992 7352 161998 7404
rect 162029 7395 162087 7401
rect 162029 7361 162041 7395
rect 162075 7392 162087 7395
rect 181530 7392 181536 7404
rect 162075 7364 181536 7392
rect 162075 7361 162087 7364
rect 162029 7355 162087 7361
rect 181530 7352 181536 7364
rect 181588 7352 181594 7404
rect 181806 7352 181812 7404
rect 181864 7352 181870 7404
rect 181993 7395 182051 7401
rect 181993 7361 182005 7395
rect 182039 7392 182051 7395
rect 182634 7392 182640 7404
rect 182039 7364 182640 7392
rect 182039 7361 182051 7364
rect 181993 7355 182051 7361
rect 182634 7352 182640 7364
rect 182692 7352 182698 7404
rect 182726 7352 182732 7404
rect 182784 7392 182790 7404
rect 188356 7392 188384 7500
rect 188798 7420 188804 7472
rect 188856 7420 188862 7472
rect 182784 7364 188384 7392
rect 182784 7352 182790 7364
rect 156046 7324 156052 7336
rect 151464 7296 156052 7324
rect 151357 7287 151415 7293
rect 141292 7228 142476 7256
rect 141292 7216 141298 7228
rect 142706 7216 142712 7268
rect 142764 7256 142770 7268
rect 144270 7256 144276 7268
rect 142764 7228 144276 7256
rect 142764 7216 142770 7228
rect 144270 7216 144276 7228
rect 144328 7216 144334 7268
rect 150342 7216 150348 7268
rect 150400 7256 150406 7268
rect 151372 7256 151400 7287
rect 156046 7284 156052 7296
rect 156104 7284 156110 7336
rect 157058 7284 157064 7336
rect 157116 7324 157122 7336
rect 161860 7324 161888 7352
rect 157116 7296 161888 7324
rect 161952 7324 161980 7352
rect 181717 7327 181775 7333
rect 181717 7324 181729 7327
rect 161952 7296 181729 7324
rect 157116 7284 157122 7296
rect 181717 7293 181729 7296
rect 181763 7293 181775 7327
rect 181824 7324 181852 7352
rect 188816 7324 188844 7420
rect 188908 7392 188936 7500
rect 189166 7420 189172 7472
rect 189224 7460 189230 7472
rect 196710 7460 196716 7472
rect 189224 7432 196716 7460
rect 189224 7420 189230 7432
rect 196710 7420 196716 7432
rect 196768 7420 196774 7472
rect 196986 7392 196992 7404
rect 188908 7364 196992 7392
rect 196986 7352 196992 7364
rect 197044 7352 197050 7404
rect 181824 7296 188844 7324
rect 181717 7287 181775 7293
rect 150400 7228 151400 7256
rect 150400 7216 150406 7228
rect 133138 7188 133144 7200
rect 130396 7160 133144 7188
rect 133138 7148 133144 7160
rect 133196 7148 133202 7200
rect 133690 7188 133696 7200
rect 133651 7160 133696 7188
rect 133690 7148 133696 7160
rect 133748 7148 133754 7200
rect 133782 7148 133788 7200
rect 133840 7188 133846 7200
rect 144641 7191 144699 7197
rect 144641 7188 144653 7191
rect 133840 7160 144653 7188
rect 133840 7148 133846 7160
rect 144641 7157 144653 7160
rect 144687 7157 144699 7191
rect 144641 7151 144699 7157
rect 1104 7098 154560 7120
rect 1104 7046 24078 7098
rect 24130 7046 64078 7098
rect 64130 7046 104078 7098
rect 104130 7046 144078 7098
rect 144130 7046 154560 7098
rect 1104 7024 154560 7046
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 17681 6987 17739 6993
rect 17681 6984 17693 6987
rect 17000 6956 17693 6984
rect 17000 6944 17006 6956
rect 17681 6953 17693 6956
rect 17727 6953 17739 6987
rect 17681 6947 17739 6953
rect 18046 6944 18052 6996
rect 18104 6984 18110 6996
rect 18693 6987 18751 6993
rect 18693 6984 18705 6987
rect 18104 6956 18705 6984
rect 18104 6944 18110 6956
rect 18693 6953 18705 6956
rect 18739 6953 18751 6987
rect 18693 6947 18751 6953
rect 25314 6944 25320 6996
rect 25372 6984 25378 6996
rect 30558 6984 30564 6996
rect 25372 6956 30564 6984
rect 25372 6944 25378 6956
rect 30558 6944 30564 6956
rect 30616 6944 30622 6996
rect 91738 6944 91744 6996
rect 91796 6984 91802 6996
rect 95878 6984 95884 6996
rect 91796 6956 95884 6984
rect 91796 6944 91802 6956
rect 95878 6944 95884 6956
rect 95936 6944 95942 6996
rect 96522 6944 96528 6996
rect 96580 6984 96586 6996
rect 99374 6984 99380 6996
rect 96580 6956 99380 6984
rect 96580 6944 96586 6956
rect 99374 6944 99380 6956
rect 99432 6944 99438 6996
rect 99466 6944 99472 6996
rect 99524 6984 99530 6996
rect 99524 6956 99569 6984
rect 99524 6944 99530 6956
rect 105630 6944 105636 6996
rect 105688 6984 105694 6996
rect 108022 6984 108028 6996
rect 105688 6956 108028 6984
rect 105688 6944 105694 6956
rect 108022 6944 108028 6956
rect 108080 6944 108086 6996
rect 120166 6944 120172 6996
rect 120224 6984 120230 6996
rect 137462 6984 137468 6996
rect 120224 6956 137468 6984
rect 120224 6944 120230 6956
rect 137462 6944 137468 6956
rect 137520 6944 137526 6996
rect 137922 6944 137928 6996
rect 137980 6984 137986 6996
rect 139578 6984 139584 6996
rect 137980 6956 139584 6984
rect 137980 6944 137986 6956
rect 139578 6944 139584 6956
rect 139636 6944 139642 6996
rect 139762 6984 139768 6996
rect 139723 6956 139768 6984
rect 139762 6944 139768 6956
rect 139820 6944 139826 6996
rect 140314 6944 140320 6996
rect 140372 6984 140378 6996
rect 143994 6984 144000 6996
rect 140372 6956 144000 6984
rect 140372 6944 140378 6956
rect 143994 6944 144000 6956
rect 144052 6944 144058 6996
rect 42426 6876 42432 6928
rect 42484 6916 42490 6928
rect 49326 6916 49332 6928
rect 42484 6888 49332 6916
rect 42484 6876 42490 6888
rect 49326 6876 49332 6888
rect 49384 6876 49390 6928
rect 52454 6876 52460 6928
rect 52512 6916 52518 6928
rect 52512 6888 53052 6916
rect 52512 6876 52518 6888
rect 2958 6848 2964 6860
rect 2919 6820 2964 6848
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6848 3111 6851
rect 5718 6848 5724 6860
rect 3099 6820 5724 6848
rect 3099 6817 3111 6820
rect 3053 6811 3111 6817
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6848 6331 6851
rect 7190 6848 7196 6860
rect 6319 6820 7196 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 7190 6808 7196 6820
rect 7248 6808 7254 6860
rect 8662 6848 8668 6860
rect 8623 6820 8668 6848
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 9732 6820 10609 6848
rect 9732 6808 9738 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 11698 6848 11704 6860
rect 11659 6820 11704 6848
rect 10597 6811 10655 6817
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6848 13047 6851
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 13035 6820 15301 6848
rect 13035 6817 13047 6820
rect 12989 6811 13047 6817
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 16574 6848 16580 6860
rect 16535 6820 16580 6848
rect 15289 6811 15347 6817
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 21269 6851 21327 6857
rect 21269 6817 21281 6851
rect 21315 6848 21327 6851
rect 21726 6848 21732 6860
rect 21315 6820 21732 6848
rect 21315 6817 21327 6820
rect 21269 6811 21327 6817
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 22370 6848 22376 6860
rect 22331 6820 22376 6848
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 23566 6808 23572 6860
rect 23624 6848 23630 6860
rect 23661 6851 23719 6857
rect 23661 6848 23673 6851
rect 23624 6820 23673 6848
rect 23624 6808 23630 6820
rect 23661 6817 23673 6820
rect 23707 6817 23719 6851
rect 24946 6848 24952 6860
rect 24907 6820 24952 6848
rect 23661 6811 23719 6817
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 27246 6848 27252 6860
rect 26559 6820 27252 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 27246 6808 27252 6820
rect 27304 6808 27310 6860
rect 27706 6848 27712 6860
rect 27667 6820 27712 6848
rect 27706 6808 27712 6820
rect 27764 6808 27770 6860
rect 28442 6808 28448 6860
rect 28500 6848 28506 6860
rect 30282 6848 30288 6860
rect 28500 6820 30288 6848
rect 28500 6808 28506 6820
rect 30282 6808 30288 6820
rect 30340 6808 30346 6860
rect 33318 6848 33324 6860
rect 33279 6820 33324 6848
rect 33318 6808 33324 6820
rect 33376 6808 33382 6860
rect 33962 6808 33968 6860
rect 34020 6848 34026 6860
rect 35894 6848 35900 6860
rect 34020 6820 35900 6848
rect 34020 6808 34026 6820
rect 35894 6808 35900 6820
rect 35952 6808 35958 6860
rect 37734 6808 37740 6860
rect 37792 6848 37798 6860
rect 38105 6851 38163 6857
rect 38105 6848 38117 6851
rect 37792 6820 38117 6848
rect 37792 6808 37798 6820
rect 38105 6817 38117 6820
rect 38151 6817 38163 6851
rect 38105 6811 38163 6817
rect 38194 6808 38200 6860
rect 38252 6848 38258 6860
rect 39942 6848 39948 6860
rect 38252 6820 39948 6848
rect 38252 6808 38258 6820
rect 39942 6808 39948 6820
rect 40000 6808 40006 6860
rect 42245 6851 42303 6857
rect 42245 6817 42257 6851
rect 42291 6848 42303 6851
rect 42886 6848 42892 6860
rect 42291 6820 42892 6848
rect 42291 6817 42303 6820
rect 42245 6811 42303 6817
rect 42886 6808 42892 6820
rect 42944 6808 42950 6860
rect 45554 6808 45560 6860
rect 45612 6848 45618 6860
rect 46385 6851 46443 6857
rect 45612 6820 45657 6848
rect 45612 6808 45618 6820
rect 46385 6817 46397 6851
rect 46431 6848 46443 6851
rect 47302 6848 47308 6860
rect 46431 6820 47308 6848
rect 46431 6817 46443 6820
rect 46385 6811 46443 6817
rect 47302 6808 47308 6820
rect 47360 6808 47366 6860
rect 47578 6848 47584 6860
rect 47539 6820 47584 6848
rect 47578 6808 47584 6820
rect 47636 6808 47642 6860
rect 48958 6848 48964 6860
rect 48919 6820 48964 6848
rect 48958 6808 48964 6820
rect 49016 6808 49022 6860
rect 49142 6808 49148 6860
rect 49200 6848 49206 6860
rect 50065 6851 50123 6857
rect 50065 6848 50077 6851
rect 49200 6820 50077 6848
rect 49200 6808 49206 6820
rect 50065 6817 50077 6820
rect 50111 6817 50123 6851
rect 50065 6811 50123 6817
rect 51813 6851 51871 6857
rect 51813 6817 51825 6851
rect 51859 6848 51871 6851
rect 52546 6848 52552 6860
rect 51859 6820 52552 6848
rect 51859 6817 51871 6820
rect 51813 6811 51871 6817
rect 52546 6808 52552 6820
rect 52604 6808 52610 6860
rect 52638 6808 52644 6860
rect 52696 6848 52702 6860
rect 52917 6851 52975 6857
rect 52917 6848 52929 6851
rect 52696 6820 52929 6848
rect 52696 6808 52702 6820
rect 52917 6817 52929 6820
rect 52963 6817 52975 6851
rect 53024 6848 53052 6888
rect 58636 6888 59216 6916
rect 58636 6860 58664 6888
rect 53024 6820 54892 6848
rect 52917 6811 52975 6817
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6730 6780 6736 6792
rect 6227 6752 6736 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 8478 6780 8484 6792
rect 7147 6752 8484 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 9766 6780 9772 6792
rect 8619 6752 9772 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 12342 6780 12348 6792
rect 12115 6752 12348 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 17954 6780 17960 6792
rect 16807 6752 17960 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 22281 6783 22339 6789
rect 22281 6780 22293 6783
rect 21968 6752 22293 6780
rect 21968 6740 21974 6752
rect 22281 6749 22293 6752
rect 22327 6749 22339 6783
rect 22281 6743 22339 6749
rect 23750 6740 23756 6792
rect 23808 6780 23814 6792
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 23808 6752 24685 6780
rect 23808 6740 23814 6752
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 26694 6740 26700 6792
rect 26752 6780 26758 6792
rect 27525 6783 27583 6789
rect 27525 6780 27537 6783
rect 26752 6752 27537 6780
rect 26752 6740 26758 6752
rect 27525 6749 27537 6752
rect 27571 6749 27583 6783
rect 27525 6743 27583 6749
rect 28626 6740 28632 6792
rect 28684 6780 28690 6792
rect 28905 6783 28963 6789
rect 28905 6780 28917 6783
rect 28684 6752 28917 6780
rect 28684 6740 28690 6752
rect 28905 6749 28917 6752
rect 28951 6749 28963 6783
rect 28905 6743 28963 6749
rect 29638 6740 29644 6792
rect 29696 6780 29702 6792
rect 31021 6783 31079 6789
rect 31021 6780 31033 6783
rect 29696 6752 31033 6780
rect 29696 6740 29702 6752
rect 31021 6749 31033 6752
rect 31067 6749 31079 6783
rect 31021 6743 31079 6749
rect 32125 6783 32183 6789
rect 32125 6749 32137 6783
rect 32171 6780 32183 6783
rect 34517 6783 34575 6789
rect 34517 6780 34529 6783
rect 32171 6752 34529 6780
rect 32171 6749 32183 6752
rect 32125 6743 32183 6749
rect 34517 6749 34529 6752
rect 34563 6749 34575 6783
rect 34517 6743 34575 6749
rect 36633 6783 36691 6789
rect 36633 6749 36645 6783
rect 36679 6780 36691 6783
rect 37826 6780 37832 6792
rect 36679 6752 37832 6780
rect 36679 6749 36691 6752
rect 36633 6743 36691 6749
rect 37826 6740 37832 6752
rect 37884 6740 37890 6792
rect 40678 6740 40684 6792
rect 40736 6780 40742 6792
rect 40736 6752 41552 6780
rect 40736 6740 40742 6752
rect 566 6672 572 6724
rect 624 6712 630 6724
rect 624 6684 3924 6712
rect 624 6672 630 6684
rect 2314 6604 2320 6656
rect 2372 6644 2378 6656
rect 3786 6644 3792 6656
rect 2372 6616 3792 6644
rect 2372 6604 2378 6616
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 3896 6644 3924 6684
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 11330 6712 11336 6724
rect 4028 6684 11336 6712
rect 4028 6672 4034 6684
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 30190 6672 30196 6724
rect 30248 6712 30254 6724
rect 33413 6715 33471 6721
rect 33413 6712 33425 6715
rect 30248 6684 33425 6712
rect 30248 6672 30254 6684
rect 33413 6681 33425 6684
rect 33459 6681 33471 6715
rect 33413 6675 33471 6681
rect 37182 6672 37188 6724
rect 37240 6712 37246 6724
rect 41414 6712 41420 6724
rect 37240 6684 41420 6712
rect 37240 6672 37246 6684
rect 41414 6672 41420 6684
rect 41472 6672 41478 6724
rect 41524 6712 41552 6752
rect 42610 6740 42616 6792
rect 42668 6780 42674 6792
rect 43993 6783 44051 6789
rect 43993 6780 44005 6783
rect 42668 6752 44005 6780
rect 42668 6740 42674 6752
rect 43993 6749 44005 6752
rect 44039 6749 44051 6783
rect 43993 6743 44051 6749
rect 45465 6783 45523 6789
rect 45465 6749 45477 6783
rect 45511 6780 45523 6783
rect 45922 6780 45928 6792
rect 45511 6752 45928 6780
rect 45511 6749 45523 6752
rect 45465 6743 45523 6749
rect 45922 6740 45928 6752
rect 45980 6740 45986 6792
rect 47397 6783 47455 6789
rect 47397 6749 47409 6783
rect 47443 6749 47455 6783
rect 47397 6743 47455 6749
rect 47412 6712 47440 6743
rect 47670 6740 47676 6792
rect 47728 6780 47734 6792
rect 49973 6783 50031 6789
rect 49973 6780 49985 6783
rect 47728 6752 49985 6780
rect 47728 6740 47734 6752
rect 49973 6749 49985 6752
rect 50019 6749 50031 6783
rect 49973 6743 50031 6749
rect 52825 6783 52883 6789
rect 52825 6749 52837 6783
rect 52871 6749 52883 6783
rect 52825 6743 52883 6749
rect 41524 6684 47440 6712
rect 7834 6644 7840 6656
rect 3896 6616 7840 6644
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 28902 6604 28908 6656
rect 28960 6644 28966 6656
rect 33226 6644 33232 6656
rect 28960 6616 33232 6644
rect 28960 6604 28966 6616
rect 33226 6604 33232 6616
rect 33284 6604 33290 6656
rect 50430 6604 50436 6656
rect 50488 6644 50494 6656
rect 52840 6644 52868 6743
rect 53006 6740 53012 6792
rect 53064 6780 53070 6792
rect 54573 6783 54631 6789
rect 54573 6780 54585 6783
rect 53064 6752 54585 6780
rect 53064 6740 53070 6752
rect 54573 6749 54585 6752
rect 54619 6749 54631 6783
rect 54573 6743 54631 6749
rect 54864 6712 54892 6820
rect 56594 6808 56600 6860
rect 56652 6848 56658 6860
rect 57241 6851 57299 6857
rect 57241 6848 57253 6851
rect 56652 6820 57253 6848
rect 56652 6808 56658 6820
rect 57241 6817 57253 6820
rect 57287 6817 57299 6851
rect 57241 6811 57299 6817
rect 58618 6808 58624 6860
rect 58676 6808 58682 6860
rect 58802 6848 58808 6860
rect 58763 6820 58808 6848
rect 58802 6808 58808 6820
rect 58860 6808 58866 6860
rect 59081 6851 59139 6857
rect 59081 6817 59093 6851
rect 59127 6817 59139 6851
rect 59188 6848 59216 6888
rect 60384 6888 60596 6916
rect 60384 6848 60412 6888
rect 59188 6820 60412 6848
rect 60461 6851 60519 6857
rect 59081 6811 59139 6817
rect 60461 6817 60473 6851
rect 60507 6817 60519 6851
rect 60568 6848 60596 6888
rect 68020 6888 68232 6916
rect 60737 6851 60795 6857
rect 60737 6848 60749 6851
rect 60568 6820 60749 6848
rect 60461 6811 60519 6817
rect 60737 6817 60749 6820
rect 60783 6817 60795 6851
rect 60737 6811 60795 6817
rect 62485 6851 62543 6857
rect 62485 6817 62497 6851
rect 62531 6848 62543 6851
rect 62574 6848 62580 6860
rect 62531 6820 62580 6848
rect 62531 6817 62543 6820
rect 62485 6811 62543 6817
rect 56137 6783 56195 6789
rect 56137 6749 56149 6783
rect 56183 6780 56195 6783
rect 57330 6780 57336 6792
rect 56183 6752 57336 6780
rect 56183 6749 56195 6752
rect 56137 6743 56195 6749
rect 57330 6740 57336 6752
rect 57388 6740 57394 6792
rect 57698 6740 57704 6792
rect 57756 6780 57762 6792
rect 59096 6780 59124 6811
rect 57756 6752 59124 6780
rect 60476 6780 60504 6811
rect 62574 6808 62580 6820
rect 62632 6808 62638 6860
rect 62945 6851 63003 6857
rect 62945 6817 62957 6851
rect 62991 6848 63003 6851
rect 63770 6848 63776 6860
rect 62991 6820 63776 6848
rect 62991 6817 63003 6820
rect 62945 6811 63003 6817
rect 63770 6808 63776 6820
rect 63828 6808 63834 6860
rect 64046 6848 64052 6860
rect 64007 6820 64052 6848
rect 64046 6808 64052 6820
rect 64104 6808 64110 6860
rect 64230 6808 64236 6860
rect 64288 6848 64294 6860
rect 64325 6851 64383 6857
rect 64325 6848 64337 6851
rect 64288 6820 64337 6848
rect 64288 6808 64294 6820
rect 64325 6817 64337 6820
rect 64371 6817 64383 6851
rect 64325 6811 64383 6817
rect 66165 6851 66223 6857
rect 66165 6817 66177 6851
rect 66211 6848 66223 6851
rect 66346 6848 66352 6860
rect 66211 6820 66352 6848
rect 66211 6817 66223 6820
rect 66165 6811 66223 6817
rect 66346 6808 66352 6820
rect 66404 6808 66410 6860
rect 66533 6851 66591 6857
rect 66533 6817 66545 6851
rect 66579 6817 66591 6851
rect 66533 6811 66591 6817
rect 61654 6780 61660 6792
rect 60476 6752 61660 6780
rect 57756 6740 57762 6752
rect 61654 6740 61660 6752
rect 61712 6740 61718 6792
rect 65518 6740 65524 6792
rect 65576 6780 65582 6792
rect 66548 6780 66576 6811
rect 67174 6808 67180 6860
rect 67232 6848 67238 6860
rect 67545 6851 67603 6857
rect 67545 6848 67557 6851
rect 67232 6820 67557 6848
rect 67232 6808 67238 6820
rect 67545 6817 67557 6820
rect 67591 6817 67603 6851
rect 67545 6811 67603 6817
rect 65576 6752 66576 6780
rect 65576 6740 65582 6752
rect 66806 6740 66812 6792
rect 66864 6780 66870 6792
rect 68020 6780 68048 6888
rect 68097 6851 68155 6857
rect 68097 6817 68109 6851
rect 68143 6817 68155 6851
rect 68097 6811 68155 6817
rect 66864 6752 68048 6780
rect 66864 6740 66870 6752
rect 57425 6715 57483 6721
rect 57425 6712 57437 6715
rect 54864 6684 57437 6712
rect 57425 6681 57437 6684
rect 57471 6681 57483 6715
rect 57425 6675 57483 6681
rect 66438 6672 66444 6724
rect 66496 6712 66502 6724
rect 68112 6712 68140 6811
rect 68204 6780 68232 6888
rect 73172 6888 73568 6916
rect 69014 6808 69020 6860
rect 69072 6848 69078 6860
rect 69109 6851 69167 6857
rect 69109 6848 69121 6851
rect 69072 6820 69121 6848
rect 69072 6808 69078 6820
rect 69109 6817 69121 6820
rect 69155 6817 69167 6851
rect 69661 6851 69719 6857
rect 69661 6848 69673 6851
rect 69109 6811 69167 6817
rect 69216 6820 69673 6848
rect 69216 6780 69244 6820
rect 69661 6817 69673 6820
rect 69707 6817 69719 6851
rect 69661 6811 69719 6817
rect 70302 6808 70308 6860
rect 70360 6848 70366 6860
rect 71409 6851 71467 6857
rect 71409 6848 71421 6851
rect 70360 6820 71421 6848
rect 70360 6808 70366 6820
rect 71409 6817 71421 6820
rect 71455 6817 71467 6851
rect 71409 6811 71467 6817
rect 71961 6851 72019 6857
rect 71961 6817 71973 6851
rect 72007 6817 72019 6851
rect 71961 6811 72019 6817
rect 69474 6780 69480 6792
rect 68204 6752 69244 6780
rect 69435 6752 69480 6780
rect 69474 6740 69480 6752
rect 69532 6740 69538 6792
rect 69842 6740 69848 6792
rect 69900 6780 69906 6792
rect 71976 6780 72004 6811
rect 69900 6752 72004 6780
rect 69900 6740 69906 6752
rect 66496 6684 68140 6712
rect 66496 6672 66502 6684
rect 70210 6672 70216 6724
rect 70268 6712 70274 6724
rect 73172 6712 73200 6888
rect 73540 6857 73568 6888
rect 75472 6888 75684 6916
rect 73249 6851 73307 6857
rect 73249 6817 73261 6851
rect 73295 6848 73307 6851
rect 73525 6851 73583 6857
rect 73295 6820 73476 6848
rect 73295 6817 73307 6820
rect 73249 6811 73307 6817
rect 73341 6783 73399 6789
rect 73341 6749 73353 6783
rect 73387 6749 73399 6783
rect 73448 6780 73476 6820
rect 73525 6817 73537 6851
rect 73571 6817 73583 6851
rect 73525 6811 73583 6817
rect 74258 6808 74264 6860
rect 74316 6848 74322 6860
rect 75472 6848 75500 6888
rect 74316 6820 75500 6848
rect 75549 6851 75607 6857
rect 74316 6808 74322 6820
rect 75549 6817 75561 6851
rect 75595 6817 75607 6851
rect 75656 6848 75684 6888
rect 77496 6888 77708 6916
rect 75917 6851 75975 6857
rect 75917 6848 75929 6851
rect 75656 6820 75929 6848
rect 75549 6811 75607 6817
rect 75917 6817 75929 6820
rect 75963 6817 75975 6851
rect 75917 6811 75975 6817
rect 74534 6780 74540 6792
rect 73448 6752 74540 6780
rect 73341 6743 73399 6749
rect 70268 6684 73200 6712
rect 70268 6672 70274 6684
rect 73246 6672 73252 6724
rect 73304 6712 73310 6724
rect 73356 6712 73384 6743
rect 74534 6740 74540 6752
rect 74592 6740 74598 6792
rect 73304 6684 73384 6712
rect 75564 6712 75592 6811
rect 76466 6808 76472 6860
rect 76524 6848 76530 6860
rect 77496 6848 77524 6888
rect 76524 6820 77524 6848
rect 77573 6851 77631 6857
rect 76524 6808 76530 6820
rect 77573 6817 77585 6851
rect 77619 6817 77631 6851
rect 77680 6848 77708 6888
rect 85316 6888 85528 6916
rect 77849 6851 77907 6857
rect 77849 6848 77861 6851
rect 77680 6820 77861 6848
rect 77573 6811 77631 6817
rect 77849 6817 77861 6820
rect 77895 6817 77907 6851
rect 79873 6851 79931 6857
rect 79873 6848 79885 6851
rect 77849 6811 77907 6817
rect 78048 6820 79885 6848
rect 77588 6780 77616 6811
rect 78048 6780 78076 6820
rect 79873 6817 79885 6820
rect 79919 6817 79931 6851
rect 79873 6811 79931 6817
rect 81161 6851 81219 6857
rect 81161 6817 81173 6851
rect 81207 6817 81219 6851
rect 81161 6811 81219 6817
rect 81621 6851 81679 6857
rect 81621 6817 81633 6851
rect 81667 6817 81679 6851
rect 82630 6848 82636 6860
rect 82591 6820 82636 6848
rect 81621 6811 81679 6817
rect 77588 6752 78076 6780
rect 78861 6783 78919 6789
rect 78861 6749 78873 6783
rect 78907 6749 78919 6783
rect 78861 6743 78919 6749
rect 78876 6712 78904 6743
rect 75564 6684 78904 6712
rect 81176 6712 81204 6811
rect 81253 6783 81311 6789
rect 81253 6749 81265 6783
rect 81299 6780 81311 6783
rect 81526 6780 81532 6792
rect 81299 6752 81532 6780
rect 81299 6749 81311 6752
rect 81253 6743 81311 6749
rect 81526 6740 81532 6752
rect 81584 6740 81590 6792
rect 81636 6780 81664 6811
rect 82630 6808 82636 6820
rect 82688 6808 82694 6860
rect 83366 6848 83372 6860
rect 82740 6820 83136 6848
rect 83327 6820 83372 6848
rect 82740 6780 82768 6820
rect 82998 6780 83004 6792
rect 81636 6752 82768 6780
rect 82959 6752 83004 6780
rect 82998 6740 83004 6752
rect 83056 6740 83062 6792
rect 83108 6780 83136 6820
rect 83366 6808 83372 6820
rect 83424 6808 83430 6860
rect 85114 6808 85120 6860
rect 85172 6848 85178 6860
rect 85316 6848 85344 6888
rect 85172 6820 85344 6848
rect 85393 6851 85451 6857
rect 85172 6808 85178 6820
rect 85393 6817 85405 6851
rect 85439 6817 85451 6851
rect 85500 6848 85528 6888
rect 86954 6876 86960 6928
rect 87012 6916 87018 6928
rect 87012 6888 88380 6916
rect 87012 6876 87018 6888
rect 85669 6851 85727 6857
rect 85669 6848 85681 6851
rect 85500 6820 85681 6848
rect 85393 6811 85451 6817
rect 85669 6817 85681 6820
rect 85715 6817 85727 6851
rect 88245 6851 88303 6857
rect 88245 6848 88257 6851
rect 85669 6811 85727 6817
rect 85776 6820 88257 6848
rect 84286 6780 84292 6792
rect 83108 6752 84292 6780
rect 84286 6740 84292 6752
rect 84344 6740 84350 6792
rect 85408 6780 85436 6811
rect 85776 6780 85804 6820
rect 88245 6817 88257 6820
rect 88291 6817 88303 6851
rect 88352 6848 88380 6888
rect 91848 6888 92060 6916
rect 89898 6848 89904 6860
rect 88352 6820 89904 6848
rect 88245 6811 88303 6817
rect 89898 6808 89904 6820
rect 89956 6808 89962 6860
rect 90358 6848 90364 6860
rect 90319 6820 90364 6848
rect 90358 6808 90364 6820
rect 90416 6808 90422 6860
rect 90821 6851 90879 6857
rect 90821 6817 90833 6851
rect 90867 6848 90879 6851
rect 91848 6848 91876 6888
rect 90867 6820 91876 6848
rect 91925 6851 91983 6857
rect 90867 6817 90879 6820
rect 90821 6811 90879 6817
rect 91925 6817 91937 6851
rect 91971 6817 91983 6851
rect 92032 6848 92060 6888
rect 94700 6888 95280 6916
rect 92106 6848 92112 6860
rect 92032 6820 92112 6848
rect 91925 6811 91983 6817
rect 85408 6752 85804 6780
rect 86681 6783 86739 6789
rect 86681 6749 86693 6783
rect 86727 6749 86739 6783
rect 86681 6743 86739 6749
rect 86696 6712 86724 6743
rect 81176 6684 86724 6712
rect 91940 6712 91968 6811
rect 92106 6808 92112 6820
rect 92164 6808 92170 6860
rect 92385 6851 92443 6857
rect 92385 6817 92397 6851
rect 92431 6848 92443 6851
rect 94700 6848 94728 6888
rect 92431 6820 94728 6848
rect 94777 6851 94835 6857
rect 92431 6817 92443 6820
rect 92385 6811 92443 6817
rect 94777 6817 94789 6851
rect 94823 6848 94835 6851
rect 95142 6848 95148 6860
rect 94823 6820 95004 6848
rect 95103 6820 95148 6848
rect 94823 6817 94835 6820
rect 94777 6811 94835 6817
rect 94976 6712 95004 6820
rect 95142 6808 95148 6820
rect 95200 6808 95206 6860
rect 95252 6848 95280 6888
rect 97902 6876 97908 6928
rect 97960 6916 97966 6928
rect 105906 6916 105912 6928
rect 97960 6888 105912 6916
rect 97960 6876 97966 6888
rect 105906 6876 105912 6888
rect 105964 6876 105970 6928
rect 106550 6916 106556 6928
rect 106384 6888 106556 6916
rect 96338 6848 96344 6860
rect 95252 6820 96344 6848
rect 96338 6808 96344 6820
rect 96396 6808 96402 6860
rect 96433 6851 96491 6857
rect 96433 6817 96445 6851
rect 96479 6848 96491 6851
rect 96706 6848 96712 6860
rect 96479 6820 96712 6848
rect 96479 6817 96491 6820
rect 96433 6811 96491 6817
rect 96706 6808 96712 6820
rect 96764 6808 96770 6860
rect 96893 6851 96951 6857
rect 96893 6817 96905 6851
rect 96939 6848 96951 6851
rect 97442 6848 97448 6860
rect 96939 6820 97448 6848
rect 96939 6817 96951 6820
rect 96893 6811 96951 6817
rect 97442 6808 97448 6820
rect 97500 6808 97506 6860
rect 97997 6851 98055 6857
rect 97997 6817 98009 6851
rect 98043 6817 98055 6851
rect 97997 6811 98055 6817
rect 98457 6851 98515 6857
rect 98457 6817 98469 6851
rect 98503 6848 98515 6851
rect 99558 6848 99564 6860
rect 98503 6820 99564 6848
rect 98503 6817 98515 6820
rect 98457 6811 98515 6817
rect 96246 6740 96252 6792
rect 96304 6780 96310 6792
rect 96525 6783 96583 6789
rect 96525 6780 96537 6783
rect 96304 6752 96537 6780
rect 96304 6740 96310 6752
rect 96525 6749 96537 6752
rect 96571 6749 96583 6783
rect 98012 6780 98040 6811
rect 99558 6808 99564 6820
rect 99616 6808 99622 6860
rect 99742 6808 99748 6860
rect 99800 6848 99806 6860
rect 103054 6848 103060 6860
rect 99800 6820 103060 6848
rect 99800 6808 99806 6820
rect 103054 6808 103060 6820
rect 103112 6808 103118 6860
rect 106384 6857 106412 6888
rect 106550 6876 106556 6888
rect 106608 6876 106614 6928
rect 110417 6919 110475 6925
rect 110417 6885 110429 6919
rect 110463 6916 110475 6919
rect 110463 6888 111380 6916
rect 110463 6885 110475 6888
rect 110417 6879 110475 6885
rect 103977 6851 104035 6857
rect 103977 6817 103989 6851
rect 104023 6848 104035 6851
rect 106369 6851 106427 6857
rect 104023 6820 106228 6848
rect 104023 6817 104035 6820
rect 103977 6811 104035 6817
rect 99282 6780 99288 6792
rect 98012 6752 99288 6780
rect 96525 6743 96583 6749
rect 99282 6740 99288 6752
rect 99340 6740 99346 6792
rect 100757 6783 100815 6789
rect 100757 6749 100769 6783
rect 100803 6780 100815 6783
rect 102413 6783 102471 6789
rect 102413 6780 102425 6783
rect 100803 6752 102425 6780
rect 100803 6749 100815 6752
rect 100757 6743 100815 6749
rect 102413 6749 102425 6752
rect 102459 6749 102471 6783
rect 102413 6743 102471 6749
rect 103885 6783 103943 6789
rect 103885 6749 103897 6783
rect 103931 6780 103943 6783
rect 104434 6780 104440 6792
rect 103931 6752 104440 6780
rect 103931 6749 103943 6752
rect 103885 6743 103943 6749
rect 104434 6740 104440 6752
rect 104492 6740 104498 6792
rect 105078 6740 105084 6792
rect 105136 6780 105142 6792
rect 105265 6783 105323 6789
rect 105265 6780 105277 6783
rect 105136 6752 105277 6780
rect 105136 6740 105142 6752
rect 105265 6749 105277 6752
rect 105311 6749 105323 6783
rect 105265 6743 105323 6749
rect 91940 6684 94728 6712
rect 94976 6684 97948 6712
rect 73304 6672 73310 6684
rect 58618 6644 58624 6656
rect 50488 6616 52868 6644
rect 58579 6616 58624 6644
rect 50488 6604 50494 6616
rect 58618 6604 58624 6616
rect 58676 6604 58682 6656
rect 58894 6604 58900 6656
rect 58952 6644 58958 6656
rect 60277 6647 60335 6653
rect 60277 6644 60289 6647
rect 58952 6616 60289 6644
rect 58952 6604 58958 6616
rect 60277 6613 60289 6616
rect 60323 6613 60335 6647
rect 62298 6644 62304 6656
rect 62259 6616 62304 6644
rect 60277 6607 60335 6613
rect 62298 6604 62304 6616
rect 62356 6604 62362 6656
rect 63494 6604 63500 6656
rect 63552 6644 63558 6656
rect 63865 6647 63923 6653
rect 63865 6644 63877 6647
rect 63552 6616 63877 6644
rect 63552 6604 63558 6616
rect 63865 6613 63877 6616
rect 63911 6613 63923 6647
rect 63865 6607 63923 6613
rect 66073 6647 66131 6653
rect 66073 6613 66085 6647
rect 66119 6644 66131 6647
rect 66254 6644 66260 6656
rect 66119 6616 66260 6644
rect 66119 6613 66131 6616
rect 66073 6607 66131 6613
rect 66254 6604 66260 6616
rect 66312 6604 66318 6656
rect 67634 6644 67640 6656
rect 67595 6616 67640 6644
rect 67634 6604 67640 6616
rect 67692 6604 67698 6656
rect 67726 6604 67732 6656
rect 67784 6644 67790 6656
rect 68830 6644 68836 6656
rect 67784 6616 68836 6644
rect 67784 6604 67790 6616
rect 68830 6604 68836 6616
rect 68888 6604 68894 6656
rect 69014 6604 69020 6656
rect 69072 6644 69078 6656
rect 70118 6644 70124 6656
rect 69072 6616 70124 6644
rect 69072 6604 69078 6616
rect 70118 6604 70124 6616
rect 70176 6604 70182 6656
rect 71498 6644 71504 6656
rect 71459 6616 71504 6644
rect 71498 6604 71504 6616
rect 71556 6604 71562 6656
rect 72786 6604 72792 6656
rect 72844 6644 72850 6656
rect 75365 6647 75423 6653
rect 75365 6644 75377 6647
rect 72844 6616 75377 6644
rect 72844 6604 72850 6616
rect 75365 6613 75377 6616
rect 75411 6613 75423 6647
rect 75365 6607 75423 6613
rect 76190 6604 76196 6656
rect 76248 6644 76254 6656
rect 77389 6647 77447 6653
rect 77389 6644 77401 6647
rect 76248 6616 77401 6644
rect 76248 6604 76254 6616
rect 77389 6613 77401 6616
rect 77435 6613 77447 6647
rect 77389 6607 77447 6613
rect 80790 6604 80796 6656
rect 80848 6644 80854 6656
rect 83458 6644 83464 6656
rect 80848 6616 83464 6644
rect 80848 6604 80854 6616
rect 83458 6604 83464 6616
rect 83516 6604 83522 6656
rect 84654 6604 84660 6656
rect 84712 6644 84718 6656
rect 85209 6647 85267 6653
rect 85209 6644 85221 6647
rect 84712 6616 85221 6644
rect 84712 6604 84718 6616
rect 85209 6613 85221 6616
rect 85255 6613 85267 6647
rect 90174 6644 90180 6656
rect 90135 6616 90180 6644
rect 85209 6607 85267 6613
rect 90174 6604 90180 6616
rect 90232 6604 90238 6656
rect 91646 6604 91652 6656
rect 91704 6644 91710 6656
rect 91741 6647 91799 6653
rect 91741 6644 91753 6647
rect 91704 6616 91753 6644
rect 91704 6604 91710 6616
rect 91741 6613 91753 6616
rect 91787 6613 91799 6647
rect 91741 6607 91799 6613
rect 93578 6604 93584 6656
rect 93636 6644 93642 6656
rect 94593 6647 94651 6653
rect 94593 6644 94605 6647
rect 93636 6616 94605 6644
rect 93636 6604 93642 6616
rect 94593 6613 94605 6616
rect 94639 6613 94651 6647
rect 94700 6644 94728 6684
rect 97626 6644 97632 6656
rect 94700 6616 97632 6644
rect 94593 6607 94651 6613
rect 97626 6604 97632 6616
rect 97684 6604 97690 6656
rect 97810 6644 97816 6656
rect 97771 6616 97816 6644
rect 97810 6604 97816 6616
rect 97868 6604 97874 6656
rect 97920 6644 97948 6684
rect 97994 6672 98000 6724
rect 98052 6712 98058 6724
rect 101674 6712 101680 6724
rect 98052 6684 101680 6712
rect 98052 6672 98058 6684
rect 101674 6672 101680 6684
rect 101732 6672 101738 6724
rect 102686 6672 102692 6724
rect 102744 6712 102750 6724
rect 106090 6712 106096 6724
rect 102744 6684 106096 6712
rect 102744 6672 102750 6684
rect 106090 6672 106096 6684
rect 106148 6672 106154 6724
rect 106200 6712 106228 6820
rect 106369 6817 106381 6851
rect 106415 6817 106427 6851
rect 106369 6811 106427 6817
rect 109221 6851 109279 6857
rect 109221 6817 109233 6851
rect 109267 6848 109279 6851
rect 110509 6851 110567 6857
rect 110509 6848 110521 6851
rect 109267 6820 110521 6848
rect 109267 6817 109279 6820
rect 109221 6811 109279 6817
rect 110509 6817 110521 6820
rect 110555 6817 110567 6851
rect 110509 6811 110567 6817
rect 110969 6851 111027 6857
rect 110969 6817 110981 6851
rect 111015 6848 111027 6851
rect 111058 6848 111064 6860
rect 111015 6820 111064 6848
rect 111015 6817 111027 6820
rect 110969 6811 111027 6817
rect 111058 6808 111064 6820
rect 111116 6808 111122 6860
rect 111245 6851 111303 6857
rect 111245 6817 111257 6851
rect 111291 6817 111303 6851
rect 111352 6848 111380 6888
rect 114940 6888 115244 6916
rect 114940 6848 114968 6888
rect 115106 6848 115112 6860
rect 111352 6820 114968 6848
rect 115067 6820 115112 6848
rect 111245 6811 111303 6817
rect 106274 6740 106280 6792
rect 106332 6780 106338 6792
rect 107657 6783 107715 6789
rect 107657 6780 107669 6783
rect 106332 6752 107669 6780
rect 106332 6740 106338 6752
rect 107657 6749 107669 6752
rect 107703 6749 107715 6783
rect 108850 6780 108856 6792
rect 108811 6752 108856 6780
rect 107657 6743 107715 6749
rect 108850 6740 108856 6752
rect 108908 6740 108914 6792
rect 109494 6740 109500 6792
rect 109552 6780 109558 6792
rect 111260 6780 111288 6811
rect 115106 6808 115112 6820
rect 115164 6808 115170 6860
rect 115216 6848 115244 6888
rect 127710 6876 127716 6928
rect 127768 6916 127774 6928
rect 127768 6888 139348 6916
rect 127768 6876 127774 6888
rect 115658 6848 115664 6860
rect 115216 6820 115664 6848
rect 115658 6808 115664 6820
rect 115716 6808 115722 6860
rect 116302 6848 116308 6860
rect 116263 6820 116308 6848
rect 116302 6808 116308 6820
rect 116360 6808 116366 6860
rect 117869 6851 117927 6857
rect 117869 6817 117881 6851
rect 117915 6848 117927 6851
rect 119798 6848 119804 6860
rect 117915 6820 119804 6848
rect 117915 6817 117927 6820
rect 117869 6811 117927 6817
rect 119798 6808 119804 6820
rect 119856 6808 119862 6860
rect 120166 6848 120172 6860
rect 120127 6820 120172 6848
rect 120166 6808 120172 6820
rect 120224 6808 120230 6860
rect 120258 6808 120264 6860
rect 120316 6848 120322 6860
rect 122009 6851 122067 6857
rect 122009 6848 122021 6851
rect 120316 6820 122021 6848
rect 120316 6808 120322 6820
rect 122009 6817 122021 6820
rect 122055 6817 122067 6851
rect 122009 6811 122067 6817
rect 123573 6851 123631 6857
rect 123573 6817 123585 6851
rect 123619 6848 123631 6851
rect 123662 6848 123668 6860
rect 123619 6820 123668 6848
rect 123619 6817 123631 6820
rect 123573 6811 123631 6817
rect 123662 6808 123668 6820
rect 123720 6808 123726 6860
rect 124582 6848 124588 6860
rect 124543 6820 124588 6848
rect 124582 6808 124588 6820
rect 124640 6808 124646 6860
rect 125502 6808 125508 6860
rect 125560 6848 125566 6860
rect 125962 6848 125968 6860
rect 125560 6820 125968 6848
rect 125560 6808 125566 6820
rect 125962 6808 125968 6820
rect 126020 6808 126026 6860
rect 126149 6851 126207 6857
rect 126149 6817 126161 6851
rect 126195 6848 126207 6851
rect 129090 6848 129096 6860
rect 126195 6820 129096 6848
rect 126195 6817 126207 6820
rect 126149 6811 126207 6817
rect 129090 6808 129096 6820
rect 129148 6808 129154 6860
rect 129274 6848 129280 6860
rect 129235 6820 129280 6848
rect 129274 6808 129280 6820
rect 129332 6808 129338 6860
rect 131298 6848 131304 6860
rect 129384 6820 131304 6848
rect 109552 6752 111288 6780
rect 112441 6783 112499 6789
rect 109552 6740 109558 6752
rect 112441 6749 112453 6783
rect 112487 6780 112499 6783
rect 113545 6783 113603 6789
rect 113545 6780 113557 6783
rect 112487 6752 113557 6780
rect 112487 6749 112499 6752
rect 112441 6743 112499 6749
rect 113545 6749 113557 6752
rect 113591 6749 113603 6783
rect 113545 6743 113603 6749
rect 114462 6740 114468 6792
rect 114520 6780 114526 6792
rect 114830 6780 114836 6792
rect 114520 6752 114836 6780
rect 114520 6740 114526 6752
rect 114830 6740 114836 6752
rect 114888 6740 114894 6792
rect 115017 6783 115075 6789
rect 115017 6749 115029 6783
rect 115063 6780 115075 6783
rect 117777 6783 117835 6789
rect 115063 6752 117728 6780
rect 115063 6749 115075 6752
rect 115017 6743 115075 6749
rect 106642 6712 106648 6724
rect 106200 6684 106648 6712
rect 106642 6672 106648 6684
rect 106700 6672 106706 6724
rect 106737 6715 106795 6721
rect 106737 6681 106749 6715
rect 106783 6681 106795 6715
rect 106737 6675 106795 6681
rect 99190 6644 99196 6656
rect 97920 6616 99196 6644
rect 99190 6604 99196 6616
rect 99248 6604 99254 6656
rect 106752 6644 106780 6675
rect 106826 6672 106832 6724
rect 106884 6712 106890 6724
rect 110417 6715 110475 6721
rect 110417 6712 110429 6715
rect 106884 6684 110429 6712
rect 106884 6672 106890 6684
rect 110417 6681 110429 6684
rect 110463 6681 110475 6715
rect 110417 6675 110475 6681
rect 110509 6715 110567 6721
rect 110509 6681 110521 6715
rect 110555 6712 110567 6715
rect 115750 6712 115756 6724
rect 110555 6684 115756 6712
rect 110555 6681 110567 6684
rect 110509 6675 110567 6681
rect 115750 6672 115756 6684
rect 115808 6672 115814 6724
rect 117700 6712 117728 6752
rect 117777 6749 117789 6783
rect 117823 6780 117835 6783
rect 118142 6780 118148 6792
rect 117823 6752 118148 6780
rect 117823 6749 117835 6752
rect 117777 6743 117835 6749
rect 118142 6740 118148 6752
rect 118200 6740 118206 6792
rect 118694 6740 118700 6792
rect 118752 6780 118758 6792
rect 118752 6752 118797 6780
rect 118752 6740 118758 6752
rect 118878 6740 118884 6792
rect 118936 6780 118942 6792
rect 122098 6780 122104 6792
rect 118936 6752 122104 6780
rect 118936 6740 118942 6752
rect 122098 6740 122104 6752
rect 122156 6740 122162 6792
rect 123481 6783 123539 6789
rect 123481 6749 123493 6783
rect 123527 6780 123539 6783
rect 124214 6780 124220 6792
rect 123527 6752 124220 6780
rect 123527 6749 123539 6752
rect 123481 6743 123539 6749
rect 124214 6740 124220 6752
rect 124272 6740 124278 6792
rect 124306 6740 124312 6792
rect 124364 6780 124370 6792
rect 124950 6780 124956 6792
rect 124364 6752 124956 6780
rect 124364 6740 124370 6752
rect 124950 6740 124956 6752
rect 125008 6740 125014 6792
rect 126057 6783 126115 6789
rect 126057 6749 126069 6783
rect 126103 6780 126115 6783
rect 127618 6780 127624 6792
rect 126103 6752 127624 6780
rect 126103 6749 126115 6752
rect 126057 6743 126115 6749
rect 127618 6740 127624 6752
rect 127676 6740 127682 6792
rect 127894 6780 127900 6792
rect 127855 6752 127900 6780
rect 127894 6740 127900 6752
rect 127952 6740 127958 6792
rect 129384 6789 129412 6820
rect 131298 6808 131304 6820
rect 131356 6808 131362 6860
rect 131482 6848 131488 6860
rect 131443 6820 131488 6848
rect 131482 6808 131488 6820
rect 131540 6808 131546 6860
rect 134058 6848 134064 6860
rect 131592 6820 134064 6848
rect 129369 6783 129427 6789
rect 129369 6749 129381 6783
rect 129415 6749 129427 6783
rect 129369 6743 129427 6749
rect 130289 6783 130347 6789
rect 130289 6749 130301 6783
rect 130335 6780 130347 6783
rect 131592 6780 131620 6820
rect 134058 6808 134064 6820
rect 134116 6808 134122 6860
rect 134153 6851 134211 6857
rect 134153 6817 134165 6851
rect 134199 6848 134211 6851
rect 134334 6848 134340 6860
rect 134199 6820 134340 6848
rect 134199 6817 134211 6820
rect 134153 6811 134211 6817
rect 134334 6808 134340 6820
rect 134392 6808 134398 6860
rect 134426 6808 134432 6860
rect 134484 6848 134490 6860
rect 135530 6848 135536 6860
rect 134484 6820 135536 6848
rect 134484 6808 134490 6820
rect 135530 6808 135536 6820
rect 135588 6808 135594 6860
rect 135714 6848 135720 6860
rect 135675 6820 135720 6848
rect 135714 6808 135720 6820
rect 135772 6808 135778 6860
rect 138753 6851 138811 6857
rect 138753 6848 138765 6851
rect 136468 6820 138765 6848
rect 131758 6780 131764 6792
rect 130335 6752 131620 6780
rect 131719 6752 131764 6780
rect 130335 6749 130347 6752
rect 130289 6743 130347 6749
rect 131758 6740 131764 6752
rect 131816 6740 131822 6792
rect 132494 6740 132500 6792
rect 132552 6780 132558 6792
rect 133141 6783 133199 6789
rect 133141 6780 133153 6783
rect 132552 6752 133153 6780
rect 132552 6740 132558 6752
rect 133141 6749 133153 6752
rect 133187 6749 133199 6783
rect 133141 6743 133199 6749
rect 133322 6740 133328 6792
rect 133380 6780 133386 6792
rect 135254 6780 135260 6792
rect 133380 6752 135260 6780
rect 133380 6740 133386 6752
rect 135254 6740 135260 6752
rect 135312 6740 135318 6792
rect 135622 6780 135628 6792
rect 135583 6752 135628 6780
rect 135622 6740 135628 6752
rect 135680 6740 135686 6792
rect 120169 6715 120227 6721
rect 117700 6684 118832 6712
rect 110598 6644 110604 6656
rect 106752 6616 110604 6644
rect 110598 6604 110604 6616
rect 110656 6604 110662 6656
rect 110782 6644 110788 6656
rect 110743 6616 110788 6644
rect 110782 6604 110788 6616
rect 110840 6604 110846 6656
rect 112254 6604 112260 6656
rect 112312 6644 112318 6656
rect 118326 6644 118332 6656
rect 112312 6616 118332 6644
rect 112312 6604 112318 6616
rect 118326 6604 118332 6616
rect 118384 6604 118390 6656
rect 118804 6644 118832 6684
rect 120169 6681 120181 6715
rect 120215 6712 120227 6715
rect 128814 6712 128820 6724
rect 120215 6684 128820 6712
rect 120215 6681 120227 6684
rect 120169 6675 120227 6681
rect 128814 6672 128820 6684
rect 128872 6672 128878 6724
rect 131206 6672 131212 6724
rect 131264 6712 131270 6724
rect 132034 6712 132040 6724
rect 131264 6684 132040 6712
rect 131264 6672 131270 6684
rect 132034 6672 132040 6684
rect 132092 6672 132098 6724
rect 132586 6672 132592 6724
rect 132644 6712 132650 6724
rect 136468 6712 136496 6820
rect 138753 6817 138765 6820
rect 138799 6817 138811 6851
rect 139320 6848 139348 6888
rect 140682 6876 140688 6928
rect 140740 6916 140746 6928
rect 147858 6916 147864 6928
rect 140740 6888 147864 6916
rect 140740 6876 140746 6888
rect 147858 6876 147864 6888
rect 147916 6876 147922 6928
rect 141050 6848 141056 6860
rect 139320 6820 141056 6848
rect 138753 6811 138811 6817
rect 141050 6808 141056 6820
rect 141108 6808 141114 6860
rect 141142 6808 141148 6860
rect 141200 6848 141206 6860
rect 141329 6851 141387 6857
rect 141329 6848 141341 6851
rect 141200 6820 141341 6848
rect 141200 6808 141206 6820
rect 141329 6817 141341 6820
rect 141375 6817 141387 6851
rect 141329 6811 141387 6817
rect 142433 6851 142491 6857
rect 142433 6817 142445 6851
rect 142479 6817 142491 6851
rect 142433 6811 142491 6817
rect 136545 6783 136603 6789
rect 136545 6749 136557 6783
rect 136591 6749 136603 6783
rect 136545 6743 136603 6749
rect 132644 6684 136496 6712
rect 136560 6712 136588 6743
rect 136634 6740 136640 6792
rect 136692 6780 136698 6792
rect 137557 6783 137615 6789
rect 137557 6780 137569 6783
rect 136692 6752 137569 6780
rect 136692 6740 136698 6752
rect 137557 6749 137569 6752
rect 137603 6749 137615 6783
rect 137557 6743 137615 6749
rect 137646 6740 137652 6792
rect 137704 6780 137710 6792
rect 137704 6752 138612 6780
rect 137704 6740 137710 6752
rect 138474 6712 138480 6724
rect 136560 6684 138480 6712
rect 132644 6672 132650 6684
rect 138474 6672 138480 6684
rect 138532 6672 138538 6724
rect 138584 6712 138612 6752
rect 139026 6740 139032 6792
rect 139084 6780 139090 6792
rect 142448 6780 142476 6811
rect 143626 6808 143632 6860
rect 143684 6848 143690 6860
rect 144365 6851 144423 6857
rect 144365 6848 144377 6851
rect 143684 6820 144377 6848
rect 143684 6808 143690 6820
rect 144365 6817 144377 6820
rect 144411 6817 144423 6851
rect 144365 6811 144423 6817
rect 146849 6851 146907 6857
rect 146849 6817 146861 6851
rect 146895 6848 146907 6851
rect 147766 6848 147772 6860
rect 146895 6820 147772 6848
rect 146895 6817 146907 6820
rect 146849 6811 146907 6817
rect 147766 6808 147772 6820
rect 147824 6808 147830 6860
rect 147950 6848 147956 6860
rect 147911 6820 147956 6848
rect 147950 6808 147956 6820
rect 148008 6808 148014 6860
rect 150710 6848 150716 6860
rect 150671 6820 150716 6848
rect 150710 6808 150716 6820
rect 150768 6808 150774 6860
rect 151078 6808 151084 6860
rect 151136 6848 151142 6860
rect 151725 6851 151783 6857
rect 151725 6848 151737 6851
rect 151136 6820 151737 6848
rect 151136 6808 151142 6820
rect 151725 6817 151737 6820
rect 151771 6817 151783 6851
rect 153010 6848 153016 6860
rect 152971 6820 153016 6848
rect 151725 6811 151783 6817
rect 153010 6808 153016 6820
rect 153068 6808 153074 6860
rect 139084 6752 142476 6780
rect 139084 6740 139090 6752
rect 144914 6740 144920 6792
rect 144972 6780 144978 6792
rect 145377 6783 145435 6789
rect 145377 6780 145389 6783
rect 144972 6752 145389 6780
rect 144972 6740 144978 6752
rect 145377 6749 145389 6752
rect 145423 6749 145435 6783
rect 152550 6780 152556 6792
rect 145377 6743 145435 6749
rect 148244 6752 152556 6780
rect 141142 6712 141148 6724
rect 138584 6684 141148 6712
rect 141142 6672 141148 6684
rect 141200 6672 141206 6724
rect 142801 6715 142859 6721
rect 142801 6681 142813 6715
rect 142847 6712 142859 6715
rect 148244 6712 148272 6752
rect 152550 6740 152556 6752
rect 152608 6740 152614 6792
rect 153102 6780 153108 6792
rect 153063 6752 153108 6780
rect 153102 6740 153108 6752
rect 153160 6740 153166 6792
rect 142847 6684 148272 6712
rect 148321 6715 148379 6721
rect 142847 6681 142859 6684
rect 142801 6675 142859 6681
rect 148321 6681 148333 6715
rect 148367 6712 148379 6715
rect 157153 6715 157211 6721
rect 157153 6712 157165 6715
rect 148367 6684 157165 6712
rect 148367 6681 148379 6684
rect 148321 6675 148379 6681
rect 157153 6681 157165 6684
rect 157199 6681 157211 6715
rect 157153 6675 157211 6681
rect 125778 6644 125784 6656
rect 118804 6616 125784 6644
rect 125778 6604 125784 6616
rect 125836 6604 125842 6656
rect 125962 6604 125968 6656
rect 126020 6644 126026 6656
rect 130194 6644 130200 6656
rect 126020 6616 130200 6644
rect 126020 6604 126026 6616
rect 130194 6604 130200 6616
rect 130252 6604 130258 6656
rect 130470 6604 130476 6656
rect 130528 6644 130534 6656
rect 154850 6644 154856 6656
rect 130528 6616 154856 6644
rect 130528 6604 130534 6616
rect 154850 6604 154856 6616
rect 154908 6604 154914 6656
rect 1104 6554 154560 6576
rect 1104 6502 4078 6554
rect 4130 6502 44078 6554
rect 44130 6502 84078 6554
rect 84130 6502 124078 6554
rect 124130 6502 154560 6554
rect 1104 6480 154560 6502
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 7282 6440 7288 6452
rect 3844 6412 7288 6440
rect 3844 6400 3850 6412
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 27154 6400 27160 6452
rect 27212 6440 27218 6452
rect 27212 6412 33088 6440
rect 27212 6400 27218 6412
rect 1854 6332 1860 6384
rect 1912 6372 1918 6384
rect 6914 6372 6920 6384
rect 1912 6344 6920 6372
rect 1912 6332 1918 6344
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 8754 6372 8760 6384
rect 7116 6344 8760 6372
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6304 3387 6307
rect 4614 6304 4620 6316
rect 3375 6276 4620 6304
rect 3375 6273 3387 6276
rect 3329 6267 3387 6273
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 7116 6304 7144 6344
rect 8754 6332 8760 6344
rect 8812 6332 8818 6384
rect 13725 6375 13783 6381
rect 13725 6341 13737 6375
rect 13771 6372 13783 6375
rect 15010 6372 15016 6384
rect 13771 6344 15016 6372
rect 13771 6341 13783 6344
rect 13725 6335 13783 6341
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 17037 6375 17095 6381
rect 17037 6341 17049 6375
rect 17083 6372 17095 6375
rect 17126 6372 17132 6384
rect 17083 6344 17132 6372
rect 17083 6341 17095 6344
rect 17037 6335 17095 6341
rect 17126 6332 17132 6344
rect 17184 6332 17190 6384
rect 19334 6332 19340 6384
rect 19392 6372 19398 6384
rect 20898 6372 20904 6384
rect 19392 6344 20904 6372
rect 19392 6332 19398 6344
rect 20898 6332 20904 6344
rect 20956 6332 20962 6384
rect 26878 6332 26884 6384
rect 26936 6372 26942 6384
rect 27614 6372 27620 6384
rect 26936 6344 27620 6372
rect 26936 6332 26942 6344
rect 27614 6332 27620 6344
rect 27672 6332 27678 6384
rect 29362 6332 29368 6384
rect 29420 6372 29426 6384
rect 29420 6344 30696 6372
rect 29420 6332 29426 6344
rect 8205 6307 8263 6313
rect 5859 6276 7144 6304
rect 7484 6276 8064 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 4341 6239 4399 6245
rect 4341 6236 4353 6239
rect 2004 6208 4353 6236
rect 2004 6196 2010 6208
rect 4341 6205 4353 6208
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 5905 6239 5963 6245
rect 5905 6205 5917 6239
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 5920 6168 5948 6199
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6788 6208 6837 6236
rect 6788 6196 6794 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7484 6236 7512 6276
rect 6972 6208 7512 6236
rect 6972 6196 6978 6208
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7616 6208 7941 6236
rect 7616 6196 7622 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 7929 6199 7987 6205
rect 7834 6168 7840 6180
rect 5920 6140 7840 6168
rect 7834 6128 7840 6140
rect 7892 6128 7898 6180
rect 8036 6168 8064 6276
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8386 6304 8392 6316
rect 8251 6276 8392 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 15562 6304 15568 6316
rect 15523 6276 15568 6304
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 18414 6264 18420 6316
rect 18472 6304 18478 6316
rect 19061 6307 19119 6313
rect 19061 6304 19073 6307
rect 18472 6276 19073 6304
rect 18472 6264 18478 6276
rect 19061 6273 19073 6276
rect 19107 6273 19119 6307
rect 19061 6267 19119 6273
rect 20622 6264 20628 6316
rect 20680 6304 20686 6316
rect 21821 6307 21879 6313
rect 21821 6304 21833 6307
rect 20680 6276 21833 6304
rect 20680 6264 20686 6276
rect 21821 6273 21833 6276
rect 21867 6273 21879 6307
rect 23658 6304 23664 6316
rect 23619 6276 23664 6304
rect 21821 6267 21879 6273
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 25038 6304 25044 6316
rect 24999 6276 25044 6304
rect 25038 6264 25044 6276
rect 25096 6264 25102 6316
rect 26326 6264 26332 6316
rect 26384 6304 26390 6316
rect 27801 6307 27859 6313
rect 27801 6304 27813 6307
rect 26384 6276 27813 6304
rect 26384 6264 26390 6276
rect 27801 6273 27813 6276
rect 27847 6273 27859 6307
rect 29638 6304 29644 6316
rect 29599 6276 29644 6304
rect 27801 6267 27859 6273
rect 29638 6264 29644 6276
rect 29696 6264 29702 6316
rect 30668 6313 30696 6344
rect 33060 6313 33088 6412
rect 36354 6400 36360 6452
rect 36412 6440 36418 6452
rect 36412 6412 38976 6440
rect 36412 6400 36418 6412
rect 35434 6332 35440 6384
rect 35492 6372 35498 6384
rect 36725 6375 36783 6381
rect 36725 6372 36737 6375
rect 35492 6344 36737 6372
rect 35492 6332 35498 6344
rect 36725 6341 36737 6344
rect 36771 6341 36783 6375
rect 36725 6335 36783 6341
rect 37642 6332 37648 6384
rect 37700 6372 37706 6384
rect 38948 6372 38976 6412
rect 50706 6400 50712 6452
rect 50764 6440 50770 6452
rect 60826 6440 60832 6452
rect 50764 6412 60832 6440
rect 50764 6400 50770 6412
rect 60826 6400 60832 6412
rect 60884 6400 60890 6452
rect 70213 6443 70271 6449
rect 70213 6440 70225 6443
rect 68664 6412 70225 6440
rect 37700 6344 38884 6372
rect 38948 6344 42748 6372
rect 37700 6332 37706 6344
rect 30653 6307 30711 6313
rect 30653 6273 30665 6307
rect 30699 6273 30711 6307
rect 30653 6267 30711 6273
rect 33045 6307 33103 6313
rect 33045 6273 33057 6307
rect 33091 6273 33103 6307
rect 37826 6304 37832 6316
rect 37787 6276 37832 6304
rect 33045 6267 33103 6273
rect 37826 6264 37832 6276
rect 37884 6264 37890 6316
rect 38856 6313 38884 6344
rect 38841 6307 38899 6313
rect 38841 6273 38853 6307
rect 38887 6273 38899 6307
rect 42610 6304 42616 6316
rect 42571 6276 42616 6304
rect 38841 6267 38899 6273
rect 42610 6264 42616 6276
rect 42668 6264 42674 6316
rect 42720 6304 42748 6344
rect 43714 6332 43720 6384
rect 43772 6372 43778 6384
rect 44634 6372 44640 6384
rect 43772 6344 44640 6372
rect 43772 6332 43778 6344
rect 44634 6332 44640 6344
rect 44692 6332 44698 6384
rect 52914 6332 52920 6384
rect 52972 6372 52978 6384
rect 52972 6344 54064 6372
rect 52972 6332 52978 6344
rect 44821 6307 44879 6313
rect 44821 6304 44833 6307
rect 42720 6276 44833 6304
rect 44821 6273 44833 6276
rect 44867 6273 44879 6307
rect 44821 6267 44879 6273
rect 47305 6307 47363 6313
rect 47305 6273 47317 6307
rect 47351 6273 47363 6307
rect 47305 6267 47363 6273
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6236 11391 6239
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 11379 6208 12449 6236
rect 11379 6205 11391 6208
rect 11333 6199 11391 6205
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 13538 6236 13544 6248
rect 13499 6208 13544 6236
rect 12437 6199 12495 6205
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 16666 6236 16672 6248
rect 16627 6208 16672 6236
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 18046 6236 18052 6248
rect 18007 6208 18052 6236
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 19426 6236 19432 6248
rect 19387 6208 19432 6236
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 20806 6236 20812 6248
rect 20767 6208 20812 6236
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 22005 6239 22063 6245
rect 22005 6236 22017 6239
rect 21928 6208 22017 6236
rect 21928 6180 21956 6208
rect 22005 6205 22017 6208
rect 22051 6205 22063 6239
rect 24854 6236 24860 6248
rect 24815 6208 24860 6236
rect 22005 6199 22063 6205
rect 24854 6196 24860 6208
rect 24912 6196 24918 6248
rect 26789 6239 26847 6245
rect 26789 6205 26801 6239
rect 26835 6236 26847 6239
rect 27614 6236 27620 6248
rect 26835 6208 27620 6236
rect 26835 6205 26847 6208
rect 26789 6199 26847 6205
rect 27614 6196 27620 6208
rect 27672 6196 27678 6248
rect 27890 6236 27896 6248
rect 27851 6208 27896 6236
rect 27890 6196 27896 6208
rect 27948 6196 27954 6248
rect 31205 6239 31263 6245
rect 31205 6205 31217 6239
rect 31251 6205 31263 6239
rect 31205 6199 31263 6205
rect 32033 6239 32091 6245
rect 32033 6205 32045 6239
rect 32079 6236 32091 6239
rect 32398 6236 32404 6248
rect 32079 6208 32404 6236
rect 32079 6205 32091 6208
rect 32033 6199 32091 6205
rect 13722 6168 13728 6180
rect 8036 6140 13728 6168
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 21910 6128 21916 6180
rect 21968 6128 21974 6180
rect 31220 6168 31248 6199
rect 32398 6196 32404 6208
rect 32456 6196 32462 6248
rect 33597 6239 33655 6245
rect 33597 6205 33609 6239
rect 33643 6236 33655 6239
rect 33870 6236 33876 6248
rect 33643 6208 33876 6236
rect 33643 6205 33655 6208
rect 33597 6199 33655 6205
rect 33870 6196 33876 6208
rect 33928 6196 33934 6248
rect 35437 6239 35495 6245
rect 35437 6205 35449 6239
rect 35483 6236 35495 6239
rect 36078 6236 36084 6248
rect 35483 6208 36084 6236
rect 35483 6205 35495 6208
rect 35437 6199 35495 6205
rect 36078 6196 36084 6208
rect 36136 6196 36142 6248
rect 36538 6236 36544 6248
rect 36499 6208 36544 6236
rect 36538 6196 36544 6208
rect 36596 6196 36602 6248
rect 39390 6236 39396 6248
rect 39351 6208 39396 6236
rect 39390 6196 39396 6208
rect 39448 6196 39454 6248
rect 43625 6239 43683 6245
rect 43625 6205 43637 6239
rect 43671 6236 43683 6239
rect 43990 6236 43996 6248
rect 43671 6208 43996 6236
rect 43671 6205 43683 6208
rect 43625 6199 43683 6205
rect 43990 6196 43996 6208
rect 44048 6196 44054 6248
rect 44266 6196 44272 6248
rect 44324 6236 44330 6248
rect 44729 6239 44787 6245
rect 44729 6236 44741 6239
rect 44324 6208 44741 6236
rect 44324 6196 44330 6208
rect 44729 6205 44741 6208
rect 44775 6205 44787 6239
rect 46106 6236 46112 6248
rect 46067 6208 46112 6236
rect 44729 6199 44787 6205
rect 46106 6196 46112 6208
rect 46164 6196 46170 6248
rect 47026 6196 47032 6248
rect 47084 6236 47090 6248
rect 47213 6239 47271 6245
rect 47213 6236 47225 6239
rect 47084 6208 47225 6236
rect 47084 6196 47090 6208
rect 47213 6205 47225 6208
rect 47259 6205 47271 6239
rect 47213 6199 47271 6205
rect 32766 6168 32772 6180
rect 31220 6140 32772 6168
rect 32766 6128 32772 6140
rect 32824 6128 32830 6180
rect 39850 6128 39856 6180
rect 39908 6168 39914 6180
rect 47320 6168 47348 6267
rect 49418 6264 49424 6316
rect 49476 6304 49482 6316
rect 49513 6307 49571 6313
rect 49513 6304 49525 6307
rect 49476 6276 49525 6304
rect 49476 6264 49482 6276
rect 49513 6273 49525 6276
rect 49559 6273 49571 6307
rect 53006 6304 53012 6316
rect 52967 6276 53012 6304
rect 49513 6267 49571 6273
rect 53006 6264 53012 6276
rect 53064 6264 53070 6316
rect 54036 6313 54064 6344
rect 57238 6332 57244 6384
rect 57296 6372 57302 6384
rect 57296 6344 60228 6372
rect 57296 6332 57302 6344
rect 54021 6307 54079 6313
rect 54021 6273 54033 6307
rect 54067 6273 54079 6307
rect 57330 6304 57336 6316
rect 57291 6276 57336 6304
rect 54021 6267 54079 6273
rect 57330 6264 57336 6276
rect 57388 6264 57394 6316
rect 60200 6313 60228 6344
rect 62114 6332 62120 6384
rect 62172 6372 62178 6384
rect 63681 6375 63739 6381
rect 63681 6372 63693 6375
rect 62172 6344 63693 6372
rect 62172 6332 62178 6344
rect 63681 6341 63693 6344
rect 63727 6341 63739 6375
rect 63681 6335 63739 6341
rect 66990 6332 66996 6384
rect 67048 6372 67054 6384
rect 68664 6372 68692 6412
rect 70213 6409 70225 6412
rect 70259 6409 70271 6443
rect 70213 6403 70271 6409
rect 73706 6400 73712 6452
rect 73764 6440 73770 6452
rect 106826 6440 106832 6452
rect 73764 6412 106832 6440
rect 73764 6400 73770 6412
rect 106826 6400 106832 6412
rect 106884 6400 106890 6452
rect 107657 6443 107715 6449
rect 107657 6409 107669 6443
rect 107703 6440 107715 6443
rect 108390 6440 108396 6452
rect 107703 6412 108396 6440
rect 107703 6409 107715 6412
rect 107657 6403 107715 6409
rect 108390 6400 108396 6412
rect 108448 6400 108454 6452
rect 110598 6400 110604 6452
rect 110656 6440 110662 6452
rect 110656 6412 119752 6440
rect 110656 6400 110662 6412
rect 67048 6344 68692 6372
rect 67048 6332 67054 6344
rect 68830 6332 68836 6384
rect 68888 6372 68894 6384
rect 68888 6344 69060 6372
rect 68888 6332 68894 6344
rect 60185 6307 60243 6313
rect 60185 6273 60197 6307
rect 60231 6273 60243 6307
rect 60185 6267 60243 6273
rect 64046 6264 64052 6316
rect 64104 6304 64110 6316
rect 66165 6307 66223 6313
rect 66165 6304 66177 6307
rect 64104 6276 66177 6304
rect 64104 6264 64110 6276
rect 66165 6273 66177 6276
rect 66211 6273 66223 6307
rect 67174 6304 67180 6316
rect 67135 6276 67180 6304
rect 66165 6267 66223 6273
rect 67174 6264 67180 6276
rect 67232 6264 67238 6316
rect 68925 6307 68983 6313
rect 68925 6304 68937 6307
rect 67284 6276 68937 6304
rect 48498 6236 48504 6248
rect 48459 6208 48504 6236
rect 48498 6196 48504 6208
rect 48556 6196 48562 6248
rect 49694 6236 49700 6248
rect 49655 6208 49700 6236
rect 49694 6196 49700 6208
rect 49752 6196 49758 6248
rect 54110 6236 54116 6248
rect 54071 6208 54116 6236
rect 54110 6196 54116 6208
rect 54168 6196 54174 6248
rect 59173 6239 59231 6245
rect 59173 6205 59185 6239
rect 59219 6205 59231 6239
rect 59173 6199 59231 6205
rect 39908 6140 47348 6168
rect 59188 6168 59216 6199
rect 59446 6196 59452 6248
rect 59504 6236 59510 6248
rect 60277 6239 60335 6245
rect 60277 6236 60289 6239
rect 59504 6208 60289 6236
rect 59504 6196 59510 6208
rect 60277 6205 60289 6208
rect 60323 6205 60335 6239
rect 63862 6236 63868 6248
rect 63823 6208 63868 6236
rect 60277 6199 60335 6205
rect 63862 6196 63868 6208
rect 63920 6196 63926 6248
rect 64325 6239 64383 6245
rect 64325 6205 64337 6239
rect 64371 6236 64383 6239
rect 64598 6236 64604 6248
rect 64371 6208 64604 6236
rect 64371 6205 64383 6208
rect 64325 6199 64383 6205
rect 64598 6196 64604 6208
rect 64656 6196 64662 6248
rect 64690 6196 64696 6248
rect 64748 6236 64754 6248
rect 65153 6239 65211 6245
rect 65153 6236 65165 6239
rect 64748 6208 65165 6236
rect 64748 6196 64754 6208
rect 65153 6205 65165 6208
rect 65199 6205 65211 6239
rect 65153 6199 65211 6205
rect 66898 6196 66904 6248
rect 66956 6236 66962 6248
rect 67284 6236 67312 6276
rect 68925 6273 68937 6276
rect 68971 6273 68983 6307
rect 69032 6304 69060 6344
rect 70946 6332 70952 6384
rect 71004 6372 71010 6384
rect 72050 6372 72056 6384
rect 71004 6344 72056 6372
rect 71004 6332 71010 6344
rect 72050 6332 72056 6344
rect 72108 6332 72114 6384
rect 72694 6332 72700 6384
rect 72752 6372 72758 6384
rect 74905 6375 74963 6381
rect 74905 6372 74917 6375
rect 72752 6344 74917 6372
rect 72752 6332 72758 6344
rect 74905 6341 74917 6344
rect 74951 6341 74963 6375
rect 78214 6372 78220 6384
rect 78175 6344 78220 6372
rect 74905 6335 74963 6341
rect 78214 6332 78220 6344
rect 78272 6332 78278 6384
rect 79318 6332 79324 6384
rect 79376 6372 79382 6384
rect 79873 6375 79931 6381
rect 79873 6372 79885 6375
rect 79376 6344 79885 6372
rect 79376 6332 79382 6344
rect 79873 6341 79885 6344
rect 79919 6341 79931 6375
rect 79873 6335 79931 6341
rect 79980 6344 80376 6372
rect 69032 6276 69152 6304
rect 68925 6267 68983 6273
rect 66956 6208 67312 6236
rect 68833 6239 68891 6245
rect 66956 6196 66962 6208
rect 68833 6205 68845 6239
rect 68879 6236 68891 6239
rect 69014 6236 69020 6248
rect 68879 6208 69020 6236
rect 68879 6205 68891 6208
rect 68833 6199 68891 6205
rect 69014 6196 69020 6208
rect 69072 6196 69078 6248
rect 69124 6245 69152 6276
rect 69566 6264 69572 6316
rect 69624 6304 69630 6316
rect 69624 6276 72280 6304
rect 69624 6264 69630 6276
rect 69109 6239 69167 6245
rect 69109 6205 69121 6239
rect 69155 6205 69167 6239
rect 69109 6199 69167 6205
rect 70394 6196 70400 6248
rect 70452 6236 70458 6248
rect 70670 6236 70676 6248
rect 70452 6208 70497 6236
rect 70631 6208 70676 6236
rect 70452 6196 70458 6208
rect 70670 6196 70676 6208
rect 70728 6196 70734 6248
rect 71774 6236 71780 6248
rect 71735 6208 71780 6236
rect 71774 6196 71780 6208
rect 71832 6196 71838 6248
rect 71866 6196 71872 6248
rect 71924 6236 71930 6248
rect 72252 6245 72280 6276
rect 73338 6264 73344 6316
rect 73396 6304 73402 6316
rect 76745 6307 76803 6313
rect 73396 6276 74948 6304
rect 73396 6264 73402 6276
rect 72053 6239 72111 6245
rect 72053 6236 72065 6239
rect 71924 6208 72065 6236
rect 71924 6196 71930 6208
rect 72053 6205 72065 6208
rect 72099 6205 72111 6239
rect 72053 6199 72111 6205
rect 72237 6239 72295 6245
rect 72237 6205 72249 6239
rect 72283 6205 72295 6239
rect 72237 6199 72295 6205
rect 74721 6239 74779 6245
rect 74721 6205 74733 6239
rect 74767 6236 74779 6239
rect 74813 6239 74871 6245
rect 74813 6236 74825 6239
rect 74767 6208 74825 6236
rect 74767 6205 74779 6208
rect 74721 6199 74779 6205
rect 74813 6205 74825 6208
rect 74859 6205 74871 6239
rect 74920 6236 74948 6276
rect 76745 6273 76757 6307
rect 76791 6304 76803 6307
rect 77294 6304 77300 6316
rect 76791 6276 77300 6304
rect 76791 6273 76803 6276
rect 76745 6267 76803 6273
rect 77294 6264 77300 6276
rect 77352 6264 77358 6316
rect 79042 6264 79048 6316
rect 79100 6304 79106 6316
rect 79980 6304 80008 6344
rect 79100 6276 80008 6304
rect 79100 6264 79106 6276
rect 75365 6239 75423 6245
rect 75365 6236 75377 6239
rect 74920 6208 75377 6236
rect 74813 6199 74871 6205
rect 75365 6205 75377 6208
rect 75411 6205 75423 6239
rect 76650 6236 76656 6248
rect 76611 6208 76656 6236
rect 75365 6199 75423 6205
rect 76650 6196 76656 6208
rect 76708 6196 76714 6248
rect 77113 6239 77171 6245
rect 77113 6205 77125 6239
rect 77159 6236 77171 6239
rect 77754 6236 77760 6248
rect 77159 6208 77760 6236
rect 77159 6205 77171 6208
rect 77113 6199 77171 6205
rect 77754 6196 77760 6208
rect 77812 6196 77818 6248
rect 78398 6236 78404 6248
rect 78359 6208 78404 6236
rect 78398 6196 78404 6208
rect 78456 6196 78462 6248
rect 78861 6239 78919 6245
rect 78861 6205 78873 6239
rect 78907 6236 78919 6239
rect 79870 6236 79876 6248
rect 78907 6208 79876 6236
rect 78907 6205 78919 6208
rect 78861 6199 78919 6205
rect 79870 6196 79876 6208
rect 79928 6196 79934 6248
rect 80054 6196 80060 6248
rect 80112 6236 80118 6248
rect 80348 6245 80376 6344
rect 81986 6332 81992 6384
rect 82044 6372 82050 6384
rect 83001 6375 83059 6381
rect 83001 6372 83013 6375
rect 82044 6344 83013 6372
rect 82044 6332 82050 6344
rect 83001 6341 83013 6344
rect 83047 6341 83059 6375
rect 83001 6335 83059 6341
rect 88426 6332 88432 6384
rect 88484 6372 88490 6384
rect 88797 6375 88855 6381
rect 88797 6372 88809 6375
rect 88484 6344 88809 6372
rect 88484 6332 88490 6344
rect 88797 6341 88809 6344
rect 88843 6341 88855 6375
rect 88797 6335 88855 6341
rect 89254 6332 89260 6384
rect 89312 6372 89318 6384
rect 91189 6375 91247 6381
rect 91189 6372 91201 6375
rect 89312 6344 91201 6372
rect 89312 6332 89318 6344
rect 91189 6341 91201 6344
rect 91235 6341 91247 6375
rect 91738 6372 91744 6384
rect 91189 6335 91247 6341
rect 91296 6344 91744 6372
rect 89806 6304 89812 6316
rect 88996 6276 89812 6304
rect 80333 6239 80391 6245
rect 80112 6208 80157 6236
rect 80112 6196 80118 6208
rect 80333 6205 80345 6239
rect 80379 6205 80391 6239
rect 81434 6236 81440 6248
rect 81395 6208 81440 6236
rect 80333 6199 80391 6205
rect 81434 6196 81440 6208
rect 81492 6196 81498 6248
rect 81710 6236 81716 6248
rect 81671 6208 81716 6236
rect 81710 6196 81716 6208
rect 81768 6196 81774 6248
rect 81894 6236 81900 6248
rect 81855 6208 81900 6236
rect 81894 6196 81900 6208
rect 81952 6196 81958 6248
rect 82906 6236 82912 6248
rect 82867 6208 82912 6236
rect 82906 6196 82912 6208
rect 82964 6196 82970 6248
rect 83458 6236 83464 6248
rect 83419 6208 83464 6236
rect 83458 6196 83464 6208
rect 83516 6196 83522 6248
rect 85206 6196 85212 6248
rect 85264 6236 85270 6248
rect 85393 6239 85451 6245
rect 85393 6236 85405 6239
rect 85264 6208 85405 6236
rect 85264 6196 85270 6208
rect 85393 6205 85405 6208
rect 85439 6205 85451 6239
rect 85758 6236 85764 6248
rect 85719 6208 85764 6236
rect 85393 6199 85451 6205
rect 85758 6196 85764 6208
rect 85816 6196 85822 6248
rect 86129 6239 86187 6245
rect 86129 6205 86141 6239
rect 86175 6236 86187 6239
rect 86862 6236 86868 6248
rect 86175 6208 86868 6236
rect 86175 6205 86187 6208
rect 86129 6199 86187 6205
rect 86862 6196 86868 6208
rect 86920 6196 86926 6248
rect 87138 6236 87144 6248
rect 87099 6208 87144 6236
rect 87138 6196 87144 6208
rect 87196 6196 87202 6248
rect 87414 6196 87420 6248
rect 87472 6236 87478 6248
rect 87509 6239 87567 6245
rect 87509 6236 87521 6239
rect 87472 6208 87521 6236
rect 87472 6196 87478 6208
rect 87509 6205 87521 6208
rect 87555 6205 87567 6239
rect 87509 6199 87567 6205
rect 87877 6239 87935 6245
rect 87877 6205 87889 6239
rect 87923 6236 87935 6239
rect 88150 6236 88156 6248
rect 87923 6208 88156 6236
rect 87923 6205 87935 6208
rect 87877 6199 87935 6205
rect 88150 6196 88156 6208
rect 88208 6196 88214 6248
rect 88996 6245 89024 6276
rect 89806 6264 89812 6276
rect 89864 6264 89870 6316
rect 88981 6239 89039 6245
rect 88981 6205 88993 6239
rect 89027 6205 89039 6239
rect 88981 6199 89039 6205
rect 89162 6196 89168 6248
rect 89220 6236 89226 6248
rect 89257 6239 89315 6245
rect 89257 6236 89269 6239
rect 89220 6208 89269 6236
rect 89220 6196 89226 6208
rect 89257 6205 89269 6208
rect 89303 6205 89315 6239
rect 89257 6199 89315 6205
rect 61565 6171 61623 6177
rect 61565 6168 61577 6171
rect 59188 6140 61577 6168
rect 39908 6128 39914 6140
rect 61565 6137 61577 6140
rect 61611 6137 61623 6171
rect 61565 6131 61623 6137
rect 61838 6128 61844 6180
rect 61896 6168 61902 6180
rect 81802 6168 81808 6180
rect 61896 6140 81808 6168
rect 61896 6128 61902 6140
rect 81802 6128 81808 6140
rect 81860 6128 81866 6180
rect 82170 6128 82176 6180
rect 82228 6168 82234 6180
rect 91296 6168 91324 6344
rect 91738 6332 91744 6344
rect 91796 6332 91802 6384
rect 95142 6332 95148 6384
rect 95200 6372 95206 6384
rect 95200 6344 99236 6372
rect 95200 6332 95206 6344
rect 97534 6304 97540 6316
rect 91388 6276 97540 6304
rect 91388 6245 91416 6276
rect 97534 6264 97540 6276
rect 97592 6264 97598 6316
rect 99208 6304 99236 6344
rect 99282 6332 99288 6384
rect 99340 6372 99346 6384
rect 99340 6344 100064 6372
rect 99340 6332 99346 6344
rect 99926 6304 99932 6316
rect 99208 6276 99932 6304
rect 99926 6264 99932 6276
rect 99984 6264 99990 6316
rect 100036 6313 100064 6344
rect 100110 6332 100116 6384
rect 100168 6372 100174 6384
rect 100168 6344 106412 6372
rect 100168 6332 100174 6344
rect 100021 6307 100079 6313
rect 100021 6273 100033 6307
rect 100067 6273 100079 6307
rect 100021 6267 100079 6273
rect 100570 6264 100576 6316
rect 100628 6304 100634 6316
rect 102597 6307 102655 6313
rect 102597 6304 102609 6307
rect 100628 6276 102609 6304
rect 100628 6264 100634 6276
rect 102597 6273 102609 6276
rect 102643 6273 102655 6307
rect 104710 6304 104716 6316
rect 102597 6267 102655 6273
rect 102980 6276 104716 6304
rect 91373 6239 91431 6245
rect 91373 6205 91385 6239
rect 91419 6205 91431 6239
rect 91373 6199 91431 6205
rect 91554 6196 91560 6248
rect 91612 6236 91618 6248
rect 91649 6239 91707 6245
rect 91649 6236 91661 6239
rect 91612 6208 91661 6236
rect 91612 6196 91618 6208
rect 91649 6205 91661 6208
rect 91695 6205 91707 6239
rect 92934 6236 92940 6248
rect 92895 6208 92940 6236
rect 91649 6199 91707 6205
rect 92934 6196 92940 6208
rect 92992 6196 92998 6248
rect 93118 6196 93124 6248
rect 93176 6236 93182 6248
rect 93305 6239 93363 6245
rect 93305 6236 93317 6239
rect 93176 6208 93317 6236
rect 93176 6196 93182 6208
rect 93305 6205 93317 6208
rect 93351 6205 93363 6239
rect 93305 6199 93363 6205
rect 93673 6239 93731 6245
rect 93673 6205 93685 6239
rect 93719 6236 93731 6239
rect 93854 6236 93860 6248
rect 93719 6208 93860 6236
rect 93719 6205 93731 6208
rect 93673 6199 93731 6205
rect 93854 6196 93860 6208
rect 93912 6196 93918 6248
rect 94958 6236 94964 6248
rect 94919 6208 94964 6236
rect 94958 6196 94964 6208
rect 95016 6196 95022 6248
rect 95142 6236 95148 6248
rect 95103 6208 95148 6236
rect 95142 6196 95148 6208
rect 95200 6196 95206 6248
rect 95513 6239 95571 6245
rect 95513 6205 95525 6239
rect 95559 6236 95571 6239
rect 96798 6236 96804 6248
rect 95559 6208 96804 6236
rect 95559 6205 95571 6208
rect 95513 6199 95571 6205
rect 96798 6196 96804 6208
rect 96856 6196 96862 6248
rect 97077 6239 97135 6245
rect 97077 6205 97089 6239
rect 97123 6205 97135 6239
rect 97077 6199 97135 6205
rect 97261 6239 97319 6245
rect 97261 6205 97273 6239
rect 97307 6236 97319 6239
rect 97350 6236 97356 6248
rect 97307 6208 97356 6236
rect 97307 6205 97319 6208
rect 97261 6199 97319 6205
rect 82228 6140 91324 6168
rect 82228 6128 82234 6140
rect 91738 6128 91744 6180
rect 91796 6168 91802 6180
rect 96890 6168 96896 6180
rect 91796 6140 96896 6168
rect 91796 6128 91802 6140
rect 96890 6128 96896 6140
rect 96948 6128 96954 6180
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 6822 6100 6828 6112
rect 3292 6072 6828 6100
rect 3292 6060 3298 6072
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 9217 6103 9275 6109
rect 9217 6100 9229 6103
rect 6972 6072 9229 6100
rect 6972 6060 6978 6072
rect 9217 6069 9229 6072
rect 9263 6069 9275 6103
rect 9217 6063 9275 6069
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 9732 6072 10241 6100
rect 9732 6060 9738 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 10229 6063 10287 6069
rect 21542 6060 21548 6112
rect 21600 6100 21606 6112
rect 22462 6100 22468 6112
rect 21600 6072 22468 6100
rect 21600 6060 21606 6072
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 29822 6060 29828 6112
rect 29880 6100 29886 6112
rect 30374 6100 30380 6112
rect 29880 6072 30380 6100
rect 29880 6060 29886 6072
rect 30374 6060 30380 6072
rect 30432 6060 30438 6112
rect 45462 6060 45468 6112
rect 45520 6100 45526 6112
rect 50430 6100 50436 6112
rect 45520 6072 50436 6100
rect 45520 6060 45526 6072
rect 50430 6060 50436 6072
rect 50488 6060 50494 6112
rect 50522 6060 50528 6112
rect 50580 6100 50586 6112
rect 51721 6103 51779 6109
rect 51721 6100 51733 6103
rect 50580 6072 51733 6100
rect 50580 6060 50586 6072
rect 51721 6069 51733 6072
rect 51767 6069 51779 6103
rect 51721 6063 51779 6069
rect 54570 6060 54576 6112
rect 54628 6100 54634 6112
rect 55401 6103 55459 6109
rect 55401 6100 55413 6103
rect 54628 6072 55413 6100
rect 54628 6060 54634 6072
rect 55401 6069 55413 6072
rect 55447 6069 55459 6103
rect 55401 6063 55459 6069
rect 56778 6060 56784 6112
rect 56836 6100 56842 6112
rect 59170 6100 59176 6112
rect 56836 6072 59176 6100
rect 56836 6060 56842 6072
rect 59170 6060 59176 6072
rect 59228 6060 59234 6112
rect 59814 6060 59820 6112
rect 59872 6100 59878 6112
rect 61930 6100 61936 6112
rect 59872 6072 61936 6100
rect 59872 6060 59878 6072
rect 61930 6060 61936 6072
rect 61988 6060 61994 6112
rect 67726 6060 67732 6112
rect 67784 6100 67790 6112
rect 69106 6100 69112 6112
rect 67784 6072 69112 6100
rect 67784 6060 67790 6072
rect 69106 6060 69112 6072
rect 69164 6060 69170 6112
rect 74721 6103 74779 6109
rect 74721 6069 74733 6103
rect 74767 6100 74779 6103
rect 77018 6100 77024 6112
rect 74767 6072 77024 6100
rect 74767 6069 74779 6072
rect 74721 6063 74779 6069
rect 77018 6060 77024 6072
rect 77076 6060 77082 6112
rect 91554 6060 91560 6112
rect 91612 6100 91618 6112
rect 96982 6100 96988 6112
rect 91612 6072 96988 6100
rect 91612 6060 91618 6072
rect 96982 6060 96988 6072
rect 97040 6060 97046 6112
rect 97092 6100 97120 6199
rect 97350 6196 97356 6208
rect 97408 6196 97414 6248
rect 97629 6239 97687 6245
rect 97629 6205 97641 6239
rect 97675 6236 97687 6239
rect 97994 6236 98000 6248
rect 97675 6208 98000 6236
rect 97675 6205 97687 6208
rect 97629 6199 97687 6205
rect 97994 6196 98000 6208
rect 98052 6196 98058 6248
rect 98638 6236 98644 6248
rect 98599 6208 98644 6236
rect 98638 6196 98644 6208
rect 98696 6196 98702 6248
rect 98822 6236 98828 6248
rect 98783 6208 98828 6236
rect 98822 6196 98828 6208
rect 98880 6196 98886 6248
rect 99193 6239 99251 6245
rect 99193 6205 99205 6239
rect 99239 6236 99251 6239
rect 99466 6236 99472 6248
rect 99239 6208 99472 6236
rect 99239 6205 99251 6208
rect 99193 6199 99251 6205
rect 99466 6196 99472 6208
rect 99524 6196 99530 6248
rect 102980 6245 103008 6276
rect 104710 6264 104716 6276
rect 104768 6264 104774 6316
rect 105265 6307 105323 6313
rect 105265 6273 105277 6307
rect 105311 6273 105323 6307
rect 106274 6304 106280 6316
rect 106235 6276 106280 6304
rect 105265 6267 105323 6273
rect 102505 6239 102563 6245
rect 102505 6205 102517 6239
rect 102551 6205 102563 6239
rect 102505 6199 102563 6205
rect 102965 6239 103023 6245
rect 102965 6205 102977 6239
rect 103011 6205 103023 6239
rect 103882 6236 103888 6248
rect 103843 6208 103888 6236
rect 102965 6199 103023 6205
rect 101033 6171 101091 6177
rect 101033 6168 101045 6171
rect 99944 6140 101045 6168
rect 99006 6100 99012 6112
rect 97092 6072 99012 6100
rect 99006 6060 99012 6072
rect 99064 6060 99070 6112
rect 99282 6060 99288 6112
rect 99340 6100 99346 6112
rect 99944 6100 99972 6140
rect 101033 6137 101045 6140
rect 101079 6137 101091 6171
rect 101033 6131 101091 6137
rect 99340 6072 99972 6100
rect 99340 6060 99346 6072
rect 100018 6060 100024 6112
rect 100076 6100 100082 6112
rect 101214 6100 101220 6112
rect 100076 6072 101220 6100
rect 100076 6060 100082 6072
rect 101214 6060 101220 6072
rect 101272 6060 101278 6112
rect 102520 6100 102548 6199
rect 103882 6196 103888 6208
rect 103940 6196 103946 6248
rect 105280 6168 105308 6267
rect 106274 6264 106280 6276
rect 106332 6264 106338 6316
rect 106384 6304 106412 6344
rect 106550 6332 106556 6384
rect 106608 6372 106614 6384
rect 108574 6372 108580 6384
rect 106608 6344 108580 6372
rect 106608 6332 106614 6344
rect 108574 6332 108580 6344
rect 108632 6332 108638 6384
rect 108666 6332 108672 6384
rect 108724 6372 108730 6384
rect 108724 6344 110000 6372
rect 108724 6332 108730 6344
rect 109862 6304 109868 6316
rect 106384 6276 109868 6304
rect 109862 6264 109868 6276
rect 109920 6264 109926 6316
rect 105354 6196 105360 6248
rect 105412 6236 105418 6248
rect 105412 6208 105457 6236
rect 105412 6196 105418 6208
rect 105538 6196 105544 6248
rect 105596 6236 105602 6248
rect 107657 6239 107715 6245
rect 107657 6236 107669 6239
rect 105596 6208 107669 6236
rect 105596 6196 105602 6208
rect 107657 6205 107669 6208
rect 107703 6205 107715 6239
rect 108022 6236 108028 6248
rect 107983 6208 108028 6236
rect 107657 6199 107715 6205
rect 108022 6196 108028 6208
rect 108080 6196 108086 6248
rect 108206 6236 108212 6248
rect 108167 6208 108212 6236
rect 108206 6196 108212 6208
rect 108264 6196 108270 6248
rect 108390 6236 108396 6248
rect 108351 6208 108396 6236
rect 108390 6196 108396 6208
rect 108448 6196 108454 6248
rect 109586 6236 109592 6248
rect 109547 6208 109592 6236
rect 109586 6196 109592 6208
rect 109644 6196 109650 6248
rect 109770 6236 109776 6248
rect 109731 6208 109776 6236
rect 109770 6196 109776 6208
rect 109828 6196 109834 6248
rect 109972 6245 110000 6344
rect 110046 6332 110052 6384
rect 110104 6372 110110 6384
rect 111061 6375 111119 6381
rect 111061 6372 111073 6375
rect 110104 6344 111073 6372
rect 110104 6332 110110 6344
rect 111061 6341 111073 6344
rect 111107 6341 111119 6375
rect 111061 6335 111119 6341
rect 111242 6332 111248 6384
rect 111300 6372 111306 6384
rect 116026 6372 116032 6384
rect 111300 6344 116032 6372
rect 111300 6332 111306 6344
rect 116026 6332 116032 6344
rect 116084 6332 116090 6384
rect 116305 6375 116363 6381
rect 116305 6341 116317 6375
rect 116351 6372 116363 6375
rect 118789 6375 118847 6381
rect 118789 6372 118801 6375
rect 116351 6344 118801 6372
rect 116351 6341 116363 6344
rect 116305 6335 116363 6341
rect 118789 6341 118801 6344
rect 118835 6341 118847 6375
rect 118789 6335 118847 6341
rect 117777 6307 117835 6313
rect 110340 6276 117636 6304
rect 109957 6239 110015 6245
rect 109957 6205 109969 6239
rect 110003 6205 110015 6239
rect 109957 6199 110015 6205
rect 110340 6168 110368 6276
rect 111245 6239 111303 6245
rect 111245 6205 111257 6239
rect 111291 6236 111303 6239
rect 111426 6236 111432 6248
rect 111291 6208 111432 6236
rect 111291 6205 111303 6208
rect 111245 6199 111303 6205
rect 111426 6196 111432 6208
rect 111484 6196 111490 6248
rect 111705 6239 111763 6245
rect 111705 6205 111717 6239
rect 111751 6236 111763 6239
rect 112530 6236 112536 6248
rect 111751 6208 112536 6236
rect 111751 6205 111763 6208
rect 111705 6199 111763 6205
rect 112530 6196 112536 6208
rect 112588 6196 112594 6248
rect 113821 6239 113879 6245
rect 113821 6205 113833 6239
rect 113867 6236 113879 6239
rect 114833 6239 114891 6245
rect 114833 6236 114845 6239
rect 113867 6208 114845 6236
rect 113867 6205 113879 6208
rect 113821 6199 113879 6205
rect 114833 6205 114845 6208
rect 114879 6205 114891 6239
rect 116394 6236 116400 6248
rect 116355 6208 116400 6236
rect 114833 6199 114891 6205
rect 116394 6196 116400 6208
rect 116452 6196 116458 6248
rect 117498 6168 117504 6180
rect 105280 6140 110368 6168
rect 110432 6140 117504 6168
rect 106550 6100 106556 6112
rect 102520 6072 106556 6100
rect 106550 6060 106556 6072
rect 106608 6060 106614 6112
rect 106642 6060 106648 6112
rect 106700 6100 106706 6112
rect 107562 6100 107568 6112
rect 106700 6072 107568 6100
rect 106700 6060 106706 6072
rect 107562 6060 107568 6072
rect 107620 6060 107626 6112
rect 107654 6060 107660 6112
rect 107712 6100 107718 6112
rect 110432 6100 110460 6140
rect 117498 6128 117504 6140
rect 117556 6128 117562 6180
rect 117608 6168 117636 6276
rect 117777 6273 117789 6307
rect 117823 6304 117835 6307
rect 118694 6304 118700 6316
rect 117823 6276 118700 6304
rect 117823 6273 117835 6276
rect 117777 6267 117835 6273
rect 118694 6264 118700 6276
rect 118752 6264 118758 6316
rect 119062 6304 119068 6316
rect 119023 6276 119068 6304
rect 119062 6264 119068 6276
rect 119120 6264 119126 6316
rect 119724 6236 119752 6412
rect 119798 6400 119804 6452
rect 119856 6440 119862 6452
rect 122006 6440 122012 6452
rect 119856 6412 122012 6440
rect 119856 6400 119862 6412
rect 122006 6400 122012 6412
rect 122064 6400 122070 6452
rect 122098 6400 122104 6452
rect 122156 6440 122162 6452
rect 122742 6440 122748 6452
rect 122156 6412 122748 6440
rect 122156 6400 122162 6412
rect 122742 6400 122748 6412
rect 122800 6400 122806 6452
rect 123110 6400 123116 6452
rect 123168 6440 123174 6452
rect 126054 6440 126060 6452
rect 123168 6412 126060 6440
rect 123168 6400 123174 6412
rect 126054 6400 126060 6412
rect 126112 6400 126118 6452
rect 126164 6412 131896 6440
rect 124398 6332 124404 6384
rect 124456 6372 124462 6384
rect 126164 6381 126192 6412
rect 126149 6375 126207 6381
rect 124456 6344 126100 6372
rect 124456 6332 124462 6344
rect 120534 6304 120540 6316
rect 120495 6276 120540 6304
rect 120534 6264 120540 6276
rect 120592 6264 120598 6316
rect 121454 6304 121460 6316
rect 121415 6276 121460 6304
rect 121454 6264 121460 6276
rect 121512 6264 121518 6316
rect 122929 6307 122987 6313
rect 122929 6273 122941 6307
rect 122975 6304 122987 6307
rect 125962 6304 125968 6316
rect 122975 6276 125968 6304
rect 122975 6273 122987 6276
rect 122929 6267 122987 6273
rect 125962 6264 125968 6276
rect 126020 6264 126026 6316
rect 126072 6304 126100 6344
rect 126149 6341 126161 6375
rect 126195 6341 126207 6375
rect 128633 6375 128691 6381
rect 126149 6335 126207 6341
rect 126256 6344 128584 6372
rect 126256 6304 126284 6344
rect 126072 6276 126284 6304
rect 127161 6307 127219 6313
rect 127161 6273 127173 6307
rect 127207 6304 127219 6307
rect 128262 6304 128268 6316
rect 127207 6276 128268 6304
rect 127207 6273 127219 6276
rect 127161 6267 127219 6273
rect 128262 6264 128268 6276
rect 128320 6264 128326 6316
rect 128556 6304 128584 6344
rect 128633 6341 128645 6375
rect 128679 6372 128691 6375
rect 131758 6372 131764 6384
rect 128679 6344 131764 6372
rect 128679 6341 128691 6344
rect 128633 6335 128691 6341
rect 131758 6332 131764 6344
rect 131816 6332 131822 6384
rect 131868 6372 131896 6412
rect 131942 6400 131948 6452
rect 132000 6440 132006 6452
rect 138290 6440 138296 6452
rect 132000 6412 138296 6440
rect 132000 6400 132006 6412
rect 138290 6400 138296 6412
rect 138348 6400 138354 6452
rect 149974 6440 149980 6452
rect 139964 6412 149980 6440
rect 139964 6381 139992 6412
rect 149974 6400 149980 6412
rect 150032 6400 150038 6452
rect 139949 6375 140007 6381
rect 131868 6344 139900 6372
rect 131393 6307 131451 6313
rect 128556 6276 131068 6304
rect 119724 6208 120212 6236
rect 120074 6168 120080 6180
rect 117608 6140 120080 6168
rect 120074 6128 120080 6140
rect 120132 6128 120138 6180
rect 120184 6168 120212 6208
rect 120626 6196 120632 6248
rect 120684 6236 120690 6248
rect 120684 6208 120729 6236
rect 120684 6196 120690 6208
rect 120810 6196 120816 6248
rect 120868 6236 120874 6248
rect 122834 6236 122840 6248
rect 120868 6208 122328 6236
rect 122795 6208 122840 6236
rect 120868 6196 120874 6208
rect 122300 6168 122328 6208
rect 122834 6196 122840 6208
rect 122892 6196 122898 6248
rect 123754 6196 123760 6248
rect 123812 6236 123818 6248
rect 124398 6236 124404 6248
rect 123812 6208 124404 6236
rect 123812 6196 123818 6208
rect 124398 6196 124404 6208
rect 124456 6196 124462 6248
rect 124674 6236 124680 6248
rect 124635 6208 124680 6236
rect 124674 6196 124680 6208
rect 124732 6196 124738 6248
rect 125778 6236 125784 6248
rect 125739 6208 125784 6236
rect 125778 6196 125784 6208
rect 125836 6196 125842 6248
rect 128725 6239 128783 6245
rect 128725 6205 128737 6239
rect 128771 6236 128783 6239
rect 130930 6236 130936 6248
rect 128771 6208 130936 6236
rect 128771 6205 128783 6208
rect 128725 6199 128783 6205
rect 130930 6196 130936 6208
rect 130988 6196 130994 6248
rect 131040 6236 131068 6276
rect 131393 6273 131405 6307
rect 131439 6304 131451 6307
rect 132586 6304 132592 6316
rect 131439 6276 132592 6304
rect 131439 6273 131451 6276
rect 131393 6267 131451 6273
rect 132586 6264 132592 6276
rect 132644 6264 132650 6316
rect 132770 6304 132776 6316
rect 132731 6276 132776 6304
rect 132770 6264 132776 6276
rect 132828 6264 132834 6316
rect 133598 6304 133604 6316
rect 132880 6276 133604 6304
rect 132218 6236 132224 6248
rect 131040 6208 132224 6236
rect 132218 6196 132224 6208
rect 132276 6196 132282 6248
rect 120184 6140 120948 6168
rect 122300 6140 127756 6168
rect 107712 6072 110460 6100
rect 107712 6060 107718 6072
rect 113542 6060 113548 6112
rect 113600 6100 113606 6112
rect 118602 6100 118608 6112
rect 113600 6072 118608 6100
rect 113600 6060 113606 6072
rect 118602 6060 118608 6072
rect 118660 6060 118666 6112
rect 118789 6103 118847 6109
rect 118789 6069 118801 6103
rect 118835 6100 118847 6103
rect 120810 6100 120816 6112
rect 118835 6072 120816 6100
rect 118835 6069 118847 6072
rect 118789 6063 118847 6069
rect 120810 6060 120816 6072
rect 120868 6060 120874 6112
rect 120920 6100 120948 6140
rect 125502 6100 125508 6112
rect 120920 6072 125508 6100
rect 125502 6060 125508 6072
rect 125560 6060 125566 6112
rect 125686 6060 125692 6112
rect 125744 6100 125750 6112
rect 127618 6100 127624 6112
rect 125744 6072 127624 6100
rect 125744 6060 125750 6072
rect 127618 6060 127624 6072
rect 127676 6060 127682 6112
rect 127728 6100 127756 6140
rect 130194 6128 130200 6180
rect 130252 6168 130258 6180
rect 130252 6140 131252 6168
rect 130252 6128 130258 6140
rect 129182 6100 129188 6112
rect 127728 6072 129188 6100
rect 129182 6060 129188 6072
rect 129240 6060 129246 6112
rect 130289 6103 130347 6109
rect 130289 6069 130301 6103
rect 130335 6100 130347 6103
rect 131114 6100 131120 6112
rect 130335 6072 131120 6100
rect 130335 6069 130347 6072
rect 130289 6063 130347 6069
rect 131114 6060 131120 6072
rect 131172 6060 131178 6112
rect 131224 6100 131252 6140
rect 131574 6128 131580 6180
rect 131632 6168 131638 6180
rect 132880 6168 132908 6276
rect 133598 6264 133604 6276
rect 133656 6264 133662 6316
rect 133966 6264 133972 6316
rect 134024 6304 134030 6316
rect 135898 6304 135904 6316
rect 134024 6276 135904 6304
rect 134024 6264 134030 6276
rect 135898 6264 135904 6276
rect 135956 6264 135962 6316
rect 136085 6307 136143 6313
rect 136085 6273 136097 6307
rect 136131 6304 136143 6307
rect 137554 6304 137560 6316
rect 136131 6276 137416 6304
rect 137515 6276 137560 6304
rect 136131 6273 136143 6276
rect 136085 6267 136143 6273
rect 132957 6239 133015 6245
rect 132957 6205 132969 6239
rect 133003 6236 133015 6239
rect 133506 6236 133512 6248
rect 133003 6208 133512 6236
rect 133003 6205 133015 6208
rect 132957 6199 133015 6205
rect 133506 6196 133512 6208
rect 133564 6196 133570 6248
rect 134426 6196 134432 6248
rect 134484 6236 134490 6248
rect 134484 6208 134932 6236
rect 134484 6196 134490 6208
rect 131632 6140 132908 6168
rect 132972 6140 133920 6168
rect 131632 6128 131638 6140
rect 132972 6100 133000 6140
rect 131224 6072 133000 6100
rect 133598 6060 133604 6112
rect 133656 6100 133662 6112
rect 133785 6103 133843 6109
rect 133785 6100 133797 6103
rect 133656 6072 133797 6100
rect 133656 6060 133662 6072
rect 133785 6069 133797 6072
rect 133831 6069 133843 6103
rect 133892 6100 133920 6140
rect 133966 6128 133972 6180
rect 134024 6168 134030 6180
rect 134797 6171 134855 6177
rect 134797 6168 134809 6171
rect 134024 6140 134809 6168
rect 134024 6128 134030 6140
rect 134797 6137 134809 6140
rect 134843 6137 134855 6171
rect 134904 6168 134932 6208
rect 134978 6196 134984 6248
rect 135036 6236 135042 6248
rect 136542 6236 136548 6248
rect 135036 6208 136548 6236
rect 135036 6196 135042 6208
rect 136542 6196 136548 6208
rect 136600 6196 136606 6248
rect 136726 6196 136732 6248
rect 136784 6236 136790 6248
rect 137189 6239 137247 6245
rect 137189 6236 137201 6239
rect 136784 6208 137201 6236
rect 136784 6196 136790 6208
rect 137189 6205 137201 6208
rect 137235 6205 137247 6239
rect 137388 6236 137416 6276
rect 137554 6264 137560 6276
rect 137612 6264 137618 6316
rect 139872 6304 139900 6344
rect 139949 6341 139961 6375
rect 139995 6341 140007 6375
rect 155310 6372 155316 6384
rect 139949 6335 140007 6341
rect 140056 6344 155316 6372
rect 140056 6304 140084 6344
rect 155310 6332 155316 6344
rect 155368 6332 155374 6384
rect 138308 6276 139716 6304
rect 139872 6276 140084 6304
rect 138308 6236 138336 6276
rect 138474 6236 138480 6248
rect 137388 6208 138336 6236
rect 138435 6208 138480 6236
rect 137189 6199 137247 6205
rect 138474 6196 138480 6208
rect 138532 6196 138538 6248
rect 139578 6236 139584 6248
rect 139539 6208 139584 6236
rect 139578 6196 139584 6208
rect 139636 6196 139642 6248
rect 139688 6236 139716 6276
rect 140498 6264 140504 6316
rect 140556 6304 140562 6316
rect 142525 6307 142583 6313
rect 142525 6304 142537 6307
rect 140556 6276 142537 6304
rect 140556 6264 140562 6276
rect 142525 6273 142537 6276
rect 142571 6273 142583 6307
rect 142525 6267 142583 6273
rect 142614 6264 142620 6316
rect 142672 6304 142678 6316
rect 145374 6304 145380 6316
rect 142672 6276 145236 6304
rect 145335 6276 145380 6304
rect 142672 6264 142678 6276
rect 141513 6239 141571 6245
rect 141513 6236 141525 6239
rect 139688 6208 141525 6236
rect 141513 6205 141525 6208
rect 141559 6205 141571 6239
rect 143902 6236 143908 6248
rect 143863 6208 143908 6236
rect 141513 6199 141571 6205
rect 143902 6196 143908 6208
rect 143960 6196 143966 6248
rect 145098 6236 145104 6248
rect 145059 6208 145104 6236
rect 145098 6196 145104 6208
rect 145156 6196 145162 6248
rect 145208 6236 145236 6276
rect 145374 6264 145380 6276
rect 145432 6264 145438 6316
rect 147125 6307 147183 6313
rect 147125 6273 147137 6307
rect 147171 6304 147183 6307
rect 147674 6304 147680 6316
rect 147171 6276 147680 6304
rect 147171 6273 147183 6276
rect 147125 6267 147183 6273
rect 147674 6264 147680 6276
rect 147732 6264 147738 6316
rect 150618 6304 150624 6316
rect 150579 6276 150624 6304
rect 150618 6264 150624 6276
rect 150676 6264 150682 6316
rect 151630 6304 151636 6316
rect 151591 6276 151636 6304
rect 151630 6264 151636 6276
rect 151688 6264 151694 6316
rect 153286 6304 153292 6316
rect 153247 6276 153292 6304
rect 153286 6264 153292 6276
rect 153344 6264 153350 6316
rect 153930 6236 153936 6248
rect 145208 6208 153936 6236
rect 153930 6196 153936 6208
rect 153988 6196 153994 6248
rect 134904 6140 135300 6168
rect 134797 6131 134855 6137
rect 134702 6100 134708 6112
rect 133892 6072 134708 6100
rect 133785 6063 133843 6069
rect 134702 6060 134708 6072
rect 134760 6060 134766 6112
rect 135272 6100 135300 6140
rect 135530 6128 135536 6180
rect 135588 6168 135594 6180
rect 152182 6168 152188 6180
rect 135588 6140 152188 6168
rect 135588 6128 135594 6140
rect 152182 6128 152188 6140
rect 152240 6128 152246 6180
rect 140406 6100 140412 6112
rect 135272 6072 140412 6100
rect 140406 6060 140412 6072
rect 140464 6060 140470 6112
rect 145098 6060 145104 6112
rect 145156 6100 145162 6112
rect 145834 6100 145840 6112
rect 145156 6072 145840 6100
rect 145156 6060 145162 6072
rect 145834 6060 145840 6072
rect 145892 6060 145898 6112
rect 1104 6010 154560 6032
rect 1104 5958 24078 6010
rect 24130 5958 64078 6010
rect 64130 5958 104078 6010
rect 104130 5958 144078 6010
rect 144130 5958 154560 6010
rect 1104 5936 154560 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 8297 5899 8355 5905
rect 8297 5896 8309 5899
rect 6788 5868 8309 5896
rect 6788 5856 6794 5868
rect 8297 5865 8309 5868
rect 8343 5865 8355 5899
rect 8297 5859 8355 5865
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 10134 5896 10140 5908
rect 8628 5868 10140 5896
rect 8628 5856 8634 5868
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 10226 5856 10232 5908
rect 10284 5896 10290 5908
rect 13446 5896 13452 5908
rect 10284 5868 13452 5896
rect 10284 5856 10290 5868
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 21082 5856 21088 5908
rect 21140 5896 21146 5908
rect 27614 5896 27620 5908
rect 21140 5868 22508 5896
rect 27575 5868 27620 5896
rect 21140 5856 21146 5868
rect 4706 5788 4712 5840
rect 4764 5828 4770 5840
rect 7285 5831 7343 5837
rect 7285 5828 7297 5831
rect 4764 5800 7297 5828
rect 4764 5788 4770 5800
rect 7285 5797 7297 5800
rect 7331 5797 7343 5831
rect 12250 5828 12256 5840
rect 7285 5791 7343 5797
rect 8680 5800 12256 5828
rect 6454 5760 6460 5772
rect 6415 5732 6460 5760
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 3007 5664 4905 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 4893 5661 4905 5664
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 7466 5692 7472 5704
rect 6411 5664 7472 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 3602 5584 3608 5636
rect 3660 5624 3666 5636
rect 8680 5624 8708 5800
rect 12250 5788 12256 5800
rect 12308 5788 12314 5840
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 9876 5732 10793 5760
rect 8938 5652 8944 5704
rect 8996 5692 9002 5704
rect 9876 5692 9904 5732
rect 10781 5729 10793 5732
rect 10827 5729 10839 5763
rect 13446 5760 13452 5772
rect 13407 5732 13452 5760
rect 10781 5723 10839 5729
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 14056 5732 15301 5760
rect 14056 5720 14062 5732
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 16393 5763 16451 5769
rect 16393 5729 16405 5763
rect 16439 5729 16451 5763
rect 19978 5760 19984 5772
rect 19939 5732 19984 5760
rect 16393 5723 16451 5729
rect 8996 5664 9904 5692
rect 8996 5652 9002 5664
rect 10594 5652 10600 5704
rect 10652 5692 10658 5704
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10652 5664 10701 5692
rect 10652 5652 10658 5664
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 12069 5695 12127 5701
rect 10928 5664 12020 5692
rect 10928 5652 10934 5664
rect 3660 5596 8708 5624
rect 3660 5584 3666 5596
rect 8754 5584 8760 5636
rect 8812 5624 8818 5636
rect 11882 5624 11888 5636
rect 8812 5596 11888 5624
rect 8812 5584 8818 5596
rect 11882 5584 11888 5596
rect 11940 5584 11946 5636
rect 11992 5624 12020 5664
rect 12069 5661 12081 5695
rect 12115 5692 12127 5695
rect 12434 5692 12440 5704
rect 12115 5664 12440 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 14090 5692 14096 5704
rect 13587 5664 14096 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14918 5652 14924 5704
rect 14976 5692 14982 5704
rect 16408 5692 16436 5723
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 21082 5720 21088 5772
rect 21140 5760 21146 5772
rect 22373 5763 22431 5769
rect 22373 5760 22385 5763
rect 21140 5732 22385 5760
rect 21140 5720 21146 5732
rect 22373 5729 22385 5732
rect 22419 5729 22431 5763
rect 22373 5723 22431 5729
rect 14976 5664 16436 5692
rect 16485 5695 16543 5701
rect 14976 5652 14982 5664
rect 16485 5661 16497 5695
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5692 18475 5695
rect 19334 5692 19340 5704
rect 18463 5664 19340 5692
rect 18463 5661 18475 5664
rect 18417 5655 18475 5661
rect 12802 5624 12808 5636
rect 11992 5596 12808 5624
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 16298 5584 16304 5636
rect 16356 5624 16362 5636
rect 16500 5624 16528 5655
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5692 19947 5695
rect 20162 5692 20168 5704
rect 19935 5664 20168 5692
rect 19935 5661 19947 5664
rect 19889 5655 19947 5661
rect 20162 5652 20168 5664
rect 20220 5652 20226 5704
rect 21266 5692 21272 5704
rect 21227 5664 21272 5692
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 22480 5701 22508 5868
rect 27614 5856 27620 5868
rect 27672 5856 27678 5908
rect 32398 5896 32404 5908
rect 32359 5868 32404 5896
rect 32398 5856 32404 5868
rect 32456 5856 32462 5908
rect 36078 5896 36084 5908
rect 36039 5868 36084 5896
rect 36078 5856 36084 5868
rect 36136 5856 36142 5908
rect 43990 5896 43996 5908
rect 43951 5868 43996 5896
rect 43990 5856 43996 5868
rect 44048 5856 44054 5908
rect 46106 5856 46112 5908
rect 46164 5896 46170 5908
rect 47397 5899 47455 5905
rect 47397 5896 47409 5899
rect 46164 5868 47409 5896
rect 46164 5856 46170 5868
rect 47397 5865 47409 5868
rect 47443 5865 47455 5899
rect 47397 5859 47455 5865
rect 53742 5856 53748 5908
rect 53800 5896 53806 5908
rect 67082 5896 67088 5908
rect 53800 5868 67088 5896
rect 53800 5856 53806 5868
rect 67082 5856 67088 5868
rect 67140 5856 67146 5908
rect 68094 5856 68100 5908
rect 68152 5896 68158 5908
rect 70670 5896 70676 5908
rect 68152 5868 70676 5896
rect 68152 5856 68158 5868
rect 70670 5856 70676 5868
rect 70728 5856 70734 5908
rect 82538 5856 82544 5908
rect 82596 5896 82602 5908
rect 83366 5896 83372 5908
rect 82596 5868 83372 5896
rect 82596 5856 82602 5868
rect 83366 5856 83372 5868
rect 83424 5856 83430 5908
rect 85206 5896 85212 5908
rect 85167 5868 85212 5896
rect 85206 5856 85212 5868
rect 85264 5856 85270 5908
rect 89714 5856 89720 5908
rect 89772 5896 89778 5908
rect 99466 5896 99472 5908
rect 89772 5868 99472 5896
rect 89772 5856 89778 5868
rect 99466 5856 99472 5868
rect 99524 5856 99530 5908
rect 99650 5856 99656 5908
rect 99708 5896 99714 5908
rect 100481 5899 100539 5905
rect 100481 5896 100493 5899
rect 99708 5868 100493 5896
rect 99708 5856 99714 5868
rect 100481 5865 100493 5868
rect 100527 5865 100539 5899
rect 100481 5859 100539 5865
rect 101861 5899 101919 5905
rect 101861 5865 101873 5899
rect 101907 5896 101919 5899
rect 103882 5896 103888 5908
rect 101907 5868 103888 5896
rect 101907 5865 101919 5868
rect 101861 5859 101919 5865
rect 103882 5856 103888 5868
rect 103940 5856 103946 5908
rect 105078 5896 105084 5908
rect 105039 5868 105084 5896
rect 105078 5856 105084 5868
rect 105136 5856 105142 5908
rect 105354 5856 105360 5908
rect 105412 5896 105418 5908
rect 108942 5896 108948 5908
rect 105412 5868 108948 5896
rect 105412 5856 105418 5868
rect 108942 5856 108948 5868
rect 109000 5856 109006 5908
rect 109126 5856 109132 5908
rect 109184 5896 109190 5908
rect 115014 5896 115020 5908
rect 109184 5868 115020 5896
rect 109184 5856 109190 5868
rect 115014 5856 115020 5868
rect 115072 5856 115078 5908
rect 115106 5856 115112 5908
rect 115164 5896 115170 5908
rect 115164 5868 119936 5896
rect 115164 5856 115170 5868
rect 24578 5788 24584 5840
rect 24636 5828 24642 5840
rect 24636 5800 29684 5828
rect 24636 5788 24642 5800
rect 25038 5760 25044 5772
rect 24999 5732 25044 5760
rect 25038 5720 25044 5732
rect 25096 5720 25102 5772
rect 28626 5760 28632 5772
rect 28587 5732 28632 5760
rect 28626 5720 28632 5732
rect 28684 5720 28690 5772
rect 29656 5701 29684 5800
rect 34330 5788 34336 5840
rect 34388 5828 34394 5840
rect 34606 5828 34612 5840
rect 34388 5800 34612 5828
rect 34388 5788 34394 5800
rect 34606 5788 34612 5800
rect 34664 5788 34670 5840
rect 46750 5788 46756 5840
rect 46808 5828 46814 5840
rect 47118 5828 47124 5840
rect 46808 5800 47124 5828
rect 46808 5788 46814 5800
rect 47118 5788 47124 5800
rect 47176 5788 47182 5840
rect 58986 5788 58992 5840
rect 59044 5828 59050 5840
rect 59044 5800 63356 5828
rect 59044 5788 59050 5800
rect 29730 5720 29736 5772
rect 29788 5760 29794 5772
rect 29788 5732 29833 5760
rect 29788 5720 29794 5732
rect 30558 5720 30564 5772
rect 30616 5760 30622 5772
rect 31938 5760 31944 5772
rect 30616 5732 31944 5760
rect 30616 5720 30622 5732
rect 31938 5720 31944 5732
rect 31996 5720 32002 5772
rect 33594 5720 33600 5772
rect 33652 5760 33658 5772
rect 34517 5763 34575 5769
rect 34517 5760 34529 5763
rect 33652 5732 34529 5760
rect 33652 5720 33658 5732
rect 34517 5729 34529 5732
rect 34563 5729 34575 5763
rect 34517 5723 34575 5729
rect 36722 5720 36728 5772
rect 36780 5760 36786 5772
rect 39114 5760 39120 5772
rect 36780 5732 38792 5760
rect 39075 5732 39120 5760
rect 36780 5720 36786 5732
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5661 22523 5695
rect 22465 5655 22523 5661
rect 23661 5695 23719 5701
rect 23661 5661 23673 5695
rect 23707 5692 23719 5695
rect 26513 5695 26571 5701
rect 26513 5692 26525 5695
rect 23707 5664 26525 5692
rect 23707 5661 23719 5664
rect 23661 5655 23719 5661
rect 26513 5661 26525 5664
rect 26559 5661 26571 5695
rect 26513 5655 26571 5661
rect 29641 5695 29699 5701
rect 29641 5661 29653 5695
rect 29687 5661 29699 5695
rect 29641 5655 29699 5661
rect 31021 5695 31079 5701
rect 31021 5661 31033 5695
rect 31067 5692 31079 5695
rect 31754 5692 31760 5704
rect 31067 5664 31760 5692
rect 31067 5661 31079 5664
rect 31021 5655 31079 5661
rect 31754 5652 31760 5664
rect 31812 5652 31818 5704
rect 33413 5695 33471 5701
rect 33413 5661 33425 5695
rect 33459 5692 33471 5695
rect 34882 5692 34888 5704
rect 33459 5664 34888 5692
rect 33459 5661 33471 5664
rect 33413 5655 33471 5661
rect 34882 5652 34888 5664
rect 34940 5652 34946 5704
rect 37734 5692 37740 5704
rect 37695 5664 37740 5692
rect 37734 5652 37740 5664
rect 37792 5652 37798 5704
rect 38764 5701 38792 5732
rect 39114 5720 39120 5732
rect 39172 5720 39178 5772
rect 46566 5760 46572 5772
rect 46527 5732 46572 5760
rect 46566 5720 46572 5732
rect 46624 5720 46630 5772
rect 48961 5763 49019 5769
rect 48961 5760 48973 5763
rect 46768 5732 48973 5760
rect 38749 5695 38807 5701
rect 38749 5661 38761 5695
rect 38795 5661 38807 5695
rect 40126 5692 40132 5704
rect 40087 5664 40132 5692
rect 38749 5655 38807 5661
rect 40126 5652 40132 5664
rect 40184 5652 40190 5704
rect 41966 5692 41972 5704
rect 41927 5664 41972 5692
rect 41966 5652 41972 5664
rect 42024 5652 42030 5704
rect 45005 5695 45063 5701
rect 45005 5661 45017 5695
rect 45051 5692 45063 5695
rect 46768 5692 46796 5732
rect 48961 5729 48973 5732
rect 49007 5729 49019 5763
rect 50522 5760 50528 5772
rect 50483 5732 50528 5760
rect 48961 5723 49019 5729
rect 50522 5720 50528 5732
rect 50580 5720 50586 5772
rect 51626 5760 51632 5772
rect 51587 5732 51632 5760
rect 51626 5720 51632 5732
rect 51684 5720 51690 5772
rect 54570 5760 54576 5772
rect 54531 5732 54576 5760
rect 54570 5720 54576 5732
rect 54628 5720 54634 5772
rect 55677 5763 55735 5769
rect 55677 5760 55689 5763
rect 54680 5732 55689 5760
rect 45051 5664 46796 5692
rect 45051 5661 45063 5664
rect 45005 5655 45063 5661
rect 50154 5652 50160 5704
rect 50212 5692 50218 5704
rect 51537 5695 51595 5701
rect 51537 5692 51549 5695
rect 50212 5664 51549 5692
rect 50212 5652 50218 5664
rect 51537 5661 51549 5664
rect 51583 5661 51595 5695
rect 52914 5692 52920 5704
rect 52875 5664 52920 5692
rect 51537 5655 51595 5661
rect 52914 5652 52920 5664
rect 52972 5652 52978 5704
rect 53834 5652 53840 5704
rect 53892 5692 53898 5704
rect 54680 5692 54708 5732
rect 55677 5729 55689 5732
rect 55723 5729 55735 5763
rect 55677 5723 55735 5729
rect 56318 5720 56324 5772
rect 56376 5760 56382 5772
rect 59262 5760 59268 5772
rect 56376 5732 59124 5760
rect 59223 5732 59268 5760
rect 56376 5720 56382 5732
rect 53892 5664 54708 5692
rect 53892 5652 53898 5664
rect 54754 5652 54760 5704
rect 54812 5692 54818 5704
rect 55585 5695 55643 5701
rect 55585 5692 55597 5695
rect 54812 5664 55597 5692
rect 54812 5652 54818 5664
rect 55585 5661 55597 5664
rect 55631 5661 55643 5695
rect 57698 5692 57704 5704
rect 57659 5664 57704 5692
rect 55585 5655 55643 5661
rect 57698 5652 57704 5664
rect 57756 5652 57762 5704
rect 59096 5692 59124 5732
rect 59262 5720 59268 5732
rect 59320 5720 59326 5772
rect 61933 5763 61991 5769
rect 61933 5729 61945 5763
rect 61979 5760 61991 5763
rect 62022 5760 62028 5772
rect 61979 5732 62028 5760
rect 61979 5729 61991 5732
rect 61933 5723 61991 5729
rect 62022 5720 62028 5732
rect 62080 5720 62086 5772
rect 63328 5769 63356 5800
rect 72878 5788 72884 5840
rect 72936 5828 72942 5840
rect 72936 5800 74396 5828
rect 72936 5788 72942 5800
rect 63037 5763 63095 5769
rect 63037 5729 63049 5763
rect 63083 5729 63095 5763
rect 63037 5723 63095 5729
rect 63313 5763 63371 5769
rect 63313 5729 63325 5763
rect 63359 5729 63371 5763
rect 68830 5760 68836 5772
rect 68791 5732 68836 5760
rect 63313 5723 63371 5729
rect 60366 5692 60372 5704
rect 59096 5664 59308 5692
rect 60327 5664 60372 5692
rect 16356 5596 16528 5624
rect 16356 5584 16362 5596
rect 23290 5584 23296 5636
rect 23348 5624 23354 5636
rect 24949 5627 25007 5633
rect 24949 5624 24961 5627
rect 23348 5596 24961 5624
rect 23348 5584 23354 5596
rect 24949 5593 24961 5596
rect 24995 5593 25007 5627
rect 24949 5587 25007 5593
rect 32858 5584 32864 5636
rect 32916 5624 32922 5636
rect 34701 5627 34759 5633
rect 34701 5624 34713 5627
rect 32916 5596 34713 5624
rect 32916 5584 32922 5596
rect 34701 5593 34713 5596
rect 34747 5593 34759 5627
rect 34701 5587 34759 5593
rect 46477 5627 46535 5633
rect 46477 5593 46489 5627
rect 46523 5624 46535 5627
rect 47210 5624 47216 5636
rect 46523 5596 47216 5624
rect 46523 5593 46535 5596
rect 46477 5587 46535 5593
rect 47210 5584 47216 5596
rect 47268 5584 47274 5636
rect 59173 5627 59231 5633
rect 59173 5593 59185 5627
rect 59219 5593 59231 5627
rect 59280 5624 59308 5664
rect 60366 5652 60372 5664
rect 60424 5652 60430 5704
rect 61838 5692 61844 5704
rect 61799 5664 61844 5692
rect 61838 5652 61844 5664
rect 61896 5652 61902 5704
rect 63052 5692 63080 5723
rect 68830 5720 68836 5732
rect 68888 5720 68894 5772
rect 72602 5760 72608 5772
rect 72563 5732 72608 5760
rect 72602 5720 72608 5732
rect 72660 5720 72666 5772
rect 73154 5720 73160 5772
rect 73212 5760 73218 5772
rect 74368 5769 74396 5800
rect 81452 5800 103928 5828
rect 73801 5763 73859 5769
rect 73801 5760 73813 5763
rect 73212 5732 73813 5760
rect 73212 5720 73218 5732
rect 73801 5729 73813 5732
rect 73847 5729 73859 5763
rect 73801 5723 73859 5729
rect 74353 5763 74411 5769
rect 74353 5729 74365 5763
rect 74399 5729 74411 5763
rect 74353 5723 74411 5729
rect 74442 5720 74448 5772
rect 74500 5760 74506 5772
rect 75365 5763 75423 5769
rect 75365 5760 75377 5763
rect 74500 5732 75377 5760
rect 74500 5720 74506 5732
rect 75365 5729 75377 5732
rect 75411 5729 75423 5763
rect 75365 5723 75423 5729
rect 76101 5763 76159 5769
rect 76101 5729 76113 5763
rect 76147 5760 76159 5763
rect 78122 5760 78128 5772
rect 76147 5732 78128 5760
rect 76147 5729 76159 5732
rect 76101 5723 76159 5729
rect 78122 5720 78128 5732
rect 78180 5720 78186 5772
rect 79134 5760 79140 5772
rect 79095 5732 79140 5760
rect 79134 5720 79140 5732
rect 79192 5720 79198 5772
rect 80974 5720 80980 5772
rect 81032 5760 81038 5772
rect 81069 5763 81127 5769
rect 81069 5760 81081 5763
rect 81032 5732 81081 5760
rect 81032 5720 81038 5732
rect 81069 5729 81081 5732
rect 81115 5729 81127 5763
rect 81069 5723 81127 5729
rect 64325 5695 64383 5701
rect 64325 5692 64337 5695
rect 63052 5664 64337 5692
rect 64325 5661 64337 5664
rect 64371 5661 64383 5695
rect 66438 5692 66444 5704
rect 66399 5664 66444 5692
rect 64325 5655 64383 5661
rect 66438 5652 66444 5664
rect 66496 5652 66502 5704
rect 67450 5692 67456 5704
rect 67411 5664 67456 5692
rect 67450 5652 67456 5664
rect 67508 5652 67514 5704
rect 68738 5692 68744 5704
rect 68699 5664 68744 5692
rect 68738 5652 68744 5664
rect 68796 5652 68802 5704
rect 70213 5695 70271 5701
rect 70213 5661 70225 5695
rect 70259 5692 70271 5695
rect 71409 5695 71467 5701
rect 71409 5692 71421 5695
rect 70259 5664 71421 5692
rect 70259 5661 70271 5664
rect 70213 5655 70271 5661
rect 71409 5661 71421 5664
rect 71455 5661 71467 5695
rect 77570 5692 77576 5704
rect 71409 5655 71467 5661
rect 72620 5664 75592 5692
rect 77531 5664 77576 5692
rect 61194 5624 61200 5636
rect 59280 5596 61200 5624
rect 59173 5587 59231 5593
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 10226 5556 10232 5568
rect 2832 5528 10232 5556
rect 2832 5516 2838 5528
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 12710 5516 12716 5568
rect 12768 5556 12774 5568
rect 14550 5556 14556 5568
rect 12768 5528 14556 5556
rect 12768 5516 12774 5528
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 18874 5516 18880 5568
rect 18932 5556 18938 5568
rect 20254 5556 20260 5568
rect 18932 5528 20260 5556
rect 18932 5516 18938 5528
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 22830 5516 22836 5568
rect 22888 5556 22894 5568
rect 25222 5556 25228 5568
rect 22888 5528 25228 5556
rect 22888 5516 22894 5528
rect 25222 5516 25228 5528
rect 25280 5516 25286 5568
rect 43254 5516 43260 5568
rect 43312 5556 43318 5568
rect 45646 5556 45652 5568
rect 43312 5528 45652 5556
rect 43312 5516 43318 5528
rect 45646 5516 45652 5528
rect 45704 5516 45710 5568
rect 59188 5556 59216 5587
rect 61194 5584 61200 5596
rect 61252 5584 61258 5636
rect 72620 5624 72648 5664
rect 61672 5596 72648 5624
rect 72881 5627 72939 5633
rect 61672 5556 61700 5596
rect 72881 5593 72893 5627
rect 72927 5624 72939 5627
rect 73706 5624 73712 5636
rect 72927 5596 73712 5624
rect 72927 5593 72939 5596
rect 72881 5587 72939 5593
rect 73706 5584 73712 5596
rect 73764 5584 73770 5636
rect 73798 5584 73804 5636
rect 73856 5624 73862 5636
rect 74718 5624 74724 5636
rect 73856 5596 74724 5624
rect 73856 5584 73862 5596
rect 74718 5584 74724 5596
rect 74776 5584 74782 5636
rect 59188 5528 61700 5556
rect 62850 5516 62856 5568
rect 62908 5556 62914 5568
rect 62908 5528 62953 5556
rect 62908 5516 62914 5528
rect 73154 5516 73160 5568
rect 73212 5556 73218 5568
rect 73893 5559 73951 5565
rect 73893 5556 73905 5559
rect 73212 5528 73905 5556
rect 73212 5516 73218 5528
rect 73893 5525 73905 5528
rect 73939 5525 73951 5559
rect 75454 5556 75460 5568
rect 75415 5528 75460 5556
rect 73893 5519 73951 5525
rect 75454 5516 75460 5528
rect 75512 5516 75518 5568
rect 75564 5556 75592 5664
rect 77570 5652 77576 5664
rect 77628 5652 77634 5704
rect 77662 5652 77668 5704
rect 77720 5692 77726 5704
rect 81452 5701 81480 5800
rect 103900 5772 103928 5800
rect 104158 5788 104164 5840
rect 104216 5828 104222 5840
rect 109586 5828 109592 5840
rect 104216 5800 109592 5828
rect 104216 5788 104222 5800
rect 109586 5788 109592 5800
rect 109644 5788 109650 5840
rect 109862 5788 109868 5840
rect 109920 5828 109926 5840
rect 114462 5828 114468 5840
rect 109920 5800 114468 5828
rect 109920 5788 109926 5800
rect 114462 5788 114468 5800
rect 114520 5788 114526 5840
rect 119908 5828 119936 5868
rect 120626 5856 120632 5908
rect 120684 5896 120690 5908
rect 126517 5899 126575 5905
rect 126517 5896 126529 5899
rect 120684 5868 126529 5896
rect 120684 5856 120690 5868
rect 126517 5865 126529 5868
rect 126563 5865 126575 5899
rect 126517 5859 126575 5865
rect 126606 5856 126612 5908
rect 126664 5896 126670 5908
rect 127066 5896 127072 5908
rect 126664 5868 127072 5896
rect 126664 5856 126670 5868
rect 127066 5856 127072 5868
rect 127124 5856 127130 5908
rect 128262 5856 128268 5908
rect 128320 5896 128326 5908
rect 133506 5896 133512 5908
rect 128320 5868 133512 5896
rect 128320 5856 128326 5868
rect 133506 5856 133512 5868
rect 133564 5856 133570 5908
rect 133598 5856 133604 5908
rect 133656 5896 133662 5908
rect 133782 5896 133788 5908
rect 133656 5868 133788 5896
rect 133656 5856 133662 5868
rect 133782 5856 133788 5868
rect 133840 5856 133846 5908
rect 134058 5856 134064 5908
rect 134116 5896 134122 5908
rect 141145 5899 141203 5905
rect 141145 5896 141157 5899
rect 134116 5868 141157 5896
rect 134116 5856 134122 5868
rect 141145 5865 141157 5868
rect 141191 5865 141203 5899
rect 142154 5896 142160 5908
rect 142115 5868 142160 5896
rect 141145 5859 141203 5865
rect 142154 5856 142160 5868
rect 142212 5856 142218 5908
rect 143258 5896 143264 5908
rect 143219 5868 143264 5896
rect 143258 5856 143264 5868
rect 143316 5856 143322 5908
rect 143902 5856 143908 5908
rect 143960 5896 143966 5908
rect 145377 5899 145435 5905
rect 145377 5896 145389 5899
rect 143960 5868 145389 5896
rect 143960 5856 143966 5868
rect 145377 5865 145389 5868
rect 145423 5865 145435 5899
rect 145377 5859 145435 5865
rect 121822 5828 121828 5840
rect 114572 5800 119844 5828
rect 119908 5800 121828 5828
rect 82817 5763 82875 5769
rect 82817 5729 82829 5763
rect 82863 5729 82875 5763
rect 83366 5760 83372 5772
rect 83327 5732 83372 5760
rect 82817 5723 82875 5729
rect 79965 5695 80023 5701
rect 79965 5692 79977 5695
rect 77720 5664 79977 5692
rect 77720 5652 77726 5664
rect 79965 5661 79977 5664
rect 80011 5661 80023 5695
rect 79965 5655 80023 5661
rect 81437 5695 81495 5701
rect 81437 5661 81449 5695
rect 81483 5661 81495 5695
rect 82832 5692 82860 5723
rect 83366 5720 83372 5732
rect 83424 5720 83430 5772
rect 89622 5760 89628 5772
rect 89583 5732 89628 5760
rect 89622 5720 89628 5732
rect 89680 5720 89686 5772
rect 91186 5720 91192 5772
rect 91244 5760 91250 5772
rect 91281 5763 91339 5769
rect 91281 5760 91293 5763
rect 91244 5732 91293 5760
rect 91244 5720 91250 5732
rect 91281 5729 91293 5732
rect 91327 5729 91339 5763
rect 91281 5723 91339 5729
rect 92017 5763 92075 5769
rect 92017 5729 92029 5763
rect 92063 5760 92075 5763
rect 94682 5760 94688 5772
rect 92063 5732 94688 5760
rect 92063 5729 92075 5732
rect 92017 5723 92075 5729
rect 94682 5720 94688 5732
rect 94740 5720 94746 5772
rect 95789 5763 95847 5769
rect 95789 5729 95801 5763
rect 95835 5760 95847 5763
rect 96798 5760 96804 5772
rect 95835 5732 96804 5760
rect 95835 5729 95847 5732
rect 95789 5723 95847 5729
rect 96798 5720 96804 5732
rect 96856 5720 96862 5772
rect 96982 5720 96988 5772
rect 97040 5760 97046 5772
rect 97718 5760 97724 5772
rect 97040 5732 97724 5760
rect 97040 5720 97046 5732
rect 97718 5720 97724 5732
rect 97776 5720 97782 5772
rect 98457 5763 98515 5769
rect 98457 5729 98469 5763
rect 98503 5760 98515 5763
rect 99098 5760 99104 5772
rect 98503 5732 99104 5760
rect 98503 5729 98515 5732
rect 98457 5723 98515 5729
rect 99098 5720 99104 5732
rect 99156 5720 99162 5772
rect 103701 5763 103759 5769
rect 103701 5729 103713 5763
rect 103747 5729 103759 5763
rect 103701 5723 103759 5729
rect 84197 5695 84255 5701
rect 84197 5692 84209 5695
rect 82832 5664 84209 5692
rect 81437 5655 81495 5661
rect 84197 5661 84209 5664
rect 84243 5661 84255 5695
rect 84197 5655 84255 5661
rect 86773 5695 86831 5701
rect 86773 5661 86785 5695
rect 86819 5692 86831 5695
rect 88245 5695 88303 5701
rect 88245 5692 88257 5695
rect 86819 5664 88257 5692
rect 86819 5661 86831 5664
rect 86773 5655 86831 5661
rect 88245 5661 88257 5664
rect 88291 5661 88303 5695
rect 94225 5695 94283 5701
rect 88245 5655 88303 5661
rect 88352 5664 93808 5692
rect 79042 5624 79048 5636
rect 79003 5596 79048 5624
rect 79042 5584 79048 5596
rect 79100 5584 79106 5636
rect 80422 5584 80428 5636
rect 80480 5624 80486 5636
rect 82725 5627 82783 5633
rect 82725 5624 82737 5627
rect 80480 5596 82737 5624
rect 80480 5584 80486 5596
rect 82725 5593 82737 5596
rect 82771 5593 82783 5627
rect 88352 5624 88380 5664
rect 82725 5587 82783 5593
rect 82832 5596 88380 5624
rect 82832 5556 82860 5596
rect 89714 5584 89720 5636
rect 89772 5624 89778 5636
rect 89772 5596 89817 5624
rect 89772 5584 89778 5596
rect 91370 5556 91376 5568
rect 75564 5528 82860 5556
rect 91331 5528 91376 5556
rect 91370 5516 91376 5528
rect 91428 5516 91434 5568
rect 93780 5556 93808 5664
rect 94225 5661 94237 5695
rect 94271 5692 94283 5695
rect 94774 5692 94780 5704
rect 94271 5664 94780 5692
rect 94271 5661 94283 5664
rect 94225 5655 94283 5661
rect 94774 5652 94780 5664
rect 94832 5652 94838 5704
rect 95694 5692 95700 5704
rect 95655 5664 95700 5692
rect 95694 5652 95700 5664
rect 95752 5652 95758 5704
rect 96893 5695 96951 5701
rect 96893 5661 96905 5695
rect 96939 5692 96951 5695
rect 98178 5692 98184 5704
rect 96939 5664 98184 5692
rect 96939 5661 96951 5664
rect 96893 5655 96951 5661
rect 98178 5652 98184 5664
rect 98236 5652 98242 5704
rect 98365 5695 98423 5701
rect 98365 5661 98377 5695
rect 98411 5692 98423 5695
rect 99282 5692 99288 5704
rect 98411 5664 99288 5692
rect 98411 5661 98423 5664
rect 98365 5655 98423 5661
rect 99282 5652 99288 5664
rect 99340 5652 99346 5704
rect 99466 5692 99472 5704
rect 99427 5664 99472 5692
rect 99466 5652 99472 5664
rect 99524 5652 99530 5704
rect 103716 5692 103744 5723
rect 103882 5720 103888 5772
rect 103940 5720 103946 5772
rect 104066 5760 104072 5772
rect 104027 5732 104072 5760
rect 104066 5720 104072 5732
rect 104124 5720 104130 5772
rect 104342 5720 104348 5772
rect 104400 5760 104406 5772
rect 107470 5760 107476 5772
rect 104400 5732 107476 5760
rect 104400 5720 104406 5732
rect 107470 5720 107476 5732
rect 107528 5720 107534 5772
rect 107749 5763 107807 5769
rect 107749 5729 107761 5763
rect 107795 5760 107807 5763
rect 107930 5760 107936 5772
rect 107795 5732 107936 5760
rect 107795 5729 107807 5732
rect 107749 5723 107807 5729
rect 107930 5720 107936 5732
rect 107988 5720 107994 5772
rect 108758 5760 108764 5772
rect 108719 5732 108764 5760
rect 108758 5720 108764 5732
rect 108816 5720 108822 5772
rect 109313 5763 109371 5769
rect 109313 5729 109325 5763
rect 109359 5760 109371 5763
rect 111610 5760 111616 5772
rect 109359 5732 111616 5760
rect 109359 5729 109371 5732
rect 109313 5723 109371 5729
rect 111610 5720 111616 5732
rect 111668 5720 111674 5772
rect 112254 5760 112260 5772
rect 112215 5732 112260 5760
rect 112254 5720 112260 5732
rect 112312 5720 112318 5772
rect 106185 5695 106243 5701
rect 103716 5664 105768 5692
rect 94498 5584 94504 5636
rect 94556 5624 94562 5636
rect 94866 5624 94872 5636
rect 94556 5596 94872 5624
rect 94556 5584 94562 5596
rect 94866 5584 94872 5596
rect 94924 5584 94930 5636
rect 95620 5596 104204 5624
rect 95620 5556 95648 5596
rect 93780 5528 95648 5556
rect 98638 5516 98644 5568
rect 98696 5556 98702 5568
rect 103054 5556 103060 5568
rect 98696 5528 103060 5556
rect 98696 5516 98702 5528
rect 103054 5516 103060 5528
rect 103112 5516 103118 5568
rect 103146 5516 103152 5568
rect 103204 5556 103210 5568
rect 103517 5559 103575 5565
rect 103517 5556 103529 5559
rect 103204 5528 103529 5556
rect 103204 5516 103210 5528
rect 103517 5525 103529 5528
rect 103563 5525 103575 5559
rect 104176 5556 104204 5596
rect 104250 5584 104256 5636
rect 104308 5624 104314 5636
rect 105630 5624 105636 5636
rect 104308 5596 105636 5624
rect 104308 5584 104314 5596
rect 105630 5584 105636 5596
rect 105688 5584 105694 5636
rect 105740 5624 105768 5664
rect 106185 5661 106197 5695
rect 106231 5692 106243 5695
rect 106366 5692 106372 5704
rect 106231 5664 106372 5692
rect 106231 5661 106243 5664
rect 106185 5655 106243 5661
rect 106366 5652 106372 5664
rect 106424 5652 106430 5704
rect 107654 5692 107660 5704
rect 107615 5664 107660 5692
rect 107654 5652 107660 5664
rect 107712 5652 107718 5704
rect 108942 5652 108948 5704
rect 109000 5692 109006 5704
rect 109862 5692 109868 5704
rect 109000 5664 109868 5692
rect 109000 5652 109006 5664
rect 109862 5652 109868 5664
rect 109920 5652 109926 5704
rect 110690 5692 110696 5704
rect 110651 5664 110696 5692
rect 110690 5652 110696 5664
rect 110748 5652 110754 5704
rect 113082 5692 113088 5704
rect 110984 5664 112300 5692
rect 113043 5664 113088 5692
rect 106734 5624 106740 5636
rect 105740 5596 106740 5624
rect 106734 5584 106740 5596
rect 106792 5584 106798 5636
rect 107930 5584 107936 5636
rect 107988 5624 107994 5636
rect 107988 5596 108804 5624
rect 107988 5584 107994 5596
rect 108390 5556 108396 5568
rect 104176 5528 108396 5556
rect 103517 5519 103575 5525
rect 108390 5516 108396 5528
rect 108448 5516 108454 5568
rect 108482 5516 108488 5568
rect 108540 5556 108546 5568
rect 108669 5559 108727 5565
rect 108669 5556 108681 5559
rect 108540 5528 108681 5556
rect 108540 5516 108546 5528
rect 108669 5525 108681 5528
rect 108715 5525 108727 5559
rect 108776 5556 108804 5596
rect 110230 5584 110236 5636
rect 110288 5624 110294 5636
rect 110874 5624 110880 5636
rect 110288 5596 110880 5624
rect 110288 5584 110294 5596
rect 110874 5584 110880 5596
rect 110932 5584 110938 5636
rect 110984 5556 111012 5664
rect 111426 5584 111432 5636
rect 111484 5624 111490 5636
rect 111610 5624 111616 5636
rect 111484 5596 111616 5624
rect 111484 5584 111490 5596
rect 111610 5584 111616 5596
rect 111668 5584 111674 5636
rect 112165 5627 112223 5633
rect 112165 5593 112177 5627
rect 112211 5593 112223 5627
rect 112272 5624 112300 5664
rect 113082 5652 113088 5664
rect 113140 5652 113146 5704
rect 114572 5701 114600 5800
rect 114649 5763 114707 5769
rect 114649 5729 114661 5763
rect 114695 5760 114707 5763
rect 117038 5760 117044 5772
rect 114695 5732 117044 5760
rect 114695 5729 114707 5732
rect 114649 5723 114707 5729
rect 117038 5720 117044 5732
rect 117096 5720 117102 5772
rect 114557 5695 114615 5701
rect 114557 5661 114569 5695
rect 114603 5661 114615 5695
rect 114557 5655 114615 5661
rect 114738 5652 114744 5704
rect 114796 5692 114802 5704
rect 116118 5692 116124 5704
rect 114796 5664 116124 5692
rect 114796 5652 114802 5664
rect 116118 5652 116124 5664
rect 116176 5652 116182 5704
rect 116302 5692 116308 5704
rect 116263 5664 116308 5692
rect 116302 5652 116308 5664
rect 116360 5652 116366 5704
rect 117317 5695 117375 5701
rect 117317 5661 117329 5695
rect 117363 5692 117375 5695
rect 118329 5695 118387 5701
rect 118329 5692 118341 5695
rect 117363 5664 118341 5692
rect 117363 5661 117375 5664
rect 117317 5655 117375 5661
rect 118329 5661 118341 5664
rect 118375 5661 118387 5695
rect 119816 5692 119844 5800
rect 121822 5788 121828 5800
rect 121880 5788 121886 5840
rect 127434 5828 127440 5840
rect 124692 5800 127440 5828
rect 119893 5763 119951 5769
rect 119893 5729 119905 5763
rect 119939 5760 119951 5763
rect 121362 5760 121368 5772
rect 119939 5732 121368 5760
rect 119939 5729 119951 5732
rect 119893 5723 119951 5729
rect 121362 5720 121368 5732
rect 121420 5720 121426 5772
rect 122650 5720 122656 5772
rect 122708 5760 122714 5772
rect 124692 5769 124720 5800
rect 127434 5788 127440 5800
rect 127492 5788 127498 5840
rect 127526 5788 127532 5840
rect 127584 5828 127590 5840
rect 154390 5828 154396 5840
rect 127584 5800 154396 5828
rect 127584 5788 127590 5800
rect 154390 5788 154396 5800
rect 154448 5788 154454 5840
rect 123113 5763 123171 5769
rect 123113 5760 123125 5763
rect 122708 5732 123125 5760
rect 122708 5720 122714 5732
rect 123113 5729 123125 5732
rect 123159 5729 123171 5763
rect 123113 5723 123171 5729
rect 124677 5763 124735 5769
rect 124677 5729 124689 5763
rect 124723 5729 124735 5763
rect 124677 5723 124735 5729
rect 124766 5720 124772 5772
rect 124824 5760 124830 5772
rect 126330 5760 126336 5772
rect 124824 5732 126336 5760
rect 124824 5720 124830 5732
rect 126330 5720 126336 5732
rect 126388 5720 126394 5772
rect 126425 5763 126483 5769
rect 126425 5729 126437 5763
rect 126471 5760 126483 5763
rect 128170 5760 128176 5772
rect 126471 5732 128176 5760
rect 126471 5729 126483 5732
rect 126425 5723 126483 5729
rect 128170 5720 128176 5732
rect 128228 5720 128234 5772
rect 128814 5760 128820 5772
rect 128775 5732 128820 5760
rect 128814 5720 128820 5732
rect 128872 5720 128878 5772
rect 129274 5720 129280 5772
rect 129332 5760 129338 5772
rect 131758 5760 131764 5772
rect 129332 5732 130792 5760
rect 131719 5732 131764 5760
rect 129332 5720 129338 5732
rect 120813 5695 120871 5701
rect 119816 5664 119936 5692
rect 118329 5655 118387 5661
rect 117682 5624 117688 5636
rect 112272 5596 117688 5624
rect 112165 5587 112223 5593
rect 108776 5528 111012 5556
rect 112180 5556 112208 5587
rect 117682 5584 117688 5596
rect 117740 5584 117746 5636
rect 119801 5627 119859 5633
rect 119801 5593 119813 5627
rect 119847 5593 119859 5627
rect 119908 5624 119936 5664
rect 120813 5661 120825 5695
rect 120859 5692 120871 5695
rect 122006 5692 122012 5704
rect 120859 5664 122012 5692
rect 120859 5661 120871 5664
rect 120813 5655 120871 5661
rect 122006 5652 122012 5664
rect 122064 5652 122070 5704
rect 122101 5695 122159 5701
rect 122101 5661 122113 5695
rect 122147 5692 122159 5695
rect 123018 5692 123024 5704
rect 122147 5664 123024 5692
rect 122147 5661 122159 5664
rect 122101 5655 122159 5661
rect 123018 5652 123024 5664
rect 123076 5652 123082 5704
rect 123478 5652 123484 5704
rect 123536 5692 123542 5704
rect 127526 5692 127532 5704
rect 123536 5664 127532 5692
rect 123536 5652 123542 5664
rect 127526 5652 127532 5664
rect 127584 5652 127590 5704
rect 127618 5652 127624 5704
rect 127676 5692 127682 5704
rect 130654 5692 130660 5704
rect 127676 5664 127721 5692
rect 130615 5664 130660 5692
rect 127676 5652 127682 5664
rect 130654 5652 130660 5664
rect 130712 5652 130718 5704
rect 130764 5692 130792 5732
rect 131758 5720 131764 5732
rect 131816 5720 131822 5772
rect 133138 5760 133144 5772
rect 133099 5732 133144 5760
rect 133138 5720 133144 5732
rect 133196 5720 133202 5772
rect 133598 5720 133604 5772
rect 133656 5760 133662 5772
rect 134610 5760 134616 5772
rect 133656 5732 134616 5760
rect 133656 5720 133662 5732
rect 134610 5720 134616 5732
rect 134668 5720 134674 5772
rect 134705 5763 134763 5769
rect 134705 5729 134717 5763
rect 134751 5760 134763 5763
rect 134886 5760 134892 5772
rect 134751 5732 134892 5760
rect 134751 5729 134763 5732
rect 134705 5723 134763 5729
rect 134886 5720 134892 5732
rect 134944 5720 134950 5772
rect 135533 5763 135591 5769
rect 135533 5729 135545 5763
rect 135579 5760 135591 5763
rect 136634 5760 136640 5772
rect 135579 5732 136640 5760
rect 135579 5729 135591 5732
rect 135533 5723 135591 5729
rect 136634 5720 136640 5732
rect 136692 5720 136698 5772
rect 137097 5763 137155 5769
rect 137097 5729 137109 5763
rect 137143 5760 137155 5763
rect 139854 5760 139860 5772
rect 137143 5732 139860 5760
rect 137143 5729 137155 5732
rect 137097 5723 137155 5729
rect 139854 5720 139860 5732
rect 139912 5720 139918 5772
rect 140317 5763 140375 5769
rect 140317 5729 140329 5763
rect 140363 5760 140375 5763
rect 140363 5732 141096 5760
rect 140363 5729 140375 5732
rect 140317 5723 140375 5729
rect 130764 5664 132080 5692
rect 123938 5624 123944 5636
rect 119908 5596 123944 5624
rect 119801 5587 119859 5593
rect 119614 5556 119620 5568
rect 112180 5528 119620 5556
rect 108669 5519 108727 5525
rect 119614 5516 119620 5528
rect 119672 5516 119678 5568
rect 119816 5556 119844 5587
rect 123938 5584 123944 5596
rect 123996 5584 124002 5636
rect 124585 5627 124643 5633
rect 124585 5593 124597 5627
rect 124631 5624 124643 5627
rect 128906 5624 128912 5636
rect 124631 5596 128676 5624
rect 128867 5596 128912 5624
rect 124631 5593 124643 5596
rect 124585 5587 124643 5593
rect 128538 5556 128544 5568
rect 119816 5528 128544 5556
rect 128538 5516 128544 5528
rect 128596 5516 128602 5568
rect 128648 5556 128676 5596
rect 128906 5584 128912 5596
rect 128964 5584 128970 5636
rect 129366 5584 129372 5636
rect 129424 5624 129430 5636
rect 131574 5624 131580 5636
rect 129424 5596 131580 5624
rect 129424 5584 129430 5596
rect 131574 5584 131580 5596
rect 131632 5584 131638 5636
rect 131942 5624 131948 5636
rect 131903 5596 131948 5624
rect 131942 5584 131948 5596
rect 132000 5584 132006 5636
rect 132052 5624 132080 5664
rect 132218 5652 132224 5704
rect 132276 5692 132282 5704
rect 132276 5664 134748 5692
rect 132276 5652 132282 5664
rect 134150 5624 134156 5636
rect 132052 5596 134156 5624
rect 134150 5584 134156 5596
rect 134208 5584 134214 5636
rect 134610 5624 134616 5636
rect 134571 5596 134616 5624
rect 134610 5584 134616 5596
rect 134668 5584 134674 5636
rect 134720 5624 134748 5664
rect 134794 5652 134800 5704
rect 134852 5692 134858 5704
rect 138750 5692 138756 5704
rect 134852 5664 137784 5692
rect 138711 5664 138756 5692
rect 134852 5652 134858 5664
rect 135530 5624 135536 5636
rect 134720 5596 135536 5624
rect 135530 5584 135536 5596
rect 135588 5584 135594 5636
rect 135898 5584 135904 5636
rect 135956 5624 135962 5636
rect 137005 5627 137063 5633
rect 135956 5596 136312 5624
rect 135956 5584 135962 5596
rect 136174 5556 136180 5568
rect 128648 5528 136180 5556
rect 136174 5516 136180 5528
rect 136232 5516 136238 5568
rect 136284 5556 136312 5596
rect 137005 5593 137017 5627
rect 137051 5624 137063 5627
rect 137646 5624 137652 5636
rect 137051 5596 137652 5624
rect 137051 5593 137063 5596
rect 137005 5587 137063 5593
rect 137646 5584 137652 5596
rect 137704 5584 137710 5636
rect 137554 5556 137560 5568
rect 136284 5528 137560 5556
rect 137554 5516 137560 5528
rect 137612 5516 137618 5568
rect 137756 5556 137784 5664
rect 138750 5652 138756 5664
rect 138808 5652 138814 5704
rect 141068 5692 141096 5732
rect 141142 5720 141148 5772
rect 141200 5760 141206 5772
rect 144365 5763 144423 5769
rect 144365 5760 144377 5763
rect 141200 5732 144377 5760
rect 141200 5720 141206 5732
rect 144365 5729 144377 5732
rect 144411 5729 144423 5763
rect 144365 5723 144423 5729
rect 153473 5763 153531 5769
rect 153473 5729 153485 5763
rect 153519 5760 153531 5763
rect 153654 5760 153660 5772
rect 153519 5732 153660 5760
rect 153519 5729 153531 5732
rect 153473 5723 153531 5729
rect 153654 5720 153660 5732
rect 153712 5720 153718 5772
rect 146110 5692 146116 5704
rect 141068 5664 146116 5692
rect 146110 5652 146116 5664
rect 146168 5652 146174 5704
rect 146386 5652 146392 5704
rect 146444 5692 146450 5704
rect 148778 5692 148784 5704
rect 146444 5664 148784 5692
rect 146444 5652 146450 5664
rect 148778 5652 148784 5664
rect 148836 5652 148842 5704
rect 151909 5695 151967 5701
rect 151909 5661 151921 5695
rect 151955 5692 151967 5695
rect 153286 5692 153292 5704
rect 151955 5664 153292 5692
rect 151955 5661 151967 5664
rect 151909 5655 151967 5661
rect 153286 5652 153292 5664
rect 153344 5652 153350 5704
rect 140225 5627 140283 5633
rect 140225 5593 140237 5627
rect 140271 5624 140283 5627
rect 151354 5624 151360 5636
rect 140271 5596 151360 5624
rect 140271 5593 140283 5596
rect 140225 5587 140283 5593
rect 151354 5584 151360 5596
rect 151412 5584 151418 5636
rect 152918 5584 152924 5636
rect 152976 5624 152982 5636
rect 153197 5627 153255 5633
rect 153197 5624 153209 5627
rect 152976 5596 153209 5624
rect 152976 5584 152982 5596
rect 153197 5593 153209 5596
rect 153243 5593 153255 5627
rect 153197 5587 153255 5593
rect 156506 5556 156512 5568
rect 137756 5528 156512 5556
rect 156506 5516 156512 5528
rect 156564 5516 156570 5568
rect 1104 5466 154560 5488
rect 1104 5414 4078 5466
rect 4130 5414 44078 5466
rect 44130 5414 84078 5466
rect 84130 5414 124078 5466
rect 124130 5414 154560 5466
rect 1104 5392 154560 5414
rect 70486 5312 70492 5364
rect 70544 5352 70550 5364
rect 94498 5352 94504 5364
rect 70544 5324 94504 5352
rect 70544 5312 70550 5324
rect 94498 5312 94504 5324
rect 94556 5312 94562 5364
rect 94682 5312 94688 5364
rect 94740 5352 94746 5364
rect 96062 5352 96068 5364
rect 94740 5324 96068 5352
rect 94740 5312 94746 5324
rect 96062 5312 96068 5324
rect 96120 5312 96126 5364
rect 96433 5355 96491 5361
rect 96433 5321 96445 5355
rect 96479 5352 96491 5355
rect 101214 5352 101220 5364
rect 96479 5324 101220 5352
rect 96479 5321 96491 5324
rect 96433 5315 96491 5321
rect 101214 5312 101220 5324
rect 101272 5312 101278 5364
rect 118510 5352 118516 5364
rect 101324 5324 118516 5352
rect 5813 5287 5871 5293
rect 5813 5253 5825 5287
rect 5859 5284 5871 5287
rect 8018 5284 8024 5296
rect 5859 5256 8024 5284
rect 5859 5253 5871 5256
rect 5813 5247 5871 5253
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 8113 5287 8171 5293
rect 8113 5253 8125 5287
rect 8159 5284 8171 5287
rect 9306 5284 9312 5296
rect 8159 5256 9312 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 37645 5287 37703 5293
rect 37645 5253 37657 5287
rect 37691 5284 37703 5287
rect 38470 5284 38476 5296
rect 37691 5256 38476 5284
rect 37691 5253 37703 5256
rect 37645 5247 37703 5253
rect 38470 5244 38476 5256
rect 38528 5244 38534 5296
rect 41969 5287 42027 5293
rect 41969 5253 41981 5287
rect 42015 5284 42027 5287
rect 43714 5284 43720 5296
rect 42015 5256 43720 5284
rect 42015 5253 42027 5256
rect 41969 5247 42027 5253
rect 43714 5244 43720 5256
rect 43772 5244 43778 5296
rect 45097 5287 45155 5293
rect 45097 5253 45109 5287
rect 45143 5284 45155 5287
rect 49602 5284 49608 5296
rect 45143 5256 49608 5284
rect 45143 5253 45155 5256
rect 45097 5247 45155 5253
rect 49602 5244 49608 5256
rect 49660 5244 49666 5296
rect 55950 5244 55956 5296
rect 56008 5284 56014 5296
rect 56137 5287 56195 5293
rect 56137 5284 56149 5287
rect 56008 5256 56149 5284
rect 56008 5244 56014 5256
rect 56137 5253 56149 5256
rect 56183 5253 56195 5287
rect 57974 5284 57980 5296
rect 57935 5256 57980 5284
rect 56137 5247 56195 5253
rect 57974 5244 57980 5256
rect 58032 5244 58038 5296
rect 59170 5244 59176 5296
rect 59228 5284 59234 5296
rect 59228 5256 60504 5284
rect 59228 5244 59234 5256
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 6914 5216 6920 5228
rect 6871 5188 6920 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 8536 5188 9229 5216
rect 8536 5176 8542 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 13630 5216 13636 5228
rect 13591 5188 13636 5216
rect 9217 5179 9275 5185
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15436 5188 15853 5216
rect 15436 5176 15442 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 20254 5216 20260 5228
rect 20215 5188 20260 5216
rect 15841 5179 15899 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20806 5176 20812 5228
rect 20864 5216 20870 5228
rect 21637 5219 21695 5225
rect 21637 5216 21649 5219
rect 20864 5188 21649 5216
rect 20864 5176 20870 5188
rect 21637 5185 21649 5188
rect 21683 5185 21695 5219
rect 21637 5179 21695 5185
rect 22462 5176 22468 5228
rect 22520 5216 22526 5228
rect 24673 5219 24731 5225
rect 24673 5216 24685 5219
rect 22520 5188 24685 5216
rect 22520 5176 22526 5188
rect 24673 5185 24685 5188
rect 24719 5185 24731 5219
rect 30374 5216 30380 5228
rect 30335 5188 30380 5216
rect 24673 5179 24731 5185
rect 30374 5176 30380 5188
rect 30432 5176 30438 5228
rect 31754 5216 31760 5228
rect 31715 5188 31760 5216
rect 31754 5176 31760 5188
rect 31812 5176 31818 5228
rect 32306 5176 32312 5228
rect 32364 5216 32370 5228
rect 32769 5219 32827 5225
rect 32769 5216 32781 5219
rect 32364 5188 32781 5216
rect 32364 5176 32370 5188
rect 32769 5185 32781 5188
rect 32815 5185 32827 5219
rect 34882 5216 34888 5228
rect 34843 5188 34888 5216
rect 32769 5179 32827 5185
rect 34882 5176 34888 5188
rect 34940 5176 34946 5228
rect 40126 5176 40132 5228
rect 40184 5216 40190 5228
rect 40497 5219 40555 5225
rect 40497 5216 40509 5219
rect 40184 5188 40509 5216
rect 40184 5176 40190 5188
rect 40497 5185 40509 5188
rect 40543 5185 40555 5219
rect 47118 5216 47124 5228
rect 47079 5188 47124 5216
rect 40497 5179 40555 5185
rect 47118 5176 47124 5188
rect 47176 5176 47182 5228
rect 48498 5176 48504 5228
rect 48556 5216 48562 5228
rect 49237 5219 49295 5225
rect 49237 5216 49249 5219
rect 48556 5188 49249 5216
rect 48556 5176 48562 5188
rect 49237 5185 49249 5188
rect 49283 5185 49295 5219
rect 49237 5179 49295 5185
rect 52273 5219 52331 5225
rect 52273 5185 52285 5219
rect 52319 5216 52331 5219
rect 52914 5216 52920 5228
rect 52319 5188 52920 5216
rect 52319 5185 52331 5188
rect 52273 5179 52331 5185
rect 52914 5176 52920 5188
rect 52972 5176 52978 5228
rect 53282 5216 53288 5228
rect 53243 5188 53288 5216
rect 53282 5176 53288 5188
rect 53340 5176 53346 5228
rect 59078 5176 59084 5228
rect 59136 5216 59142 5228
rect 60476 5225 60504 5256
rect 62206 5244 62212 5296
rect 62264 5284 62270 5296
rect 63037 5287 63095 5293
rect 63037 5284 63049 5287
rect 62264 5256 63049 5284
rect 62264 5244 62270 5256
rect 63037 5253 63049 5256
rect 63083 5253 63095 5287
rect 63037 5247 63095 5253
rect 66530 5244 66536 5296
rect 66588 5284 66594 5296
rect 66993 5287 67051 5293
rect 66993 5284 67005 5287
rect 66588 5256 67005 5284
rect 66588 5244 66594 5256
rect 66993 5253 67005 5256
rect 67039 5253 67051 5287
rect 66993 5247 67051 5253
rect 72234 5244 72240 5296
rect 72292 5284 72298 5296
rect 72292 5256 78260 5284
rect 72292 5244 72298 5256
rect 60461 5219 60519 5225
rect 59136 5188 59584 5216
rect 59136 5176 59142 5188
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5148 3387 5151
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 3375 5120 4353 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5148 5963 5151
rect 7466 5148 7472 5160
rect 5951 5120 7472 5148
rect 5951 5117 5963 5120
rect 5905 5111 5963 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 7926 5148 7932 5160
rect 7887 5120 7932 5148
rect 7926 5108 7932 5120
rect 7984 5108 7990 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 13354 5148 13360 5160
rect 12483 5120 13360 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 13814 5148 13820 5160
rect 13775 5120 13820 5148
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 15286 5148 15292 5160
rect 14875 5120 15292 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 15930 5148 15936 5160
rect 15891 5120 15936 5148
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 19245 5151 19303 5157
rect 19245 5117 19257 5151
rect 19291 5148 19303 5151
rect 20438 5148 20444 5160
rect 19291 5120 20444 5148
rect 19291 5117 19303 5120
rect 19245 5111 19303 5117
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 20714 5148 20720 5160
rect 20675 5120 20720 5148
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 23474 5108 23480 5160
rect 23532 5148 23538 5160
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 23532 5120 23673 5148
rect 23532 5108 23538 5120
rect 23661 5117 23673 5120
rect 23707 5117 23719 5151
rect 23661 5111 23719 5117
rect 23750 5108 23756 5160
rect 23808 5148 23814 5160
rect 24765 5151 24823 5157
rect 24765 5148 24777 5151
rect 23808 5120 24777 5148
rect 23808 5108 23814 5120
rect 24765 5117 24777 5120
rect 24811 5117 24823 5151
rect 29362 5148 29368 5160
rect 29323 5120 29368 5148
rect 24765 5111 24823 5117
rect 29362 5108 29368 5120
rect 29420 5108 29426 5160
rect 30466 5148 30472 5160
rect 30427 5120 30472 5148
rect 30466 5108 30472 5120
rect 30524 5108 30530 5160
rect 32950 5148 32956 5160
rect 32911 5120 32956 5148
rect 32950 5108 32956 5120
rect 33008 5108 33014 5160
rect 36078 5108 36084 5160
rect 36136 5148 36142 5160
rect 36173 5151 36231 5157
rect 36173 5148 36185 5151
rect 36136 5120 36185 5148
rect 36136 5108 36142 5120
rect 36173 5117 36185 5120
rect 36219 5117 36231 5151
rect 36173 5111 36231 5117
rect 37737 5151 37795 5157
rect 37737 5117 37749 5151
rect 37783 5148 37795 5151
rect 41138 5148 41144 5160
rect 37783 5120 41144 5148
rect 37783 5117 37795 5120
rect 37737 5111 37795 5117
rect 41138 5108 41144 5120
rect 41196 5108 41202 5160
rect 42061 5151 42119 5157
rect 42061 5117 42073 5151
rect 42107 5148 42119 5151
rect 42334 5148 42340 5160
rect 42107 5120 42340 5148
rect 42107 5117 42119 5120
rect 42061 5111 42119 5117
rect 42334 5108 42340 5120
rect 42392 5108 42398 5160
rect 43625 5151 43683 5157
rect 43625 5117 43637 5151
rect 43671 5148 43683 5151
rect 44542 5148 44548 5160
rect 43671 5120 44548 5148
rect 43671 5117 43683 5120
rect 43625 5111 43683 5117
rect 44542 5108 44548 5120
rect 44600 5108 44606 5160
rect 45189 5151 45247 5157
rect 45189 5117 45201 5151
rect 45235 5117 45247 5151
rect 46106 5148 46112 5160
rect 46067 5120 46112 5148
rect 45189 5111 45247 5117
rect 45204 5080 45232 5111
rect 46106 5108 46112 5120
rect 46164 5108 46170 5160
rect 47210 5148 47216 5160
rect 47171 5120 47216 5148
rect 47210 5108 47216 5120
rect 47268 5108 47274 5160
rect 53558 5148 53564 5160
rect 53519 5120 53564 5148
rect 53558 5108 53564 5120
rect 53616 5108 53622 5160
rect 54846 5148 54852 5160
rect 54807 5120 54852 5148
rect 54846 5108 54852 5120
rect 54904 5108 54910 5160
rect 55950 5148 55956 5160
rect 55911 5120 55956 5148
rect 55950 5108 55956 5120
rect 56008 5108 56014 5160
rect 57977 5151 58035 5157
rect 57977 5117 57989 5151
rect 58023 5117 58035 5151
rect 57977 5111 58035 5117
rect 47762 5080 47768 5092
rect 45204 5052 47768 5080
rect 47762 5040 47768 5052
rect 47820 5040 47826 5092
rect 57992 5080 58020 5111
rect 58066 5108 58072 5160
rect 58124 5148 58130 5160
rect 58437 5151 58495 5157
rect 58437 5148 58449 5151
rect 58124 5120 58449 5148
rect 58124 5108 58130 5120
rect 58437 5117 58449 5120
rect 58483 5117 58495 5151
rect 58437 5111 58495 5117
rect 59449 5151 59507 5157
rect 59449 5117 59461 5151
rect 59495 5117 59507 5151
rect 59556 5148 59584 5188
rect 60461 5185 60473 5219
rect 60507 5185 60519 5219
rect 60461 5179 60519 5185
rect 61930 5176 61936 5228
rect 61988 5216 61994 5228
rect 61988 5188 63540 5216
rect 61988 5176 61994 5188
rect 60645 5151 60703 5157
rect 60645 5148 60657 5151
rect 59556 5120 60657 5148
rect 59449 5111 59507 5117
rect 60645 5117 60657 5120
rect 60691 5117 60703 5151
rect 63218 5148 63224 5160
rect 63179 5120 63224 5148
rect 60645 5111 60703 5117
rect 59354 5080 59360 5092
rect 57992 5052 59360 5080
rect 59354 5040 59360 5052
rect 59412 5040 59418 5092
rect 59464 5080 59492 5111
rect 63218 5108 63224 5120
rect 63276 5108 63282 5160
rect 63512 5157 63540 5188
rect 63862 5176 63868 5228
rect 63920 5216 63926 5228
rect 64509 5219 64567 5225
rect 64509 5216 64521 5219
rect 63920 5188 64521 5216
rect 63920 5176 63926 5188
rect 64509 5185 64521 5188
rect 64555 5185 64567 5219
rect 64509 5179 64567 5185
rect 69293 5219 69351 5225
rect 69293 5185 69305 5219
rect 69339 5216 69351 5219
rect 70578 5216 70584 5228
rect 69339 5188 70584 5216
rect 69339 5185 69351 5188
rect 69293 5179 69351 5185
rect 70578 5176 70584 5188
rect 70636 5176 70642 5228
rect 70762 5176 70768 5228
rect 70820 5216 70826 5228
rect 76101 5219 76159 5225
rect 70820 5188 71084 5216
rect 70820 5176 70826 5188
rect 63497 5151 63555 5157
rect 63497 5117 63509 5151
rect 63543 5117 63555 5151
rect 63497 5111 63555 5117
rect 66438 5108 66444 5160
rect 66496 5148 66502 5160
rect 66901 5151 66959 5157
rect 66901 5148 66913 5151
rect 66496 5120 66913 5148
rect 66496 5108 66502 5120
rect 66901 5117 66913 5120
rect 66947 5117 66959 5151
rect 66901 5111 66959 5117
rect 67545 5151 67603 5157
rect 67545 5117 67557 5151
rect 67591 5148 67603 5151
rect 67726 5148 67732 5160
rect 67591 5120 67732 5148
rect 67591 5117 67603 5120
rect 67545 5111 67603 5117
rect 67726 5108 67732 5120
rect 67784 5108 67790 5160
rect 69014 5148 69020 5160
rect 68975 5120 69020 5148
rect 69014 5108 69020 5120
rect 69072 5108 69078 5160
rect 69661 5151 69719 5157
rect 69661 5117 69673 5151
rect 69707 5117 69719 5151
rect 69661 5111 69719 5117
rect 61841 5083 61899 5089
rect 61841 5080 61853 5083
rect 59464 5052 61853 5080
rect 61841 5049 61853 5052
rect 61887 5049 61899 5083
rect 69676 5080 69704 5111
rect 69934 5108 69940 5160
rect 69992 5148 69998 5160
rect 70489 5151 70547 5157
rect 70489 5148 70501 5151
rect 69992 5120 70501 5148
rect 69992 5108 69998 5120
rect 70489 5117 70501 5120
rect 70535 5117 70547 5151
rect 70854 5148 70860 5160
rect 70815 5120 70860 5148
rect 70489 5111 70547 5117
rect 70854 5108 70860 5120
rect 70912 5108 70918 5160
rect 71056 5157 71084 5188
rect 76101 5185 76113 5219
rect 76147 5216 76159 5219
rect 77570 5216 77576 5228
rect 76147 5188 77576 5216
rect 76147 5185 76159 5188
rect 76101 5179 76159 5185
rect 77570 5176 77576 5188
rect 77628 5176 77634 5228
rect 71041 5151 71099 5157
rect 71041 5117 71053 5151
rect 71087 5117 71099 5151
rect 71041 5111 71099 5117
rect 72053 5151 72111 5157
rect 72053 5117 72065 5151
rect 72099 5117 72111 5151
rect 72418 5148 72424 5160
rect 72379 5120 72424 5148
rect 72053 5111 72111 5117
rect 71222 5080 71228 5092
rect 69676 5052 71228 5080
rect 61841 5043 61899 5049
rect 71222 5040 71228 5052
rect 71280 5040 71286 5092
rect 2317 5015 2375 5021
rect 2317 4981 2329 5015
rect 2363 5012 2375 5015
rect 7006 5012 7012 5024
rect 2363 4984 7012 5012
rect 2363 4981 2375 4984
rect 2317 4975 2375 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 10873 5015 10931 5021
rect 10873 4981 10885 5015
rect 10919 5012 10931 5015
rect 10962 5012 10968 5024
rect 10919 4984 10968 5012
rect 10919 4981 10931 4984
rect 10873 4975 10931 4981
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 50617 5015 50675 5021
rect 50617 4981 50629 5015
rect 50663 5012 50675 5015
rect 51718 5012 51724 5024
rect 50663 4984 51724 5012
rect 50663 4981 50675 4984
rect 50617 4975 50675 4981
rect 51718 4972 51724 4984
rect 51776 4972 51782 5024
rect 65889 5015 65947 5021
rect 65889 4981 65901 5015
rect 65935 5012 65947 5015
rect 67542 5012 67548 5024
rect 65935 4984 67548 5012
rect 65935 4981 65947 4984
rect 65889 4975 65947 4981
rect 67542 4972 67548 4984
rect 67600 4972 67606 5024
rect 67726 4972 67732 5024
rect 67784 5012 67790 5024
rect 72068 5012 72096 5111
rect 72418 5108 72424 5120
rect 72476 5108 72482 5160
rect 72510 5108 72516 5160
rect 72568 5148 72574 5160
rect 72605 5151 72663 5157
rect 72605 5148 72617 5151
rect 72568 5120 72617 5148
rect 72568 5108 72574 5120
rect 72605 5117 72617 5120
rect 72651 5117 72663 5151
rect 74166 5148 74172 5160
rect 74127 5120 74172 5148
rect 72605 5111 72663 5117
rect 74166 5108 74172 5120
rect 74224 5108 74230 5160
rect 74534 5148 74540 5160
rect 74495 5120 74540 5148
rect 74534 5108 74540 5120
rect 74592 5108 74598 5160
rect 74718 5148 74724 5160
rect 74679 5120 74724 5148
rect 74718 5108 74724 5120
rect 74776 5108 74782 5160
rect 77113 5151 77171 5157
rect 77113 5117 77125 5151
rect 77159 5148 77171 5151
rect 77662 5148 77668 5160
rect 77159 5120 77668 5148
rect 77159 5117 77171 5120
rect 77113 5111 77171 5117
rect 77662 5108 77668 5120
rect 77720 5108 77726 5160
rect 78232 5157 78260 5256
rect 78766 5244 78772 5296
rect 78824 5284 78830 5296
rect 81437 5287 81495 5293
rect 81437 5284 81449 5287
rect 78824 5256 81449 5284
rect 78824 5244 78830 5256
rect 81437 5253 81449 5256
rect 81483 5253 81495 5287
rect 81437 5247 81495 5253
rect 81618 5244 81624 5296
rect 81676 5244 81682 5296
rect 89990 5284 89996 5296
rect 89951 5256 89996 5284
rect 89990 5244 89996 5256
rect 90048 5244 90054 5296
rect 99561 5287 99619 5293
rect 99561 5284 99573 5287
rect 94516 5256 99573 5284
rect 81636 5216 81664 5244
rect 80532 5188 81664 5216
rect 86865 5219 86923 5225
rect 78217 5151 78275 5157
rect 78217 5117 78229 5151
rect 78263 5117 78275 5151
rect 79778 5148 79784 5160
rect 79739 5120 79784 5148
rect 78217 5111 78275 5117
rect 79778 5108 79784 5120
rect 79836 5108 79842 5160
rect 80146 5148 80152 5160
rect 80107 5120 80152 5148
rect 80146 5108 80152 5120
rect 80204 5108 80210 5160
rect 80532 5157 80560 5188
rect 86865 5185 86877 5219
rect 86911 5216 86923 5219
rect 94516 5216 94544 5256
rect 99561 5253 99573 5256
rect 99607 5253 99619 5287
rect 99561 5247 99619 5253
rect 101125 5287 101183 5293
rect 101125 5253 101137 5287
rect 101171 5284 101183 5287
rect 101324 5284 101352 5324
rect 118510 5312 118516 5324
rect 118568 5312 118574 5364
rect 118602 5312 118608 5364
rect 118660 5352 118666 5364
rect 119522 5352 119528 5364
rect 118660 5324 119528 5352
rect 118660 5312 118666 5324
rect 119522 5312 119528 5324
rect 119580 5312 119586 5364
rect 123478 5352 123484 5364
rect 121840 5324 123484 5352
rect 117409 5287 117467 5293
rect 101171 5256 101352 5284
rect 103992 5256 116440 5284
rect 101171 5253 101183 5256
rect 101125 5247 101183 5253
rect 86911 5188 94544 5216
rect 94777 5219 94835 5225
rect 86911 5185 86923 5188
rect 86865 5179 86923 5185
rect 94777 5185 94789 5219
rect 94823 5216 94835 5219
rect 94823 5188 99420 5216
rect 94823 5185 94835 5188
rect 94777 5179 94835 5185
rect 80517 5151 80575 5157
rect 80517 5117 80529 5151
rect 80563 5117 80575 5151
rect 81618 5148 81624 5160
rect 81579 5120 81624 5148
rect 80517 5111 80575 5117
rect 81618 5108 81624 5120
rect 81676 5108 81682 5160
rect 82078 5148 82084 5160
rect 82039 5120 82084 5148
rect 82078 5108 82084 5120
rect 82136 5108 82142 5160
rect 84289 5151 84347 5157
rect 84289 5117 84301 5151
rect 84335 5148 84347 5151
rect 85393 5151 85451 5157
rect 85393 5148 85405 5151
rect 84335 5120 85405 5148
rect 84335 5117 84347 5120
rect 84289 5111 84347 5117
rect 85393 5117 85405 5120
rect 85439 5117 85451 5151
rect 86770 5148 86776 5160
rect 86731 5120 86776 5148
rect 85393 5111 85451 5117
rect 86770 5108 86776 5120
rect 86828 5108 86834 5160
rect 88518 5148 88524 5160
rect 88479 5120 88524 5148
rect 88518 5108 88524 5120
rect 88576 5108 88582 5160
rect 90085 5151 90143 5157
rect 90085 5117 90097 5151
rect 90131 5148 90143 5151
rect 90266 5148 90272 5160
rect 90131 5120 90272 5148
rect 90131 5117 90143 5120
rect 90085 5111 90143 5117
rect 90266 5108 90272 5120
rect 90324 5108 90330 5160
rect 91646 5148 91652 5160
rect 91607 5120 91652 5148
rect 91646 5108 91652 5120
rect 91704 5108 91710 5160
rect 91741 5151 91799 5157
rect 91741 5117 91753 5151
rect 91787 5148 91799 5151
rect 92750 5148 92756 5160
rect 91787 5120 92756 5148
rect 91787 5117 91799 5120
rect 91741 5111 91799 5117
rect 92750 5108 92756 5120
rect 92808 5108 92814 5160
rect 93305 5151 93363 5157
rect 93305 5117 93317 5151
rect 93351 5148 93363 5151
rect 93854 5148 93860 5160
rect 93351 5120 93860 5148
rect 93351 5117 93363 5120
rect 93305 5111 93363 5117
rect 93854 5108 93860 5120
rect 93912 5108 93918 5160
rect 94869 5151 94927 5157
rect 94869 5117 94881 5151
rect 94915 5148 94927 5151
rect 96433 5151 96491 5157
rect 96433 5148 96445 5151
rect 94915 5120 96445 5148
rect 94915 5117 94927 5120
rect 94869 5111 94927 5117
rect 96433 5117 96445 5120
rect 96479 5117 96491 5151
rect 96433 5111 96491 5117
rect 96522 5108 96528 5160
rect 96580 5148 96586 5160
rect 96617 5151 96675 5157
rect 96617 5148 96629 5151
rect 96580 5120 96629 5148
rect 96580 5108 96586 5120
rect 96617 5117 96629 5120
rect 96663 5117 96675 5151
rect 96617 5111 96675 5117
rect 96706 5108 96712 5160
rect 96764 5148 96770 5160
rect 98178 5148 98184 5160
rect 96764 5120 96809 5148
rect 98139 5120 98184 5148
rect 96764 5108 96770 5120
rect 98178 5108 98184 5120
rect 98236 5108 98242 5160
rect 99392 5148 99420 5188
rect 99466 5176 99472 5228
rect 99524 5216 99530 5228
rect 99653 5219 99711 5225
rect 99653 5216 99665 5219
rect 99524 5188 99665 5216
rect 99524 5176 99530 5188
rect 99653 5185 99665 5188
rect 99699 5185 99711 5219
rect 103992 5216 104020 5256
rect 105446 5216 105452 5228
rect 99653 5179 99711 5185
rect 99760 5188 104020 5216
rect 105407 5188 105452 5216
rect 99760 5148 99788 5188
rect 105446 5176 105452 5188
rect 105504 5176 105510 5228
rect 106366 5216 106372 5228
rect 106327 5188 106372 5216
rect 106366 5176 106372 5188
rect 106424 5176 106430 5228
rect 106550 5176 106556 5228
rect 106608 5216 106614 5228
rect 111794 5216 111800 5228
rect 106608 5188 111800 5216
rect 106608 5176 106614 5188
rect 111794 5176 111800 5188
rect 111852 5176 111858 5228
rect 112349 5219 112407 5225
rect 112349 5185 112361 5219
rect 112395 5216 112407 5219
rect 113082 5216 113088 5228
rect 112395 5188 113088 5216
rect 112395 5185 112407 5188
rect 112349 5179 112407 5185
rect 113082 5176 113088 5188
rect 113140 5176 113146 5228
rect 114925 5219 114983 5225
rect 114925 5185 114937 5219
rect 114971 5185 114983 5219
rect 114925 5179 114983 5185
rect 115937 5219 115995 5225
rect 115937 5185 115949 5219
rect 115983 5216 115995 5219
rect 116302 5216 116308 5228
rect 115983 5188 116308 5216
rect 115983 5185 115995 5188
rect 115937 5179 115995 5185
rect 99392 5120 99788 5148
rect 101217 5151 101275 5157
rect 101217 5117 101229 5151
rect 101263 5148 101275 5151
rect 102870 5148 102876 5160
rect 101263 5120 102876 5148
rect 101263 5117 101275 5120
rect 101217 5111 101275 5117
rect 102870 5108 102876 5120
rect 102928 5108 102934 5160
rect 102965 5151 103023 5157
rect 102965 5117 102977 5151
rect 103011 5148 103023 5151
rect 103977 5151 104035 5157
rect 103977 5148 103989 5151
rect 103011 5120 103989 5148
rect 103011 5117 103023 5120
rect 102965 5111 103023 5117
rect 103977 5117 103989 5120
rect 104023 5117 104035 5151
rect 105078 5148 105084 5160
rect 105039 5120 105084 5148
rect 103977 5111 104035 5117
rect 105078 5108 105084 5120
rect 105136 5108 105142 5160
rect 105170 5108 105176 5160
rect 105228 5148 105234 5160
rect 106274 5148 106280 5160
rect 105228 5120 106280 5148
rect 105228 5108 105234 5120
rect 106274 5108 106280 5120
rect 106332 5108 106338 5160
rect 108114 5148 108120 5160
rect 106384 5120 106688 5148
rect 108075 5120 108120 5148
rect 72878 5040 72884 5092
rect 72936 5080 72942 5092
rect 106384 5080 106412 5120
rect 72936 5052 106412 5080
rect 106660 5080 106688 5120
rect 108114 5108 108120 5120
rect 108172 5108 108178 5160
rect 108209 5151 108267 5157
rect 108209 5117 108221 5151
rect 108255 5148 108267 5151
rect 108390 5148 108396 5160
rect 108255 5120 108396 5148
rect 108255 5117 108267 5120
rect 108209 5111 108267 5117
rect 108390 5108 108396 5120
rect 108448 5108 108454 5160
rect 108577 5151 108635 5157
rect 108577 5117 108589 5151
rect 108623 5148 108635 5151
rect 110230 5148 110236 5160
rect 108623 5120 110236 5148
rect 108623 5117 108635 5120
rect 108577 5111 108635 5117
rect 110230 5108 110236 5120
rect 110288 5108 110294 5160
rect 110414 5148 110420 5160
rect 110375 5120 110420 5148
rect 110414 5108 110420 5120
rect 110472 5108 110478 5160
rect 110598 5148 110604 5160
rect 110559 5120 110604 5148
rect 110598 5108 110604 5120
rect 110656 5108 110662 5160
rect 110969 5151 111027 5157
rect 110969 5117 110981 5151
rect 111015 5117 111027 5151
rect 110969 5111 111027 5117
rect 110874 5080 110880 5092
rect 106660 5052 110880 5080
rect 72936 5040 72942 5052
rect 110874 5040 110880 5052
rect 110932 5040 110938 5092
rect 110984 5080 111012 5111
rect 111426 5108 111432 5160
rect 111484 5148 111490 5160
rect 113453 5151 113511 5157
rect 113453 5148 113465 5151
rect 111484 5120 113465 5148
rect 111484 5108 111490 5120
rect 113453 5117 113465 5120
rect 113499 5117 113511 5151
rect 113453 5111 113511 5117
rect 112990 5080 112996 5092
rect 110984 5052 112996 5080
rect 112990 5040 112996 5052
rect 113048 5040 113054 5092
rect 113082 5040 113088 5092
rect 113140 5080 113146 5092
rect 114830 5080 114836 5092
rect 113140 5052 114836 5080
rect 113140 5040 113146 5052
rect 114830 5040 114836 5052
rect 114888 5040 114894 5092
rect 67784 4984 72096 5012
rect 67784 4972 67790 4984
rect 77018 4972 77024 5024
rect 77076 5012 77082 5024
rect 78401 5015 78459 5021
rect 78401 5012 78413 5015
rect 77076 4984 78413 5012
rect 77076 4972 77082 4984
rect 78401 4981 78413 4984
rect 78447 4981 78459 5015
rect 78401 4975 78459 4981
rect 81434 4972 81440 5024
rect 81492 5012 81498 5024
rect 82909 5015 82967 5021
rect 82909 5012 82921 5015
rect 81492 4984 82921 5012
rect 81492 4972 81498 4984
rect 82909 4981 82921 4984
rect 82955 4981 82967 5015
rect 82909 4975 82967 4981
rect 88702 4972 88708 5024
rect 88760 5012 88766 5024
rect 94682 5012 94688 5024
rect 88760 4984 94688 5012
rect 88760 4972 88766 4984
rect 94682 4972 94688 4984
rect 94740 4972 94746 5024
rect 95050 4972 95056 5024
rect 95108 5012 95114 5024
rect 96614 5012 96620 5024
rect 95108 4984 96620 5012
rect 95108 4972 95114 4984
rect 96614 4972 96620 4984
rect 96672 4972 96678 5024
rect 99561 5015 99619 5021
rect 99561 4981 99573 5015
rect 99607 5012 99619 5015
rect 106366 5012 106372 5024
rect 99607 4984 106372 5012
rect 99607 4981 99619 4984
rect 99561 4975 99619 4981
rect 106366 4972 106372 4984
rect 106424 4972 106430 5024
rect 106550 4972 106556 5024
rect 106608 5012 106614 5024
rect 113818 5012 113824 5024
rect 106608 4984 113824 5012
rect 106608 4972 106614 4984
rect 113818 4972 113824 4984
rect 113876 4972 113882 5024
rect 114940 5012 114968 5179
rect 116302 5176 116308 5188
rect 116360 5176 116366 5228
rect 116412 5216 116440 5256
rect 117409 5253 117421 5287
rect 117455 5284 117467 5287
rect 121840 5284 121868 5324
rect 123478 5312 123484 5324
rect 123536 5312 123542 5364
rect 123570 5312 123576 5364
rect 123628 5352 123634 5364
rect 124766 5352 124772 5364
rect 123628 5324 124772 5352
rect 123628 5312 123634 5324
rect 124766 5312 124772 5324
rect 124824 5312 124830 5364
rect 129366 5352 129372 5364
rect 126164 5324 129372 5352
rect 117455 5256 121868 5284
rect 117455 5253 117467 5256
rect 117409 5247 117467 5253
rect 122006 5244 122012 5296
rect 122064 5284 122070 5296
rect 124674 5284 124680 5296
rect 122064 5256 124680 5284
rect 122064 5244 122070 5256
rect 124674 5244 124680 5256
rect 124732 5244 124738 5296
rect 126164 5293 126192 5324
rect 129366 5312 129372 5324
rect 129424 5312 129430 5364
rect 129734 5312 129740 5364
rect 129792 5352 129798 5364
rect 131206 5352 131212 5364
rect 129792 5324 131212 5352
rect 129792 5312 129798 5324
rect 131206 5312 131212 5324
rect 131264 5312 131270 5364
rect 131298 5312 131304 5364
rect 131356 5352 131362 5364
rect 138198 5352 138204 5364
rect 131356 5324 138204 5352
rect 131356 5312 131362 5324
rect 138198 5312 138204 5324
rect 138256 5312 138262 5364
rect 144822 5352 144828 5364
rect 139688 5324 144828 5352
rect 126149 5287 126207 5293
rect 126149 5253 126161 5287
rect 126195 5253 126207 5287
rect 126149 5247 126207 5253
rect 126238 5244 126244 5296
rect 126296 5284 126302 5296
rect 128725 5287 128783 5293
rect 126296 5256 128676 5284
rect 126296 5244 126302 5256
rect 118510 5216 118516 5228
rect 116412 5188 118516 5216
rect 118510 5176 118516 5188
rect 118568 5176 118574 5228
rect 121733 5219 121791 5225
rect 121733 5185 121745 5219
rect 121779 5216 121791 5219
rect 128170 5216 128176 5228
rect 121779 5188 128176 5216
rect 121779 5185 121791 5188
rect 121733 5179 121791 5185
rect 128170 5176 128176 5188
rect 128228 5176 128234 5228
rect 128648 5216 128676 5256
rect 128725 5253 128737 5287
rect 128771 5284 128783 5287
rect 131022 5284 131028 5296
rect 128771 5256 131028 5284
rect 128771 5253 128783 5256
rect 128725 5247 128783 5253
rect 131022 5244 131028 5256
rect 131080 5244 131086 5296
rect 137278 5284 137284 5296
rect 131224 5256 137284 5284
rect 131114 5216 131120 5228
rect 128648 5188 130424 5216
rect 131075 5188 131120 5216
rect 115017 5151 115075 5157
rect 115017 5117 115029 5151
rect 115063 5117 115075 5151
rect 115017 5111 115075 5117
rect 115032 5080 115060 5111
rect 115106 5108 115112 5160
rect 115164 5148 115170 5160
rect 117222 5148 117228 5160
rect 115164 5120 117228 5148
rect 115164 5108 115170 5120
rect 117222 5108 117228 5120
rect 117280 5108 117286 5160
rect 117501 5151 117559 5157
rect 117501 5117 117513 5151
rect 117547 5148 117559 5151
rect 119249 5151 119307 5157
rect 117547 5120 119200 5148
rect 117547 5117 117559 5120
rect 117501 5111 117559 5117
rect 118786 5080 118792 5092
rect 115032 5052 118792 5080
rect 118786 5040 118792 5052
rect 118844 5040 118850 5092
rect 119172 5080 119200 5120
rect 119249 5117 119261 5151
rect 119295 5148 119307 5151
rect 120261 5151 120319 5157
rect 120261 5148 120273 5151
rect 119295 5120 120273 5148
rect 119295 5117 119307 5120
rect 119249 5111 119307 5117
rect 120261 5117 120273 5120
rect 120307 5117 120319 5151
rect 120261 5111 120319 5117
rect 121825 5151 121883 5157
rect 121825 5117 121837 5151
rect 121871 5148 121883 5151
rect 123294 5148 123300 5160
rect 121871 5120 123300 5148
rect 121871 5117 121883 5120
rect 121825 5111 121883 5117
rect 123294 5108 123300 5120
rect 123352 5108 123358 5160
rect 123565 5151 123623 5157
rect 123565 5117 123577 5151
rect 123611 5117 123623 5151
rect 124674 5148 124680 5160
rect 124635 5120 124680 5148
rect 123565 5111 123623 5117
rect 123478 5080 123484 5092
rect 119172 5052 123484 5080
rect 123478 5040 123484 5052
rect 123536 5040 123542 5092
rect 123588 5080 123616 5111
rect 124674 5108 124680 5120
rect 124732 5108 124738 5160
rect 126238 5148 126244 5160
rect 126199 5120 126244 5148
rect 126238 5108 126244 5120
rect 126296 5108 126302 5160
rect 127253 5151 127311 5157
rect 127253 5117 127265 5151
rect 127299 5148 127311 5151
rect 128630 5148 128636 5160
rect 127299 5120 128636 5148
rect 127299 5117 127311 5120
rect 127253 5111 127311 5117
rect 128630 5108 128636 5120
rect 128688 5108 128694 5160
rect 128817 5151 128875 5157
rect 128817 5117 128829 5151
rect 128863 5148 128875 5151
rect 130194 5148 130200 5160
rect 128863 5120 130200 5148
rect 128863 5117 128875 5120
rect 128817 5111 128875 5117
rect 130194 5108 130200 5120
rect 130252 5108 130258 5160
rect 130396 5080 130424 5188
rect 131114 5176 131120 5188
rect 131172 5176 131178 5228
rect 130470 5108 130476 5160
rect 130528 5148 130534 5160
rect 131224 5148 131252 5256
rect 137278 5244 137284 5256
rect 137336 5244 137342 5296
rect 137373 5287 137431 5293
rect 137373 5253 137385 5287
rect 137419 5284 137431 5287
rect 139688 5284 139716 5324
rect 144822 5312 144828 5324
rect 144880 5312 144886 5364
rect 145374 5312 145380 5364
rect 145432 5352 145438 5364
rect 155954 5352 155960 5364
rect 145432 5324 155960 5352
rect 145432 5312 145438 5324
rect 155954 5312 155960 5324
rect 156012 5312 156018 5364
rect 137419 5256 139716 5284
rect 139765 5287 139823 5293
rect 137419 5253 137431 5256
rect 137373 5247 137431 5253
rect 139765 5253 139777 5287
rect 139811 5284 139823 5287
rect 149606 5284 149612 5296
rect 139811 5256 149612 5284
rect 139811 5253 139823 5256
rect 139765 5247 139823 5253
rect 149606 5244 149612 5256
rect 149664 5244 149670 5296
rect 131482 5176 131488 5228
rect 131540 5216 131546 5228
rect 131540 5188 132356 5216
rect 131540 5176 131546 5188
rect 132218 5148 132224 5160
rect 130528 5120 131252 5148
rect 132179 5120 132224 5148
rect 130528 5108 130534 5120
rect 132218 5108 132224 5120
rect 132276 5108 132282 5160
rect 132328 5148 132356 5188
rect 132402 5176 132408 5228
rect 132460 5216 132466 5228
rect 132460 5188 132505 5216
rect 132460 5176 132466 5188
rect 132586 5176 132592 5228
rect 132644 5216 132650 5228
rect 133322 5216 133328 5228
rect 132644 5188 133328 5216
rect 132644 5176 132650 5188
rect 133322 5176 133328 5188
rect 133380 5176 133386 5228
rect 133506 5216 133512 5228
rect 133467 5188 133512 5216
rect 133506 5176 133512 5188
rect 133564 5176 133570 5228
rect 133966 5176 133972 5228
rect 134024 5216 134030 5228
rect 135070 5216 135076 5228
rect 134024 5188 135076 5216
rect 134024 5176 134030 5188
rect 135070 5176 135076 5188
rect 135128 5176 135134 5228
rect 135346 5176 135352 5228
rect 135404 5216 135410 5228
rect 135901 5219 135959 5225
rect 135901 5216 135913 5219
rect 135404 5188 135913 5216
rect 135404 5176 135410 5188
rect 135901 5185 135913 5188
rect 135947 5185 135959 5219
rect 135901 5179 135959 5185
rect 136174 5176 136180 5228
rect 136232 5216 136238 5228
rect 137186 5216 137192 5228
rect 136232 5188 137192 5216
rect 136232 5176 136238 5188
rect 137186 5176 137192 5188
rect 137244 5176 137250 5228
rect 137388 5188 137600 5216
rect 137388 5160 137416 5188
rect 137002 5148 137008 5160
rect 132328 5120 137008 5148
rect 137002 5108 137008 5120
rect 137060 5108 137066 5160
rect 137370 5108 137376 5160
rect 137428 5108 137434 5160
rect 137465 5151 137523 5157
rect 137465 5117 137477 5151
rect 137511 5117 137523 5151
rect 137572 5148 137600 5188
rect 137646 5176 137652 5228
rect 137704 5216 137710 5228
rect 142614 5216 142620 5228
rect 137704 5188 142620 5216
rect 137704 5176 137710 5188
rect 142614 5176 142620 5188
rect 142672 5176 142678 5228
rect 143169 5219 143227 5225
rect 143169 5185 143181 5219
rect 143215 5216 143227 5219
rect 143258 5216 143264 5228
rect 143215 5188 143264 5216
rect 143215 5185 143227 5188
rect 143169 5179 143227 5185
rect 143258 5176 143264 5188
rect 143316 5176 143322 5228
rect 144362 5216 144368 5228
rect 144323 5188 144368 5216
rect 144362 5176 144368 5188
rect 144420 5176 144426 5228
rect 144472 5188 144776 5216
rect 138293 5151 138351 5157
rect 138293 5148 138305 5151
rect 137572 5120 138305 5148
rect 137465 5111 137523 5117
rect 138293 5117 138305 5120
rect 138339 5117 138351 5151
rect 138293 5111 138351 5117
rect 139857 5151 139915 5157
rect 139857 5117 139869 5151
rect 139903 5148 139915 5151
rect 143350 5148 143356 5160
rect 139903 5120 143356 5148
rect 139903 5117 139915 5120
rect 139857 5111 139915 5117
rect 131114 5080 131120 5092
rect 123588 5052 128492 5080
rect 130396 5052 131120 5080
rect 121270 5012 121276 5024
rect 114940 4984 121276 5012
rect 121270 4972 121276 4984
rect 121328 4972 121334 5024
rect 121362 4972 121368 5024
rect 121420 5012 121426 5024
rect 123665 5015 123723 5021
rect 123665 5012 123677 5015
rect 121420 4984 123677 5012
rect 121420 4972 121426 4984
rect 123665 4981 123677 4984
rect 123711 4981 123723 5015
rect 123665 4975 123723 4981
rect 123754 4972 123760 5024
rect 123812 5012 123818 5024
rect 126054 5012 126060 5024
rect 123812 4984 126060 5012
rect 123812 4972 123818 4984
rect 126054 4972 126060 4984
rect 126112 4972 126118 5024
rect 126698 4972 126704 5024
rect 126756 5012 126762 5024
rect 128078 5012 128084 5024
rect 126756 4984 128084 5012
rect 126756 4972 126762 4984
rect 128078 4972 128084 4984
rect 128136 4972 128142 5024
rect 128464 5012 128492 5052
rect 131114 5040 131120 5052
rect 131172 5040 131178 5092
rect 131206 5040 131212 5092
rect 131264 5080 131270 5092
rect 136818 5080 136824 5092
rect 131264 5052 136824 5080
rect 131264 5040 131270 5052
rect 136818 5040 136824 5052
rect 136876 5040 136882 5092
rect 137480 5080 137508 5111
rect 143350 5108 143356 5120
rect 143408 5108 143414 5160
rect 138842 5080 138848 5092
rect 137480 5052 138848 5080
rect 138842 5040 138848 5052
rect 138900 5040 138906 5092
rect 144472 5080 144500 5188
rect 144549 5151 144607 5157
rect 144549 5117 144561 5151
rect 144595 5117 144607 5151
rect 144549 5111 144607 5117
rect 138952 5052 144500 5080
rect 132586 5012 132592 5024
rect 128464 4984 132592 5012
rect 132586 4972 132592 4984
rect 132644 4972 132650 5024
rect 132678 4972 132684 5024
rect 132736 5012 132742 5024
rect 133598 5012 133604 5024
rect 132736 4984 133604 5012
rect 132736 4972 132742 4984
rect 133598 4972 133604 4984
rect 133656 4972 133662 5024
rect 133782 4972 133788 5024
rect 133840 5012 133846 5024
rect 134334 5012 134340 5024
rect 133840 4984 134340 5012
rect 133840 4972 133846 4984
rect 134334 4972 134340 4984
rect 134392 4972 134398 5024
rect 134518 5012 134524 5024
rect 134479 4984 134524 5012
rect 134518 4972 134524 4984
rect 134576 4972 134582 5024
rect 134610 4972 134616 5024
rect 134668 5012 134674 5024
rect 138952 5012 138980 5052
rect 134668 4984 138980 5012
rect 134668 4972 134674 4984
rect 140774 4972 140780 5024
rect 140832 5012 140838 5024
rect 141513 5015 141571 5021
rect 141513 5012 141525 5015
rect 140832 4984 141525 5012
rect 140832 4972 140838 4984
rect 141513 4981 141525 4984
rect 141559 4981 141571 5015
rect 144564 5012 144592 5111
rect 144748 5080 144776 5188
rect 144822 5176 144828 5228
rect 144880 5216 144886 5228
rect 146386 5216 146392 5228
rect 144880 5188 146392 5216
rect 144880 5176 144886 5188
rect 146386 5176 146392 5188
rect 146444 5176 146450 5228
rect 153286 5216 153292 5228
rect 153247 5188 153292 5216
rect 153286 5176 153292 5188
rect 153344 5176 153350 5228
rect 156506 5080 156512 5092
rect 144748 5052 156512 5080
rect 156506 5040 156512 5052
rect 156564 5040 156570 5092
rect 144822 5012 144828 5024
rect 144564 4984 144828 5012
rect 141513 4975 141571 4981
rect 144822 4972 144828 4984
rect 144880 4972 144886 5024
rect 1104 4922 154560 4944
rect 1104 4870 24078 4922
rect 24130 4870 64078 4922
rect 64130 4870 104078 4922
rect 104130 4870 144078 4922
rect 144130 4870 154560 4922
rect 1104 4848 154560 4870
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 15286 4808 15292 4820
rect 15247 4780 15292 4808
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 18046 4808 18052 4820
rect 16807 4780 18052 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 19334 4808 19340 4820
rect 19295 4780 19340 4808
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 20438 4768 20444 4820
rect 20496 4808 20502 4820
rect 20901 4811 20959 4817
rect 20901 4808 20913 4811
rect 20496 4780 20913 4808
rect 20496 4768 20502 4780
rect 20901 4777 20913 4780
rect 20947 4777 20959 4811
rect 20901 4771 20959 4777
rect 21266 4768 21272 4820
rect 21324 4808 21330 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 21324 4780 21925 4808
rect 21324 4768 21330 4780
rect 21913 4777 21925 4780
rect 21959 4777 21971 4811
rect 36078 4808 36084 4820
rect 36039 4780 36084 4808
rect 21913 4771 21971 4777
rect 36078 4768 36084 4780
rect 36136 4768 36142 4820
rect 37734 4808 37740 4820
rect 37695 4780 37740 4808
rect 37734 4768 37740 4780
rect 37792 4768 37798 4820
rect 43441 4811 43499 4817
rect 43441 4777 43453 4811
rect 43487 4808 43499 4811
rect 43622 4808 43628 4820
rect 43487 4780 43628 4808
rect 43487 4777 43499 4780
rect 43441 4771 43499 4777
rect 43622 4768 43628 4780
rect 43680 4768 43686 4820
rect 46106 4768 46112 4820
rect 46164 4808 46170 4820
rect 47489 4811 47547 4817
rect 47489 4808 47501 4811
rect 46164 4780 47501 4808
rect 46164 4768 46170 4780
rect 47489 4777 47501 4780
rect 47535 4777 47547 4811
rect 47489 4771 47547 4777
rect 54846 4768 54852 4820
rect 54904 4808 54910 4820
rect 57057 4811 57115 4817
rect 57057 4808 57069 4811
rect 54904 4780 57069 4808
rect 54904 4768 54910 4780
rect 57057 4777 57069 4780
rect 57103 4777 57115 4811
rect 57057 4771 57115 4777
rect 61654 4768 61660 4820
rect 61712 4808 61718 4820
rect 62577 4811 62635 4817
rect 62577 4808 62589 4811
rect 61712 4780 62589 4808
rect 61712 4768 61718 4780
rect 62577 4777 62589 4780
rect 62623 4777 62635 4811
rect 62577 4771 62635 4777
rect 63218 4768 63224 4820
rect 63276 4808 63282 4820
rect 63589 4811 63647 4817
rect 63589 4808 63601 4811
rect 63276 4780 63601 4808
rect 63276 4768 63282 4780
rect 63589 4777 63601 4780
rect 63635 4777 63647 4811
rect 63589 4771 63647 4777
rect 66901 4811 66959 4817
rect 66901 4777 66913 4811
rect 66947 4808 66959 4811
rect 67450 4808 67456 4820
rect 66947 4780 67456 4808
rect 66947 4777 66959 4780
rect 66901 4771 66959 4777
rect 67450 4768 67456 4780
rect 67508 4768 67514 4820
rect 71314 4768 71320 4820
rect 71372 4808 71378 4820
rect 82633 4811 82691 4817
rect 71372 4780 77524 4808
rect 71372 4768 71378 4780
rect 52730 4740 52736 4752
rect 50540 4712 52736 4740
rect 5718 4672 5724 4684
rect 5679 4644 5724 4672
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 7006 4672 7012 4684
rect 6967 4644 7012 4672
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 10962 4672 10968 4684
rect 10923 4644 10968 4672
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 12526 4672 12532 4684
rect 12487 4644 12532 4672
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 23566 4632 23572 4684
rect 23624 4672 23630 4684
rect 24213 4675 24271 4681
rect 24213 4672 24225 4675
rect 23624 4644 24225 4672
rect 23624 4632 23630 4644
rect 24213 4641 24225 4644
rect 24259 4641 24271 4675
rect 24213 4635 24271 4641
rect 29825 4675 29883 4681
rect 29825 4641 29837 4675
rect 29871 4672 29883 4675
rect 32306 4672 32312 4684
rect 29871 4644 32312 4672
rect 29871 4641 29883 4644
rect 29825 4635 29883 4641
rect 32306 4632 32312 4644
rect 32364 4632 32370 4684
rect 34241 4675 34299 4681
rect 34241 4641 34253 4675
rect 34287 4672 34299 4675
rect 34974 4672 34980 4684
rect 34287 4644 34980 4672
rect 34287 4641 34299 4644
rect 34241 4635 34299 4641
rect 34974 4632 34980 4644
rect 35032 4632 35038 4684
rect 42337 4675 42395 4681
rect 42337 4641 42349 4675
rect 42383 4641 42395 4675
rect 42337 4635 42395 4641
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 3007 4576 4629 4604
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 4617 4573 4629 4576
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6270 4604 6276 4616
rect 6135 4576 6276 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 8570 4604 8576 4616
rect 8527 4576 8576 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 9674 4604 9680 4616
rect 9635 4576 9680 4604
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 13262 4604 13268 4616
rect 12483 4576 13268 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 23109 4607 23167 4613
rect 23109 4573 23121 4607
rect 23155 4604 23167 4607
rect 23842 4604 23848 4616
rect 23155 4576 23848 4604
rect 23155 4573 23167 4576
rect 23109 4567 23167 4573
rect 23842 4564 23848 4576
rect 23900 4564 23906 4616
rect 24121 4607 24179 4613
rect 24121 4573 24133 4607
rect 24167 4573 24179 4607
rect 26970 4604 26976 4616
rect 26931 4576 26976 4604
rect 24121 4567 24179 4573
rect 20898 4496 20904 4548
rect 20956 4536 20962 4548
rect 24136 4536 24164 4567
rect 26970 4564 26976 4576
rect 27028 4564 27034 4616
rect 28258 4604 28264 4616
rect 28219 4576 28264 4604
rect 28258 4564 28264 4576
rect 28316 4564 28322 4616
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4604 29791 4607
rect 30558 4604 30564 4616
rect 29779 4576 30564 4604
rect 29779 4573 29791 4576
rect 29733 4567 29791 4573
rect 30558 4564 30564 4576
rect 30616 4564 30622 4616
rect 30742 4604 30748 4616
rect 30703 4576 30748 4604
rect 30742 4564 30748 4576
rect 30800 4564 30806 4616
rect 32677 4607 32735 4613
rect 32677 4573 32689 4607
rect 32723 4604 32735 4607
rect 33502 4604 33508 4616
rect 32723 4576 33508 4604
rect 32723 4573 32735 4576
rect 32677 4567 32735 4573
rect 33502 4564 33508 4576
rect 33560 4564 33566 4616
rect 33686 4604 33692 4616
rect 33647 4576 33692 4604
rect 33686 4564 33692 4576
rect 33744 4564 33750 4616
rect 33778 4564 33784 4616
rect 33836 4604 33842 4616
rect 35069 4607 35127 4613
rect 35069 4604 35081 4607
rect 33836 4576 35081 4604
rect 33836 4564 33842 4576
rect 35069 4573 35081 4576
rect 35115 4573 35127 4607
rect 40770 4604 40776 4616
rect 40731 4576 40776 4604
rect 35069 4567 35127 4573
rect 40770 4564 40776 4576
rect 40828 4564 40834 4616
rect 42058 4604 42064 4616
rect 42019 4576 42064 4604
rect 42058 4564 42064 4576
rect 42116 4564 42122 4616
rect 42352 4604 42380 4635
rect 42794 4632 42800 4684
rect 42852 4672 42858 4684
rect 43349 4675 43407 4681
rect 43349 4672 43361 4675
rect 42852 4644 43361 4672
rect 42852 4632 42858 4644
rect 43349 4641 43361 4644
rect 43395 4641 43407 4675
rect 43349 4635 43407 4641
rect 46661 4675 46719 4681
rect 46661 4641 46673 4675
rect 46707 4672 46719 4675
rect 47302 4672 47308 4684
rect 46707 4644 47308 4672
rect 46707 4641 46719 4644
rect 46661 4635 46719 4641
rect 47302 4632 47308 4644
rect 47360 4632 47366 4684
rect 50540 4681 50568 4712
rect 52730 4700 52736 4712
rect 52788 4700 52794 4752
rect 77386 4740 77392 4752
rect 72988 4712 77392 4740
rect 50525 4675 50583 4681
rect 50525 4641 50537 4675
rect 50571 4641 50583 4675
rect 51718 4672 51724 4684
rect 51679 4644 51724 4672
rect 50525 4635 50583 4641
rect 51718 4632 51724 4644
rect 51776 4632 51782 4684
rect 53285 4675 53343 4681
rect 53285 4641 53297 4675
rect 53331 4672 53343 4675
rect 54754 4672 54760 4684
rect 53331 4644 54760 4672
rect 53331 4641 53343 4644
rect 53285 4635 53343 4641
rect 54754 4632 54760 4644
rect 54812 4632 54818 4684
rect 56226 4672 56232 4684
rect 56187 4644 56232 4672
rect 56226 4632 56232 4644
rect 56284 4632 56290 4684
rect 59538 4632 59544 4684
rect 59596 4672 59602 4684
rect 61289 4675 61347 4681
rect 61289 4672 61301 4675
rect 59596 4644 61301 4672
rect 59596 4632 59602 4644
rect 61289 4641 61301 4644
rect 61335 4641 61347 4675
rect 70486 4672 70492 4684
rect 70447 4644 70492 4672
rect 61289 4635 61347 4641
rect 70486 4632 70492 4644
rect 70544 4632 70550 4684
rect 72988 4681 73016 4712
rect 77386 4700 77392 4712
rect 77444 4700 77450 4752
rect 72973 4675 73031 4681
rect 72973 4641 72985 4675
rect 73019 4641 73031 4675
rect 72973 4635 73031 4641
rect 73062 4632 73068 4684
rect 73120 4672 73126 4684
rect 77496 4681 77524 4780
rect 82633 4777 82645 4811
rect 82679 4808 82691 4811
rect 82906 4808 82912 4820
rect 82679 4780 82912 4808
rect 82679 4777 82691 4780
rect 82633 4771 82691 4777
rect 82906 4768 82912 4780
rect 82964 4768 82970 4820
rect 87141 4811 87199 4817
rect 87141 4777 87153 4811
rect 87187 4808 87199 4811
rect 88518 4808 88524 4820
rect 87187 4780 88524 4808
rect 87187 4777 87199 4780
rect 87141 4771 87199 4777
rect 88518 4768 88524 4780
rect 88576 4768 88582 4820
rect 88702 4808 88708 4820
rect 88663 4780 88708 4808
rect 88702 4768 88708 4780
rect 88760 4768 88766 4820
rect 88978 4768 88984 4820
rect 89036 4808 89042 4820
rect 102594 4808 102600 4820
rect 89036 4780 102600 4808
rect 89036 4768 89042 4780
rect 102594 4768 102600 4780
rect 102652 4768 102658 4820
rect 106090 4808 106096 4820
rect 103716 4780 106096 4808
rect 79962 4700 79968 4752
rect 80020 4740 80026 4752
rect 99282 4740 99288 4752
rect 80020 4712 86540 4740
rect 80020 4700 80026 4712
rect 74537 4675 74595 4681
rect 74537 4672 74549 4675
rect 73120 4644 74549 4672
rect 73120 4632 73126 4644
rect 74537 4641 74549 4644
rect 74583 4641 74595 4675
rect 74537 4635 74595 4641
rect 77481 4675 77539 4681
rect 77481 4641 77493 4675
rect 77527 4641 77539 4675
rect 81066 4672 81072 4684
rect 81027 4644 81072 4672
rect 77481 4635 77539 4641
rect 81066 4632 81072 4644
rect 81124 4632 81130 4684
rect 83918 4672 83924 4684
rect 83879 4644 83924 4672
rect 83918 4632 83924 4644
rect 83976 4632 83982 4684
rect 84378 4672 84384 4684
rect 84339 4644 84384 4672
rect 84378 4632 84384 4644
rect 84436 4632 84442 4684
rect 85574 4672 85580 4684
rect 85535 4644 85580 4672
rect 85574 4632 85580 4644
rect 85632 4632 85638 4684
rect 86221 4675 86279 4681
rect 86221 4641 86233 4675
rect 86267 4672 86279 4675
rect 86402 4672 86408 4684
rect 86267 4644 86408 4672
rect 86267 4641 86279 4644
rect 86221 4635 86279 4641
rect 86402 4632 86408 4644
rect 86460 4632 86466 4684
rect 86512 4672 86540 4712
rect 89364 4712 97304 4740
rect 87049 4675 87107 4681
rect 87049 4672 87061 4675
rect 86512 4644 87061 4672
rect 87049 4641 87061 4644
rect 87095 4641 87107 4675
rect 87049 4635 87107 4641
rect 88889 4675 88947 4681
rect 88889 4641 88901 4675
rect 88935 4672 88947 4675
rect 89254 4672 89260 4684
rect 88935 4644 89260 4672
rect 88935 4641 88947 4644
rect 88889 4635 88947 4641
rect 89254 4632 89260 4644
rect 89312 4632 89318 4684
rect 44358 4604 44364 4616
rect 42352 4576 44364 4604
rect 44358 4564 44364 4576
rect 44416 4564 44422 4616
rect 45094 4604 45100 4616
rect 45055 4576 45100 4604
rect 45094 4564 45100 4576
rect 45152 4564 45158 4616
rect 46569 4607 46627 4613
rect 46569 4573 46581 4607
rect 46615 4604 46627 4607
rect 48130 4604 48136 4616
rect 46615 4576 48136 4604
rect 46615 4573 46627 4576
rect 46569 4567 46627 4573
rect 48130 4564 48136 4576
rect 48188 4564 48194 4616
rect 48958 4604 48964 4616
rect 48919 4576 48964 4604
rect 48958 4564 48964 4576
rect 49016 4564 49022 4616
rect 50433 4607 50491 4613
rect 50433 4573 50445 4607
rect 50479 4604 50491 4607
rect 51994 4604 52000 4616
rect 50479 4576 52000 4604
rect 50479 4573 50491 4576
rect 50433 4567 50491 4573
rect 51994 4564 52000 4576
rect 52052 4564 52058 4616
rect 53193 4607 53251 4613
rect 53193 4573 53205 4607
rect 53239 4604 53251 4607
rect 54202 4604 54208 4616
rect 53239 4576 54208 4604
rect 53239 4573 53251 4576
rect 53193 4567 53251 4573
rect 54202 4564 54208 4576
rect 54260 4564 54266 4616
rect 54665 4607 54723 4613
rect 54665 4573 54677 4607
rect 54711 4573 54723 4607
rect 58066 4604 58072 4616
rect 58027 4576 58072 4604
rect 54665 4567 54723 4573
rect 20956 4508 24164 4536
rect 20956 4496 20962 4508
rect 52362 4496 52368 4548
rect 52420 4536 52426 4548
rect 54680 4536 54708 4567
rect 58066 4564 58072 4576
rect 58124 4564 58130 4616
rect 59081 4607 59139 4613
rect 59081 4573 59093 4607
rect 59127 4604 59139 4607
rect 60185 4607 60243 4613
rect 60185 4604 60197 4607
rect 59127 4576 60197 4604
rect 59127 4573 59139 4576
rect 59081 4567 59139 4573
rect 60185 4573 60197 4576
rect 60231 4573 60243 4607
rect 61194 4604 61200 4616
rect 61155 4576 61200 4604
rect 60185 4567 60243 4573
rect 61194 4564 61200 4576
rect 61252 4564 61258 4616
rect 67913 4607 67971 4613
rect 67913 4573 67925 4607
rect 67959 4604 67971 4607
rect 68925 4607 68983 4613
rect 68925 4604 68937 4607
rect 67959 4576 68937 4604
rect 67959 4573 67971 4576
rect 67913 4567 67971 4573
rect 68925 4573 68937 4576
rect 68971 4573 68983 4607
rect 70302 4604 70308 4616
rect 70263 4576 70308 4604
rect 68925 4567 68983 4573
rect 70302 4564 70308 4576
rect 70360 4564 70366 4616
rect 71406 4604 71412 4616
rect 71367 4576 71412 4604
rect 71406 4564 71412 4576
rect 71464 4564 71470 4616
rect 72878 4604 72884 4616
rect 72839 4576 72884 4604
rect 72878 4564 72884 4576
rect 72936 4564 72942 4616
rect 74626 4564 74632 4616
rect 74684 4604 74690 4616
rect 77021 4607 77079 4613
rect 77021 4604 77033 4607
rect 74684 4576 77033 4604
rect 74684 4564 74690 4576
rect 77021 4573 77033 4576
rect 77067 4573 77079 4607
rect 79502 4604 79508 4616
rect 79463 4576 79508 4604
rect 77021 4567 77079 4573
rect 79502 4564 79508 4576
rect 79560 4564 79566 4616
rect 80977 4607 81035 4613
rect 80977 4573 80989 4607
rect 81023 4604 81035 4607
rect 88978 4604 88984 4616
rect 81023 4576 88984 4604
rect 81023 4573 81035 4576
rect 80977 4567 81035 4573
rect 88978 4564 88984 4576
rect 89036 4564 89042 4616
rect 52420 4508 54708 4536
rect 56137 4539 56195 4545
rect 52420 4496 52426 4508
rect 56137 4505 56149 4539
rect 56183 4536 56195 4539
rect 87049 4539 87107 4545
rect 56183 4508 75040 4536
rect 56183 4505 56195 4508
rect 56137 4499 56195 4505
rect 74718 4468 74724 4480
rect 74679 4440 74724 4468
rect 74718 4428 74724 4440
rect 74776 4428 74782 4480
rect 75012 4468 75040 4508
rect 80072 4508 85804 4536
rect 80072 4468 80100 4508
rect 75012 4440 80100 4468
rect 85577 4471 85635 4477
rect 85577 4437 85589 4471
rect 85623 4468 85635 4471
rect 85666 4468 85672 4480
rect 85623 4440 85672 4468
rect 85623 4437 85635 4440
rect 85577 4431 85635 4437
rect 85666 4428 85672 4440
rect 85724 4428 85730 4480
rect 85776 4468 85804 4508
rect 87049 4505 87061 4539
rect 87095 4536 87107 4539
rect 89364 4536 89392 4712
rect 92014 4672 92020 4684
rect 91975 4644 92020 4672
rect 92014 4632 92020 4644
rect 92072 4632 92078 4684
rect 92106 4632 92112 4684
rect 92164 4672 92170 4684
rect 93949 4675 94007 4681
rect 93949 4672 93961 4675
rect 92164 4644 93961 4672
rect 92164 4632 92170 4644
rect 93949 4641 93961 4644
rect 93995 4641 94007 4675
rect 96706 4672 96712 4684
rect 93949 4635 94007 4641
rect 94056 4644 96712 4672
rect 90450 4604 90456 4616
rect 90411 4576 90456 4604
rect 90450 4564 90456 4576
rect 90508 4564 90514 4616
rect 91922 4604 91928 4616
rect 91883 4576 91928 4604
rect 91922 4564 91928 4576
rect 91980 4564 91986 4616
rect 93026 4564 93032 4616
rect 93084 4604 93090 4616
rect 93857 4607 93915 4613
rect 93857 4604 93869 4607
rect 93084 4576 93869 4604
rect 93084 4564 93090 4576
rect 93857 4573 93869 4576
rect 93903 4573 93915 4607
rect 94056 4604 94084 4644
rect 96706 4632 96712 4644
rect 96764 4632 96770 4684
rect 95786 4604 95792 4616
rect 93857 4567 93915 4573
rect 93964 4576 94084 4604
rect 95747 4576 95792 4604
rect 87095 4508 89392 4536
rect 87095 4505 87107 4508
rect 87049 4499 87107 4505
rect 91830 4496 91836 4548
rect 91888 4536 91894 4548
rect 93964 4536 93992 4576
rect 95786 4564 95792 4576
rect 95844 4564 95850 4616
rect 97276 4604 97304 4712
rect 97368 4712 99288 4740
rect 97368 4681 97396 4712
rect 99282 4700 99288 4712
rect 99340 4700 99346 4752
rect 103606 4740 103612 4752
rect 99760 4712 103612 4740
rect 97353 4675 97411 4681
rect 97353 4641 97365 4675
rect 97399 4641 97411 4675
rect 99760 4672 99788 4712
rect 103606 4700 103612 4712
rect 103664 4700 103670 4752
rect 97353 4635 97411 4641
rect 97460 4644 99788 4672
rect 101033 4675 101091 4681
rect 97460 4604 97488 4644
rect 101033 4641 101045 4675
rect 101079 4672 101091 4675
rect 102134 4672 102140 4684
rect 101079 4644 102140 4672
rect 101079 4641 101091 4644
rect 101033 4635 101091 4641
rect 102134 4632 102140 4644
rect 102192 4632 102198 4684
rect 103716 4672 103744 4780
rect 106090 4768 106096 4780
rect 106148 4768 106154 4820
rect 106182 4768 106188 4820
rect 106240 4808 106246 4820
rect 111242 4808 111248 4820
rect 106240 4780 111248 4808
rect 106240 4768 106246 4780
rect 111242 4768 111248 4780
rect 111300 4768 111306 4820
rect 111426 4808 111432 4820
rect 111387 4780 111432 4808
rect 111426 4768 111432 4780
rect 111484 4768 111490 4820
rect 118602 4808 118608 4820
rect 111536 4780 118608 4808
rect 106550 4740 106556 4752
rect 102336 4644 103744 4672
rect 103900 4712 106556 4740
rect 97276 4576 97488 4604
rect 98365 4607 98423 4613
rect 98365 4573 98377 4607
rect 98411 4604 98423 4607
rect 99469 4607 99527 4613
rect 99469 4604 99481 4607
rect 98411 4576 99481 4604
rect 98411 4573 98423 4576
rect 98365 4567 98423 4573
rect 99469 4573 99481 4576
rect 99515 4573 99527 4607
rect 99469 4567 99527 4573
rect 100941 4607 100999 4613
rect 100941 4573 100953 4607
rect 100987 4604 100999 4607
rect 102336 4604 102364 4644
rect 102502 4604 102508 4616
rect 100987 4576 102364 4604
rect 102463 4576 102508 4604
rect 100987 4573 100999 4576
rect 100941 4567 100999 4573
rect 102502 4564 102508 4576
rect 102560 4564 102566 4616
rect 103900 4613 103928 4712
rect 106550 4700 106556 4712
rect 106608 4700 106614 4752
rect 106645 4743 106703 4749
rect 106645 4709 106657 4743
rect 106691 4740 106703 4743
rect 108022 4740 108028 4752
rect 106691 4712 108028 4740
rect 106691 4709 106703 4712
rect 106645 4703 106703 4709
rect 108022 4700 108028 4712
rect 108080 4700 108086 4752
rect 111536 4740 111564 4780
rect 118602 4768 118608 4780
rect 118660 4768 118666 4820
rect 118878 4768 118884 4820
rect 118936 4808 118942 4820
rect 124950 4808 124956 4820
rect 118936 4780 124956 4808
rect 118936 4768 118942 4780
rect 124950 4768 124956 4780
rect 125008 4768 125014 4820
rect 126238 4768 126244 4820
rect 126296 4808 126302 4820
rect 130841 4811 130899 4817
rect 130841 4808 130853 4811
rect 126296 4780 130853 4808
rect 126296 4768 126302 4780
rect 130841 4777 130853 4780
rect 130887 4777 130899 4811
rect 130841 4771 130899 4777
rect 130930 4768 130936 4820
rect 130988 4808 130994 4820
rect 131853 4811 131911 4817
rect 131853 4808 131865 4811
rect 130988 4780 131865 4808
rect 130988 4768 130994 4780
rect 131853 4777 131865 4780
rect 131899 4777 131911 4811
rect 137554 4808 137560 4820
rect 131853 4771 131911 4777
rect 132696 4780 137560 4808
rect 108132 4712 111564 4740
rect 104069 4675 104127 4681
rect 104069 4641 104081 4675
rect 104115 4672 104127 4675
rect 104894 4672 104900 4684
rect 104115 4644 104900 4672
rect 104115 4641 104127 4644
rect 104069 4635 104127 4641
rect 104894 4632 104900 4644
rect 104952 4632 104958 4684
rect 105354 4672 105360 4684
rect 105315 4644 105360 4672
rect 105354 4632 105360 4644
rect 105412 4632 105418 4684
rect 105630 4672 105636 4684
rect 105591 4644 105636 4672
rect 105630 4632 105636 4644
rect 105688 4632 105694 4684
rect 105740 4644 106136 4672
rect 103885 4607 103943 4613
rect 103885 4573 103897 4607
rect 103931 4573 103943 4607
rect 103885 4567 103943 4573
rect 104158 4564 104164 4616
rect 104216 4604 104222 4616
rect 105740 4604 105768 4644
rect 104216 4576 105768 4604
rect 106108 4604 106136 4644
rect 106182 4632 106188 4684
rect 106240 4672 106246 4684
rect 108132 4672 108160 4712
rect 113818 4700 113824 4752
rect 113876 4740 113882 4752
rect 119893 4743 119951 4749
rect 119893 4740 119905 4743
rect 113876 4712 119905 4740
rect 113876 4700 113882 4712
rect 119893 4709 119905 4712
rect 119939 4709 119951 4743
rect 119893 4703 119951 4709
rect 120000 4712 126284 4740
rect 106240 4644 108160 4672
rect 109313 4675 109371 4681
rect 106240 4632 106246 4644
rect 109313 4641 109325 4675
rect 109359 4672 109371 4675
rect 113082 4672 113088 4684
rect 109359 4644 113088 4672
rect 109359 4641 109371 4644
rect 109313 4635 109371 4641
rect 113082 4632 113088 4644
rect 113140 4632 113146 4684
rect 113545 4675 113603 4681
rect 113545 4641 113557 4675
rect 113591 4641 113603 4675
rect 113545 4635 113603 4641
rect 106645 4607 106703 4613
rect 106645 4604 106657 4607
rect 106108 4576 106657 4604
rect 104216 4564 104222 4576
rect 106645 4573 106657 4576
rect 106691 4573 106703 4607
rect 106645 4567 106703 4573
rect 106737 4607 106795 4613
rect 106737 4573 106749 4607
rect 106783 4604 106795 4607
rect 107749 4607 107807 4613
rect 107749 4604 107761 4607
rect 106783 4576 107761 4604
rect 106783 4573 106795 4576
rect 106737 4567 106795 4573
rect 107749 4573 107761 4576
rect 107795 4573 107807 4607
rect 107749 4567 107807 4573
rect 107930 4564 107936 4616
rect 107988 4604 107994 4616
rect 108850 4604 108856 4616
rect 107988 4576 108856 4604
rect 107988 4564 107994 4576
rect 108850 4564 108856 4576
rect 108908 4564 108914 4616
rect 112438 4604 112444 4616
rect 112399 4576 112444 4604
rect 112438 4564 112444 4576
rect 112496 4564 112502 4616
rect 113560 4604 113588 4635
rect 113634 4632 113640 4684
rect 113692 4672 113698 4684
rect 118418 4672 118424 4684
rect 113692 4644 118424 4672
rect 113692 4632 113698 4644
rect 118418 4632 118424 4644
rect 118476 4632 118482 4684
rect 118697 4675 118755 4681
rect 118697 4641 118709 4675
rect 118743 4672 118755 4675
rect 119798 4672 119804 4684
rect 118743 4644 119804 4672
rect 118743 4641 118755 4644
rect 118697 4635 118755 4641
rect 119798 4632 119804 4644
rect 119856 4632 119862 4684
rect 120000 4681 120028 4712
rect 119985 4675 120043 4681
rect 119985 4641 119997 4675
rect 120031 4641 120043 4675
rect 119985 4635 120043 4641
rect 120077 4675 120135 4681
rect 120077 4641 120089 4675
rect 120123 4672 120135 4675
rect 120166 4672 120172 4684
rect 120123 4644 120172 4672
rect 120123 4641 120135 4644
rect 120077 4635 120135 4641
rect 120166 4632 120172 4644
rect 120224 4632 120230 4684
rect 120534 4632 120540 4684
rect 120592 4672 120598 4684
rect 123846 4672 123852 4684
rect 120592 4644 122880 4672
rect 123807 4644 123852 4672
rect 120592 4632 120598 4644
rect 114738 4604 114744 4616
rect 113560 4576 114744 4604
rect 114738 4564 114744 4576
rect 114796 4564 114802 4616
rect 114833 4607 114891 4613
rect 114833 4573 114845 4607
rect 114879 4604 114891 4607
rect 114922 4604 114928 4616
rect 114879 4576 114928 4604
rect 114879 4573 114891 4576
rect 114833 4567 114891 4573
rect 114922 4564 114928 4576
rect 114980 4564 114986 4616
rect 117130 4604 117136 4616
rect 117091 4576 117136 4604
rect 117130 4564 117136 4576
rect 117188 4564 117194 4616
rect 118513 4607 118571 4613
rect 118513 4573 118525 4607
rect 118559 4604 118571 4607
rect 119338 4604 119344 4616
rect 118559 4576 119344 4604
rect 118559 4573 118571 4576
rect 118513 4567 118571 4573
rect 119338 4564 119344 4576
rect 119396 4564 119402 4616
rect 122653 4607 122711 4613
rect 122653 4573 122665 4607
rect 122699 4573 122711 4607
rect 122852 4604 122880 4644
rect 123846 4632 123852 4644
rect 123904 4632 123910 4684
rect 125042 4672 125048 4684
rect 123956 4644 124260 4672
rect 125003 4644 125048 4672
rect 123956 4604 123984 4644
rect 124122 4604 124128 4616
rect 122852 4576 123984 4604
rect 124083 4576 124128 4604
rect 122653 4567 122711 4573
rect 91888 4508 93992 4536
rect 94056 4508 94268 4536
rect 91888 4496 91894 4508
rect 94056 4468 94084 4508
rect 85776 4440 94084 4468
rect 94240 4468 94268 4508
rect 94314 4496 94320 4548
rect 94372 4536 94378 4548
rect 96522 4536 96528 4548
rect 94372 4508 96528 4536
rect 94372 4496 94378 4508
rect 96522 4496 96528 4508
rect 96580 4496 96586 4548
rect 97261 4539 97319 4545
rect 97261 4505 97273 4539
rect 97307 4536 97319 4539
rect 106182 4536 106188 4548
rect 97307 4508 106188 4536
rect 97307 4505 97319 4508
rect 97261 4499 97319 4505
rect 106182 4496 106188 4508
rect 106240 4496 106246 4548
rect 106550 4536 106556 4548
rect 106292 4508 106556 4536
rect 102410 4468 102416 4480
rect 94240 4440 102416 4468
rect 102410 4428 102416 4440
rect 102468 4428 102474 4480
rect 102594 4428 102600 4480
rect 102652 4468 102658 4480
rect 104158 4468 104164 4480
rect 102652 4440 104164 4468
rect 102652 4428 102658 4440
rect 104158 4428 104164 4440
rect 104216 4428 104222 4480
rect 104342 4428 104348 4480
rect 104400 4468 104406 4480
rect 105173 4471 105231 4477
rect 105173 4468 105185 4471
rect 104400 4440 105185 4468
rect 104400 4428 104406 4440
rect 105173 4437 105185 4440
rect 105219 4437 105231 4471
rect 105173 4431 105231 4437
rect 105998 4428 106004 4480
rect 106056 4468 106062 4480
rect 106292 4468 106320 4508
rect 106550 4496 106556 4508
rect 106608 4496 106614 4548
rect 109221 4539 109279 4545
rect 109221 4505 109233 4539
rect 109267 4505 109279 4539
rect 109221 4499 109279 4505
rect 106056 4440 106320 4468
rect 106056 4428 106062 4440
rect 108022 4428 108028 4480
rect 108080 4468 108086 4480
rect 109126 4468 109132 4480
rect 108080 4440 109132 4468
rect 108080 4428 108086 4440
rect 109126 4428 109132 4440
rect 109184 4428 109190 4480
rect 109236 4468 109264 4499
rect 109310 4496 109316 4548
rect 109368 4536 109374 4548
rect 112254 4536 112260 4548
rect 109368 4508 112260 4536
rect 109368 4496 109374 4508
rect 112254 4496 112260 4508
rect 112312 4496 112318 4548
rect 113542 4496 113548 4548
rect 113600 4536 113606 4548
rect 113729 4539 113787 4545
rect 113729 4536 113741 4539
rect 113600 4508 113741 4536
rect 113600 4496 113606 4508
rect 113729 4505 113741 4508
rect 113775 4505 113787 4539
rect 119614 4536 119620 4548
rect 113729 4499 113787 4505
rect 114020 4508 119620 4536
rect 113818 4468 113824 4480
rect 109236 4440 113824 4468
rect 113818 4428 113824 4440
rect 113876 4428 113882 4480
rect 113910 4428 113916 4480
rect 113968 4468 113974 4480
rect 114020 4468 114048 4508
rect 119614 4496 119620 4508
rect 119672 4496 119678 4548
rect 121638 4536 121644 4548
rect 119724 4508 121644 4536
rect 113968 4440 114048 4468
rect 113968 4428 113974 4440
rect 114738 4428 114744 4480
rect 114796 4468 114802 4480
rect 116946 4468 116952 4480
rect 114796 4440 116952 4468
rect 114796 4428 114802 4440
rect 116946 4428 116952 4440
rect 117004 4428 117010 4480
rect 118326 4428 118332 4480
rect 118384 4468 118390 4480
rect 119724 4468 119752 4508
rect 121638 4496 121644 4508
rect 121696 4496 121702 4548
rect 122668 4536 122696 4567
rect 124122 4564 124128 4576
rect 124180 4564 124186 4616
rect 124232 4604 124260 4644
rect 125042 4632 125048 4644
rect 125100 4632 125106 4684
rect 126146 4672 126152 4684
rect 126107 4644 126152 4672
rect 126146 4632 126152 4644
rect 126204 4632 126210 4684
rect 126256 4672 126284 4712
rect 126330 4700 126336 4752
rect 126388 4740 126394 4752
rect 132696 4740 132724 4780
rect 137554 4768 137560 4780
rect 137612 4768 137618 4820
rect 137646 4768 137652 4820
rect 137704 4808 137710 4820
rect 138750 4808 138756 4820
rect 137704 4780 138612 4808
rect 138711 4780 138756 4808
rect 137704 4768 137710 4780
rect 138290 4740 138296 4752
rect 126388 4712 132724 4740
rect 134260 4712 138296 4740
rect 126388 4700 126394 4712
rect 127986 4672 127992 4684
rect 126256 4644 127992 4672
rect 127986 4632 127992 4644
rect 128044 4632 128050 4684
rect 129918 4672 129924 4684
rect 129879 4644 129924 4672
rect 129918 4632 129924 4644
rect 129976 4632 129982 4684
rect 130749 4675 130807 4681
rect 130749 4641 130761 4675
rect 130795 4672 130807 4675
rect 131666 4672 131672 4684
rect 130795 4644 131672 4672
rect 130795 4641 130807 4644
rect 130749 4635 130807 4641
rect 131666 4632 131672 4644
rect 131724 4632 131730 4684
rect 131761 4675 131819 4681
rect 131761 4641 131773 4675
rect 131807 4672 131819 4675
rect 133506 4672 133512 4684
rect 131807 4644 133512 4672
rect 131807 4641 131819 4644
rect 131761 4635 131819 4641
rect 133506 4632 133512 4644
rect 133564 4632 133570 4684
rect 133901 4675 133959 4681
rect 133901 4641 133913 4675
rect 133947 4672 133959 4675
rect 134260 4672 134288 4712
rect 138290 4700 138296 4712
rect 138348 4700 138354 4752
rect 138584 4740 138612 4780
rect 138750 4768 138756 4780
rect 138808 4768 138814 4820
rect 141050 4808 141056 4820
rect 139772 4780 141056 4808
rect 139670 4740 139676 4752
rect 138584 4712 139676 4740
rect 139670 4700 139676 4712
rect 139728 4700 139734 4752
rect 133947 4644 134288 4672
rect 133947 4641 133959 4644
rect 133901 4635 133959 4641
rect 134334 4632 134340 4684
rect 134392 4672 134398 4684
rect 134981 4675 135039 4681
rect 134981 4672 134993 4675
rect 134392 4644 134993 4672
rect 134392 4632 134398 4644
rect 134981 4641 134993 4644
rect 135027 4641 135039 4675
rect 136082 4672 136088 4684
rect 136043 4644 136088 4672
rect 134981 4635 135039 4641
rect 136082 4632 136088 4644
rect 136140 4632 136146 4684
rect 137204 4644 137508 4672
rect 124232 4576 126744 4604
rect 126330 4536 126336 4548
rect 122668 4508 126336 4536
rect 126330 4496 126336 4508
rect 126388 4496 126394 4548
rect 126514 4536 126520 4548
rect 126475 4508 126520 4536
rect 126514 4496 126520 4508
rect 126572 4496 126578 4548
rect 126716 4536 126744 4576
rect 126790 4564 126796 4616
rect 126848 4604 126854 4616
rect 128357 4607 128415 4613
rect 128357 4604 128369 4607
rect 126848 4576 128369 4604
rect 126848 4564 126854 4576
rect 128357 4573 128369 4576
rect 128403 4573 128415 4607
rect 128357 4567 128415 4573
rect 129829 4607 129887 4613
rect 129829 4573 129841 4607
rect 129875 4604 129887 4607
rect 131298 4604 131304 4616
rect 129875 4576 131304 4604
rect 129875 4573 129887 4576
rect 129829 4567 129887 4573
rect 131298 4564 131304 4576
rect 131356 4564 131362 4616
rect 137204 4604 137232 4644
rect 137370 4604 137376 4616
rect 131408 4576 137232 4604
rect 137331 4576 137376 4604
rect 126716 4508 126928 4536
rect 118384 4440 119752 4468
rect 119893 4471 119951 4477
rect 118384 4428 118390 4440
rect 119893 4437 119905 4471
rect 119939 4468 119951 4471
rect 123386 4468 123392 4480
rect 119939 4440 123392 4468
rect 119939 4437 119951 4440
rect 119893 4431 119951 4437
rect 123386 4428 123392 4440
rect 123444 4428 123450 4480
rect 125226 4428 125232 4480
rect 125284 4468 125290 4480
rect 126790 4468 126796 4480
rect 125284 4440 126796 4468
rect 125284 4428 125290 4440
rect 126790 4428 126796 4440
rect 126848 4428 126854 4480
rect 126900 4468 126928 4508
rect 127894 4496 127900 4548
rect 127952 4536 127958 4548
rect 131408 4536 131436 4576
rect 137370 4564 137376 4576
rect 137428 4564 137434 4616
rect 137480 4604 137508 4644
rect 137554 4632 137560 4684
rect 137612 4672 137618 4684
rect 139772 4672 139800 4780
rect 141050 4768 141056 4780
rect 141108 4768 141114 4820
rect 148318 4768 148324 4820
rect 148376 4808 148382 4820
rect 155494 4808 155500 4820
rect 148376 4780 155500 4808
rect 148376 4768 148382 4780
rect 155494 4768 155500 4780
rect 155552 4768 155558 4820
rect 144181 4743 144239 4749
rect 144181 4740 144193 4743
rect 140148 4712 144193 4740
rect 140148 4672 140176 4712
rect 144181 4709 144193 4712
rect 144227 4709 144239 4743
rect 144181 4703 144239 4709
rect 141602 4672 141608 4684
rect 137612 4644 139800 4672
rect 139872 4644 140176 4672
rect 141563 4644 141608 4672
rect 137612 4632 137618 4644
rect 139872 4604 139900 4644
rect 141602 4632 141608 4644
rect 141660 4632 141666 4684
rect 140038 4604 140044 4616
rect 137480 4576 139900 4604
rect 139999 4576 140044 4604
rect 140038 4564 140044 4576
rect 140096 4564 140102 4616
rect 142430 4604 142436 4616
rect 142391 4576 142436 4604
rect 142430 4564 142436 4576
rect 142488 4564 142494 4616
rect 144181 4607 144239 4613
rect 144181 4573 144193 4607
rect 144227 4604 144239 4607
rect 148318 4604 148324 4616
rect 144227 4576 148324 4604
rect 144227 4573 144239 4576
rect 144181 4567 144239 4573
rect 148318 4564 148324 4576
rect 148376 4564 148382 4616
rect 127952 4508 131436 4536
rect 127952 4496 127958 4508
rect 133506 4496 133512 4548
rect 133564 4536 133570 4548
rect 136358 4536 136364 4548
rect 133564 4508 136364 4536
rect 133564 4496 133570 4508
rect 136358 4496 136364 4508
rect 136416 4496 136422 4548
rect 136453 4539 136511 4545
rect 136453 4505 136465 4539
rect 136499 4505 136511 4539
rect 136453 4499 136511 4505
rect 128630 4468 128636 4480
rect 126900 4440 128636 4468
rect 128630 4428 128636 4440
rect 128688 4428 128694 4480
rect 132034 4428 132040 4480
rect 132092 4468 132098 4480
rect 133969 4471 134027 4477
rect 133969 4468 133981 4471
rect 132092 4440 133981 4468
rect 132092 4428 132098 4440
rect 133969 4437 133981 4440
rect 134015 4437 134027 4471
rect 133969 4431 134027 4437
rect 134702 4428 134708 4480
rect 134760 4468 134766 4480
rect 136174 4468 136180 4480
rect 134760 4440 136180 4468
rect 134760 4428 134766 4440
rect 136174 4428 136180 4440
rect 136232 4428 136238 4480
rect 136468 4468 136496 4499
rect 136634 4496 136640 4548
rect 136692 4536 136698 4548
rect 140682 4536 140688 4548
rect 136692 4508 140688 4536
rect 136692 4496 136698 4508
rect 140682 4496 140688 4508
rect 140740 4496 140746 4548
rect 141510 4536 141516 4548
rect 141471 4508 141516 4536
rect 141510 4496 141516 4508
rect 141568 4496 141574 4548
rect 137738 4468 137744 4480
rect 136468 4440 137744 4468
rect 137738 4428 137744 4440
rect 137796 4428 137802 4480
rect 137830 4428 137836 4480
rect 137888 4468 137894 4480
rect 145374 4468 145380 4480
rect 137888 4440 145380 4468
rect 137888 4428 137894 4440
rect 145374 4428 145380 4440
rect 145432 4428 145438 4480
rect 1104 4378 154560 4400
rect 1104 4326 4078 4378
rect 4130 4326 44078 4378
rect 44130 4326 84078 4378
rect 84130 4326 124078 4378
rect 124130 4326 154560 4378
rect 1104 4304 154560 4326
rect 56226 4224 56232 4276
rect 56284 4264 56290 4276
rect 75914 4264 75920 4276
rect 56284 4236 75920 4264
rect 56284 4224 56290 4236
rect 75914 4224 75920 4236
rect 75972 4224 75978 4276
rect 88886 4224 88892 4276
rect 88944 4264 88950 4276
rect 92106 4264 92112 4276
rect 88944 4236 92112 4264
rect 88944 4224 88950 4236
rect 92106 4224 92112 4236
rect 92164 4224 92170 4276
rect 94498 4224 94504 4276
rect 94556 4264 94562 4276
rect 100202 4264 100208 4276
rect 94556 4236 100208 4264
rect 94556 4224 94562 4236
rect 100202 4224 100208 4236
rect 100260 4224 100266 4276
rect 107654 4264 107660 4276
rect 102336 4236 107660 4264
rect 27985 4199 28043 4205
rect 27985 4165 27997 4199
rect 28031 4196 28043 4199
rect 30282 4196 30288 4208
rect 28031 4168 30288 4196
rect 28031 4165 28043 4168
rect 27985 4159 28043 4165
rect 30282 4156 30288 4168
rect 30340 4156 30346 4208
rect 32585 4199 32643 4205
rect 32585 4165 32597 4199
rect 32631 4196 32643 4199
rect 34330 4196 34336 4208
rect 32631 4168 34336 4196
rect 32631 4165 32643 4168
rect 32585 4159 32643 4165
rect 34330 4156 34336 4168
rect 34388 4156 34394 4208
rect 43717 4199 43775 4205
rect 43717 4165 43729 4199
rect 43763 4196 43775 4199
rect 45002 4196 45008 4208
rect 43763 4168 45008 4196
rect 43763 4165 43775 4168
rect 43717 4159 43775 4165
rect 45002 4156 45008 4168
rect 45060 4156 45066 4208
rect 53193 4199 53251 4205
rect 46308 4168 46612 4196
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 5353 4131 5411 4137
rect 4212 4100 5304 4128
rect 4212 4088 4218 4100
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4060 3295 4063
rect 3602 4060 3608 4072
rect 3283 4032 3608 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 5276 4069 5304 4100
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 5534 4128 5540 4140
rect 5399 4100 5540 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 8754 4128 8760 4140
rect 8715 4100 8760 4128
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9674 4128 9680 4140
rect 9635 4100 9680 4128
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 10870 4128 10876 4140
rect 10831 4100 10876 4128
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 20993 4131 21051 4137
rect 12492 4100 12537 4128
rect 12492 4088 12498 4100
rect 20993 4097 21005 4131
rect 21039 4097 21051 4131
rect 20993 4091 21051 4097
rect 22557 4131 22615 4137
rect 22557 4097 22569 4131
rect 22603 4128 22615 4131
rect 23474 4128 23480 4140
rect 22603 4100 23480 4128
rect 22603 4097 22615 4100
rect 22557 4091 22615 4097
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4029 5319 4063
rect 5261 4023 5319 4029
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4060 8907 4063
rect 9950 4060 9956 4072
rect 8895 4032 9956 4060
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 4264 3992 4292 4023
rect 3252 3964 4292 3992
rect 4341 3995 4399 4001
rect 3252 3936 3280 3964
rect 4341 3961 4353 3995
rect 4387 3992 4399 3995
rect 5626 3992 5632 4004
rect 4387 3964 5632 3992
rect 4387 3961 4399 3964
rect 4341 3955 4399 3961
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 7300 3992 7328 4023
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 11146 4060 11152 4072
rect 11107 4032 11152 4060
rect 11146 4020 11152 4032
rect 11204 4020 11210 4072
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 19794 4060 19800 4072
rect 19567 4032 19800 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 19794 4020 19800 4032
rect 19852 4020 19858 4072
rect 9674 3992 9680 4004
rect 7300 3964 9680 3992
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 11238 3952 11244 4004
rect 11296 3992 11302 4004
rect 13449 3995 13507 4001
rect 13449 3992 13461 3995
rect 11296 3964 13461 3992
rect 11296 3952 11302 3964
rect 13449 3961 13461 3964
rect 13495 3961 13507 3995
rect 13449 3955 13507 3961
rect 3234 3884 3240 3936
rect 3292 3884 3298 3936
rect 3329 3927 3387 3933
rect 3329 3893 3341 3927
rect 3375 3924 3387 3927
rect 6086 3924 6092 3936
rect 3375 3896 6092 3924
rect 3375 3893 3387 3896
rect 3329 3887 3387 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 21008 3924 21036 4091
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 25133 4131 25191 4137
rect 25133 4097 25145 4131
rect 25179 4128 25191 4131
rect 25222 4128 25228 4140
rect 25179 4100 25228 4128
rect 25179 4097 25191 4100
rect 25133 4091 25191 4097
rect 25222 4088 25228 4100
rect 25280 4088 25286 4140
rect 26513 4131 26571 4137
rect 26513 4097 26525 4131
rect 26559 4128 26571 4131
rect 26970 4128 26976 4140
rect 26559 4100 26976 4128
rect 26559 4097 26571 4100
rect 26513 4091 26571 4097
rect 26970 4088 26976 4100
rect 27028 4088 27034 4140
rect 29362 4088 29368 4140
rect 29420 4128 29426 4140
rect 29641 4131 29699 4137
rect 29641 4128 29653 4131
rect 29420 4100 29653 4128
rect 29420 4088 29426 4100
rect 29641 4097 29653 4100
rect 29687 4097 29699 4131
rect 29641 4091 29699 4097
rect 30742 4088 30748 4140
rect 30800 4128 30806 4140
rect 31113 4131 31171 4137
rect 31113 4128 31125 4131
rect 30800 4100 31125 4128
rect 30800 4088 30806 4100
rect 31113 4097 31125 4100
rect 31159 4097 31171 4131
rect 33502 4128 33508 4140
rect 33463 4100 33508 4128
rect 31113 4091 31171 4097
rect 33502 4088 33508 4100
rect 33560 4088 33566 4140
rect 40497 4131 40555 4137
rect 40497 4097 40509 4131
rect 40543 4128 40555 4131
rect 40770 4128 40776 4140
rect 40543 4100 40776 4128
rect 40543 4097 40555 4100
rect 40497 4091 40555 4097
rect 40770 4088 40776 4100
rect 40828 4088 40834 4140
rect 41966 4088 41972 4140
rect 42024 4128 42030 4140
rect 42245 4131 42303 4137
rect 42245 4128 42257 4131
rect 42024 4100 42257 4128
rect 42024 4088 42030 4100
rect 42245 4097 42257 4100
rect 42291 4097 42303 4131
rect 42245 4091 42303 4097
rect 44542 4088 44548 4140
rect 44600 4128 44606 4140
rect 46308 4128 46336 4168
rect 46474 4128 46480 4140
rect 44600 4100 46336 4128
rect 46435 4100 46480 4128
rect 44600 4088 44606 4100
rect 46474 4088 46480 4100
rect 46532 4088 46538 4140
rect 46584 4128 46612 4168
rect 53193 4165 53205 4199
rect 53239 4196 53251 4199
rect 55122 4196 55128 4208
rect 53239 4168 55128 4196
rect 53239 4165 53251 4168
rect 53193 4159 53251 4165
rect 55122 4156 55128 4168
rect 55180 4156 55186 4208
rect 60476 4168 60780 4196
rect 47397 4131 47455 4137
rect 47397 4128 47409 4131
rect 46584 4100 47409 4128
rect 47397 4097 47409 4100
rect 47443 4097 47455 4131
rect 47397 4091 47455 4097
rect 48593 4131 48651 4137
rect 48593 4097 48605 4131
rect 48639 4128 48651 4131
rect 48958 4128 48964 4140
rect 48639 4100 48964 4128
rect 48639 4097 48651 4100
rect 48593 4091 48651 4097
rect 48958 4088 48964 4100
rect 49016 4088 49022 4140
rect 51994 4088 52000 4140
rect 52052 4128 52058 4140
rect 52052 4100 56180 4128
rect 52052 4088 52058 4100
rect 21085 4063 21143 4069
rect 21085 4029 21097 4063
rect 21131 4060 21143 4063
rect 22738 4060 22744 4072
rect 21131 4032 22744 4060
rect 21131 4029 21143 4032
rect 21085 4023 21143 4029
rect 22738 4020 22744 4032
rect 22796 4020 22802 4072
rect 22830 4020 22836 4072
rect 22888 4060 22894 4072
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 22888 4032 23673 4060
rect 22888 4020 22894 4032
rect 23661 4029 23673 4032
rect 23707 4029 23719 4063
rect 24762 4060 24768 4072
rect 24723 4032 24768 4060
rect 23661 4023 23719 4029
rect 24762 4020 24768 4032
rect 24820 4020 24826 4072
rect 28077 4063 28135 4069
rect 28077 4029 28089 4063
rect 28123 4060 28135 4063
rect 30190 4060 30196 4072
rect 28123 4032 30196 4060
rect 28123 4029 28135 4032
rect 28077 4023 28135 4029
rect 30190 4020 30196 4032
rect 30248 4020 30254 4072
rect 32677 4063 32735 4069
rect 32677 4029 32689 4063
rect 32723 4060 32735 4063
rect 33410 4060 33416 4072
rect 32723 4032 33416 4060
rect 32723 4029 32735 4032
rect 32677 4023 32735 4029
rect 33410 4020 33416 4032
rect 33468 4020 33474 4072
rect 43346 4060 43352 4072
rect 43307 4032 43352 4060
rect 43346 4020 43352 4032
rect 43404 4020 43410 4072
rect 44726 4020 44732 4072
rect 44784 4060 44790 4072
rect 46385 4063 46443 4069
rect 46385 4060 46397 4063
rect 44784 4032 46397 4060
rect 44784 4020 44790 4032
rect 46385 4029 46397 4032
rect 46431 4029 46443 4063
rect 46385 4023 46443 4029
rect 50617 4063 50675 4069
rect 50617 4029 50629 4063
rect 50663 4060 50675 4063
rect 51721 4063 51779 4069
rect 51721 4060 51733 4063
rect 50663 4032 51733 4060
rect 50663 4029 50675 4032
rect 50617 4023 50675 4029
rect 51721 4029 51733 4032
rect 51767 4029 51779 4063
rect 52822 4060 52828 4072
rect 52783 4032 52828 4060
rect 51721 4023 51779 4029
rect 52822 4020 52828 4032
rect 52880 4020 52886 4072
rect 54113 4063 54171 4069
rect 54113 4060 54125 4063
rect 52932 4032 54125 4060
rect 48958 3952 48964 4004
rect 49016 3992 49022 4004
rect 52932 3992 52960 4032
rect 54113 4029 54125 4032
rect 54159 4029 54171 4063
rect 54113 4023 54171 4029
rect 55125 4063 55183 4069
rect 55125 4029 55137 4063
rect 55171 4029 55183 4063
rect 55125 4023 55183 4029
rect 55140 3992 55168 4023
rect 55214 4020 55220 4072
rect 55272 4060 55278 4072
rect 56152 4069 56180 4100
rect 58066 4088 58072 4140
rect 58124 4128 58130 4140
rect 59265 4131 59323 4137
rect 59265 4128 59277 4131
rect 58124 4100 59277 4128
rect 58124 4088 58130 4100
rect 59265 4097 59277 4100
rect 59311 4097 59323 4131
rect 60476 4128 60504 4168
rect 60642 4128 60648 4140
rect 59265 4091 59323 4097
rect 60292 4100 60504 4128
rect 60603 4100 60648 4128
rect 56137 4063 56195 4069
rect 55272 4032 55317 4060
rect 55272 4020 55278 4032
rect 56137 4029 56149 4063
rect 56183 4029 56195 4063
rect 58250 4060 58256 4072
rect 58211 4032 58256 4060
rect 56137 4023 56195 4029
rect 58250 4020 58256 4032
rect 58308 4020 58314 4072
rect 60292 4060 60320 4100
rect 60642 4088 60648 4100
rect 60700 4088 60706 4140
rect 60752 4128 60780 4168
rect 68830 4156 68836 4208
rect 68888 4196 68894 4208
rect 102336 4196 102364 4236
rect 107654 4224 107660 4236
rect 107712 4224 107718 4276
rect 109678 4224 109684 4276
rect 109736 4264 109742 4276
rect 118510 4264 118516 4276
rect 109736 4236 118516 4264
rect 109736 4224 109742 4236
rect 118510 4224 118516 4236
rect 118568 4224 118574 4276
rect 118602 4224 118608 4276
rect 118660 4264 118666 4276
rect 118878 4264 118884 4276
rect 118660 4236 118884 4264
rect 118660 4224 118666 4236
rect 118878 4224 118884 4236
rect 118936 4224 118942 4276
rect 119890 4264 119896 4276
rect 118988 4236 119896 4264
rect 68888 4168 102364 4196
rect 68888 4156 68894 4168
rect 102410 4156 102416 4208
rect 102468 4196 102474 4208
rect 108298 4196 108304 4208
rect 102468 4168 108304 4196
rect 102468 4156 102474 4168
rect 108298 4156 108304 4168
rect 108356 4156 108362 4208
rect 109126 4156 109132 4208
rect 109184 4196 109190 4208
rect 118988 4196 119016 4236
rect 119890 4224 119896 4236
rect 119948 4224 119954 4276
rect 119982 4224 119988 4276
rect 120040 4264 120046 4276
rect 122466 4264 122472 4276
rect 120040 4236 122472 4264
rect 120040 4224 120046 4236
rect 122466 4224 122472 4236
rect 122524 4224 122530 4276
rect 123478 4224 123484 4276
rect 123536 4264 123542 4276
rect 123573 4267 123631 4273
rect 123573 4264 123585 4267
rect 123536 4236 123585 4264
rect 123536 4224 123542 4236
rect 123573 4233 123585 4236
rect 123619 4233 123631 4267
rect 125045 4267 125103 4273
rect 125045 4264 125057 4267
rect 123573 4227 123631 4233
rect 123680 4236 125057 4264
rect 121917 4199 121975 4205
rect 109184 4168 119016 4196
rect 119080 4168 120672 4196
rect 109184 4156 109190 4168
rect 63678 4128 63684 4140
rect 60752 4100 63684 4128
rect 63678 4088 63684 4100
rect 63736 4088 63742 4140
rect 67542 4088 67548 4140
rect 67600 4128 67606 4140
rect 67600 4100 70164 4128
rect 67600 4088 67606 4100
rect 60458 4060 60464 4072
rect 58360 4032 60320 4060
rect 60419 4032 60464 4060
rect 49016 3964 52960 3992
rect 53116 3964 55168 3992
rect 56229 3995 56287 4001
rect 49016 3952 49022 3964
rect 26878 3924 26884 3936
rect 21008 3896 26884 3924
rect 26878 3884 26884 3896
rect 26936 3884 26942 3936
rect 44634 3884 44640 3936
rect 44692 3924 44698 3936
rect 44729 3927 44787 3933
rect 44729 3924 44741 3927
rect 44692 3896 44741 3924
rect 44692 3884 44698 3896
rect 44729 3893 44741 3896
rect 44775 3893 44787 3927
rect 44729 3887 44787 3893
rect 49418 3884 49424 3936
rect 49476 3924 49482 3936
rect 53116 3924 53144 3964
rect 56229 3961 56241 3995
rect 56275 3992 56287 3995
rect 58360 3992 58388 4032
rect 60458 4020 60464 4032
rect 60516 4020 60522 4072
rect 63310 4020 63316 4072
rect 63368 4060 63374 4072
rect 63405 4063 63463 4069
rect 63405 4060 63417 4063
rect 63368 4032 63417 4060
rect 63368 4020 63374 4032
rect 63405 4029 63417 4032
rect 63451 4029 63463 4063
rect 63405 4023 63463 4029
rect 67453 4063 67511 4069
rect 67453 4029 67465 4063
rect 67499 4060 67511 4063
rect 67726 4060 67732 4072
rect 67499 4032 67732 4060
rect 67499 4029 67511 4032
rect 67453 4023 67511 4029
rect 67726 4020 67732 4032
rect 67784 4020 67790 4072
rect 67910 4020 67916 4072
rect 67968 4060 67974 4072
rect 70136 4069 70164 4100
rect 70394 4088 70400 4140
rect 70452 4128 70458 4140
rect 71685 4131 71743 4137
rect 71685 4128 71697 4131
rect 70452 4100 71697 4128
rect 70452 4088 70458 4100
rect 71685 4097 71697 4100
rect 71731 4097 71743 4131
rect 71685 4091 71743 4097
rect 71774 4088 71780 4140
rect 71832 4128 71838 4140
rect 72697 4131 72755 4137
rect 72697 4128 72709 4131
rect 71832 4100 72709 4128
rect 71832 4088 71838 4100
rect 72697 4097 72709 4100
rect 72743 4097 72755 4131
rect 72697 4091 72755 4097
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75917 4131 75975 4137
rect 75917 4128 75929 4131
rect 73856 4100 75929 4128
rect 73856 4088 73862 4100
rect 75917 4097 75929 4100
rect 75963 4097 75975 4131
rect 75917 4091 75975 4097
rect 79502 4088 79508 4140
rect 79560 4128 79566 4140
rect 79781 4131 79839 4137
rect 79781 4128 79793 4131
rect 79560 4100 79793 4128
rect 79560 4088 79566 4100
rect 79781 4097 79793 4100
rect 79827 4097 79839 4131
rect 79781 4091 79839 4097
rect 80054 4088 80060 4140
rect 80112 4128 80118 4140
rect 80977 4131 81035 4137
rect 80977 4128 80989 4131
rect 80112 4100 80989 4128
rect 80112 4088 80118 4100
rect 80977 4097 80989 4100
rect 81023 4097 81035 4131
rect 80977 4091 81035 4097
rect 81618 4088 81624 4140
rect 81676 4128 81682 4140
rect 81989 4131 82047 4137
rect 81989 4128 82001 4131
rect 81676 4100 82001 4128
rect 81676 4088 81682 4100
rect 81989 4097 82001 4100
rect 82035 4097 82047 4131
rect 81989 4091 82047 4097
rect 82262 4088 82268 4140
rect 82320 4128 82326 4140
rect 84286 4128 84292 4140
rect 82320 4100 84292 4128
rect 82320 4088 82326 4100
rect 84286 4088 84292 4100
rect 84344 4088 84350 4140
rect 85393 4131 85451 4137
rect 85393 4097 85405 4131
rect 85439 4128 85451 4131
rect 85574 4128 85580 4140
rect 85439 4100 85580 4128
rect 85439 4097 85451 4100
rect 85393 4091 85451 4097
rect 85574 4088 85580 4100
rect 85632 4088 85638 4140
rect 86126 4088 86132 4140
rect 86184 4128 86190 4140
rect 86184 4100 89024 4128
rect 86184 4088 86190 4100
rect 68649 4063 68707 4069
rect 68649 4060 68661 4063
rect 67968 4032 68661 4060
rect 67968 4020 67974 4032
rect 68649 4029 68661 4032
rect 68695 4029 68707 4063
rect 68649 4023 68707 4029
rect 70121 4063 70179 4069
rect 70121 4029 70133 4063
rect 70167 4029 70179 4063
rect 70121 4023 70179 4029
rect 70489 4063 70547 4069
rect 70489 4029 70501 4063
rect 70535 4029 70547 4063
rect 70489 4023 70547 4029
rect 70857 4063 70915 4069
rect 70857 4029 70869 4063
rect 70903 4060 70915 4063
rect 70946 4060 70952 4072
rect 70903 4032 70952 4060
rect 70903 4029 70915 4032
rect 70857 4023 70915 4029
rect 56275 3964 58388 3992
rect 58437 3995 58495 4001
rect 56275 3961 56287 3964
rect 56229 3955 56287 3961
rect 58437 3961 58449 3995
rect 58483 3992 58495 3995
rect 58986 3992 58992 4004
rect 58483 3964 58992 3992
rect 58483 3961 58495 3964
rect 58437 3955 58495 3961
rect 58986 3952 58992 3964
rect 59044 3952 59050 4004
rect 59354 3952 59360 4004
rect 59412 3992 59418 4004
rect 61657 3995 61715 4001
rect 61657 3992 61669 3995
rect 59412 3964 61669 3992
rect 59412 3952 59418 3964
rect 61657 3961 61669 3964
rect 61703 3961 61715 3995
rect 61657 3955 61715 3961
rect 65518 3952 65524 4004
rect 65576 3992 65582 4004
rect 68557 3995 68615 4001
rect 68557 3992 68569 3995
rect 65576 3964 68569 3992
rect 65576 3952 65582 3964
rect 68557 3961 68569 3964
rect 68603 3961 68615 3995
rect 70504 3992 70532 4023
rect 70946 4020 70952 4032
rect 71004 4020 71010 4072
rect 72970 4020 72976 4072
rect 73028 4060 73034 4072
rect 74261 4063 74319 4069
rect 74261 4060 74273 4063
rect 73028 4032 74273 4060
rect 73028 4020 73034 4032
rect 74261 4029 74273 4032
rect 74307 4029 74319 4063
rect 76009 4063 76067 4069
rect 76009 4060 76021 4063
rect 74261 4023 74319 4029
rect 74368 4032 76021 4060
rect 72602 3992 72608 4004
rect 70504 3964 72608 3992
rect 68557 3955 68615 3961
rect 72602 3952 72608 3964
rect 72660 3952 72666 4004
rect 72878 3952 72884 4004
rect 72936 3992 72942 4004
rect 74169 3995 74227 4001
rect 74169 3992 74181 3995
rect 72936 3964 74181 3992
rect 72936 3952 72942 3964
rect 74169 3961 74181 3964
rect 74215 3961 74227 3995
rect 74169 3955 74227 3961
rect 49476 3896 53144 3924
rect 54205 3927 54263 3933
rect 49476 3884 49482 3896
rect 54205 3893 54217 3927
rect 54251 3924 54263 3927
rect 59630 3924 59636 3936
rect 54251 3896 59636 3924
rect 54251 3893 54263 3896
rect 54205 3887 54263 3893
rect 59630 3884 59636 3896
rect 59688 3884 59694 3936
rect 61194 3884 61200 3936
rect 61252 3924 61258 3936
rect 63589 3927 63647 3933
rect 63589 3924 63601 3927
rect 61252 3896 63601 3924
rect 61252 3884 61258 3896
rect 63589 3893 63601 3896
rect 63635 3893 63647 3927
rect 63589 3887 63647 3893
rect 71958 3884 71964 3936
rect 72016 3924 72022 3936
rect 74368 3924 74396 4032
rect 76009 4029 76021 4032
rect 76055 4029 76067 4063
rect 76009 4023 76067 4029
rect 78585 4063 78643 4069
rect 78585 4029 78597 4063
rect 78631 4060 78643 4063
rect 78766 4060 78772 4072
rect 78631 4032 78772 4060
rect 78631 4029 78643 4032
rect 78585 4023 78643 4029
rect 78766 4020 78772 4032
rect 78824 4020 78830 4072
rect 78861 4063 78919 4069
rect 78861 4029 78873 4063
rect 78907 4060 78919 4063
rect 80330 4060 80336 4072
rect 78907 4032 80336 4060
rect 78907 4029 78919 4032
rect 78861 4023 78919 4029
rect 80330 4020 80336 4032
rect 80388 4020 80394 4072
rect 80882 4020 80888 4072
rect 80940 4060 80946 4072
rect 83553 4063 83611 4069
rect 83553 4060 83565 4063
rect 80940 4032 83565 4060
rect 80940 4020 80946 4032
rect 83553 4029 83565 4032
rect 83599 4029 83611 4063
rect 83553 4023 83611 4029
rect 83826 4020 83832 4072
rect 83884 4060 83890 4072
rect 86034 4060 86040 4072
rect 83884 4032 86040 4060
rect 83884 4020 83890 4032
rect 86034 4020 86040 4032
rect 86092 4020 86098 4072
rect 86862 4020 86868 4072
rect 86920 4060 86926 4072
rect 87325 4063 87383 4069
rect 87325 4060 87337 4063
rect 86920 4032 87337 4060
rect 86920 4020 86926 4032
rect 87325 4029 87337 4032
rect 87371 4029 87383 4063
rect 87325 4023 87383 4029
rect 87417 4063 87475 4069
rect 87417 4029 87429 4063
rect 87463 4029 87475 4063
rect 87417 4023 87475 4029
rect 75914 3952 75920 4004
rect 75972 3992 75978 4004
rect 87230 3992 87236 4004
rect 75972 3964 87236 3992
rect 75972 3952 75978 3964
rect 87230 3952 87236 3964
rect 87288 3952 87294 4004
rect 72016 3896 74396 3924
rect 72016 3884 72022 3896
rect 77386 3884 77392 3936
rect 77444 3924 77450 3936
rect 83734 3924 83740 3936
rect 77444 3896 83740 3924
rect 77444 3884 77450 3896
rect 83734 3884 83740 3896
rect 83792 3884 83798 3936
rect 83826 3884 83832 3936
rect 83884 3924 83890 3936
rect 83921 3927 83979 3933
rect 83921 3924 83933 3927
rect 83884 3896 83933 3924
rect 83884 3884 83890 3896
rect 83921 3893 83933 3896
rect 83967 3893 83979 3927
rect 83921 3887 83979 3893
rect 84102 3884 84108 3936
rect 84160 3924 84166 3936
rect 87432 3924 87460 4023
rect 87782 4020 87788 4072
rect 87840 4060 87846 4072
rect 88996 4069 89024 4100
rect 90450 4088 90456 4140
rect 90508 4128 90514 4140
rect 91005 4131 91063 4137
rect 91005 4128 91017 4131
rect 90508 4100 91017 4128
rect 90508 4088 90514 4100
rect 91005 4097 91017 4100
rect 91051 4097 91063 4131
rect 91005 4091 91063 4097
rect 92566 4088 92572 4140
rect 92624 4128 92630 4140
rect 92624 4100 94452 4128
rect 92624 4088 92630 4100
rect 88889 4063 88947 4069
rect 88889 4060 88901 4063
rect 87840 4032 88901 4060
rect 87840 4020 87846 4032
rect 88889 4029 88901 4032
rect 88935 4029 88947 4063
rect 88889 4023 88947 4029
rect 88981 4063 89039 4069
rect 88981 4029 88993 4063
rect 89027 4029 89039 4063
rect 88981 4023 89039 4029
rect 91094 4020 91100 4072
rect 91152 4060 91158 4072
rect 92477 4063 92535 4069
rect 92477 4060 92489 4063
rect 91152 4032 92489 4060
rect 91152 4020 91158 4032
rect 92477 4029 92489 4032
rect 92523 4029 92535 4063
rect 92477 4023 92535 4029
rect 93394 4020 93400 4072
rect 93452 4060 93458 4072
rect 94314 4060 94320 4072
rect 93452 4032 94320 4060
rect 93452 4020 93458 4032
rect 94314 4020 94320 4032
rect 94372 4020 94378 4072
rect 94424 4060 94452 4100
rect 94774 4088 94780 4140
rect 94832 4128 94838 4140
rect 94961 4131 95019 4137
rect 94961 4128 94973 4131
rect 94832 4100 94973 4128
rect 94832 4088 94838 4100
rect 94961 4097 94973 4100
rect 95007 4097 95019 4131
rect 94961 4091 95019 4097
rect 95602 4088 95608 4140
rect 95660 4128 95666 4140
rect 99009 4131 99067 4137
rect 99009 4128 99021 4131
rect 95660 4100 99021 4128
rect 95660 4088 95666 4100
rect 99009 4097 99021 4100
rect 99055 4097 99067 4131
rect 99009 4091 99067 4097
rect 99190 4088 99196 4140
rect 99248 4128 99254 4140
rect 100110 4128 100116 4140
rect 99248 4100 100116 4128
rect 99248 4088 99254 4100
rect 100110 4088 100116 4100
rect 100168 4088 100174 4140
rect 102229 4131 102287 4137
rect 102229 4097 102241 4131
rect 102275 4128 102287 4131
rect 102502 4128 102508 4140
rect 102275 4100 102508 4128
rect 102275 4097 102287 4100
rect 102229 4091 102287 4097
rect 102502 4088 102508 4100
rect 102560 4088 102566 4140
rect 105538 4128 105544 4140
rect 105499 4100 105544 4128
rect 105538 4088 105544 4100
rect 105596 4088 105602 4140
rect 105722 4088 105728 4140
rect 105780 4128 105786 4140
rect 107841 4131 107899 4137
rect 107841 4128 107853 4131
rect 105780 4100 107853 4128
rect 105780 4088 105786 4100
rect 107841 4097 107853 4100
rect 107887 4097 107899 4131
rect 107841 4091 107899 4097
rect 109405 4131 109463 4137
rect 109405 4097 109417 4131
rect 109451 4128 109463 4131
rect 110690 4128 110696 4140
rect 109451 4100 110696 4128
rect 109451 4097 109463 4100
rect 109405 4091 109463 4097
rect 110690 4088 110696 4100
rect 110748 4088 110754 4140
rect 111981 4131 112039 4137
rect 111981 4097 111993 4131
rect 112027 4128 112039 4131
rect 112438 4128 112444 4140
rect 112027 4100 112444 4128
rect 112027 4097 112039 4100
rect 111981 4091 112039 4097
rect 112438 4088 112444 4100
rect 112496 4088 112502 4140
rect 115934 4128 115940 4140
rect 113376 4100 115940 4128
rect 96985 4063 97043 4069
rect 96985 4060 96997 4063
rect 94424 4032 96997 4060
rect 96985 4029 96997 4032
rect 97031 4029 97043 4063
rect 96985 4023 97043 4029
rect 98546 4020 98552 4072
rect 98604 4060 98610 4072
rect 99101 4063 99159 4069
rect 99101 4060 99113 4063
rect 98604 4032 99113 4060
rect 98604 4020 98610 4032
rect 99101 4029 99113 4032
rect 99147 4029 99159 4063
rect 100754 4060 100760 4072
rect 100715 4032 100760 4060
rect 99101 4023 99159 4029
rect 100754 4020 100760 4032
rect 100812 4020 100818 4072
rect 103333 4063 103391 4069
rect 103333 4029 103345 4063
rect 103379 4060 103391 4063
rect 104345 4063 104403 4069
rect 104345 4060 104357 4063
rect 103379 4032 104357 4060
rect 103379 4029 103391 4032
rect 103333 4023 103391 4029
rect 104345 4029 104357 4032
rect 104391 4029 104403 4063
rect 104345 4023 104403 4029
rect 105817 4063 105875 4069
rect 105817 4029 105829 4063
rect 105863 4029 105875 4063
rect 106734 4060 106740 4072
rect 106695 4032 106740 4060
rect 105817 4023 105875 4029
rect 90818 3952 90824 4004
rect 90876 3992 90882 4004
rect 92385 3995 92443 4001
rect 92385 3992 92397 3995
rect 90876 3964 92397 3992
rect 90876 3952 90882 3964
rect 92385 3961 92397 3964
rect 92431 3961 92443 3995
rect 92385 3955 92443 3961
rect 93762 3952 93768 4004
rect 93820 3992 93826 4004
rect 93949 3995 94007 4001
rect 93949 3992 93961 3995
rect 93820 3964 93961 3992
rect 93820 3952 93826 3964
rect 93949 3961 93961 3964
rect 93995 3961 94007 3995
rect 93949 3955 94007 3961
rect 94130 3952 94136 4004
rect 94188 3992 94194 4004
rect 96893 3995 96951 4001
rect 96893 3992 96905 3995
rect 94188 3964 96905 3992
rect 94188 3952 94194 3964
rect 96893 3961 96905 3964
rect 96939 3961 96951 3995
rect 96893 3955 96951 3961
rect 98638 3952 98644 4004
rect 98696 3992 98702 4004
rect 100573 3995 100631 4001
rect 100573 3992 100585 3995
rect 98696 3964 100585 3992
rect 98696 3952 98702 3964
rect 100573 3961 100585 3964
rect 100619 3961 100631 3995
rect 105832 3992 105860 4023
rect 106734 4020 106740 4032
rect 106792 4020 106798 4072
rect 107746 4020 107752 4072
rect 107804 4060 107810 4072
rect 107933 4063 107991 4069
rect 107933 4060 107945 4063
rect 107804 4032 107945 4060
rect 107804 4020 107810 4032
rect 107933 4029 107945 4032
rect 107979 4029 107991 4063
rect 110414 4060 110420 4072
rect 110375 4032 110420 4060
rect 107933 4023 107991 4029
rect 110414 4020 110420 4032
rect 110472 4020 110478 4072
rect 113376 3992 113404 4100
rect 115934 4088 115940 4100
rect 115992 4088 115998 4140
rect 116029 4131 116087 4137
rect 116029 4097 116041 4131
rect 116075 4097 116087 4131
rect 116029 4091 116087 4097
rect 113453 4063 113511 4069
rect 113453 4029 113465 4063
rect 113499 4060 113511 4063
rect 114465 4063 114523 4069
rect 114465 4060 114477 4063
rect 113499 4032 114477 4060
rect 113499 4029 113511 4032
rect 113453 4023 113511 4029
rect 114465 4029 114477 4032
rect 114511 4029 114523 4063
rect 114465 4023 114523 4029
rect 114557 4063 114615 4069
rect 114557 4029 114569 4063
rect 114603 4060 114615 4063
rect 114922 4060 114928 4072
rect 114603 4032 114928 4060
rect 114603 4029 114615 4032
rect 114557 4023 114615 4029
rect 114922 4020 114928 4032
rect 114980 4020 114986 4072
rect 115934 3992 115940 4004
rect 105832 3964 113404 3992
rect 115216 3964 115940 3992
rect 100573 3955 100631 3961
rect 84160 3896 87460 3924
rect 84160 3884 84166 3896
rect 92750 3884 92756 3936
rect 92808 3924 92814 3936
rect 94682 3924 94688 3936
rect 92808 3896 94688 3924
rect 92808 3884 92814 3896
rect 94682 3884 94688 3896
rect 94740 3884 94746 3936
rect 98914 3884 98920 3936
rect 98972 3924 98978 3936
rect 101490 3924 101496 3936
rect 98972 3896 101496 3924
rect 98972 3884 98978 3896
rect 101490 3884 101496 3896
rect 101548 3884 101554 3936
rect 102134 3884 102140 3936
rect 102192 3924 102198 3936
rect 113358 3924 113364 3936
rect 102192 3896 113364 3924
rect 102192 3884 102198 3896
rect 113358 3884 113364 3896
rect 113416 3884 113422 3936
rect 113450 3884 113456 3936
rect 113508 3924 113514 3936
rect 113545 3927 113603 3933
rect 113545 3924 113557 3927
rect 113508 3896 113557 3924
rect 113508 3884 113514 3896
rect 113545 3893 113557 3896
rect 113591 3893 113603 3927
rect 113545 3887 113603 3893
rect 114465 3927 114523 3933
rect 114465 3893 114477 3927
rect 114511 3924 114523 3927
rect 115216 3924 115244 3964
rect 115934 3952 115940 3964
rect 115992 3952 115998 4004
rect 116044 3992 116072 4091
rect 117130 4088 117136 4140
rect 117188 4128 117194 4140
rect 117961 4131 118019 4137
rect 117961 4128 117973 4131
rect 117188 4100 117973 4128
rect 117188 4088 117194 4100
rect 117961 4097 117973 4100
rect 118007 4097 118019 4131
rect 117961 4091 118019 4097
rect 118142 4088 118148 4140
rect 118200 4128 118206 4140
rect 119080 4128 119108 4168
rect 118200 4100 119108 4128
rect 120644 4128 120672 4168
rect 121917 4165 121929 4199
rect 121963 4196 121975 4199
rect 123110 4196 123116 4208
rect 121963 4168 123116 4196
rect 121963 4165 121975 4168
rect 121917 4159 121975 4165
rect 123110 4156 123116 4168
rect 123168 4156 123174 4208
rect 123294 4156 123300 4208
rect 123352 4196 123358 4208
rect 123680 4196 123708 4236
rect 125045 4233 125057 4236
rect 125091 4233 125103 4267
rect 125045 4227 125103 4233
rect 126514 4224 126520 4276
rect 126572 4264 126578 4276
rect 126572 4236 131068 4264
rect 126572 4224 126578 4236
rect 123352 4168 123708 4196
rect 124493 4199 124551 4205
rect 123352 4156 123358 4168
rect 124493 4165 124505 4199
rect 124539 4196 124551 4199
rect 126330 4196 126336 4208
rect 124539 4168 126336 4196
rect 124539 4165 124551 4168
rect 124493 4159 124551 4165
rect 126330 4156 126336 4168
rect 126388 4156 126394 4208
rect 126422 4156 126428 4208
rect 126480 4196 126486 4208
rect 126882 4196 126888 4208
rect 126480 4168 126888 4196
rect 126480 4156 126486 4168
rect 126882 4156 126888 4168
rect 126940 4156 126946 4208
rect 128446 4196 128452 4208
rect 128407 4168 128452 4196
rect 128446 4156 128452 4168
rect 128504 4156 128510 4208
rect 128630 4156 128636 4208
rect 128688 4196 128694 4208
rect 130378 4196 130384 4208
rect 128688 4168 130384 4196
rect 128688 4156 128694 4168
rect 130378 4156 130384 4168
rect 130436 4156 130442 4208
rect 131040 4196 131068 4236
rect 131114 4224 131120 4276
rect 131172 4264 131178 4276
rect 133966 4264 133972 4276
rect 131172 4236 133972 4264
rect 131172 4224 131178 4236
rect 133966 4224 133972 4236
rect 134024 4224 134030 4276
rect 135993 4267 136051 4273
rect 135993 4233 136005 4267
rect 136039 4264 136051 4267
rect 136082 4264 136088 4276
rect 136039 4236 136088 4264
rect 136039 4233 136051 4236
rect 135993 4227 136051 4233
rect 136082 4224 136088 4236
rect 136140 4224 136146 4276
rect 136542 4224 136548 4276
rect 136600 4264 136606 4276
rect 137830 4264 137836 4276
rect 136600 4236 137836 4264
rect 136600 4224 136606 4236
rect 137830 4224 137836 4236
rect 137888 4224 137894 4276
rect 145650 4264 145656 4276
rect 138032 4236 145656 4264
rect 131574 4196 131580 4208
rect 131040 4168 131580 4196
rect 131574 4156 131580 4168
rect 131632 4156 131638 4208
rect 131945 4199 132003 4205
rect 131945 4165 131957 4199
rect 131991 4196 132003 4199
rect 137186 4196 137192 4208
rect 131991 4168 137192 4196
rect 131991 4165 132003 4168
rect 131945 4159 132003 4165
rect 137186 4156 137192 4168
rect 137244 4156 137250 4208
rect 137278 4156 137284 4208
rect 137336 4196 137342 4208
rect 138032 4196 138060 4236
rect 145650 4224 145656 4236
rect 145708 4224 145714 4276
rect 137336 4168 138060 4196
rect 137336 4156 137342 4168
rect 138198 4156 138204 4208
rect 138256 4196 138262 4208
rect 139118 4196 139124 4208
rect 138256 4168 139124 4196
rect 138256 4156 138262 4168
rect 139118 4156 139124 4168
rect 139176 4156 139182 4208
rect 139964 4168 140544 4196
rect 121546 4128 121552 4140
rect 120644 4100 121552 4128
rect 118200 4088 118206 4100
rect 121546 4088 121552 4100
rect 121604 4088 121610 4140
rect 122006 4088 122012 4140
rect 122064 4128 122070 4140
rect 127437 4131 127495 4137
rect 122064 4100 127388 4128
rect 122064 4088 122070 4100
rect 116121 4063 116179 4069
rect 116121 4029 116133 4063
rect 116167 4060 116179 4063
rect 116670 4060 116676 4072
rect 116167 4032 116676 4060
rect 116167 4029 116179 4032
rect 116121 4023 116179 4029
rect 116670 4020 116676 4032
rect 116728 4020 116734 4072
rect 116949 4063 117007 4069
rect 116949 4029 116961 4063
rect 116995 4060 117007 4063
rect 119338 4060 119344 4072
rect 116995 4032 119344 4060
rect 116995 4029 117007 4032
rect 116949 4023 117007 4029
rect 119338 4020 119344 4032
rect 119396 4020 119402 4072
rect 119433 4063 119491 4069
rect 119433 4029 119445 4063
rect 119479 4060 119491 4063
rect 120445 4063 120503 4069
rect 120445 4060 120457 4063
rect 119479 4032 120457 4060
rect 119479 4029 119491 4032
rect 119433 4023 119491 4029
rect 120445 4029 120457 4032
rect 120491 4029 120503 4063
rect 120445 4023 120503 4029
rect 121917 4063 121975 4069
rect 121917 4029 121929 4063
rect 121963 4060 121975 4063
rect 123386 4060 123392 4072
rect 121963 4032 123392 4060
rect 121963 4029 121975 4032
rect 121917 4023 121975 4029
rect 123386 4020 123392 4032
rect 123444 4020 123450 4072
rect 123481 4063 123539 4069
rect 123481 4029 123493 4063
rect 123527 4060 123539 4063
rect 124493 4063 124551 4069
rect 124493 4060 124505 4063
rect 123527 4032 124505 4060
rect 123527 4029 123539 4032
rect 123481 4023 123539 4029
rect 124493 4029 124505 4032
rect 124539 4029 124551 4063
rect 124493 4023 124551 4029
rect 124953 4063 125011 4069
rect 124953 4029 124965 4063
rect 124999 4060 125011 4063
rect 125870 4060 125876 4072
rect 124999 4032 125876 4060
rect 124999 4029 125011 4032
rect 124953 4023 125011 4029
rect 125870 4020 125876 4032
rect 125928 4020 125934 4072
rect 125965 4063 126023 4069
rect 125965 4029 125977 4063
rect 126011 4029 126023 4063
rect 127158 4060 127164 4072
rect 127119 4032 127164 4060
rect 125965 4023 126023 4029
rect 125686 3992 125692 4004
rect 116044 3964 125692 3992
rect 125686 3952 125692 3964
rect 125744 3952 125750 4004
rect 125980 3992 126008 4023
rect 127158 4020 127164 4032
rect 127216 4020 127222 4072
rect 127360 4060 127388 4100
rect 127437 4097 127449 4131
rect 127483 4128 127495 4131
rect 131022 4128 131028 4140
rect 127483 4100 131028 4128
rect 127483 4097 127495 4100
rect 127437 4091 127495 4097
rect 131022 4088 131028 4100
rect 131080 4088 131086 4140
rect 132494 4128 132500 4140
rect 131868 4100 132500 4128
rect 128170 4060 128176 4072
rect 127360 4032 128176 4060
rect 128170 4020 128176 4032
rect 128228 4020 128234 4072
rect 128357 4063 128415 4069
rect 128357 4029 128369 4063
rect 128403 4060 128415 4063
rect 130381 4063 130439 4069
rect 130381 4060 130393 4063
rect 128403 4032 130393 4060
rect 128403 4029 128415 4032
rect 128357 4023 128415 4029
rect 130381 4029 130393 4032
rect 130427 4029 130439 4063
rect 130381 4023 130439 4029
rect 130473 4063 130531 4069
rect 130473 4029 130485 4063
rect 130519 4060 130531 4063
rect 131868 4060 131896 4100
rect 132494 4088 132500 4100
rect 132552 4088 132558 4140
rect 132865 4131 132923 4137
rect 132865 4097 132877 4131
rect 132911 4128 132923 4131
rect 133690 4128 133696 4140
rect 132911 4100 133696 4128
rect 132911 4097 132923 4100
rect 132865 4091 132923 4097
rect 133690 4088 133696 4100
rect 133748 4088 133754 4140
rect 134242 4128 134248 4140
rect 134203 4100 134248 4128
rect 134242 4088 134248 4100
rect 134300 4088 134306 4140
rect 135714 4128 135720 4140
rect 134352 4100 135720 4128
rect 132034 4060 132040 4072
rect 130519 4032 131896 4060
rect 131995 4032 132040 4060
rect 130519 4029 130531 4032
rect 130473 4023 130531 4029
rect 132034 4020 132040 4032
rect 132092 4020 132098 4072
rect 132402 4020 132408 4072
rect 132460 4060 132466 4072
rect 134352 4060 134380 4100
rect 135714 4088 135720 4100
rect 135772 4088 135778 4140
rect 136542 4128 136548 4140
rect 135824 4100 136548 4128
rect 132460 4032 134380 4060
rect 134429 4063 134487 4069
rect 132460 4020 132466 4032
rect 134429 4029 134441 4063
rect 134475 4060 134487 4063
rect 134610 4060 134616 4072
rect 134475 4032 134616 4060
rect 134475 4029 134487 4032
rect 134429 4023 134487 4029
rect 134610 4020 134616 4032
rect 134668 4020 134674 4072
rect 134978 4020 134984 4072
rect 135036 4060 135042 4072
rect 135824 4060 135852 4100
rect 136542 4088 136548 4100
rect 136600 4088 136606 4140
rect 136634 4088 136640 4140
rect 136692 4128 136698 4140
rect 139305 4131 139363 4137
rect 136692 4100 139164 4128
rect 136692 4088 136698 4100
rect 139136 4072 139164 4100
rect 139305 4097 139317 4131
rect 139351 4128 139363 4131
rect 139964 4128 139992 4168
rect 139351 4100 139992 4128
rect 139351 4097 139363 4100
rect 139305 4091 139363 4097
rect 140038 4088 140044 4140
rect 140096 4128 140102 4140
rect 140409 4131 140467 4137
rect 140409 4128 140421 4131
rect 140096 4100 140421 4128
rect 140096 4088 140102 4100
rect 140409 4097 140421 4100
rect 140455 4097 140467 4131
rect 140516 4128 140544 4168
rect 140590 4156 140596 4208
rect 140648 4196 140654 4208
rect 143534 4196 143540 4208
rect 140648 4168 143540 4196
rect 140648 4156 140654 4168
rect 143534 4156 143540 4168
rect 143592 4156 143598 4208
rect 140866 4128 140872 4140
rect 140516 4100 140872 4128
rect 140409 4091 140467 4097
rect 140866 4088 140872 4100
rect 140924 4088 140930 4140
rect 141510 4128 141516 4140
rect 141471 4100 141516 4128
rect 141510 4088 141516 4100
rect 141568 4088 141574 4140
rect 135036 4032 135852 4060
rect 135901 4063 135959 4069
rect 135036 4020 135042 4032
rect 135901 4029 135913 4063
rect 135947 4060 135959 4063
rect 136818 4060 136824 4072
rect 135947 4032 136824 4060
rect 135947 4029 135959 4032
rect 135901 4023 135959 4029
rect 136818 4020 136824 4032
rect 136876 4020 136882 4072
rect 136913 4063 136971 4069
rect 136913 4029 136925 4063
rect 136959 4060 136971 4063
rect 138017 4063 138075 4069
rect 138017 4060 138029 4063
rect 136959 4032 138029 4060
rect 136959 4029 136971 4032
rect 136913 4023 136971 4029
rect 138017 4029 138029 4032
rect 138063 4029 138075 4063
rect 138017 4023 138075 4029
rect 138106 4020 138112 4072
rect 138164 4060 138170 4072
rect 138164 4032 138796 4060
rect 138164 4020 138170 4032
rect 133690 3992 133696 4004
rect 125980 3964 128216 3992
rect 114511 3896 115244 3924
rect 114511 3893 114523 3896
rect 114465 3887 114523 3893
rect 115290 3884 115296 3936
rect 115348 3924 115354 3936
rect 117041 3927 117099 3933
rect 117041 3924 117053 3927
rect 115348 3896 117053 3924
rect 115348 3884 115354 3896
rect 117041 3893 117053 3896
rect 117087 3893 117099 3927
rect 117041 3887 117099 3893
rect 119522 3884 119528 3936
rect 119580 3924 119586 3936
rect 125962 3924 125968 3936
rect 119580 3896 125968 3924
rect 119580 3884 119586 3896
rect 125962 3884 125968 3896
rect 126020 3884 126026 3936
rect 128188 3924 128216 3964
rect 128556 3964 133696 3992
rect 128556 3924 128584 3964
rect 133690 3952 133696 3964
rect 133748 3952 133754 4004
rect 134242 3952 134248 4004
rect 134300 3992 134306 4004
rect 135438 3992 135444 4004
rect 134300 3964 135444 3992
rect 134300 3952 134306 3964
rect 135438 3952 135444 3964
rect 135496 3952 135502 4004
rect 136542 3952 136548 4004
rect 136600 3992 136606 4004
rect 136600 3964 137508 3992
rect 136600 3952 136606 3964
rect 128188 3896 128584 3924
rect 130381 3927 130439 3933
rect 130381 3893 130393 3927
rect 130427 3924 130439 3927
rect 131574 3924 131580 3936
rect 130427 3896 131580 3924
rect 130427 3893 130439 3896
rect 130381 3887 130439 3893
rect 131574 3884 131580 3896
rect 131632 3884 131638 3936
rect 131666 3884 131672 3936
rect 131724 3924 131730 3936
rect 134334 3924 134340 3936
rect 131724 3896 134340 3924
rect 131724 3884 131730 3896
rect 134334 3884 134340 3896
rect 134392 3884 134398 3936
rect 134702 3884 134708 3936
rect 134760 3924 134766 3936
rect 137370 3924 137376 3936
rect 134760 3896 137376 3924
rect 134760 3884 134766 3896
rect 137370 3884 137376 3896
rect 137428 3884 137434 3936
rect 137480 3924 137508 3964
rect 137738 3952 137744 4004
rect 137796 3992 137802 4004
rect 138658 3992 138664 4004
rect 137796 3964 138664 3992
rect 137796 3952 137802 3964
rect 138658 3952 138664 3964
rect 138716 3952 138722 4004
rect 138768 3992 138796 4032
rect 139118 4020 139124 4072
rect 139176 4020 139182 4072
rect 139210 4020 139216 4072
rect 139268 4060 139274 4072
rect 139268 4032 139313 4060
rect 139268 4020 139274 4032
rect 139394 4020 139400 4072
rect 139452 4060 139458 4072
rect 152366 4060 152372 4072
rect 139452 4032 152372 4060
rect 139452 4020 139458 4032
rect 152366 4020 152372 4032
rect 152424 4020 152430 4072
rect 142525 3995 142583 4001
rect 142525 3992 142537 3995
rect 138768 3964 142537 3992
rect 142525 3961 142537 3964
rect 142571 3961 142583 3995
rect 142525 3955 142583 3961
rect 138934 3924 138940 3936
rect 137480 3896 138940 3924
rect 138934 3884 138940 3896
rect 138992 3884 138998 3936
rect 140314 3884 140320 3936
rect 140372 3924 140378 3936
rect 151722 3924 151728 3936
rect 140372 3896 151728 3924
rect 140372 3884 140378 3896
rect 151722 3884 151728 3896
rect 151780 3884 151786 3936
rect 1104 3834 154560 3856
rect 1104 3782 24078 3834
rect 24130 3782 64078 3834
rect 64130 3782 104078 3834
rect 104130 3782 144078 3834
rect 144130 3782 154560 3834
rect 1104 3760 154560 3782
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 8294 3720 8300 3732
rect 7975 3692 8300 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 9674 3720 9680 3732
rect 9635 3692 9680 3720
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 18877 3723 18935 3729
rect 18877 3689 18889 3723
rect 18923 3720 18935 3723
rect 18966 3720 18972 3732
rect 18923 3692 18972 3720
rect 18923 3689 18935 3692
rect 18877 3683 18935 3689
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 19794 3720 19800 3732
rect 19755 3692 19800 3720
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 22830 3720 22836 3732
rect 22791 3692 22836 3720
rect 22830 3680 22836 3692
rect 22888 3680 22894 3732
rect 23842 3720 23848 3732
rect 23803 3692 23848 3720
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 24949 3723 25007 3729
rect 24949 3689 24961 3723
rect 24995 3720 25007 3723
rect 26050 3720 26056 3732
rect 24995 3692 26056 3720
rect 24995 3689 25007 3692
rect 24949 3683 25007 3689
rect 26050 3680 26056 3692
rect 26108 3680 26114 3732
rect 28258 3680 28264 3732
rect 28316 3720 28322 3732
rect 28353 3723 28411 3729
rect 28353 3720 28365 3723
rect 28316 3692 28365 3720
rect 28316 3680 28322 3692
rect 28353 3689 28365 3692
rect 28399 3689 28411 3723
rect 28353 3683 28411 3689
rect 37829 3723 37887 3729
rect 37829 3689 37841 3723
rect 37875 3720 37887 3723
rect 38286 3720 38292 3732
rect 37875 3692 38292 3720
rect 37875 3689 37887 3692
rect 37829 3683 37887 3689
rect 38286 3680 38292 3692
rect 38344 3680 38350 3732
rect 43438 3720 43444 3732
rect 43399 3692 43444 3720
rect 43438 3680 43444 3692
rect 43496 3680 43502 3732
rect 50893 3723 50951 3729
rect 50893 3689 50905 3723
rect 50939 3720 50951 3723
rect 52362 3720 52368 3732
rect 50939 3692 52368 3720
rect 50939 3689 50951 3692
rect 50893 3683 50951 3689
rect 52362 3680 52368 3692
rect 52420 3680 52426 3732
rect 53009 3723 53067 3729
rect 53009 3689 53021 3723
rect 53055 3720 53067 3723
rect 53098 3720 53104 3732
rect 53055 3692 53104 3720
rect 53055 3689 53067 3692
rect 53009 3683 53067 3689
rect 53098 3680 53104 3692
rect 53156 3680 53162 3732
rect 55582 3720 55588 3732
rect 55543 3692 55588 3720
rect 55582 3680 55588 3692
rect 55640 3680 55646 3732
rect 57149 3723 57207 3729
rect 57149 3689 57161 3723
rect 57195 3720 57207 3723
rect 57698 3720 57704 3732
rect 57195 3692 57704 3720
rect 57195 3689 57207 3692
rect 57149 3683 57207 3689
rect 57698 3680 57704 3692
rect 57756 3680 57762 3732
rect 58802 3680 58808 3732
rect 58860 3720 58866 3732
rect 59081 3723 59139 3729
rect 59081 3720 59093 3723
rect 58860 3692 59093 3720
rect 58860 3680 58866 3692
rect 59081 3689 59093 3692
rect 59127 3689 59139 3723
rect 59081 3683 59139 3689
rect 60185 3723 60243 3729
rect 60185 3689 60197 3723
rect 60231 3720 60243 3723
rect 60366 3720 60372 3732
rect 60231 3692 60372 3720
rect 60231 3689 60243 3692
rect 60185 3683 60243 3689
rect 60366 3680 60372 3692
rect 60424 3680 60430 3732
rect 68833 3723 68891 3729
rect 68833 3689 68845 3723
rect 68879 3720 68891 3723
rect 69014 3720 69020 3732
rect 68879 3692 69020 3720
rect 68879 3689 68891 3692
rect 68833 3683 68891 3689
rect 69014 3680 69020 3692
rect 69072 3680 69078 3732
rect 69845 3723 69903 3729
rect 69845 3689 69857 3723
rect 69891 3720 69903 3723
rect 71406 3720 71412 3732
rect 69891 3692 71412 3720
rect 69891 3689 69903 3692
rect 69845 3683 69903 3689
rect 71406 3680 71412 3692
rect 71464 3680 71470 3732
rect 73617 3723 73675 3729
rect 73617 3689 73629 3723
rect 73663 3720 73675 3723
rect 74166 3720 74172 3732
rect 73663 3692 74172 3720
rect 73663 3689 73675 3692
rect 73617 3683 73675 3689
rect 74166 3680 74172 3692
rect 74224 3680 74230 3732
rect 76650 3680 76656 3732
rect 76708 3720 76714 3732
rect 77021 3723 77079 3729
rect 77021 3720 77033 3723
rect 76708 3692 77033 3720
rect 76708 3680 76714 3692
rect 77021 3689 77033 3692
rect 77067 3689 77079 3723
rect 77021 3683 77079 3689
rect 83185 3723 83243 3729
rect 83185 3689 83197 3723
rect 83231 3720 83243 3723
rect 83274 3720 83280 3732
rect 83231 3692 83280 3720
rect 83231 3689 83243 3692
rect 83185 3683 83243 3689
rect 83274 3680 83280 3692
rect 83332 3680 83338 3732
rect 83734 3680 83740 3732
rect 83792 3720 83798 3732
rect 94498 3720 94504 3732
rect 83792 3692 94504 3720
rect 83792 3680 83798 3692
rect 94498 3680 94504 3692
rect 94556 3680 94562 3732
rect 95421 3723 95479 3729
rect 95421 3689 95433 3723
rect 95467 3720 95479 3723
rect 95786 3720 95792 3732
rect 95467 3692 95792 3720
rect 95467 3689 95479 3692
rect 95421 3683 95479 3689
rect 95786 3680 95792 3692
rect 95844 3680 95850 3732
rect 96154 3680 96160 3732
rect 96212 3720 96218 3732
rect 96212 3692 97948 3720
rect 96212 3680 96218 3692
rect 4617 3655 4675 3661
rect 4617 3621 4629 3655
rect 4663 3652 4675 3655
rect 17034 3652 17040 3664
rect 4663 3624 17040 3652
rect 4663 3621 4675 3624
rect 4617 3615 4675 3621
rect 17034 3612 17040 3624
rect 17092 3612 17098 3664
rect 27249 3655 27307 3661
rect 27249 3621 27261 3655
rect 27295 3652 27307 3655
rect 33042 3652 33048 3664
rect 27295 3624 33048 3652
rect 27295 3621 27307 3624
rect 27249 3615 27307 3621
rect 33042 3612 33048 3624
rect 33100 3612 33106 3664
rect 41417 3655 41475 3661
rect 41417 3621 41429 3655
rect 41463 3652 41475 3655
rect 47394 3652 47400 3664
rect 41463 3624 47400 3652
rect 41463 3621 41475 3624
rect 41417 3615 41475 3621
rect 47394 3612 47400 3624
rect 47452 3612 47458 3664
rect 51997 3655 52055 3661
rect 51997 3621 52009 3655
rect 52043 3652 52055 3655
rect 52086 3652 52092 3664
rect 52043 3624 52092 3652
rect 52043 3621 52055 3624
rect 51997 3615 52055 3621
rect 52086 3612 52092 3624
rect 52144 3612 52150 3664
rect 55214 3612 55220 3664
rect 55272 3652 55278 3664
rect 61286 3652 61292 3664
rect 55272 3624 61292 3652
rect 55272 3612 55278 3624
rect 61286 3612 61292 3624
rect 61344 3612 61350 3664
rect 73338 3612 73344 3664
rect 73396 3652 73402 3664
rect 74718 3652 74724 3664
rect 73396 3624 74724 3652
rect 73396 3612 73402 3624
rect 74718 3612 74724 3624
rect 74776 3612 74782 3664
rect 97626 3652 97632 3664
rect 74828 3624 97632 3652
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 2372 3556 4537 3584
rect 2372 3544 2378 3556
rect 4525 3553 4537 3556
rect 4571 3553 4583 3587
rect 4525 3547 4583 3553
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3553 5595 3587
rect 6549 3587 6607 3593
rect 6549 3584 6561 3587
rect 5537 3547 5595 3553
rect 5644 3556 6561 3584
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 5552 3516 5580 3547
rect 624 3488 5580 3516
rect 624 3476 630 3488
rect 2774 3408 2780 3460
rect 2832 3448 2838 3460
rect 5644 3448 5672 3556
rect 6549 3553 6561 3556
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3584 7895 3587
rect 8386 3584 8392 3596
rect 7883 3556 8392 3584
rect 7883 3553 7895 3556
rect 7837 3547 7895 3553
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 13906 3584 13912 3596
rect 12851 3556 13912 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 18046 3544 18052 3596
rect 18104 3584 18110 3596
rect 18785 3587 18843 3593
rect 18785 3584 18797 3587
rect 18104 3556 18797 3584
rect 18104 3544 18110 3556
rect 18785 3553 18797 3556
rect 18831 3553 18843 3587
rect 18785 3547 18843 3553
rect 24857 3587 24915 3593
rect 24857 3553 24869 3587
rect 24903 3584 24915 3587
rect 26326 3584 26332 3596
rect 24903 3556 26332 3584
rect 24903 3553 24915 3556
rect 24857 3547 24915 3553
rect 26326 3544 26332 3556
rect 26384 3544 26390 3596
rect 27154 3584 27160 3596
rect 27115 3556 27160 3584
rect 27154 3544 27160 3556
rect 27212 3544 27218 3596
rect 32493 3587 32551 3593
rect 32493 3553 32505 3587
rect 32539 3584 32551 3587
rect 33778 3584 33784 3596
rect 32539 3556 33784 3584
rect 32539 3553 32551 3556
rect 32493 3547 32551 3553
rect 33778 3544 33784 3556
rect 33836 3544 33842 3596
rect 34057 3587 34115 3593
rect 34057 3553 34069 3587
rect 34103 3584 34115 3587
rect 34514 3584 34520 3596
rect 34103 3556 34520 3584
rect 34103 3553 34115 3556
rect 34057 3547 34115 3553
rect 34514 3544 34520 3556
rect 34572 3544 34578 3596
rect 37642 3544 37648 3596
rect 37700 3584 37706 3596
rect 37737 3587 37795 3593
rect 37737 3584 37749 3587
rect 37700 3556 37749 3584
rect 37700 3544 37706 3556
rect 37737 3553 37749 3556
rect 37783 3553 37795 3587
rect 37737 3547 37795 3553
rect 39850 3544 39856 3596
rect 39908 3584 39914 3596
rect 41325 3587 41383 3593
rect 41325 3584 41337 3587
rect 39908 3556 41337 3584
rect 39908 3544 39914 3556
rect 41325 3553 41337 3556
rect 41371 3553 41383 3587
rect 41325 3547 41383 3553
rect 43349 3587 43407 3593
rect 43349 3553 43361 3587
rect 43395 3553 43407 3587
rect 44634 3584 44640 3596
rect 44595 3556 44640 3584
rect 43349 3547 43407 3553
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3516 6699 3519
rect 11606 3516 11612 3528
rect 6687 3488 11612 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 12710 3516 12716 3528
rect 12671 3488 12716 3516
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 33962 3516 33968 3528
rect 33923 3488 33968 3516
rect 33962 3476 33968 3488
rect 34020 3476 34026 3528
rect 41230 3476 41236 3528
rect 41288 3516 41294 3528
rect 43364 3516 43392 3547
rect 44634 3544 44640 3556
rect 44692 3544 44698 3596
rect 46198 3584 46204 3596
rect 46159 3556 46204 3584
rect 46198 3544 46204 3556
rect 46256 3544 46262 3596
rect 46750 3544 46756 3596
rect 46808 3584 46814 3596
rect 51905 3587 51963 3593
rect 51905 3584 51917 3587
rect 46808 3556 51917 3584
rect 46808 3544 46814 3556
rect 51905 3553 51917 3556
rect 51951 3553 51963 3587
rect 51905 3547 51963 3553
rect 52917 3587 52975 3593
rect 52917 3553 52929 3587
rect 52963 3553 52975 3587
rect 52917 3547 52975 3553
rect 45646 3516 45652 3528
rect 41288 3488 43392 3516
rect 45607 3488 45652 3516
rect 41288 3476 41294 3488
rect 45646 3476 45652 3488
rect 45704 3476 45710 3528
rect 47394 3476 47400 3528
rect 47452 3516 47458 3528
rect 52932 3516 52960 3547
rect 53282 3544 53288 3596
rect 53340 3584 53346 3596
rect 55493 3587 55551 3593
rect 55493 3584 55505 3587
rect 53340 3556 55505 3584
rect 53340 3544 53346 3556
rect 55493 3553 55505 3556
rect 55539 3553 55551 3587
rect 61562 3584 61568 3596
rect 61523 3556 61568 3584
rect 55493 3547 55551 3553
rect 61562 3544 61568 3556
rect 61620 3544 61626 3596
rect 66530 3584 66536 3596
rect 66491 3556 66536 3584
rect 66530 3544 66536 3556
rect 66588 3544 66594 3596
rect 72697 3587 72755 3593
rect 72697 3553 72709 3587
rect 72743 3584 72755 3587
rect 72786 3584 72792 3596
rect 72743 3556 72792 3584
rect 72743 3553 72755 3556
rect 72697 3547 72755 3553
rect 72786 3544 72792 3556
rect 72844 3544 72850 3596
rect 74258 3544 74264 3596
rect 74316 3584 74322 3596
rect 74626 3584 74632 3596
rect 74316 3556 74632 3584
rect 74316 3544 74322 3556
rect 74626 3544 74632 3556
rect 74684 3544 74690 3596
rect 47452 3488 52960 3516
rect 47452 3476 47458 3488
rect 60734 3476 60740 3528
rect 60792 3516 60798 3528
rect 61473 3519 61531 3525
rect 61473 3516 61485 3519
rect 60792 3488 61485 3516
rect 60792 3476 60798 3488
rect 61473 3485 61485 3488
rect 61519 3485 61531 3519
rect 61473 3479 61531 3485
rect 66625 3519 66683 3525
rect 66625 3485 66637 3519
rect 66671 3516 66683 3519
rect 67266 3516 67272 3528
rect 66671 3488 67272 3516
rect 66671 3485 66683 3488
rect 66625 3479 66683 3485
rect 67266 3476 67272 3488
rect 67324 3476 67330 3528
rect 72510 3476 72516 3528
rect 72568 3516 72574 3528
rect 74828 3516 74856 3624
rect 97626 3612 97632 3624
rect 97684 3612 97690 3664
rect 74902 3544 74908 3596
rect 74960 3584 74966 3596
rect 75457 3587 75515 3593
rect 75457 3584 75469 3587
rect 74960 3556 75469 3584
rect 74960 3544 74966 3556
rect 75457 3553 75469 3556
rect 75503 3553 75515 3587
rect 75457 3547 75515 3553
rect 75546 3544 75552 3596
rect 75604 3584 75610 3596
rect 77018 3584 77024 3596
rect 75604 3556 77024 3584
rect 75604 3544 75610 3556
rect 77018 3544 77024 3556
rect 77076 3544 77082 3596
rect 79318 3584 79324 3596
rect 77312 3556 78812 3584
rect 79279 3556 79324 3584
rect 72568 3488 74856 3516
rect 72568 3476 72574 3488
rect 75086 3476 75092 3528
rect 75144 3516 75150 3528
rect 75365 3519 75423 3525
rect 75365 3516 75377 3519
rect 75144 3488 75377 3516
rect 75144 3476 75150 3488
rect 75365 3485 75377 3488
rect 75411 3485 75423 3519
rect 75365 3479 75423 3485
rect 75822 3476 75828 3528
rect 75880 3516 75886 3528
rect 77312 3516 77340 3556
rect 75880 3488 77340 3516
rect 75880 3476 75886 3488
rect 77386 3476 77392 3528
rect 77444 3516 77450 3528
rect 78677 3519 78735 3525
rect 78677 3516 78689 3519
rect 77444 3488 78689 3516
rect 77444 3476 77450 3488
rect 78677 3485 78689 3488
rect 78723 3485 78735 3519
rect 78784 3516 78812 3556
rect 79318 3544 79324 3556
rect 79376 3544 79382 3596
rect 80238 3544 80244 3596
rect 80296 3584 80302 3596
rect 80333 3587 80391 3593
rect 80333 3584 80345 3587
rect 80296 3556 80345 3584
rect 80296 3544 80302 3556
rect 80333 3553 80345 3556
rect 80379 3553 80391 3587
rect 80333 3547 80391 3553
rect 82078 3544 82084 3596
rect 82136 3584 82142 3596
rect 83918 3584 83924 3596
rect 82136 3556 83924 3584
rect 82136 3544 82142 3556
rect 83918 3544 83924 3556
rect 83976 3544 83982 3596
rect 84286 3584 84292 3596
rect 84247 3556 84292 3584
rect 84286 3544 84292 3556
rect 84344 3544 84350 3596
rect 85853 3587 85911 3593
rect 85853 3553 85865 3587
rect 85899 3553 85911 3587
rect 85853 3547 85911 3553
rect 80882 3516 80888 3528
rect 78784 3488 80888 3516
rect 78677 3479 78735 3485
rect 80882 3476 80888 3488
rect 80940 3476 80946 3528
rect 80977 3519 81035 3525
rect 80977 3485 80989 3519
rect 81023 3516 81035 3519
rect 81158 3516 81164 3528
rect 81023 3488 81164 3516
rect 81023 3485 81035 3488
rect 80977 3479 81035 3485
rect 81158 3476 81164 3488
rect 81216 3476 81222 3528
rect 83182 3476 83188 3528
rect 83240 3516 83246 3528
rect 85868 3516 85896 3547
rect 86034 3544 86040 3596
rect 86092 3584 86098 3596
rect 89073 3587 89131 3593
rect 89073 3584 89085 3587
rect 86092 3556 89085 3584
rect 86092 3544 86098 3556
rect 89073 3553 89085 3556
rect 89119 3553 89131 3587
rect 89073 3547 89131 3553
rect 89346 3544 89352 3596
rect 89404 3584 89410 3596
rect 91557 3587 91615 3593
rect 91557 3584 91569 3587
rect 89404 3556 91569 3584
rect 89404 3544 89410 3556
rect 91557 3553 91569 3556
rect 91603 3553 91615 3587
rect 91557 3547 91615 3553
rect 91646 3544 91652 3596
rect 91704 3584 91710 3596
rect 93026 3584 93032 3596
rect 91704 3556 93032 3584
rect 91704 3544 91710 3556
rect 93026 3544 93032 3556
rect 93084 3544 93090 3596
rect 93949 3587 94007 3593
rect 93949 3553 93961 3587
rect 93995 3553 94007 3587
rect 93949 3547 94007 3553
rect 83240 3488 85896 3516
rect 83240 3476 83246 3488
rect 88150 3476 88156 3528
rect 88208 3516 88214 3528
rect 88981 3519 89039 3525
rect 88981 3516 88993 3519
rect 88208 3488 88993 3516
rect 88208 3476 88214 3488
rect 88981 3485 88993 3488
rect 89027 3485 89039 3519
rect 88981 3479 89039 3485
rect 91278 3476 91284 3528
rect 91336 3516 91342 3528
rect 91465 3519 91523 3525
rect 91465 3516 91477 3519
rect 91336 3488 91477 3516
rect 91336 3476 91342 3488
rect 91465 3485 91477 3488
rect 91511 3485 91523 3519
rect 91465 3479 91523 3485
rect 11790 3448 11796 3460
rect 2832 3420 5672 3448
rect 6564 3420 11796 3448
rect 2832 3408 2838 3420
rect 5629 3383 5687 3389
rect 5629 3349 5641 3383
rect 5675 3380 5687 3383
rect 6564 3380 6592 3420
rect 11790 3408 11796 3420
rect 11848 3408 11854 3460
rect 26510 3408 26516 3460
rect 26568 3448 26574 3460
rect 29086 3448 29092 3460
rect 26568 3420 29092 3448
rect 26568 3408 26574 3420
rect 29086 3408 29092 3420
rect 29144 3408 29150 3460
rect 34606 3408 34612 3460
rect 34664 3448 34670 3460
rect 41414 3448 41420 3460
rect 34664 3420 41420 3448
rect 34664 3408 34670 3420
rect 41414 3408 41420 3420
rect 41472 3408 41478 3460
rect 59262 3408 59268 3460
rect 59320 3448 59326 3460
rect 92474 3448 92480 3460
rect 59320 3420 92480 3448
rect 59320 3408 59326 3420
rect 92474 3408 92480 3420
rect 92532 3408 92538 3460
rect 5675 3352 6592 3380
rect 5675 3349 5687 3352
rect 5629 3343 5687 3349
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 45186 3380 45192 3392
rect 40736 3352 45192 3380
rect 40736 3340 40742 3352
rect 45186 3340 45192 3352
rect 45244 3340 45250 3392
rect 53926 3340 53932 3392
rect 53984 3380 53990 3392
rect 57238 3380 57244 3392
rect 53984 3352 57244 3380
rect 53984 3340 53990 3352
rect 57238 3340 57244 3352
rect 57296 3340 57302 3392
rect 72510 3380 72516 3392
rect 72471 3352 72516 3380
rect 72510 3340 72516 3352
rect 72568 3340 72574 3392
rect 84286 3340 84292 3392
rect 84344 3380 84350 3392
rect 84473 3383 84531 3389
rect 84473 3380 84485 3383
rect 84344 3352 84485 3380
rect 84344 3340 84350 3352
rect 84473 3349 84485 3352
rect 84519 3349 84531 3383
rect 86034 3380 86040 3392
rect 85995 3352 86040 3380
rect 84473 3343 84531 3349
rect 86034 3340 86040 3352
rect 86092 3340 86098 3392
rect 91002 3340 91008 3392
rect 91060 3380 91066 3392
rect 93964 3380 93992 3547
rect 94958 3544 94964 3596
rect 95016 3584 95022 3596
rect 96433 3587 96491 3593
rect 96433 3584 96445 3587
rect 95016 3556 96445 3584
rect 95016 3544 95022 3556
rect 96433 3553 96445 3556
rect 96479 3553 96491 3587
rect 97718 3584 97724 3596
rect 97679 3556 97724 3584
rect 96433 3547 96491 3553
rect 97718 3544 97724 3556
rect 97776 3544 97782 3596
rect 97920 3584 97948 3692
rect 99006 3680 99012 3732
rect 99064 3720 99070 3732
rect 101033 3723 101091 3729
rect 101033 3720 101045 3723
rect 99064 3692 101045 3720
rect 99064 3680 99070 3692
rect 101033 3689 101045 3692
rect 101079 3689 101091 3723
rect 103054 3720 103060 3732
rect 103015 3692 103060 3720
rect 101033 3683 101091 3689
rect 103054 3680 103060 3692
rect 103112 3680 103118 3732
rect 104894 3680 104900 3732
rect 104952 3720 104958 3732
rect 104952 3692 109816 3720
rect 104952 3680 104958 3692
rect 105170 3612 105176 3664
rect 105228 3652 105234 3664
rect 106737 3655 106795 3661
rect 106737 3652 106749 3655
rect 105228 3624 106749 3652
rect 105228 3612 105234 3624
rect 106737 3621 106749 3624
rect 106783 3621 106795 3655
rect 108206 3652 108212 3664
rect 106737 3615 106795 3621
rect 106844 3624 108212 3652
rect 99561 3587 99619 3593
rect 99561 3584 99573 3587
rect 97920 3556 99573 3584
rect 99561 3553 99573 3556
rect 99607 3553 99619 3587
rect 99561 3547 99619 3553
rect 99742 3544 99748 3596
rect 99800 3584 99806 3596
rect 102045 3587 102103 3593
rect 102045 3584 102057 3587
rect 99800 3556 102057 3584
rect 99800 3544 99806 3556
rect 102045 3553 102057 3556
rect 102091 3553 102103 3587
rect 102045 3547 102103 3553
rect 105817 3587 105875 3593
rect 105817 3553 105829 3587
rect 105863 3584 105875 3587
rect 106844 3584 106872 3624
rect 108206 3612 108212 3624
rect 108264 3612 108270 3664
rect 107286 3584 107292 3596
rect 105863 3556 106872 3584
rect 107247 3556 107292 3584
rect 105863 3553 105875 3556
rect 105817 3547 105875 3553
rect 107286 3544 107292 3556
rect 107344 3544 107350 3596
rect 108945 3587 109003 3593
rect 108945 3553 108957 3587
rect 108991 3584 109003 3587
rect 109034 3584 109040 3596
rect 108991 3556 109040 3584
rect 108991 3553 109003 3556
rect 108945 3547 109003 3553
rect 109034 3544 109040 3556
rect 109092 3544 109098 3596
rect 97350 3476 97356 3528
rect 97408 3516 97414 3528
rect 99469 3519 99527 3525
rect 99469 3516 99481 3519
rect 97408 3488 99481 3516
rect 97408 3476 97414 3488
rect 99469 3485 99481 3488
rect 99515 3485 99527 3519
rect 99469 3479 99527 3485
rect 103422 3476 103428 3528
rect 103480 3516 103486 3528
rect 105173 3519 105231 3525
rect 105173 3516 105185 3519
rect 103480 3488 105185 3516
rect 103480 3476 103486 3488
rect 105173 3485 105185 3488
rect 105219 3485 105231 3519
rect 105173 3479 105231 3485
rect 105998 3476 106004 3528
rect 106056 3516 106062 3528
rect 108301 3519 108359 3525
rect 108301 3516 108313 3519
rect 106056 3488 108313 3516
rect 106056 3476 106062 3488
rect 108301 3485 108313 3488
rect 108347 3485 108359 3519
rect 108301 3479 108359 3485
rect 94498 3408 94504 3460
rect 94556 3448 94562 3460
rect 94556 3420 102548 3448
rect 94556 3408 94562 3420
rect 91060 3352 93992 3380
rect 94317 3383 94375 3389
rect 91060 3340 91066 3352
rect 94317 3349 94329 3383
rect 94363 3380 94375 3383
rect 97718 3380 97724 3392
rect 94363 3352 97724 3380
rect 94363 3349 94375 3352
rect 94317 3343 94375 3349
rect 97718 3340 97724 3352
rect 97776 3340 97782 3392
rect 97997 3383 98055 3389
rect 97997 3349 98009 3383
rect 98043 3380 98055 3383
rect 101674 3380 101680 3392
rect 98043 3352 101680 3380
rect 98043 3349 98055 3352
rect 97997 3343 98055 3349
rect 101674 3340 101680 3352
rect 101732 3340 101738 3392
rect 102520 3380 102548 3420
rect 104158 3408 104164 3460
rect 104216 3448 104222 3460
rect 109218 3448 109224 3460
rect 104216 3420 109224 3448
rect 104216 3408 104222 3420
rect 109218 3408 109224 3420
rect 109276 3408 109282 3460
rect 105722 3380 105728 3392
rect 102520 3352 105728 3380
rect 105722 3340 105728 3352
rect 105780 3340 105786 3392
rect 106550 3340 106556 3392
rect 106608 3380 106614 3392
rect 107102 3380 107108 3392
rect 106608 3352 107108 3380
rect 106608 3340 106614 3352
rect 107102 3340 107108 3352
rect 107160 3340 107166 3392
rect 109788 3380 109816 3692
rect 110506 3680 110512 3732
rect 110564 3720 110570 3732
rect 113821 3723 113879 3729
rect 113821 3720 113833 3723
rect 110564 3692 113833 3720
rect 110564 3680 110570 3692
rect 113821 3689 113833 3692
rect 113867 3689 113879 3723
rect 115198 3720 115204 3732
rect 115159 3692 115204 3720
rect 113821 3683 113879 3689
rect 115198 3680 115204 3692
rect 115256 3680 115262 3732
rect 115382 3680 115388 3732
rect 115440 3720 115446 3732
rect 117133 3723 117191 3729
rect 117133 3720 117145 3723
rect 115440 3692 117145 3720
rect 115440 3680 115446 3692
rect 117133 3689 117145 3692
rect 117179 3689 117191 3723
rect 117133 3683 117191 3689
rect 117222 3680 117228 3732
rect 117280 3720 117286 3732
rect 119341 3723 119399 3729
rect 119341 3720 119353 3723
rect 117280 3692 119353 3720
rect 117280 3680 117286 3692
rect 119341 3689 119353 3692
rect 119387 3689 119399 3723
rect 122190 3720 122196 3732
rect 122151 3692 122196 3720
rect 119341 3683 119399 3689
rect 122190 3680 122196 3692
rect 122248 3680 122254 3732
rect 122300 3692 128216 3720
rect 111705 3655 111763 3661
rect 111705 3621 111717 3655
rect 111751 3652 111763 3655
rect 111794 3652 111800 3664
rect 111751 3624 111800 3652
rect 111751 3621 111763 3624
rect 111705 3615 111763 3621
rect 111794 3612 111800 3624
rect 111852 3612 111858 3664
rect 121917 3655 121975 3661
rect 121917 3652 121929 3655
rect 112640 3624 116992 3652
rect 110693 3587 110751 3593
rect 110693 3553 110705 3587
rect 110739 3584 110751 3587
rect 112640 3584 112668 3624
rect 110739 3556 112668 3584
rect 112709 3587 112767 3593
rect 110739 3553 110751 3556
rect 110693 3547 110751 3553
rect 112709 3553 112721 3587
rect 112755 3553 112767 3587
rect 112709 3547 112767 3553
rect 113729 3587 113787 3593
rect 113729 3553 113741 3587
rect 113775 3584 113787 3587
rect 116854 3584 116860 3596
rect 113775 3556 116860 3584
rect 113775 3553 113787 3556
rect 113729 3547 113787 3553
rect 109862 3476 109868 3528
rect 109920 3516 109926 3528
rect 110785 3519 110843 3525
rect 110785 3516 110797 3519
rect 109920 3488 110797 3516
rect 109920 3476 109926 3488
rect 110785 3485 110797 3488
rect 110831 3485 110843 3519
rect 110785 3479 110843 3485
rect 112732 3448 112760 3547
rect 116854 3544 116860 3556
rect 116912 3544 116918 3596
rect 112806 3476 112812 3528
rect 112864 3516 112870 3528
rect 112864 3488 112909 3516
rect 112864 3476 112870 3488
rect 113358 3476 113364 3528
rect 113416 3516 113422 3528
rect 116578 3516 116584 3528
rect 113416 3488 116584 3516
rect 113416 3476 113422 3488
rect 116578 3476 116584 3488
rect 116636 3476 116642 3528
rect 116964 3516 116992 3624
rect 120184 3624 121929 3652
rect 117041 3587 117099 3593
rect 117041 3553 117053 3587
rect 117087 3584 117099 3587
rect 117958 3584 117964 3596
rect 117087 3556 117964 3584
rect 117087 3553 117099 3556
rect 117041 3547 117099 3553
rect 117958 3544 117964 3556
rect 118016 3544 118022 3596
rect 118053 3587 118111 3593
rect 118053 3553 118065 3587
rect 118099 3584 118111 3587
rect 119249 3587 119307 3593
rect 118099 3556 119200 3584
rect 118099 3553 118111 3556
rect 118053 3547 118111 3553
rect 118510 3516 118516 3528
rect 116964 3488 118516 3516
rect 118510 3476 118516 3488
rect 118568 3476 118574 3528
rect 119172 3516 119200 3556
rect 119249 3553 119261 3587
rect 119295 3584 119307 3587
rect 120184 3584 120212 3624
rect 121917 3621 121929 3624
rect 121963 3621 121975 3655
rect 121917 3615 121975 3621
rect 119295 3556 120212 3584
rect 120261 3587 120319 3593
rect 119295 3553 119307 3556
rect 119249 3547 119307 3553
rect 120261 3553 120273 3587
rect 120307 3584 120319 3587
rect 122006 3584 122012 3596
rect 120307 3556 122012 3584
rect 120307 3553 120319 3556
rect 120261 3547 120319 3553
rect 122006 3544 122012 3556
rect 122064 3544 122070 3596
rect 122098 3544 122104 3596
rect 122156 3584 122162 3596
rect 122156 3556 122201 3584
rect 122156 3544 122162 3556
rect 122300 3516 122328 3692
rect 126238 3652 126244 3664
rect 124968 3624 126244 3652
rect 123018 3544 123024 3596
rect 123076 3584 123082 3596
rect 123481 3587 123539 3593
rect 123481 3584 123493 3587
rect 123076 3556 123493 3584
rect 123076 3544 123082 3556
rect 123481 3553 123493 3556
rect 123527 3553 123539 3587
rect 123481 3547 123539 3553
rect 124968 3525 124996 3624
rect 126238 3612 126244 3624
rect 126296 3612 126302 3664
rect 128188 3652 128216 3692
rect 128262 3680 128268 3732
rect 128320 3720 128326 3732
rect 128541 3723 128599 3729
rect 128541 3720 128553 3723
rect 128320 3692 128553 3720
rect 128320 3680 128326 3692
rect 128541 3689 128553 3692
rect 128587 3689 128599 3723
rect 128541 3683 128599 3689
rect 128630 3680 128636 3732
rect 128688 3720 128694 3732
rect 131298 3720 131304 3732
rect 128688 3692 131304 3720
rect 128688 3680 128694 3692
rect 131298 3680 131304 3692
rect 131356 3680 131362 3732
rect 132310 3680 132316 3732
rect 132368 3720 132374 3732
rect 133233 3723 133291 3729
rect 133233 3720 133245 3723
rect 132368 3692 133245 3720
rect 132368 3680 132374 3692
rect 133233 3689 133245 3692
rect 133279 3689 133291 3723
rect 137830 3720 137836 3732
rect 133233 3683 133291 3689
rect 133616 3692 137836 3720
rect 132402 3652 132408 3664
rect 128188 3624 132408 3652
rect 132402 3612 132408 3624
rect 132460 3612 132466 3664
rect 133046 3612 133052 3664
rect 133104 3652 133110 3664
rect 133616 3652 133644 3692
rect 137830 3680 137836 3692
rect 137888 3680 137894 3732
rect 138198 3680 138204 3732
rect 138256 3720 138262 3732
rect 140314 3720 140320 3732
rect 138256 3692 140320 3720
rect 138256 3680 138262 3692
rect 140314 3680 140320 3692
rect 140372 3680 140378 3732
rect 140777 3723 140835 3729
rect 140777 3689 140789 3723
rect 140823 3720 140835 3723
rect 140958 3720 140964 3732
rect 140823 3692 140964 3720
rect 140823 3689 140835 3692
rect 140777 3683 140835 3689
rect 140958 3680 140964 3692
rect 141016 3680 141022 3732
rect 142249 3723 142307 3729
rect 142249 3689 142261 3723
rect 142295 3720 142307 3723
rect 145466 3720 145472 3732
rect 142295 3692 145472 3720
rect 142295 3689 142307 3692
rect 142249 3683 142307 3689
rect 145466 3680 145472 3692
rect 145524 3680 145530 3732
rect 148965 3723 149023 3729
rect 148965 3689 148977 3723
rect 149011 3720 149023 3723
rect 150434 3720 150440 3732
rect 149011 3692 150440 3720
rect 149011 3689 149023 3692
rect 148965 3683 149023 3689
rect 150434 3680 150440 3692
rect 150492 3680 150498 3732
rect 133104 3624 133644 3652
rect 133104 3612 133110 3624
rect 133690 3612 133696 3664
rect 133748 3652 133754 3664
rect 137922 3652 137928 3664
rect 133748 3624 137928 3652
rect 133748 3612 133754 3624
rect 137922 3612 137928 3624
rect 137980 3612 137986 3664
rect 138382 3612 138388 3664
rect 138440 3652 138446 3664
rect 138569 3655 138627 3661
rect 138569 3652 138581 3655
rect 138440 3624 138581 3652
rect 138440 3612 138446 3624
rect 138569 3621 138581 3624
rect 138615 3621 138627 3655
rect 138569 3615 138627 3621
rect 138658 3612 138664 3664
rect 138716 3652 138722 3664
rect 139210 3652 139216 3664
rect 138716 3624 139216 3652
rect 138716 3612 138722 3624
rect 139210 3612 139216 3624
rect 139268 3612 139274 3664
rect 139762 3652 139768 3664
rect 139723 3624 139768 3652
rect 139762 3612 139768 3624
rect 139820 3612 139826 3664
rect 141326 3652 141332 3664
rect 140884 3624 141332 3652
rect 125045 3587 125103 3593
rect 125045 3553 125057 3587
rect 125091 3584 125103 3587
rect 125594 3584 125600 3596
rect 125091 3556 125600 3584
rect 125091 3553 125103 3556
rect 125045 3547 125103 3553
rect 125594 3544 125600 3556
rect 125652 3544 125658 3596
rect 125873 3587 125931 3593
rect 125873 3553 125885 3587
rect 125919 3584 125931 3587
rect 125962 3584 125968 3596
rect 125919 3556 125968 3584
rect 125919 3553 125931 3556
rect 125873 3547 125931 3553
rect 125962 3544 125968 3556
rect 126020 3544 126026 3596
rect 126054 3544 126060 3596
rect 126112 3584 126118 3596
rect 126112 3556 126157 3584
rect 126112 3544 126118 3556
rect 127434 3544 127440 3596
rect 127492 3584 127498 3596
rect 128449 3587 128507 3593
rect 127492 3556 128400 3584
rect 127492 3544 127498 3556
rect 119172 3488 122328 3516
rect 124953 3519 125011 3525
rect 124953 3485 124965 3519
rect 124999 3485 125011 3519
rect 128262 3516 128268 3528
rect 124953 3479 125011 3485
rect 125060 3488 128268 3516
rect 125060 3448 125088 3488
rect 128262 3476 128268 3488
rect 128320 3476 128326 3528
rect 128372 3516 128400 3556
rect 128449 3553 128461 3587
rect 128495 3584 128507 3587
rect 128998 3584 129004 3596
rect 128495 3556 129004 3584
rect 128495 3553 128507 3556
rect 128449 3547 128507 3553
rect 128998 3544 129004 3556
rect 129056 3544 129062 3596
rect 129829 3587 129887 3593
rect 129829 3553 129841 3587
rect 129875 3584 129887 3587
rect 130286 3584 130292 3596
rect 129875 3556 130292 3584
rect 129875 3553 129887 3556
rect 129829 3547 129887 3553
rect 130286 3544 130292 3556
rect 130344 3544 130350 3596
rect 131114 3584 131120 3596
rect 131075 3556 131120 3584
rect 131114 3544 131120 3556
rect 131172 3544 131178 3596
rect 133138 3584 133144 3596
rect 133099 3556 133144 3584
rect 133138 3544 133144 3556
rect 133196 3544 133202 3596
rect 133782 3584 133788 3596
rect 133248 3556 133788 3584
rect 133248 3516 133276 3556
rect 133782 3544 133788 3556
rect 133840 3544 133846 3596
rect 134058 3544 134064 3596
rect 134116 3584 134122 3596
rect 134153 3587 134211 3593
rect 134153 3584 134165 3587
rect 134116 3556 134165 3584
rect 134116 3544 134122 3556
rect 134153 3553 134165 3556
rect 134199 3553 134211 3587
rect 134153 3547 134211 3553
rect 134518 3544 134524 3596
rect 134576 3584 134582 3596
rect 135165 3587 135223 3593
rect 135165 3584 135177 3587
rect 134576 3556 135177 3584
rect 134576 3544 134582 3556
rect 135165 3553 135177 3556
rect 135211 3553 135223 3587
rect 136358 3584 136364 3596
rect 136319 3556 136364 3584
rect 135165 3547 135223 3553
rect 136358 3544 136364 3556
rect 136416 3544 136422 3596
rect 137462 3544 137468 3596
rect 137520 3584 137526 3596
rect 137557 3587 137615 3593
rect 137557 3584 137569 3587
rect 137520 3556 137569 3584
rect 137520 3544 137526 3556
rect 137557 3553 137569 3556
rect 137603 3553 137615 3587
rect 140884 3584 140912 3624
rect 141326 3612 141332 3624
rect 141384 3612 141390 3664
rect 151814 3652 151820 3664
rect 141988 3624 148824 3652
rect 137557 3547 137615 3553
rect 137848 3556 140912 3584
rect 137848 3528 137876 3556
rect 141142 3544 141148 3596
rect 141200 3584 141206 3596
rect 141988 3584 142016 3624
rect 142154 3584 142160 3596
rect 141200 3556 142016 3584
rect 142115 3556 142160 3584
rect 141200 3544 141206 3556
rect 142154 3544 142160 3556
rect 142212 3544 142218 3596
rect 142246 3544 142252 3596
rect 142304 3584 142310 3596
rect 144365 3587 144423 3593
rect 142304 3556 144224 3584
rect 142304 3544 142310 3556
rect 136542 3516 136548 3528
rect 128372 3488 133276 3516
rect 133340 3488 136548 3516
rect 112732 3420 125088 3448
rect 128446 3408 128452 3460
rect 128504 3448 128510 3460
rect 131117 3451 131175 3457
rect 128504 3420 130608 3448
rect 128504 3408 128510 3420
rect 116486 3380 116492 3392
rect 109788 3352 116492 3380
rect 116486 3340 116492 3352
rect 116544 3340 116550 3392
rect 118142 3380 118148 3392
rect 118103 3352 118148 3380
rect 118142 3340 118148 3352
rect 118200 3340 118206 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119522 3380 119528 3392
rect 118752 3352 119528 3380
rect 118752 3340 118758 3352
rect 119522 3340 119528 3352
rect 119580 3340 119586 3392
rect 120350 3380 120356 3392
rect 120311 3352 120356 3380
rect 120350 3340 120356 3352
rect 120408 3340 120414 3392
rect 121917 3383 121975 3389
rect 121917 3349 121929 3383
rect 121963 3380 121975 3383
rect 124582 3380 124588 3392
rect 121963 3352 124588 3380
rect 121963 3349 121975 3352
rect 121917 3343 121975 3349
rect 124582 3340 124588 3352
rect 124640 3340 124646 3392
rect 125502 3340 125508 3392
rect 125560 3380 125566 3392
rect 125962 3380 125968 3392
rect 125560 3352 125968 3380
rect 125560 3340 125566 3352
rect 125962 3340 125968 3352
rect 126020 3340 126026 3392
rect 126146 3340 126152 3392
rect 126204 3380 126210 3392
rect 130470 3380 130476 3392
rect 126204 3352 130476 3380
rect 126204 3340 126210 3352
rect 130470 3340 130476 3352
rect 130528 3340 130534 3392
rect 130580 3380 130608 3420
rect 131117 3417 131129 3451
rect 131163 3448 131175 3451
rect 131206 3448 131212 3460
rect 131163 3420 131212 3448
rect 131163 3417 131175 3420
rect 131117 3411 131175 3417
rect 131206 3408 131212 3420
rect 131264 3408 131270 3460
rect 131482 3408 131488 3460
rect 131540 3448 131546 3460
rect 133340 3448 133368 3488
rect 136542 3476 136548 3488
rect 136600 3476 136606 3528
rect 136637 3519 136695 3525
rect 136637 3485 136649 3519
rect 136683 3516 136695 3519
rect 137094 3516 137100 3528
rect 136683 3488 137100 3516
rect 136683 3485 136695 3488
rect 136637 3479 136695 3485
rect 137094 3476 137100 3488
rect 137152 3476 137158 3528
rect 137830 3476 137836 3528
rect 137888 3476 137894 3528
rect 138753 3519 138811 3525
rect 138753 3516 138765 3519
rect 137940 3488 138765 3516
rect 131540 3420 133368 3448
rect 131540 3408 131546 3420
rect 134058 3408 134064 3460
rect 134116 3448 134122 3460
rect 137278 3448 137284 3460
rect 134116 3420 137284 3448
rect 134116 3408 134122 3420
rect 137278 3408 137284 3420
rect 137336 3408 137342 3460
rect 137370 3408 137376 3460
rect 137428 3448 137434 3460
rect 137940 3448 137968 3488
rect 138753 3485 138765 3488
rect 138799 3485 138811 3519
rect 138753 3479 138811 3485
rect 138934 3476 138940 3528
rect 138992 3516 138998 3528
rect 143994 3516 144000 3528
rect 138992 3488 144000 3516
rect 138992 3476 138998 3488
rect 143994 3476 144000 3488
rect 144052 3476 144058 3528
rect 138569 3451 138627 3457
rect 138569 3448 138581 3451
rect 137428 3420 137968 3448
rect 138032 3420 138581 3448
rect 137428 3408 137434 3420
rect 131574 3380 131580 3392
rect 130580 3352 131580 3380
rect 131574 3340 131580 3352
rect 131632 3340 131638 3392
rect 131666 3340 131672 3392
rect 131724 3380 131730 3392
rect 133690 3380 133696 3392
rect 131724 3352 133696 3380
rect 131724 3340 131730 3352
rect 133690 3340 133696 3352
rect 133748 3340 133754 3392
rect 133782 3340 133788 3392
rect 133840 3380 133846 3392
rect 134245 3383 134303 3389
rect 134245 3380 134257 3383
rect 133840 3352 134257 3380
rect 133840 3340 133846 3352
rect 134245 3349 134257 3352
rect 134291 3349 134303 3383
rect 134245 3343 134303 3349
rect 134794 3340 134800 3392
rect 134852 3380 134858 3392
rect 135438 3380 135444 3392
rect 134852 3352 135444 3380
rect 134852 3340 134858 3352
rect 135438 3340 135444 3352
rect 135496 3340 135502 3392
rect 137462 3380 137468 3392
rect 137423 3352 137468 3380
rect 137462 3340 137468 3352
rect 137520 3340 137526 3392
rect 137649 3383 137707 3389
rect 137649 3349 137661 3383
rect 137695 3380 137707 3383
rect 138032 3380 138060 3420
rect 138569 3417 138581 3420
rect 138615 3417 138627 3451
rect 144196 3448 144224 3556
rect 144365 3553 144377 3587
rect 144411 3584 144423 3587
rect 144730 3584 144736 3596
rect 144411 3556 144736 3584
rect 144411 3553 144423 3556
rect 144365 3547 144423 3553
rect 144730 3544 144736 3556
rect 144788 3544 144794 3596
rect 147582 3584 147588 3596
rect 144840 3556 147588 3584
rect 144270 3476 144276 3528
rect 144328 3516 144334 3528
rect 144840 3516 144868 3556
rect 147582 3544 147588 3556
rect 147640 3544 147646 3596
rect 144328 3488 144868 3516
rect 144328 3476 144334 3488
rect 144914 3476 144920 3528
rect 144972 3516 144978 3528
rect 145742 3516 145748 3528
rect 144972 3488 145748 3516
rect 144972 3476 144978 3488
rect 145742 3476 145748 3488
rect 145800 3476 145806 3528
rect 148796 3516 148824 3624
rect 148888 3624 151820 3652
rect 148888 3593 148916 3624
rect 151814 3612 151820 3624
rect 151872 3612 151878 3664
rect 148873 3587 148931 3593
rect 148873 3553 148885 3587
rect 148919 3553 148931 3587
rect 156874 3584 156880 3596
rect 148873 3547 148931 3553
rect 148980 3556 156880 3584
rect 148980 3516 149008 3556
rect 156874 3544 156880 3556
rect 156932 3544 156938 3596
rect 148796 3488 149008 3516
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 157150 3516 157156 3528
rect 151872 3488 157156 3516
rect 151872 3476 151878 3488
rect 157150 3476 157156 3488
rect 157208 3476 157214 3528
rect 197262 3476 197268 3528
rect 197320 3516 197326 3528
rect 197998 3516 198004 3528
rect 197320 3488 198004 3516
rect 197320 3476 197326 3488
rect 197998 3476 198004 3488
rect 198056 3476 198062 3528
rect 146018 3448 146024 3460
rect 144196 3420 146024 3448
rect 138569 3411 138627 3417
rect 146018 3408 146024 3420
rect 146076 3408 146082 3460
rect 152642 3448 152648 3460
rect 148888 3420 152648 3448
rect 137695 3352 138060 3380
rect 137695 3349 137707 3352
rect 137649 3343 137707 3349
rect 138382 3340 138388 3392
rect 138440 3380 138446 3392
rect 138750 3380 138756 3392
rect 138440 3352 138756 3380
rect 138440 3340 138446 3352
rect 138750 3340 138756 3352
rect 138808 3340 138814 3392
rect 138934 3340 138940 3392
rect 138992 3380 138998 3392
rect 144270 3380 144276 3392
rect 138992 3352 144276 3380
rect 138992 3340 138998 3352
rect 144270 3340 144276 3352
rect 144328 3340 144334 3392
rect 144454 3380 144460 3392
rect 144415 3352 144460 3380
rect 144454 3340 144460 3352
rect 144512 3340 144518 3392
rect 144730 3380 144736 3392
rect 144691 3352 144736 3380
rect 144730 3340 144736 3352
rect 144788 3340 144794 3392
rect 144822 3340 144828 3392
rect 144880 3380 144886 3392
rect 148888 3380 148916 3420
rect 152642 3408 152648 3420
rect 152700 3408 152706 3460
rect 144880 3352 148916 3380
rect 144880 3340 144886 3352
rect 149698 3340 149704 3392
rect 149756 3380 149762 3392
rect 156969 3383 157027 3389
rect 156969 3380 156981 3383
rect 149756 3352 156981 3380
rect 149756 3340 149762 3352
rect 156969 3349 156981 3352
rect 157015 3349 157027 3383
rect 156969 3343 157027 3349
rect 1104 3290 154560 3312
rect 1104 3238 4078 3290
rect 4130 3238 44078 3290
rect 44130 3238 84078 3290
rect 84130 3238 124078 3290
rect 124130 3238 154560 3290
rect 1104 3216 154560 3238
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 4663 3148 7788 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 7760 3040 7788 3148
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 7929 3179 7987 3185
rect 7929 3176 7941 3179
rect 7892 3148 7941 3176
rect 7892 3136 7898 3148
rect 7929 3145 7941 3148
rect 7975 3145 7987 3179
rect 8938 3176 8944 3188
rect 8899 3148 8944 3176
rect 7929 3139 7987 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 11422 3176 11428 3188
rect 11383 3148 11428 3176
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 12526 3176 12532 3188
rect 12487 3148 12532 3176
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 13504 3148 13553 3176
rect 13504 3136 13510 3148
rect 13541 3145 13553 3148
rect 13587 3145 13599 3179
rect 14918 3176 14924 3188
rect 14879 3148 14924 3176
rect 13541 3139 13599 3145
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 19978 3176 19984 3188
rect 19939 3148 19984 3176
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 21082 3176 21088 3188
rect 21043 3148 21088 3176
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 27062 3176 27068 3188
rect 24412 3148 26924 3176
rect 27023 3148 27068 3176
rect 14182 3040 14188 3052
rect 4479 3012 6868 3040
rect 7760 3012 14188 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 6840 2981 6868 3012
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 4525 2975 4583 2981
rect 4525 2972 4537 2975
rect 1544 2944 4537 2972
rect 1544 2932 1550 2944
rect 4525 2941 4537 2944
rect 4571 2941 4583 2975
rect 4525 2935 4583 2941
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 198 2864 204 2916
rect 256 2904 262 2916
rect 5552 2904 5580 2935
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 7156 2944 7849 2972
rect 7156 2932 7162 2944
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 8846 2972 8852 2984
rect 8807 2944 8852 2972
rect 7837 2935 7895 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 11333 2975 11391 2981
rect 11333 2972 11345 2975
rect 9824 2944 11345 2972
rect 9824 2932 9830 2944
rect 11333 2941 11345 2944
rect 11379 2941 11391 2975
rect 11333 2935 11391 2941
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 11572 2944 12449 2972
rect 11572 2932 11578 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 13449 2975 13507 2981
rect 13449 2941 13461 2975
rect 13495 2941 13507 2975
rect 13449 2935 13507 2941
rect 256 2876 5580 2904
rect 6917 2907 6975 2913
rect 256 2864 262 2876
rect 6917 2873 6929 2907
rect 6963 2904 6975 2907
rect 6963 2876 11560 2904
rect 6963 2873 6975 2876
rect 6917 2867 6975 2873
rect 1854 2796 1860 2848
rect 1912 2836 1918 2848
rect 4433 2839 4491 2845
rect 4433 2836 4445 2839
rect 1912 2808 4445 2836
rect 1912 2796 1918 2808
rect 4433 2805 4445 2808
rect 4479 2805 4491 2839
rect 4433 2799 4491 2805
rect 5629 2839 5687 2845
rect 5629 2805 5641 2839
rect 5675 2836 5687 2839
rect 11054 2836 11060 2848
rect 5675 2808 11060 2836
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11532 2836 11560 2876
rect 12342 2864 12348 2916
rect 12400 2904 12406 2916
rect 13464 2904 13492 2935
rect 14550 2932 14556 2984
rect 14608 2972 14614 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14608 2944 14841 2972
rect 14608 2932 14614 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 24412 2981 24440 3148
rect 25406 3068 25412 3120
rect 25464 3108 25470 3120
rect 26896 3108 26924 3148
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 29365 3179 29423 3185
rect 29365 3145 29377 3179
rect 29411 3176 29423 3179
rect 29546 3176 29552 3188
rect 29411 3148 29552 3176
rect 29411 3145 29423 3148
rect 29365 3139 29423 3145
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 32309 3179 32367 3185
rect 32309 3145 32321 3179
rect 32355 3176 32367 3179
rect 32582 3176 32588 3188
rect 32355 3148 32588 3176
rect 32355 3145 32367 3148
rect 32309 3139 32367 3145
rect 32582 3136 32588 3148
rect 32640 3136 32646 3188
rect 33321 3179 33379 3185
rect 33321 3145 33333 3179
rect 33367 3176 33379 3179
rect 33594 3176 33600 3188
rect 33367 3148 33600 3176
rect 33367 3145 33379 3148
rect 33321 3139 33379 3145
rect 33594 3136 33600 3148
rect 33652 3136 33658 3188
rect 41233 3179 41291 3185
rect 41233 3145 41245 3179
rect 41279 3176 41291 3179
rect 41322 3176 41328 3188
rect 41279 3148 41328 3176
rect 41279 3145 41291 3148
rect 41233 3139 41291 3145
rect 41322 3136 41328 3148
rect 41380 3136 41386 3188
rect 42797 3179 42855 3185
rect 42797 3145 42809 3179
rect 42843 3176 42855 3179
rect 43070 3176 43076 3188
rect 42843 3148 43076 3176
rect 42843 3145 42855 3148
rect 42797 3139 42855 3145
rect 43070 3136 43076 3148
rect 43128 3136 43134 3188
rect 43806 3176 43812 3188
rect 43767 3148 43812 3176
rect 43806 3136 43812 3148
rect 43864 3136 43870 3188
rect 46201 3179 46259 3185
rect 46201 3145 46213 3179
rect 46247 3176 46259 3179
rect 47210 3176 47216 3188
rect 46247 3148 47216 3176
rect 46247 3145 46259 3148
rect 46201 3139 46259 3145
rect 47210 3136 47216 3148
rect 47268 3136 47274 3188
rect 48593 3179 48651 3185
rect 48593 3145 48605 3179
rect 48639 3176 48651 3179
rect 49142 3176 49148 3188
rect 48639 3148 49148 3176
rect 48639 3145 48651 3148
rect 48593 3139 48651 3145
rect 49142 3136 49148 3148
rect 49200 3136 49206 3188
rect 50709 3179 50767 3185
rect 50709 3145 50721 3179
rect 50755 3176 50767 3179
rect 52822 3176 52828 3188
rect 50755 3148 52828 3176
rect 50755 3145 50767 3148
rect 50709 3139 50767 3145
rect 52822 3136 52828 3148
rect 52880 3136 52886 3188
rect 53558 3176 53564 3188
rect 53519 3148 53564 3176
rect 53558 3136 53564 3148
rect 53616 3136 53622 3188
rect 54573 3179 54631 3185
rect 54573 3145 54585 3179
rect 54619 3176 54631 3179
rect 55950 3176 55956 3188
rect 54619 3148 55956 3176
rect 54619 3145 54631 3148
rect 54573 3139 54631 3145
rect 55950 3136 55956 3148
rect 56008 3136 56014 3188
rect 57885 3179 57943 3185
rect 57885 3145 57897 3179
rect 57931 3176 57943 3179
rect 59078 3176 59084 3188
rect 57931 3148 59084 3176
rect 57931 3145 57943 3148
rect 57885 3139 57943 3145
rect 59078 3136 59084 3148
rect 59136 3136 59142 3188
rect 92474 3136 92480 3188
rect 92532 3176 92538 3188
rect 95234 3176 95240 3188
rect 92532 3148 95240 3176
rect 92532 3136 92538 3148
rect 95234 3136 95240 3148
rect 95292 3136 95298 3188
rect 96798 3136 96804 3188
rect 96856 3176 96862 3188
rect 104158 3176 104164 3188
rect 96856 3148 104164 3176
rect 96856 3136 96862 3148
rect 104158 3136 104164 3148
rect 104216 3136 104222 3188
rect 104526 3136 104532 3188
rect 104584 3176 104590 3188
rect 104713 3179 104771 3185
rect 104713 3176 104725 3179
rect 104584 3148 104725 3176
rect 104584 3136 104590 3148
rect 104713 3145 104725 3148
rect 104759 3145 104771 3179
rect 104713 3139 104771 3145
rect 106185 3179 106243 3185
rect 106185 3145 106197 3179
rect 106231 3176 106243 3179
rect 109126 3176 109132 3188
rect 106231 3148 109132 3176
rect 106231 3145 106243 3148
rect 106185 3139 106243 3145
rect 109126 3136 109132 3148
rect 109184 3136 109190 3188
rect 111058 3176 111064 3188
rect 111019 3148 111064 3176
rect 111058 3136 111064 3148
rect 111116 3136 111122 3188
rect 116302 3176 116308 3188
rect 111904 3148 116308 3176
rect 29822 3108 29828 3120
rect 25464 3080 26648 3108
rect 26896 3080 29828 3108
rect 25464 3068 25470 3080
rect 24489 3043 24547 3049
rect 24489 3009 24501 3043
rect 24535 3040 24547 3043
rect 26510 3040 26516 3052
rect 24535 3012 26516 3040
rect 24535 3009 24547 3012
rect 24489 3003 24547 3009
rect 26510 3000 26516 3012
rect 26568 3000 26574 3052
rect 19889 2975 19947 2981
rect 19889 2972 19901 2975
rect 18472 2944 19901 2972
rect 18472 2932 18478 2944
rect 19889 2941 19901 2944
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 24397 2975 24455 2981
rect 24397 2941 24409 2975
rect 24443 2941 24455 2975
rect 24397 2935 24455 2941
rect 25409 2975 25467 2981
rect 25409 2941 25421 2975
rect 25455 2972 25467 2975
rect 25866 2972 25872 2984
rect 25455 2944 25872 2972
rect 25455 2941 25467 2944
rect 25409 2935 25467 2941
rect 12400 2876 13492 2904
rect 12400 2864 12406 2876
rect 19334 2864 19340 2916
rect 19392 2904 19398 2916
rect 21008 2904 21036 2935
rect 25866 2932 25872 2944
rect 25924 2932 25930 2984
rect 19392 2876 21036 2904
rect 19392 2864 19398 2876
rect 22738 2864 22744 2916
rect 22796 2904 22802 2916
rect 25501 2907 25559 2913
rect 25501 2904 25513 2907
rect 22796 2876 25513 2904
rect 22796 2864 22802 2876
rect 25501 2873 25513 2876
rect 25547 2873 25559 2907
rect 25501 2867 25559 2873
rect 15194 2836 15200 2848
rect 11532 2808 15200 2836
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 26620 2836 26648 3080
rect 29822 3068 29828 3080
rect 29880 3068 29886 3120
rect 37182 3068 37188 3120
rect 37240 3108 37246 3120
rect 43438 3108 43444 3120
rect 37240 3080 43444 3108
rect 37240 3068 37246 3080
rect 43438 3068 43444 3080
rect 43496 3068 43502 3120
rect 62850 3108 62856 3120
rect 52380 3080 62856 3108
rect 26694 3000 26700 3052
rect 26752 3040 26758 3052
rect 26752 3012 29316 3040
rect 26752 3000 26758 3012
rect 29288 2981 29316 3012
rect 31570 3000 31576 3052
rect 31628 3040 31634 3052
rect 31628 3012 33364 3040
rect 31628 3000 31634 3012
rect 26973 2975 27031 2981
rect 26973 2941 26985 2975
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 29273 2975 29331 2981
rect 29273 2941 29285 2975
rect 29319 2941 29331 2975
rect 29273 2935 29331 2941
rect 32217 2975 32275 2981
rect 32217 2941 32229 2975
rect 32263 2972 32275 2975
rect 33134 2972 33140 2984
rect 32263 2944 33140 2972
rect 32263 2941 32275 2944
rect 32217 2935 32275 2941
rect 26988 2904 27016 2935
rect 33134 2932 33140 2944
rect 33192 2932 33198 2984
rect 33229 2975 33287 2981
rect 33229 2941 33241 2975
rect 33275 2941 33287 2975
rect 33229 2935 33287 2941
rect 29362 2904 29368 2916
rect 26988 2876 29368 2904
rect 29362 2864 29368 2876
rect 29420 2864 29426 2916
rect 31110 2864 31116 2916
rect 31168 2904 31174 2916
rect 33244 2904 33272 2935
rect 31168 2876 33272 2904
rect 33336 2904 33364 3012
rect 35434 3000 35440 3052
rect 35492 3040 35498 3052
rect 35492 3012 36308 3040
rect 35492 3000 35498 3012
rect 36280 2972 36308 3012
rect 36354 3000 36360 3052
rect 36412 3040 36418 3052
rect 43070 3040 43076 3052
rect 36412 3012 43076 3040
rect 36412 3000 36418 3012
rect 43070 3000 43076 3012
rect 43128 3000 43134 3052
rect 44729 3043 44787 3049
rect 44729 3009 44741 3043
rect 44775 3040 44787 3043
rect 45094 3040 45100 3052
rect 44775 3012 45100 3040
rect 44775 3009 44787 3012
rect 44729 3003 44787 3009
rect 45094 3000 45100 3012
rect 45152 3000 45158 3052
rect 45186 3000 45192 3052
rect 45244 3040 45250 3052
rect 47486 3040 47492 3052
rect 45244 3012 47492 3040
rect 45244 3000 45250 3012
rect 47486 3000 47492 3012
rect 47544 3000 47550 3052
rect 36280 2944 37872 2972
rect 37734 2904 37740 2916
rect 33336 2876 37740 2904
rect 31168 2864 31174 2876
rect 37734 2864 37740 2876
rect 37792 2864 37798 2916
rect 33042 2836 33048 2848
rect 26620 2808 33048 2836
rect 33042 2796 33048 2808
rect 33100 2796 33106 2848
rect 37844 2836 37872 2944
rect 38470 2932 38476 2984
rect 38528 2972 38534 2984
rect 41141 2975 41199 2981
rect 41141 2972 41153 2975
rect 38528 2944 41153 2972
rect 38528 2932 38534 2944
rect 41141 2941 41153 2944
rect 41187 2941 41199 2975
rect 42705 2975 42763 2981
rect 42705 2972 42717 2975
rect 41141 2935 41199 2941
rect 41248 2944 42717 2972
rect 39482 2864 39488 2916
rect 39540 2904 39546 2916
rect 41248 2904 41276 2944
rect 42705 2941 42717 2944
rect 42751 2941 42763 2975
rect 42705 2935 42763 2941
rect 43717 2975 43775 2981
rect 43717 2941 43729 2975
rect 43763 2941 43775 2975
rect 43717 2935 43775 2941
rect 39540 2876 41276 2904
rect 39540 2864 39546 2876
rect 42426 2864 42432 2916
rect 42484 2904 42490 2916
rect 43732 2904 43760 2935
rect 45002 2932 45008 2984
rect 45060 2972 45066 2984
rect 52380 2981 52408 3080
rect 62850 3068 62856 3080
rect 62908 3068 62914 3120
rect 87230 3068 87236 3120
rect 87288 3108 87294 3120
rect 99190 3108 99196 3120
rect 87288 3080 99196 3108
rect 87288 3068 87294 3080
rect 99190 3068 99196 3080
rect 99248 3068 99254 3120
rect 99282 3068 99288 3120
rect 99340 3108 99346 3120
rect 99340 3080 103284 3108
rect 99340 3068 99346 3080
rect 52641 3043 52699 3049
rect 52641 3009 52653 3043
rect 52687 3040 52699 3043
rect 53926 3040 53932 3052
rect 52687 3012 53932 3040
rect 52687 3009 52699 3012
rect 52641 3003 52699 3009
rect 53926 3000 53932 3012
rect 53984 3000 53990 3052
rect 54018 3000 54024 3052
rect 54076 3040 54082 3052
rect 58066 3040 58072 3052
rect 54076 3012 58072 3040
rect 54076 3000 54082 3012
rect 58066 3000 58072 3012
rect 58124 3000 58130 3052
rect 60274 3000 60280 3052
rect 60332 3040 60338 3052
rect 62945 3043 63003 3049
rect 62945 3040 62957 3043
rect 60332 3012 62957 3040
rect 60332 3000 60338 3012
rect 62945 3009 62957 3012
rect 62991 3009 63003 3043
rect 73246 3040 73252 3052
rect 62945 3003 63003 3009
rect 69216 3012 73252 3040
rect 46109 2975 46167 2981
rect 46109 2972 46121 2975
rect 45060 2944 46121 2972
rect 45060 2932 45066 2944
rect 46109 2941 46121 2944
rect 46155 2941 46167 2975
rect 46109 2935 46167 2941
rect 48501 2975 48559 2981
rect 48501 2941 48513 2975
rect 48547 2941 48559 2975
rect 48501 2935 48559 2941
rect 50617 2975 50675 2981
rect 50617 2941 50629 2975
rect 50663 2941 50675 2975
rect 50617 2935 50675 2941
rect 52365 2975 52423 2981
rect 52365 2941 52377 2975
rect 52411 2941 52423 2975
rect 53469 2975 53527 2981
rect 53469 2972 53481 2975
rect 52365 2935 52423 2941
rect 52472 2944 53481 2972
rect 42484 2876 43760 2904
rect 43824 2876 45876 2904
rect 42484 2864 42490 2876
rect 41598 2836 41604 2848
rect 37844 2808 41604 2836
rect 41598 2796 41604 2808
rect 41656 2796 41662 2848
rect 41966 2796 41972 2848
rect 42024 2836 42030 2848
rect 42794 2836 42800 2848
rect 42024 2808 42800 2836
rect 42024 2796 42030 2808
rect 42794 2796 42800 2808
rect 42852 2796 42858 2848
rect 43714 2796 43720 2848
rect 43772 2836 43778 2848
rect 43824 2836 43852 2876
rect 43772 2808 43852 2836
rect 43772 2796 43778 2808
rect 44174 2796 44180 2848
rect 44232 2836 44238 2848
rect 45646 2836 45652 2848
rect 44232 2808 45652 2836
rect 44232 2796 44238 2808
rect 45646 2796 45652 2808
rect 45704 2796 45710 2848
rect 45848 2836 45876 2876
rect 45922 2864 45928 2916
rect 45980 2904 45986 2916
rect 48516 2904 48544 2935
rect 45980 2876 48544 2904
rect 45980 2864 45986 2876
rect 49878 2836 49884 2848
rect 45848 2808 49884 2836
rect 49878 2796 49884 2808
rect 49936 2796 49942 2848
rect 50632 2836 50660 2935
rect 51534 2864 51540 2916
rect 51592 2904 51598 2916
rect 52472 2904 52500 2944
rect 53469 2941 53481 2944
rect 53515 2941 53527 2975
rect 53469 2935 53527 2941
rect 54202 2932 54208 2984
rect 54260 2972 54266 2984
rect 54481 2975 54539 2981
rect 54481 2972 54493 2975
rect 54260 2944 54493 2972
rect 54260 2932 54266 2944
rect 54481 2941 54493 2944
rect 54527 2941 54539 2975
rect 54481 2935 54539 2941
rect 55030 2932 55036 2984
rect 55088 2972 55094 2984
rect 57793 2975 57851 2981
rect 57793 2972 57805 2975
rect 55088 2944 57805 2972
rect 55088 2932 55094 2944
rect 57793 2941 57805 2944
rect 57839 2941 57851 2975
rect 57793 2935 57851 2941
rect 58434 2932 58440 2984
rect 58492 2972 58498 2984
rect 60369 2975 60427 2981
rect 60369 2972 60381 2975
rect 58492 2944 60381 2972
rect 58492 2932 58498 2944
rect 60369 2941 60381 2944
rect 60415 2941 60427 2975
rect 63034 2972 63040 2984
rect 62995 2944 63040 2972
rect 60369 2935 60427 2941
rect 63034 2932 63040 2944
rect 63092 2932 63098 2984
rect 64506 2932 64512 2984
rect 64564 2972 64570 2984
rect 64877 2975 64935 2981
rect 64877 2972 64889 2975
rect 64564 2944 64889 2972
rect 64564 2932 64570 2944
rect 64877 2941 64889 2944
rect 64923 2941 64935 2975
rect 66990 2972 66996 2984
rect 66951 2944 66996 2972
rect 64877 2935 64935 2941
rect 66990 2932 66996 2944
rect 67048 2932 67054 2984
rect 69216 2981 69244 3012
rect 73246 3000 73252 3012
rect 73304 3000 73310 3052
rect 74169 3043 74227 3049
rect 74169 3009 74181 3043
rect 74215 3040 74227 3043
rect 74442 3040 74448 3052
rect 74215 3012 74448 3040
rect 74215 3009 74227 3012
rect 74169 3003 74227 3009
rect 74442 3000 74448 3012
rect 74500 3000 74506 3052
rect 78677 3043 78735 3049
rect 78677 3009 78689 3043
rect 78723 3040 78735 3043
rect 79778 3040 79784 3052
rect 78723 3012 79784 3040
rect 78723 3009 78735 3012
rect 78677 3003 78735 3009
rect 79778 3000 79784 3012
rect 79836 3000 79842 3052
rect 81342 3040 81348 3052
rect 81303 3012 81348 3040
rect 81342 3000 81348 3012
rect 81400 3000 81406 3052
rect 87138 3040 87144 3052
rect 87099 3012 87144 3040
rect 87138 3000 87144 3012
rect 87196 3000 87202 3052
rect 89717 3043 89775 3049
rect 89717 3009 89729 3043
rect 89763 3040 89775 3043
rect 89806 3040 89812 3052
rect 89763 3012 89812 3040
rect 89763 3009 89775 3012
rect 89717 3003 89775 3009
rect 89806 3000 89812 3012
rect 89864 3000 89870 3052
rect 93673 3043 93731 3049
rect 93673 3009 93685 3043
rect 93719 3040 93731 3043
rect 99466 3040 99472 3052
rect 93719 3012 99472 3040
rect 93719 3009 93731 3012
rect 93673 3003 93731 3009
rect 99466 3000 99472 3012
rect 99524 3000 99530 3052
rect 101214 3040 101220 3052
rect 99760 3012 101220 3040
rect 69201 2975 69259 2981
rect 69201 2941 69213 2975
rect 69247 2941 69259 2975
rect 70854 2972 70860 2984
rect 70815 2944 70860 2972
rect 69201 2935 69259 2941
rect 70854 2932 70860 2944
rect 70912 2932 70918 2984
rect 72694 2972 72700 2984
rect 72655 2944 72700 2972
rect 72694 2932 72700 2944
rect 72752 2932 72758 2984
rect 76190 2972 76196 2984
rect 76151 2944 76196 2972
rect 76190 2932 76196 2944
rect 76248 2932 76254 2984
rect 77757 2975 77815 2981
rect 77757 2941 77769 2975
rect 77803 2972 77815 2975
rect 77938 2972 77944 2984
rect 77803 2944 77944 2972
rect 77803 2941 77815 2944
rect 77757 2935 77815 2941
rect 77938 2932 77944 2944
rect 77996 2932 78002 2984
rect 80422 2972 80428 2984
rect 80383 2944 80428 2972
rect 80422 2932 80428 2944
rect 80480 2932 80486 2984
rect 80606 2932 80612 2984
rect 80664 2972 80670 2984
rect 83369 2975 83427 2981
rect 83369 2972 83381 2975
rect 80664 2944 83381 2972
rect 80664 2932 80670 2944
rect 83369 2941 83381 2944
rect 83415 2941 83427 2975
rect 85758 2972 85764 2984
rect 85719 2944 85764 2972
rect 83369 2935 83427 2941
rect 85758 2932 85764 2944
rect 85816 2932 85822 2984
rect 87322 2932 87328 2984
rect 87380 2972 87386 2984
rect 88245 2975 88303 2981
rect 88245 2972 88257 2975
rect 87380 2944 88257 2972
rect 87380 2932 87386 2944
rect 88245 2941 88257 2944
rect 88291 2941 88303 2975
rect 91462 2972 91468 2984
rect 91423 2944 91468 2972
rect 88245 2935 88303 2941
rect 91462 2932 91468 2944
rect 91520 2932 91526 2984
rect 93578 2972 93584 2984
rect 93539 2944 93584 2972
rect 93578 2932 93584 2944
rect 93636 2932 93642 2984
rect 94590 2972 94596 2984
rect 94551 2944 94596 2972
rect 94590 2932 94596 2944
rect 94648 2932 94654 2984
rect 95878 2932 95884 2984
rect 95936 2972 95942 2984
rect 98822 2972 98828 2984
rect 95936 2944 97028 2972
rect 98783 2944 98828 2972
rect 95936 2932 95942 2944
rect 51592 2876 52500 2904
rect 51592 2864 51598 2876
rect 52546 2864 52552 2916
rect 52604 2904 52610 2916
rect 54662 2904 54668 2916
rect 52604 2876 54668 2904
rect 52604 2864 52610 2876
rect 54662 2864 54668 2876
rect 54720 2864 54726 2916
rect 58526 2864 58532 2916
rect 58584 2904 58590 2916
rect 60277 2907 60335 2913
rect 60277 2904 60289 2907
rect 58584 2876 60289 2904
rect 58584 2864 58590 2876
rect 60277 2873 60289 2876
rect 60323 2873 60335 2907
rect 60277 2867 60335 2873
rect 61562 2864 61568 2916
rect 61620 2904 61626 2916
rect 64785 2907 64843 2913
rect 64785 2904 64797 2907
rect 61620 2876 64797 2904
rect 61620 2864 61626 2876
rect 64785 2873 64797 2876
rect 64831 2873 64843 2907
rect 66346 2904 66352 2916
rect 66307 2876 66352 2904
rect 64785 2867 64843 2873
rect 66346 2864 66352 2876
rect 66404 2864 66410 2916
rect 68554 2904 68560 2916
rect 68515 2876 68560 2904
rect 68554 2864 68560 2876
rect 68612 2864 68618 2916
rect 69014 2864 69020 2916
rect 69072 2904 69078 2916
rect 70489 2907 70547 2913
rect 70489 2904 70501 2907
rect 69072 2876 70501 2904
rect 69072 2864 69078 2876
rect 70489 2873 70501 2876
rect 70535 2873 70547 2907
rect 70489 2867 70547 2873
rect 71590 2864 71596 2916
rect 71648 2904 71654 2916
rect 72053 2907 72111 2913
rect 72053 2904 72065 2907
rect 71648 2876 72065 2904
rect 71648 2864 71654 2876
rect 72053 2873 72065 2876
rect 72099 2873 72111 2907
rect 72053 2867 72111 2873
rect 74626 2864 74632 2916
rect 74684 2904 74690 2916
rect 75549 2907 75607 2913
rect 75549 2904 75561 2907
rect 74684 2876 75561 2904
rect 74684 2864 74690 2876
rect 75549 2873 75561 2876
rect 75595 2873 75607 2907
rect 75549 2867 75607 2873
rect 76834 2864 76840 2916
rect 76892 2904 76898 2916
rect 77113 2907 77171 2913
rect 77113 2904 77125 2907
rect 76892 2876 77125 2904
rect 76892 2864 76898 2876
rect 77113 2873 77125 2876
rect 77159 2873 77171 2907
rect 77113 2867 77171 2873
rect 80517 2907 80575 2913
rect 80517 2873 80529 2907
rect 80563 2904 80575 2907
rect 80790 2904 80796 2916
rect 80563 2876 80796 2904
rect 80563 2873 80575 2876
rect 80517 2867 80575 2873
rect 80790 2864 80796 2876
rect 80848 2864 80854 2916
rect 82906 2864 82912 2916
rect 82964 2904 82970 2916
rect 83277 2907 83335 2913
rect 83277 2904 83289 2907
rect 82964 2876 83289 2904
rect 82964 2864 82970 2876
rect 83277 2873 83289 2876
rect 83323 2873 83335 2907
rect 83277 2867 83335 2873
rect 85114 2864 85120 2916
rect 85172 2904 85178 2916
rect 85393 2907 85451 2913
rect 85393 2904 85405 2907
rect 85172 2876 85405 2904
rect 85172 2864 85178 2876
rect 85393 2873 85405 2876
rect 85439 2873 85451 2907
rect 85393 2867 85451 2873
rect 88889 2907 88947 2913
rect 88889 2873 88901 2907
rect 88935 2904 88947 2907
rect 89438 2904 89444 2916
rect 88935 2876 89444 2904
rect 88935 2873 88947 2876
rect 88889 2867 88947 2873
rect 89438 2864 89444 2876
rect 89496 2864 89502 2916
rect 91741 2907 91799 2913
rect 91741 2873 91753 2907
rect 91787 2904 91799 2907
rect 94314 2904 94320 2916
rect 91787 2876 94320 2904
rect 91787 2873 91799 2876
rect 91741 2867 91799 2873
rect 94314 2864 94320 2876
rect 94372 2864 94378 2916
rect 95237 2907 95295 2913
rect 95237 2873 95249 2907
rect 95283 2904 95295 2907
rect 96890 2904 96896 2916
rect 95283 2876 96896 2904
rect 95283 2873 95295 2876
rect 95237 2867 95295 2873
rect 96890 2864 96896 2876
rect 96948 2864 96954 2916
rect 53466 2836 53472 2848
rect 50632 2808 53472 2836
rect 53466 2796 53472 2808
rect 53524 2796 53530 2848
rect 53558 2796 53564 2848
rect 53616 2836 53622 2848
rect 56778 2836 56784 2848
rect 53616 2808 56784 2836
rect 53616 2796 53622 2808
rect 56778 2796 56784 2808
rect 56836 2796 56842 2848
rect 90910 2796 90916 2848
rect 90968 2836 90974 2848
rect 96617 2839 96675 2845
rect 96617 2836 96629 2839
rect 90968 2808 96629 2836
rect 90968 2796 90974 2808
rect 96617 2805 96629 2808
rect 96663 2805 96675 2839
rect 97000 2836 97028 2944
rect 98822 2932 98828 2944
rect 98880 2932 98886 2984
rect 98917 2907 98975 2913
rect 98917 2873 98929 2907
rect 98963 2904 98975 2907
rect 99760 2904 99788 3012
rect 101214 3000 101220 3012
rect 101272 3000 101278 3052
rect 100570 2972 100576 2984
rect 100531 2944 100576 2972
rect 100570 2932 100576 2944
rect 100628 2932 100634 2984
rect 100665 2975 100723 2981
rect 100665 2941 100677 2975
rect 100711 2972 100723 2975
rect 102962 2972 102968 2984
rect 100711 2944 102968 2972
rect 100711 2941 100723 2944
rect 100665 2935 100723 2941
rect 102962 2932 102968 2944
rect 103020 2932 103026 2984
rect 103146 2972 103152 2984
rect 103107 2944 103152 2972
rect 103146 2932 103152 2944
rect 103204 2932 103210 2984
rect 100386 2904 100392 2916
rect 98963 2876 99788 2904
rect 99852 2876 100392 2904
rect 98963 2873 98975 2876
rect 98917 2867 98975 2873
rect 99852 2836 99880 2876
rect 100386 2864 100392 2876
rect 100444 2864 100450 2916
rect 102134 2864 102140 2916
rect 102192 2904 102198 2916
rect 102505 2907 102563 2913
rect 102505 2904 102517 2907
rect 102192 2876 102517 2904
rect 102192 2864 102198 2876
rect 102505 2873 102517 2876
rect 102551 2873 102563 2907
rect 103256 2904 103284 3080
rect 104250 3068 104256 3120
rect 104308 3108 104314 3120
rect 108114 3108 108120 3120
rect 104308 3080 108120 3108
rect 104308 3068 104314 3080
rect 108114 3068 108120 3080
rect 108172 3068 108178 3120
rect 111426 3108 111432 3120
rect 108316 3080 111432 3108
rect 108022 3040 108028 3052
rect 104636 3012 108028 3040
rect 104636 2981 104664 3012
rect 108022 3000 108028 3012
rect 108080 3000 108086 3052
rect 104621 2975 104679 2981
rect 104621 2941 104633 2975
rect 104667 2941 104679 2975
rect 104621 2935 104679 2941
rect 106185 2975 106243 2981
rect 106185 2941 106197 2975
rect 106231 2972 106243 2975
rect 106918 2972 106924 2984
rect 106231 2944 106924 2972
rect 106231 2941 106243 2944
rect 106185 2935 106243 2941
rect 106918 2932 106924 2944
rect 106976 2932 106982 2984
rect 108316 2972 108344 3080
rect 111426 3068 111432 3080
rect 111484 3068 111490 3120
rect 107028 2944 108344 2972
rect 108485 2975 108543 2981
rect 107028 2904 107056 2944
rect 108485 2941 108497 2975
rect 108531 2972 108543 2975
rect 109218 2972 109224 2984
rect 108531 2944 109224 2972
rect 108531 2941 108543 2944
rect 108485 2935 108543 2941
rect 109218 2932 109224 2944
rect 109276 2932 109282 2984
rect 109770 2972 109776 2984
rect 109328 2944 109540 2972
rect 109731 2944 109776 2972
rect 103256 2876 107056 2904
rect 102505 2867 102563 2873
rect 107102 2864 107108 2916
rect 107160 2904 107166 2916
rect 107841 2907 107899 2913
rect 107841 2904 107853 2907
rect 107160 2876 107853 2904
rect 107160 2864 107166 2876
rect 107841 2873 107853 2876
rect 107887 2873 107899 2907
rect 107841 2867 107899 2873
rect 108298 2864 108304 2916
rect 108356 2904 108362 2916
rect 109328 2904 109356 2944
rect 108356 2876 109356 2904
rect 109405 2907 109463 2913
rect 108356 2864 108362 2876
rect 109405 2873 109417 2907
rect 109451 2873 109463 2907
rect 109512 2904 109540 2944
rect 109770 2932 109776 2944
rect 109828 2932 109834 2984
rect 110969 2975 111027 2981
rect 110969 2941 110981 2975
rect 111015 2972 111027 2975
rect 111904 2972 111932 3148
rect 116302 3136 116308 3148
rect 116360 3136 116366 3188
rect 116394 3136 116400 3188
rect 116452 3176 116458 3188
rect 116489 3179 116547 3185
rect 116489 3176 116501 3179
rect 116452 3148 116501 3176
rect 116452 3136 116458 3148
rect 116489 3145 116501 3148
rect 116535 3145 116547 3179
rect 116489 3139 116547 3145
rect 116578 3136 116584 3188
rect 116636 3176 116642 3188
rect 117777 3179 117835 3185
rect 117777 3176 117789 3179
rect 116636 3148 117789 3176
rect 116636 3136 116642 3148
rect 117777 3145 117789 3148
rect 117823 3145 117835 3179
rect 117777 3139 117835 3145
rect 117958 3136 117964 3188
rect 118016 3176 118022 3188
rect 123294 3176 123300 3188
rect 118016 3148 123300 3176
rect 118016 3136 118022 3148
rect 123294 3136 123300 3148
rect 123352 3136 123358 3188
rect 123938 3136 123944 3188
rect 123996 3176 124002 3188
rect 126238 3176 126244 3188
rect 123996 3148 126244 3176
rect 123996 3136 124002 3148
rect 126238 3136 126244 3148
rect 126296 3136 126302 3188
rect 126330 3136 126336 3188
rect 126388 3176 126394 3188
rect 128262 3176 128268 3188
rect 126388 3148 128268 3176
rect 126388 3136 126394 3148
rect 128262 3136 128268 3148
rect 128320 3136 128326 3188
rect 128722 3176 128728 3188
rect 128683 3148 128728 3176
rect 128722 3136 128728 3148
rect 128780 3136 128786 3188
rect 128909 3179 128967 3185
rect 128909 3145 128921 3179
rect 128955 3176 128967 3179
rect 129090 3176 129096 3188
rect 128955 3148 129096 3176
rect 128955 3145 128967 3148
rect 128909 3139 128967 3145
rect 129090 3136 129096 3148
rect 129148 3136 129154 3188
rect 129274 3136 129280 3188
rect 129332 3176 129338 3188
rect 130102 3176 130108 3188
rect 129332 3148 130108 3176
rect 129332 3136 129338 3148
rect 130102 3136 130108 3148
rect 130160 3136 130166 3188
rect 130838 3136 130844 3188
rect 130896 3176 130902 3188
rect 131301 3179 131359 3185
rect 131301 3176 131313 3179
rect 130896 3148 131313 3176
rect 130896 3136 130902 3148
rect 131301 3145 131313 3148
rect 131347 3145 131359 3179
rect 134702 3176 134708 3188
rect 131301 3139 131359 3145
rect 132420 3148 134708 3176
rect 117498 3108 117504 3120
rect 111988 3080 117504 3108
rect 111988 2981 112016 3080
rect 117498 3068 117504 3080
rect 117556 3068 117562 3120
rect 118786 3068 118792 3120
rect 118844 3108 118850 3120
rect 121638 3108 121644 3120
rect 118844 3080 120488 3108
rect 121599 3080 121644 3108
rect 118844 3068 118850 3080
rect 112070 3000 112076 3052
rect 112128 3040 112134 3052
rect 113818 3040 113824 3052
rect 112128 3012 112173 3040
rect 113468 3012 113824 3040
rect 112128 3000 112134 3012
rect 113468 2981 113496 3012
rect 113818 3000 113824 3012
rect 113876 3000 113882 3052
rect 118602 3000 118608 3052
rect 118660 3040 118666 3052
rect 120350 3040 120356 3052
rect 118660 3012 120356 3040
rect 118660 3000 118666 3012
rect 120350 3000 120356 3012
rect 120408 3000 120414 3052
rect 120460 3040 120488 3080
rect 121638 3068 121644 3080
rect 121696 3068 121702 3120
rect 126054 3108 126060 3120
rect 125152 3080 126060 3108
rect 120629 3043 120687 3049
rect 120629 3040 120641 3043
rect 120460 3012 120641 3040
rect 120629 3009 120641 3012
rect 120675 3009 120687 3043
rect 120629 3003 120687 3009
rect 123570 3000 123576 3052
rect 123628 3040 123634 3052
rect 123628 3012 123673 3040
rect 123628 3000 123634 3012
rect 111015 2944 111932 2972
rect 111981 2975 112039 2981
rect 111015 2941 111027 2944
rect 110969 2935 111027 2941
rect 111981 2941 111993 2975
rect 112027 2941 112039 2975
rect 111981 2935 112039 2941
rect 113453 2975 113511 2981
rect 113453 2941 113465 2975
rect 113499 2941 113511 2975
rect 113453 2935 113511 2941
rect 115109 2975 115167 2981
rect 115109 2941 115121 2975
rect 115155 2941 115167 2975
rect 115109 2935 115167 2941
rect 116397 2975 116455 2981
rect 116397 2941 116409 2975
rect 116443 2972 116455 2975
rect 117709 2975 117767 2981
rect 116443 2944 117636 2972
rect 116443 2941 116455 2944
rect 116397 2935 116455 2941
rect 112990 2904 112996 2916
rect 109512 2876 112996 2904
rect 109405 2867 109463 2873
rect 97000 2808 99880 2836
rect 96617 2799 96675 2805
rect 100662 2796 100668 2848
rect 100720 2836 100726 2848
rect 103882 2836 103888 2848
rect 100720 2808 103888 2836
rect 100720 2796 100726 2808
rect 103882 2796 103888 2808
rect 103940 2796 103946 2848
rect 106918 2796 106924 2848
rect 106976 2836 106982 2848
rect 109420 2836 109448 2867
rect 112990 2864 112996 2876
rect 113048 2864 113054 2916
rect 113542 2904 113548 2916
rect 113503 2876 113548 2904
rect 113542 2864 113548 2876
rect 113600 2864 113606 2916
rect 115124 2904 115152 2935
rect 116854 2904 116860 2916
rect 115124 2876 116860 2904
rect 116854 2864 116860 2876
rect 116912 2864 116918 2916
rect 117314 2864 117320 2916
rect 117372 2864 117378 2916
rect 117608 2904 117636 2944
rect 117709 2941 117721 2975
rect 117755 2972 117767 2975
rect 119338 2972 119344 2984
rect 117755 2944 119344 2972
rect 117755 2941 117767 2944
rect 117709 2935 117767 2941
rect 119338 2932 119344 2944
rect 119396 2932 119402 2984
rect 119549 2975 119607 2981
rect 119549 2941 119561 2975
rect 119595 2972 119607 2975
rect 120534 2972 120540 2984
rect 119595 2944 120396 2972
rect 120495 2944 120540 2972
rect 119595 2941 119607 2944
rect 119549 2935 119607 2941
rect 120166 2904 120172 2916
rect 117608 2876 120172 2904
rect 120166 2864 120172 2876
rect 120224 2864 120230 2916
rect 106976 2808 109448 2836
rect 106976 2796 106982 2808
rect 109494 2796 109500 2848
rect 109552 2836 109558 2848
rect 111242 2836 111248 2848
rect 109552 2808 111248 2836
rect 109552 2796 109558 2808
rect 111242 2796 111248 2808
rect 111300 2796 111306 2848
rect 111426 2796 111432 2848
rect 111484 2836 111490 2848
rect 115201 2839 115259 2845
rect 115201 2836 115213 2839
rect 111484 2808 115213 2836
rect 111484 2796 111490 2808
rect 115201 2805 115213 2808
rect 115247 2805 115259 2839
rect 115201 2799 115259 2805
rect 116302 2796 116308 2848
rect 116360 2836 116366 2848
rect 116946 2836 116952 2848
rect 116360 2808 116952 2836
rect 116360 2796 116366 2808
rect 116946 2796 116952 2808
rect 117004 2796 117010 2848
rect 117332 2836 117360 2864
rect 119617 2839 119675 2845
rect 119617 2836 119629 2839
rect 117332 2808 119629 2836
rect 119617 2805 119629 2808
rect 119663 2805 119675 2839
rect 120368 2836 120396 2944
rect 120534 2932 120540 2944
rect 120592 2932 120598 2984
rect 121549 2975 121607 2981
rect 121549 2941 121561 2975
rect 121595 2941 121607 2975
rect 121549 2935 121607 2941
rect 123481 2975 123539 2981
rect 123481 2941 123493 2975
rect 123527 2972 123539 2975
rect 125152 2972 125180 3080
rect 126054 3068 126060 3080
rect 126112 3068 126118 3120
rect 127894 3108 127900 3120
rect 127855 3080 127900 3108
rect 127894 3068 127900 3080
rect 127952 3068 127958 3120
rect 125594 3000 125600 3052
rect 125652 3000 125658 3052
rect 126422 3040 126428 3052
rect 126383 3012 126428 3040
rect 126422 3000 126428 3012
rect 126480 3000 126486 3052
rect 123527 2944 125180 2972
rect 125413 2975 125471 2981
rect 123527 2941 123539 2944
rect 123481 2935 123539 2941
rect 125413 2941 125425 2975
rect 125459 2941 125471 2975
rect 125413 2935 125471 2941
rect 125505 2975 125563 2981
rect 125505 2941 125517 2975
rect 125551 2972 125563 2975
rect 125612 2972 125640 3000
rect 125551 2944 125640 2972
rect 125551 2941 125563 2944
rect 125505 2935 125563 2941
rect 121564 2904 121592 2935
rect 125318 2904 125324 2916
rect 121564 2876 125324 2904
rect 125318 2864 125324 2876
rect 125376 2864 125382 2916
rect 125436 2904 125464 2935
rect 126974 2932 126980 2984
rect 127032 2972 127038 2984
rect 127529 2975 127587 2981
rect 127529 2972 127541 2975
rect 127032 2944 127541 2972
rect 127032 2932 127038 2944
rect 127529 2941 127541 2944
rect 127575 2941 127587 2975
rect 128630 2972 128636 2984
rect 127529 2935 127587 2941
rect 128372 2944 128636 2972
rect 126882 2904 126888 2916
rect 125436 2876 126888 2904
rect 126882 2864 126888 2876
rect 126940 2864 126946 2916
rect 128372 2904 128400 2944
rect 128630 2932 128636 2944
rect 128688 2932 128694 2984
rect 128740 2972 128768 3136
rect 130654 3068 130660 3120
rect 130712 3108 130718 3120
rect 132420 3108 132448 3148
rect 134702 3136 134708 3148
rect 134760 3136 134766 3188
rect 134889 3179 134947 3185
rect 134889 3145 134901 3179
rect 134935 3176 134947 3179
rect 135070 3176 135076 3188
rect 134935 3148 135076 3176
rect 134935 3145 134947 3148
rect 134889 3139 134947 3145
rect 135070 3136 135076 3148
rect 135128 3136 135134 3188
rect 135622 3136 135628 3188
rect 135680 3176 135686 3188
rect 135680 3148 138060 3176
rect 135680 3136 135686 3148
rect 130712 3080 132448 3108
rect 130712 3068 130718 3080
rect 132494 3068 132500 3120
rect 132552 3108 132558 3120
rect 133877 3111 133935 3117
rect 132552 3080 133736 3108
rect 132552 3068 132558 3080
rect 129274 3000 129280 3052
rect 129332 3040 129338 3052
rect 129332 3012 130976 3040
rect 129332 3000 129338 3012
rect 128817 2975 128875 2981
rect 128817 2972 128829 2975
rect 128740 2944 128829 2972
rect 128817 2941 128829 2944
rect 128863 2941 128875 2975
rect 128817 2935 128875 2941
rect 129642 2932 129648 2984
rect 129700 2972 129706 2984
rect 129918 2972 129924 2984
rect 129700 2944 129924 2972
rect 129700 2932 129706 2944
rect 129918 2932 129924 2944
rect 129976 2932 129982 2984
rect 127176 2876 128400 2904
rect 121546 2836 121552 2848
rect 120368 2808 121552 2836
rect 119617 2799 119675 2805
rect 121546 2796 121552 2808
rect 121604 2796 121610 2848
rect 123294 2796 123300 2848
rect 123352 2836 123358 2848
rect 125134 2836 125140 2848
rect 123352 2808 125140 2836
rect 123352 2796 123358 2808
rect 125134 2796 125140 2808
rect 125192 2796 125198 2848
rect 125410 2796 125416 2848
rect 125468 2836 125474 2848
rect 127176 2836 127204 2876
rect 128446 2864 128452 2916
rect 128504 2904 128510 2916
rect 130838 2904 130844 2916
rect 128504 2876 130844 2904
rect 128504 2864 128510 2876
rect 130838 2864 130844 2876
rect 130896 2864 130902 2916
rect 130948 2904 130976 3012
rect 131114 3000 131120 3052
rect 131172 3040 131178 3052
rect 133598 3040 133604 3052
rect 131172 3012 133604 3040
rect 131172 3000 131178 3012
rect 133598 3000 133604 3012
rect 133656 3000 133662 3052
rect 133708 3040 133736 3080
rect 133877 3077 133889 3111
rect 133923 3108 133935 3111
rect 136266 3108 136272 3120
rect 133923 3080 136272 3108
rect 133923 3077 133935 3080
rect 133877 3071 133935 3077
rect 136266 3068 136272 3080
rect 136324 3068 136330 3120
rect 137002 3068 137008 3120
rect 137060 3108 137066 3120
rect 137922 3108 137928 3120
rect 137060 3080 137928 3108
rect 137060 3068 137066 3080
rect 137922 3068 137928 3080
rect 137980 3068 137986 3120
rect 138032 3108 138060 3148
rect 138106 3136 138112 3188
rect 138164 3176 138170 3188
rect 138477 3179 138535 3185
rect 138477 3176 138489 3179
rect 138164 3148 138489 3176
rect 138164 3136 138170 3148
rect 138477 3145 138489 3148
rect 138523 3145 138535 3179
rect 138477 3139 138535 3145
rect 138750 3136 138756 3188
rect 138808 3176 138814 3188
rect 141694 3176 141700 3188
rect 138808 3148 141700 3176
rect 138808 3136 138814 3148
rect 141694 3136 141700 3148
rect 141752 3136 141758 3188
rect 142154 3136 142160 3188
rect 142212 3176 142218 3188
rect 157245 3179 157303 3185
rect 157245 3176 157257 3179
rect 142212 3148 157257 3176
rect 142212 3136 142218 3148
rect 157245 3145 157257 3148
rect 157291 3145 157303 3179
rect 157245 3139 157303 3145
rect 144822 3108 144828 3120
rect 138032 3080 144828 3108
rect 144822 3068 144828 3080
rect 144880 3068 144886 3120
rect 145193 3111 145251 3117
rect 145193 3077 145205 3111
rect 145239 3108 145251 3111
rect 145558 3108 145564 3120
rect 145239 3080 145564 3108
rect 145239 3077 145251 3080
rect 145193 3071 145251 3077
rect 145558 3068 145564 3080
rect 145616 3068 145622 3120
rect 146110 3068 146116 3120
rect 146168 3108 146174 3120
rect 147122 3108 147128 3120
rect 146168 3080 147128 3108
rect 146168 3068 146174 3080
rect 147122 3068 147128 3080
rect 147180 3068 147186 3120
rect 147582 3068 147588 3120
rect 147640 3108 147646 3120
rect 151354 3108 151360 3120
rect 147640 3080 151360 3108
rect 147640 3068 147646 3080
rect 151354 3068 151360 3080
rect 151412 3068 151418 3120
rect 151449 3111 151507 3117
rect 151449 3077 151461 3111
rect 151495 3108 151507 3111
rect 156690 3108 156696 3120
rect 151495 3080 156696 3108
rect 151495 3077 151507 3080
rect 151449 3071 151507 3077
rect 156690 3068 156696 3080
rect 156748 3068 156754 3120
rect 156966 3068 156972 3120
rect 157024 3108 157030 3120
rect 157024 3080 157196 3108
rect 157024 3068 157030 3080
rect 134058 3040 134064 3052
rect 133708 3012 134064 3040
rect 134058 3000 134064 3012
rect 134116 3000 134122 3052
rect 134812 3012 137140 3040
rect 131206 2972 131212 2984
rect 131167 2944 131212 2972
rect 131206 2932 131212 2944
rect 131264 2932 131270 2984
rect 132405 2975 132463 2981
rect 132405 2941 132417 2975
rect 132451 2972 132463 2975
rect 133874 2972 133880 2984
rect 132451 2944 133880 2972
rect 132451 2941 132463 2944
rect 132405 2935 132463 2941
rect 133874 2932 133880 2944
rect 133932 2932 133938 2984
rect 133969 2975 134027 2981
rect 133969 2941 133981 2975
rect 134015 2972 134027 2975
rect 134426 2972 134432 2984
rect 134015 2944 134432 2972
rect 134015 2941 134027 2944
rect 133969 2935 134027 2941
rect 134426 2932 134432 2944
rect 134484 2932 134490 2984
rect 134812 2981 134840 3012
rect 134797 2975 134855 2981
rect 134797 2941 134809 2975
rect 134843 2941 134855 2975
rect 135898 2972 135904 2984
rect 135859 2944 135904 2972
rect 134797 2935 134855 2941
rect 135898 2932 135904 2944
rect 135956 2932 135962 2984
rect 135990 2932 135996 2984
rect 136048 2972 136054 2984
rect 136048 2944 136093 2972
rect 136048 2932 136054 2944
rect 137002 2904 137008 2916
rect 130948 2876 137008 2904
rect 137002 2864 137008 2876
rect 137060 2864 137066 2916
rect 137112 2904 137140 3012
rect 137186 3000 137192 3052
rect 137244 3040 137250 3052
rect 138014 3040 138020 3052
rect 137244 3012 137289 3040
rect 137480 3012 138020 3040
rect 137244 3000 137250 3012
rect 137204 2972 137232 3000
rect 137480 2981 137508 3012
rect 138014 3000 138020 3012
rect 138072 3000 138078 3052
rect 157061 3043 157119 3049
rect 157061 3040 157073 3043
rect 138400 3012 157073 3040
rect 137365 2975 137423 2981
rect 137365 2972 137377 2975
rect 137204 2944 137377 2972
rect 137365 2941 137377 2944
rect 137411 2941 137423 2975
rect 137365 2935 137423 2941
rect 137465 2975 137523 2981
rect 137465 2941 137477 2975
rect 137511 2941 137523 2975
rect 138198 2972 138204 2984
rect 137465 2935 137523 2941
rect 137572 2944 138204 2972
rect 137572 2904 137600 2944
rect 138198 2932 138204 2944
rect 138256 2932 138262 2984
rect 138400 2981 138428 3012
rect 157061 3009 157073 3012
rect 157107 3009 157119 3043
rect 157168 3040 157196 3080
rect 157168 3012 162716 3040
rect 157061 3003 157119 3009
rect 162688 2984 162716 3012
rect 162872 3012 167132 3040
rect 138385 2975 138443 2981
rect 138385 2941 138397 2975
rect 138431 2941 138443 2975
rect 143718 2972 143724 2984
rect 138385 2935 138443 2941
rect 138584 2944 143724 2972
rect 138584 2904 138612 2944
rect 143718 2932 143724 2944
rect 143776 2932 143782 2984
rect 145009 2975 145067 2981
rect 145009 2941 145021 2975
rect 145055 2972 145067 2975
rect 145101 2975 145159 2981
rect 145101 2972 145113 2975
rect 145055 2944 145113 2972
rect 145055 2941 145067 2944
rect 145009 2935 145067 2941
rect 145101 2941 145113 2944
rect 145147 2972 145159 2975
rect 145190 2972 145196 2984
rect 145147 2944 145196 2972
rect 145147 2941 145159 2944
rect 145101 2935 145159 2941
rect 145190 2932 145196 2944
rect 145248 2932 145254 2984
rect 145282 2932 145288 2984
rect 145340 2972 145346 2984
rect 148318 2972 148324 2984
rect 145340 2944 148324 2972
rect 145340 2932 145346 2944
rect 148318 2932 148324 2944
rect 148376 2932 148382 2984
rect 151357 2975 151415 2981
rect 151357 2941 151369 2975
rect 151403 2972 151415 2975
rect 151446 2972 151452 2984
rect 151403 2944 151452 2972
rect 151403 2941 151415 2944
rect 151357 2935 151415 2941
rect 151446 2932 151452 2944
rect 151504 2932 151510 2984
rect 151538 2932 151544 2984
rect 151596 2972 151602 2984
rect 156414 2972 156420 2984
rect 151596 2944 156420 2972
rect 151596 2932 151602 2944
rect 156414 2932 156420 2944
rect 156472 2932 156478 2984
rect 157429 2975 157487 2981
rect 157429 2941 157441 2975
rect 157475 2941 157487 2975
rect 157429 2935 157487 2941
rect 157613 2975 157671 2981
rect 157613 2941 157625 2975
rect 157659 2972 157671 2975
rect 161198 2972 161204 2984
rect 157659 2944 161204 2972
rect 157659 2941 157671 2944
rect 157613 2935 157671 2941
rect 137112 2876 137600 2904
rect 137664 2876 138612 2904
rect 125468 2808 127204 2836
rect 125468 2796 125474 2808
rect 128538 2796 128544 2848
rect 128596 2836 128602 2848
rect 137664 2836 137692 2876
rect 138658 2864 138664 2916
rect 138716 2904 138722 2916
rect 144362 2904 144368 2916
rect 138716 2876 144368 2904
rect 138716 2864 138722 2876
rect 144362 2864 144368 2876
rect 144420 2864 144426 2916
rect 144546 2864 144552 2916
rect 144604 2904 144610 2916
rect 144604 2876 145328 2904
rect 144604 2864 144610 2876
rect 128596 2808 137692 2836
rect 128596 2796 128602 2808
rect 137922 2796 137928 2848
rect 137980 2836 137986 2848
rect 138474 2836 138480 2848
rect 137980 2808 138480 2836
rect 137980 2796 137986 2808
rect 138474 2796 138480 2808
rect 138532 2796 138538 2848
rect 138566 2796 138572 2848
rect 138624 2836 138630 2848
rect 139397 2839 139455 2845
rect 139397 2836 139409 2839
rect 138624 2808 139409 2836
rect 138624 2796 138630 2808
rect 139397 2805 139409 2808
rect 139443 2805 139455 2839
rect 140406 2836 140412 2848
rect 140367 2808 140412 2836
rect 139397 2799 139455 2805
rect 140406 2796 140412 2808
rect 140464 2796 140470 2848
rect 141050 2796 141056 2848
rect 141108 2836 141114 2848
rect 141513 2839 141571 2845
rect 141513 2836 141525 2839
rect 141108 2808 141525 2836
rect 141108 2796 141114 2808
rect 141513 2805 141525 2808
rect 141559 2805 141571 2839
rect 141513 2799 141571 2805
rect 141786 2796 141792 2848
rect 141844 2836 141850 2848
rect 144454 2836 144460 2848
rect 141844 2808 144460 2836
rect 141844 2796 141850 2808
rect 144454 2796 144460 2808
rect 144512 2796 144518 2848
rect 145300 2836 145328 2876
rect 146110 2864 146116 2916
rect 146168 2904 146174 2916
rect 156138 2904 156144 2916
rect 146168 2876 156144 2904
rect 146168 2864 146174 2876
rect 156138 2864 156144 2876
rect 156196 2864 156202 2916
rect 156969 2907 157027 2913
rect 156969 2873 156981 2907
rect 157015 2873 157027 2907
rect 156969 2867 157027 2873
rect 157061 2907 157119 2913
rect 157061 2873 157073 2907
rect 157107 2904 157119 2907
rect 157337 2907 157395 2913
rect 157337 2904 157349 2907
rect 157107 2876 157349 2904
rect 157107 2873 157119 2876
rect 157061 2867 157119 2873
rect 157337 2873 157349 2876
rect 157383 2873 157395 2907
rect 157444 2904 157472 2935
rect 161198 2932 161204 2944
rect 161256 2932 161262 2984
rect 161293 2975 161351 2981
rect 161293 2941 161305 2975
rect 161339 2972 161351 2975
rect 162581 2975 162639 2981
rect 162581 2972 162593 2975
rect 161339 2944 162593 2972
rect 161339 2941 161351 2944
rect 161293 2935 161351 2941
rect 162581 2941 162593 2944
rect 162627 2941 162639 2975
rect 162581 2935 162639 2941
rect 162670 2932 162676 2984
rect 162728 2932 162734 2984
rect 162762 2932 162768 2984
rect 162820 2972 162826 2984
rect 162872 2972 162900 3012
rect 162820 2944 162900 2972
rect 162949 2975 163007 2981
rect 162820 2932 162826 2944
rect 162949 2941 162961 2975
rect 162995 2972 163007 2975
rect 166718 2972 166724 2984
rect 162995 2944 166724 2972
rect 162995 2941 163007 2944
rect 162949 2935 163007 2941
rect 166718 2932 166724 2944
rect 166776 2932 166782 2984
rect 164513 2907 164571 2913
rect 164513 2904 164525 2907
rect 157444 2876 164525 2904
rect 157337 2867 157395 2873
rect 164513 2873 164525 2876
rect 164559 2873 164571 2907
rect 166258 2904 166264 2916
rect 164513 2867 164571 2873
rect 164620 2876 166264 2904
rect 147030 2836 147036 2848
rect 145300 2808 147036 2836
rect 147030 2796 147036 2808
rect 147088 2796 147094 2848
rect 149238 2796 149244 2848
rect 149296 2836 149302 2848
rect 156877 2839 156935 2845
rect 156877 2836 156889 2839
rect 149296 2808 156889 2836
rect 149296 2796 149302 2808
rect 156877 2805 156889 2808
rect 156923 2805 156935 2839
rect 156984 2836 157012 2867
rect 157426 2836 157432 2848
rect 156984 2808 157432 2836
rect 156877 2799 156935 2805
rect 157426 2796 157432 2808
rect 157484 2796 157490 2848
rect 157521 2839 157579 2845
rect 157521 2805 157533 2839
rect 157567 2836 157579 2839
rect 158346 2836 158352 2848
rect 157567 2808 158352 2836
rect 157567 2805 157579 2808
rect 157521 2799 157579 2805
rect 158346 2796 158352 2808
rect 158404 2796 158410 2848
rect 158530 2796 158536 2848
rect 158588 2836 158594 2848
rect 161293 2839 161351 2845
rect 161293 2836 161305 2839
rect 158588 2808 161305 2836
rect 158588 2796 158594 2808
rect 161293 2805 161305 2808
rect 161339 2805 161351 2839
rect 161293 2799 161351 2805
rect 161474 2796 161480 2848
rect 161532 2836 161538 2848
rect 164620 2836 164648 2876
rect 166258 2864 166264 2876
rect 166316 2864 166322 2916
rect 167104 2904 167132 3012
rect 173802 2932 173808 2984
rect 173860 2972 173866 2984
rect 180150 2972 180156 2984
rect 173860 2944 180156 2972
rect 173860 2932 173866 2944
rect 180150 2932 180156 2944
rect 180208 2932 180214 2984
rect 180334 2932 180340 2984
rect 180392 2972 180398 2984
rect 187050 2972 187056 2984
rect 180392 2944 187056 2972
rect 180392 2932 180398 2944
rect 187050 2932 187056 2944
rect 187108 2932 187114 2984
rect 193582 2932 193588 2984
rect 193640 2972 193646 2984
rect 196894 2972 196900 2984
rect 193640 2944 196900 2972
rect 193640 2932 193646 2944
rect 196894 2932 196900 2944
rect 196952 2932 196958 2984
rect 171778 2904 171784 2916
rect 167104 2876 171784 2904
rect 171778 2864 171784 2876
rect 171836 2864 171842 2916
rect 176470 2864 176476 2916
rect 176528 2904 176534 2916
rect 176654 2904 176660 2916
rect 176528 2876 176660 2904
rect 176528 2864 176534 2876
rect 176654 2864 176660 2876
rect 176712 2864 176718 2916
rect 180426 2864 180432 2916
rect 180484 2904 180490 2916
rect 184198 2904 184204 2916
rect 180484 2876 184204 2904
rect 180484 2864 180490 2876
rect 184198 2864 184204 2876
rect 184256 2864 184262 2916
rect 195882 2864 195888 2916
rect 195940 2904 195946 2916
rect 199746 2904 199752 2916
rect 195940 2876 199752 2904
rect 195940 2864 195946 2876
rect 199746 2864 199752 2876
rect 199804 2864 199810 2916
rect 161532 2808 164648 2836
rect 164789 2839 164847 2845
rect 161532 2796 161538 2808
rect 164789 2805 164801 2839
rect 164835 2836 164847 2839
rect 165062 2836 165068 2848
rect 164835 2808 165068 2836
rect 164835 2805 164847 2808
rect 164789 2799 164847 2805
rect 165062 2796 165068 2808
rect 165120 2796 165126 2848
rect 165338 2796 165344 2848
rect 165396 2836 165402 2848
rect 167086 2836 167092 2848
rect 165396 2808 167092 2836
rect 165396 2796 165402 2808
rect 167086 2796 167092 2808
rect 167144 2796 167150 2848
rect 173342 2796 173348 2848
rect 173400 2836 173406 2848
rect 179230 2836 179236 2848
rect 173400 2808 179236 2836
rect 173400 2796 173406 2808
rect 179230 2796 179236 2808
rect 179288 2796 179294 2848
rect 190454 2796 190460 2848
rect 190512 2836 190518 2848
rect 192294 2836 192300 2848
rect 190512 2808 192300 2836
rect 190512 2796 190518 2808
rect 192294 2796 192300 2808
rect 192352 2796 192358 2848
rect 194686 2796 194692 2848
rect 194744 2836 194750 2848
rect 199286 2836 199292 2848
rect 194744 2808 199292 2836
rect 194744 2796 194750 2808
rect 199286 2796 199292 2808
rect 199344 2796 199350 2848
rect 1104 2746 198812 2768
rect 1104 2694 24078 2746
rect 24130 2694 64078 2746
rect 64130 2694 104078 2746
rect 104130 2694 144078 2746
rect 144130 2694 184078 2746
rect 184130 2694 198812 2746
rect 1104 2672 198812 2694
rect 6454 2592 6460 2644
rect 6512 2632 6518 2644
rect 6549 2635 6607 2641
rect 6549 2632 6561 2635
rect 6512 2604 6561 2632
rect 6512 2592 6518 2604
rect 6549 2601 6561 2604
rect 6595 2601 6607 2635
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 6549 2595 6607 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 8662 2632 8668 2644
rect 8619 2604 8668 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2632 11667 2635
rect 11698 2632 11704 2644
rect 11655 2604 11704 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 13906 2632 13912 2644
rect 13867 2604 13912 2632
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 15381 2635 15439 2641
rect 15381 2601 15393 2635
rect 15427 2632 15439 2635
rect 15930 2632 15936 2644
rect 15427 2604 15936 2632
rect 15427 2601 15439 2604
rect 15381 2595 15439 2601
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 17218 2632 17224 2644
rect 17179 2604 17224 2632
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 20993 2635 21051 2641
rect 20993 2632 21005 2635
rect 20772 2604 21005 2632
rect 20772 2592 20778 2604
rect 20993 2601 21005 2604
rect 21039 2601 21051 2635
rect 20993 2595 21051 2601
rect 22005 2635 22063 2641
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 22370 2632 22376 2644
rect 22051 2604 22376 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 22370 2592 22376 2604
rect 22428 2592 22434 2644
rect 23937 2635 23995 2641
rect 23937 2601 23949 2635
rect 23983 2632 23995 2635
rect 24854 2632 24860 2644
rect 23983 2604 24860 2632
rect 23983 2601 23995 2604
rect 23937 2595 23995 2601
rect 24854 2592 24860 2604
rect 24912 2592 24918 2644
rect 25130 2632 25136 2644
rect 25091 2604 25136 2632
rect 25130 2592 25136 2604
rect 25188 2592 25194 2644
rect 26605 2635 26663 2641
rect 26605 2601 26617 2635
rect 26651 2632 26663 2635
rect 27706 2632 27712 2644
rect 26651 2604 27712 2632
rect 26651 2601 26663 2604
rect 26605 2595 26663 2601
rect 27706 2592 27712 2604
rect 27764 2592 27770 2644
rect 33318 2632 33324 2644
rect 33279 2604 33324 2632
rect 33318 2592 33324 2604
rect 33376 2592 33382 2644
rect 35897 2635 35955 2641
rect 35897 2601 35909 2635
rect 35943 2632 35955 2635
rect 36538 2632 36544 2644
rect 35943 2604 36544 2632
rect 35943 2601 35955 2604
rect 35897 2595 35955 2601
rect 36538 2592 36544 2604
rect 36596 2592 36602 2644
rect 42337 2635 42395 2641
rect 42337 2601 42349 2635
rect 42383 2632 42395 2635
rect 43346 2632 43352 2644
rect 42383 2604 43352 2632
rect 42383 2601 42395 2604
rect 42337 2595 42395 2601
rect 43346 2592 43352 2604
rect 43404 2592 43410 2644
rect 44358 2592 44364 2644
rect 44416 2632 44422 2644
rect 44729 2635 44787 2641
rect 44729 2632 44741 2635
rect 44416 2604 44741 2632
rect 44416 2592 44422 2604
rect 44729 2601 44741 2604
rect 44775 2601 44787 2635
rect 44729 2595 44787 2601
rect 45554 2592 45560 2644
rect 45612 2632 45618 2644
rect 45741 2635 45799 2641
rect 45741 2632 45753 2635
rect 45612 2604 45753 2632
rect 45612 2592 45618 2604
rect 45741 2601 45753 2604
rect 45787 2601 45799 2635
rect 45741 2595 45799 2601
rect 46566 2592 46572 2644
rect 46624 2632 46630 2644
rect 46753 2635 46811 2641
rect 46753 2632 46765 2635
rect 46624 2604 46765 2632
rect 46624 2592 46630 2604
rect 46753 2601 46765 2604
rect 46799 2601 46811 2635
rect 47762 2632 47768 2644
rect 47723 2604 47768 2632
rect 46753 2595 46811 2601
rect 47762 2592 47768 2604
rect 47820 2592 47826 2644
rect 50433 2635 50491 2641
rect 50433 2601 50445 2635
rect 50479 2632 50491 2635
rect 51626 2632 51632 2644
rect 50479 2604 51632 2632
rect 50479 2601 50491 2604
rect 50433 2595 50491 2601
rect 51626 2592 51632 2604
rect 51684 2592 51690 2644
rect 51810 2632 51816 2644
rect 51771 2604 51816 2632
rect 51810 2592 51816 2604
rect 51868 2592 51874 2644
rect 52730 2592 52736 2644
rect 52788 2632 52794 2644
rect 52825 2635 52883 2641
rect 52825 2632 52837 2635
rect 52788 2604 52837 2632
rect 52788 2592 52794 2604
rect 52825 2601 52837 2604
rect 52871 2601 52883 2635
rect 54754 2632 54760 2644
rect 54715 2604 54760 2632
rect 52825 2595 52883 2601
rect 54754 2592 54760 2604
rect 54812 2592 54818 2644
rect 55214 2592 55220 2644
rect 55272 2632 55278 2644
rect 55674 2632 55680 2644
rect 55272 2604 55680 2632
rect 55272 2592 55278 2604
rect 55674 2592 55680 2604
rect 55732 2592 55738 2644
rect 55769 2635 55827 2641
rect 55769 2601 55781 2635
rect 55815 2632 55827 2635
rect 59446 2632 59452 2644
rect 55815 2604 59452 2632
rect 55815 2601 55827 2604
rect 55769 2595 55827 2601
rect 59446 2592 59452 2604
rect 59504 2592 59510 2644
rect 75270 2592 75276 2644
rect 75328 2632 75334 2644
rect 75457 2635 75515 2641
rect 75457 2632 75469 2635
rect 75328 2604 75469 2632
rect 75328 2592 75334 2604
rect 75457 2601 75469 2604
rect 75503 2601 75515 2635
rect 75457 2595 75515 2601
rect 83001 2635 83059 2641
rect 83001 2601 83013 2635
rect 83047 2632 83059 2635
rect 83090 2632 83096 2644
rect 83047 2604 83096 2632
rect 83047 2601 83059 2604
rect 83001 2595 83059 2601
rect 83090 2592 83096 2604
rect 83148 2592 83154 2644
rect 88245 2635 88303 2641
rect 88245 2601 88257 2635
rect 88291 2632 88303 2635
rect 88334 2632 88340 2644
rect 88291 2604 88340 2632
rect 88291 2601 88303 2604
rect 88245 2595 88303 2601
rect 88334 2592 88340 2604
rect 88392 2592 88398 2644
rect 92569 2635 92627 2641
rect 92569 2601 92581 2635
rect 92615 2632 92627 2635
rect 92934 2632 92940 2644
rect 92615 2604 92940 2632
rect 92615 2601 92627 2604
rect 92569 2595 92627 2601
rect 92934 2592 92940 2604
rect 92992 2592 92998 2644
rect 103057 2635 103115 2641
rect 94516 2604 101812 2632
rect 34514 2524 34520 2576
rect 34572 2564 34578 2576
rect 37921 2567 37979 2573
rect 37921 2564 37933 2567
rect 34572 2536 37933 2564
rect 34572 2524 34578 2536
rect 37921 2533 37933 2536
rect 37967 2533 37979 2567
rect 37921 2527 37979 2533
rect 43441 2567 43499 2573
rect 43441 2533 43453 2567
rect 43487 2564 43499 2567
rect 47578 2564 47584 2576
rect 43487 2536 47584 2564
rect 43487 2533 43499 2536
rect 43441 2527 43499 2533
rect 47578 2524 47584 2536
rect 47636 2524 47642 2576
rect 62022 2524 62028 2576
rect 62080 2564 62086 2576
rect 69658 2564 69664 2576
rect 62080 2536 69664 2564
rect 62080 2524 62086 2536
rect 69658 2524 69664 2536
rect 69716 2524 69722 2576
rect 85942 2524 85948 2576
rect 86000 2564 86006 2576
rect 86000 2536 89576 2564
rect 86000 2524 86006 2536
rect 1026 2456 1032 2508
rect 1084 2496 1090 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 1084 2468 5457 2496
rect 1084 2456 1090 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 5445 2459 5503 2465
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6457 2499 6515 2505
rect 6457 2496 6469 2499
rect 5868 2468 6469 2496
rect 5868 2456 5874 2468
rect 6457 2465 6469 2468
rect 6503 2465 6515 2499
rect 6457 2459 6515 2465
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 6788 2468 7481 2496
rect 6788 2456 6794 2468
rect 7469 2465 7481 2468
rect 7515 2465 7527 2499
rect 7469 2459 7527 2465
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8076 2468 8493 2496
rect 8076 2456 8082 2468
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 10594 2456 10600 2508
rect 10652 2496 10658 2508
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 10652 2468 11529 2496
rect 10652 2456 10658 2468
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11517 2459 11575 2465
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 12860 2468 13829 2496
rect 12860 2456 12866 2468
rect 13817 2465 13829 2468
rect 13863 2465 13875 2499
rect 13817 2459 13875 2465
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 17121 2499 17179 2505
rect 17121 2465 17133 2499
rect 17167 2465 17179 2499
rect 17121 2459 17179 2465
rect 13630 2388 13636 2440
rect 13688 2428 13694 2440
rect 15304 2428 15332 2459
rect 13688 2400 15332 2428
rect 13688 2388 13694 2400
rect 5537 2363 5595 2369
rect 5537 2329 5549 2363
rect 5583 2360 5595 2363
rect 12986 2360 12992 2372
rect 5583 2332 12992 2360
rect 5583 2329 5595 2332
rect 5537 2323 5595 2329
rect 12986 2320 12992 2332
rect 13044 2320 13050 2372
rect 15010 2320 15016 2372
rect 15068 2360 15074 2372
rect 17144 2360 17172 2459
rect 17218 2456 17224 2508
rect 17276 2496 17282 2508
rect 20901 2499 20959 2505
rect 20901 2496 20913 2499
rect 17276 2468 20913 2496
rect 17276 2456 17282 2468
rect 20901 2465 20913 2468
rect 20947 2465 20959 2499
rect 20901 2459 20959 2465
rect 21913 2499 21971 2505
rect 21913 2465 21925 2499
rect 21959 2465 21971 2499
rect 21913 2459 21971 2465
rect 20162 2388 20168 2440
rect 20220 2428 20226 2440
rect 21928 2428 21956 2459
rect 23290 2456 23296 2508
rect 23348 2496 23354 2508
rect 23845 2499 23903 2505
rect 23845 2496 23857 2499
rect 23348 2468 23857 2496
rect 23348 2456 23354 2468
rect 23845 2465 23857 2468
rect 23891 2465 23903 2499
rect 23845 2459 23903 2465
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24268 2468 25053 2496
rect 24268 2456 24274 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 25130 2456 25136 2508
rect 25188 2496 25194 2508
rect 26513 2499 26571 2505
rect 26513 2496 26525 2499
rect 25188 2468 26525 2496
rect 25188 2456 25194 2468
rect 26513 2465 26525 2468
rect 26559 2465 26571 2499
rect 26513 2459 26571 2465
rect 28442 2456 28448 2508
rect 28500 2496 28506 2508
rect 33229 2499 33287 2505
rect 33229 2496 33241 2499
rect 28500 2468 33241 2496
rect 28500 2456 28506 2468
rect 33229 2465 33241 2468
rect 33275 2465 33287 2499
rect 33229 2459 33287 2465
rect 33686 2456 33692 2508
rect 33744 2496 33750 2508
rect 35805 2499 35863 2505
rect 35805 2496 35817 2499
rect 33744 2468 35817 2496
rect 33744 2456 33750 2468
rect 35805 2465 35817 2468
rect 35851 2465 35863 2499
rect 35805 2459 35863 2465
rect 37829 2499 37887 2505
rect 37829 2465 37841 2499
rect 37875 2465 37887 2499
rect 37829 2459 37887 2465
rect 42245 2499 42303 2505
rect 42245 2465 42257 2499
rect 42291 2496 42303 2499
rect 43254 2496 43260 2508
rect 42291 2468 43260 2496
rect 42291 2465 42303 2468
rect 42245 2459 42303 2465
rect 20220 2400 21956 2428
rect 20220 2388 20226 2400
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 37844 2428 37872 2459
rect 43254 2456 43260 2468
rect 43312 2456 43318 2508
rect 43349 2499 43407 2505
rect 43349 2465 43361 2499
rect 43395 2465 43407 2499
rect 43349 2459 43407 2465
rect 44637 2499 44695 2505
rect 44637 2465 44649 2499
rect 44683 2465 44695 2499
rect 45646 2496 45652 2508
rect 45607 2468 45652 2496
rect 44637 2459 44695 2465
rect 34204 2400 37872 2428
rect 34204 2388 34210 2400
rect 38930 2388 38936 2440
rect 38988 2428 38994 2440
rect 43364 2428 43392 2459
rect 38988 2400 43392 2428
rect 38988 2388 38994 2400
rect 15068 2332 17172 2360
rect 15068 2320 15074 2332
rect 40218 2320 40224 2372
rect 40276 2360 40282 2372
rect 44652 2360 44680 2459
rect 45646 2456 45652 2468
rect 45704 2456 45710 2508
rect 46661 2499 46719 2505
rect 46661 2465 46673 2499
rect 46707 2465 46719 2499
rect 46661 2459 46719 2465
rect 47673 2499 47731 2505
rect 47673 2465 47685 2499
rect 47719 2496 47731 2499
rect 48130 2496 48136 2508
rect 47719 2468 48136 2496
rect 47719 2465 47731 2468
rect 47673 2459 47731 2465
rect 45462 2388 45468 2440
rect 45520 2428 45526 2440
rect 46676 2428 46704 2459
rect 48130 2456 48136 2468
rect 48188 2456 48194 2508
rect 48498 2456 48504 2508
rect 48556 2496 48562 2508
rect 50341 2499 50399 2505
rect 50341 2496 50353 2499
rect 48556 2468 50353 2496
rect 48556 2456 48562 2468
rect 50341 2465 50353 2468
rect 50387 2465 50399 2499
rect 50341 2459 50399 2465
rect 51721 2499 51779 2505
rect 51721 2465 51733 2499
rect 51767 2465 51779 2499
rect 51721 2459 51779 2465
rect 52733 2499 52791 2505
rect 52733 2465 52745 2499
rect 52779 2465 52791 2499
rect 54662 2496 54668 2508
rect 54623 2468 54668 2496
rect 52733 2459 52791 2465
rect 45520 2400 46704 2428
rect 45520 2388 45526 2400
rect 49786 2388 49792 2440
rect 49844 2428 49850 2440
rect 51736 2428 51764 2459
rect 49844 2400 51764 2428
rect 49844 2388 49850 2400
rect 40276 2332 44680 2360
rect 40276 2320 40282 2332
rect 50246 2320 50252 2372
rect 50304 2360 50310 2372
rect 52748 2360 52776 2459
rect 54662 2456 54668 2468
rect 54720 2456 54726 2508
rect 55490 2456 55496 2508
rect 55548 2496 55554 2508
rect 55677 2499 55735 2505
rect 55677 2496 55689 2499
rect 55548 2468 55689 2496
rect 55548 2456 55554 2468
rect 55677 2465 55689 2468
rect 55723 2465 55735 2499
rect 55677 2459 55735 2465
rect 57793 2499 57851 2505
rect 57793 2465 57805 2499
rect 57839 2496 57851 2499
rect 57974 2496 57980 2508
rect 57839 2468 57980 2496
rect 57839 2465 57851 2468
rect 57793 2459 57851 2465
rect 57974 2456 57980 2468
rect 58032 2456 58038 2508
rect 60550 2456 60556 2508
rect 60608 2496 60614 2508
rect 60645 2499 60703 2505
rect 60645 2496 60657 2499
rect 60608 2468 60657 2496
rect 60608 2456 60614 2468
rect 60645 2465 60657 2468
rect 60691 2465 60703 2499
rect 63402 2496 63408 2508
rect 63363 2468 63408 2496
rect 60645 2459 60703 2465
rect 63402 2456 63408 2468
rect 63460 2456 63466 2508
rect 67085 2499 67143 2505
rect 67085 2465 67097 2499
rect 67131 2496 67143 2499
rect 67634 2496 67640 2508
rect 67131 2468 67640 2496
rect 67131 2465 67143 2468
rect 67085 2459 67143 2465
rect 67634 2456 67640 2468
rect 67692 2456 67698 2508
rect 68649 2499 68707 2505
rect 68649 2465 68661 2499
rect 68695 2496 68707 2499
rect 68738 2496 68744 2508
rect 68695 2468 68744 2496
rect 68695 2465 68707 2468
rect 68649 2459 68707 2465
rect 68738 2456 68744 2468
rect 68796 2456 68802 2508
rect 70305 2499 70363 2505
rect 70305 2465 70317 2499
rect 70351 2496 70363 2499
rect 71498 2496 71504 2508
rect 70351 2468 71504 2496
rect 70351 2465 70363 2468
rect 70305 2459 70363 2465
rect 71498 2456 71504 2468
rect 71556 2456 71562 2508
rect 72697 2499 72755 2505
rect 72697 2465 72709 2499
rect 72743 2496 72755 2499
rect 73154 2496 73160 2508
rect 72743 2468 73160 2496
rect 72743 2465 72755 2468
rect 72697 2459 72755 2465
rect 73154 2456 73160 2468
rect 73212 2456 73218 2508
rect 74445 2499 74503 2505
rect 74445 2465 74457 2499
rect 74491 2496 74503 2499
rect 74534 2496 74540 2508
rect 74491 2468 74540 2496
rect 74491 2465 74503 2468
rect 74445 2459 74503 2465
rect 74534 2456 74540 2468
rect 74592 2456 74598 2508
rect 77294 2496 77300 2508
rect 77255 2468 77300 2496
rect 77294 2456 77300 2468
rect 77352 2456 77358 2508
rect 78490 2456 78496 2508
rect 78548 2496 78554 2508
rect 78769 2499 78827 2505
rect 78769 2496 78781 2499
rect 78548 2468 78781 2496
rect 78548 2456 78554 2468
rect 78769 2465 78781 2468
rect 78815 2465 78827 2499
rect 80698 2496 80704 2508
rect 80659 2468 80704 2496
rect 78769 2459 78827 2465
rect 80698 2456 80704 2468
rect 80756 2456 80762 2508
rect 81526 2456 81532 2508
rect 81584 2496 81590 2508
rect 84105 2499 84163 2505
rect 84105 2496 84117 2499
rect 81584 2468 84117 2496
rect 81584 2456 81590 2468
rect 84105 2465 84117 2468
rect 84151 2465 84163 2499
rect 84105 2459 84163 2465
rect 85298 2456 85304 2508
rect 85356 2496 85362 2508
rect 89548 2505 89576 2536
rect 89622 2524 89628 2576
rect 89680 2564 89686 2576
rect 94516 2564 94544 2604
rect 95050 2564 95056 2576
rect 89680 2536 94544 2564
rect 94608 2536 95056 2564
rect 89680 2524 89686 2536
rect 86221 2499 86279 2505
rect 86221 2496 86233 2499
rect 85356 2468 86233 2496
rect 85356 2456 85362 2468
rect 86221 2465 86233 2468
rect 86267 2465 86279 2499
rect 86221 2459 86279 2465
rect 89533 2499 89591 2505
rect 89533 2465 89545 2499
rect 89579 2465 89591 2499
rect 89533 2459 89591 2465
rect 90082 2456 90088 2508
rect 90140 2496 90146 2508
rect 91097 2499 91155 2505
rect 91097 2496 91109 2499
rect 90140 2468 91109 2496
rect 90140 2456 90146 2468
rect 91097 2465 91109 2468
rect 91143 2465 91155 2499
rect 94608 2496 94636 2536
rect 95050 2524 95056 2536
rect 95108 2524 95114 2576
rect 95237 2567 95295 2573
rect 95237 2533 95249 2567
rect 95283 2564 95295 2567
rect 95878 2564 95884 2576
rect 95283 2536 95884 2564
rect 95283 2533 95295 2536
rect 95237 2527 95295 2533
rect 95878 2524 95884 2536
rect 95936 2524 95942 2576
rect 96065 2567 96123 2573
rect 96065 2533 96077 2567
rect 96111 2564 96123 2567
rect 96338 2564 96344 2576
rect 96111 2536 96344 2564
rect 96111 2533 96123 2536
rect 96065 2527 96123 2533
rect 96338 2524 96344 2536
rect 96396 2524 96402 2576
rect 97813 2567 97871 2573
rect 97813 2533 97825 2567
rect 97859 2564 97871 2567
rect 99926 2564 99932 2576
rect 97859 2536 99932 2564
rect 97859 2533 97871 2536
rect 97813 2527 97871 2533
rect 99926 2524 99932 2536
rect 99984 2524 99990 2576
rect 101784 2564 101812 2604
rect 103057 2601 103069 2635
rect 103103 2632 103115 2635
rect 110414 2632 110420 2644
rect 103103 2604 110420 2632
rect 103103 2601 103115 2604
rect 103057 2595 103115 2601
rect 110414 2592 110420 2604
rect 110472 2592 110478 2644
rect 110506 2592 110512 2644
rect 110564 2632 110570 2644
rect 114186 2632 114192 2644
rect 110564 2604 113312 2632
rect 114147 2604 114192 2632
rect 110564 2592 110570 2604
rect 104250 2564 104256 2576
rect 101784 2536 104256 2564
rect 104250 2524 104256 2536
rect 104308 2524 104314 2576
rect 105538 2524 105544 2576
rect 105596 2564 105602 2576
rect 109494 2564 109500 2576
rect 105596 2536 109500 2564
rect 105596 2524 105602 2536
rect 109494 2524 109500 2536
rect 109552 2524 109558 2576
rect 111886 2564 111892 2576
rect 109604 2536 111892 2564
rect 94866 2496 94872 2508
rect 91097 2459 91155 2465
rect 91204 2468 94636 2496
rect 94827 2468 94872 2496
rect 56318 2388 56324 2440
rect 56376 2428 56382 2440
rect 57149 2431 57207 2437
rect 57149 2428 57161 2431
rect 56376 2400 57161 2428
rect 56376 2388 56382 2400
rect 57149 2397 57161 2400
rect 57195 2397 57207 2431
rect 57149 2391 57207 2397
rect 57330 2388 57336 2440
rect 57388 2428 57394 2440
rect 62206 2428 62212 2440
rect 57388 2400 62212 2428
rect 57388 2388 57394 2400
rect 62206 2388 62212 2400
rect 62264 2388 62270 2440
rect 64598 2388 64604 2440
rect 64656 2428 64662 2440
rect 66441 2431 66499 2437
rect 66441 2428 66453 2431
rect 64656 2400 66453 2428
rect 64656 2388 64662 2400
rect 66441 2397 66453 2400
rect 66487 2397 66499 2431
rect 66441 2391 66499 2397
rect 66806 2388 66812 2440
rect 66864 2428 66870 2440
rect 68005 2431 68063 2437
rect 68005 2428 68017 2431
rect 66864 2400 68017 2428
rect 66864 2388 66870 2400
rect 68005 2397 68017 2400
rect 68051 2397 68063 2431
rect 68005 2391 68063 2397
rect 68094 2388 68100 2440
rect 68152 2428 68158 2440
rect 69753 2431 69811 2437
rect 69753 2428 69765 2431
rect 68152 2400 69765 2428
rect 68152 2388 68158 2400
rect 69753 2397 69765 2400
rect 69799 2397 69811 2431
rect 69753 2391 69811 2397
rect 71222 2388 71228 2440
rect 71280 2428 71286 2440
rect 72053 2431 72111 2437
rect 72053 2428 72065 2431
rect 71280 2400 72065 2428
rect 71280 2388 71286 2400
rect 72053 2397 72065 2400
rect 72099 2397 72111 2431
rect 72053 2391 72111 2397
rect 72142 2388 72148 2440
rect 72200 2428 72206 2440
rect 73893 2431 73951 2437
rect 73893 2428 73905 2431
rect 72200 2400 73905 2428
rect 72200 2388 72206 2400
rect 73893 2397 73905 2400
rect 73939 2397 73951 2431
rect 73893 2391 73951 2397
rect 76006 2388 76012 2440
rect 76064 2428 76070 2440
rect 77113 2431 77171 2437
rect 77113 2428 77125 2431
rect 76064 2400 77125 2428
rect 76064 2388 76070 2400
rect 77113 2397 77125 2400
rect 77159 2397 77171 2431
rect 77113 2391 77171 2397
rect 78582 2388 78588 2440
rect 78640 2428 78646 2440
rect 78677 2431 78735 2437
rect 78677 2428 78689 2431
rect 78640 2400 78689 2428
rect 78640 2388 78646 2400
rect 78677 2397 78689 2400
rect 78723 2397 78735 2431
rect 78677 2391 78735 2397
rect 79502 2388 79508 2440
rect 79560 2428 79566 2440
rect 80241 2431 80299 2437
rect 80241 2428 80253 2431
rect 79560 2400 80253 2428
rect 79560 2388 79566 2400
rect 80241 2397 80253 2400
rect 80287 2397 80299 2431
rect 80241 2391 80299 2397
rect 82538 2388 82544 2440
rect 82596 2428 82602 2440
rect 84013 2431 84071 2437
rect 84013 2428 84025 2431
rect 82596 2400 84025 2428
rect 82596 2388 82602 2400
rect 84013 2397 84025 2400
rect 84059 2397 84071 2431
rect 84013 2391 84071 2397
rect 86865 2431 86923 2437
rect 86865 2397 86877 2431
rect 86911 2428 86923 2431
rect 88610 2428 88616 2440
rect 86911 2400 88616 2428
rect 86911 2397 86923 2400
rect 86865 2391 86923 2397
rect 88610 2388 88616 2400
rect 88668 2388 88674 2440
rect 89070 2388 89076 2440
rect 89128 2428 89134 2440
rect 89441 2431 89499 2437
rect 89441 2428 89453 2431
rect 89128 2400 89453 2428
rect 89128 2388 89134 2400
rect 89441 2397 89453 2400
rect 89487 2397 89499 2431
rect 89441 2391 89499 2397
rect 89714 2388 89720 2440
rect 89772 2428 89778 2440
rect 91204 2428 91232 2468
rect 94866 2456 94872 2468
rect 94924 2456 94930 2508
rect 97258 2496 97264 2508
rect 97219 2468 97264 2496
rect 97258 2456 97264 2468
rect 97316 2456 97322 2508
rect 98086 2456 98092 2508
rect 98144 2496 98150 2508
rect 99561 2499 99619 2505
rect 99561 2496 99573 2499
rect 98144 2468 99573 2496
rect 98144 2456 98150 2468
rect 99561 2465 99573 2468
rect 99607 2465 99619 2499
rect 99561 2459 99619 2465
rect 101677 2499 101735 2505
rect 101677 2465 101689 2499
rect 101723 2496 101735 2499
rect 103241 2499 103299 2505
rect 101723 2468 102732 2496
rect 101723 2465 101735 2468
rect 101677 2459 101735 2465
rect 89772 2400 91232 2428
rect 91741 2431 91799 2437
rect 89772 2388 89778 2400
rect 91741 2397 91753 2431
rect 91787 2428 91799 2431
rect 92566 2428 92572 2440
rect 91787 2400 92572 2428
rect 91787 2397 91799 2400
rect 91741 2391 91799 2397
rect 92566 2388 92572 2400
rect 92624 2388 92630 2440
rect 92750 2388 92756 2440
rect 92808 2428 92814 2440
rect 92808 2400 94636 2428
rect 92808 2388 92814 2400
rect 50304 2332 52776 2360
rect 50304 2320 50310 2332
rect 60458 2320 60464 2372
rect 60516 2360 60522 2372
rect 94498 2360 94504 2372
rect 60516 2332 94504 2360
rect 60516 2320 60522 2332
rect 94498 2320 94504 2332
rect 94556 2320 94562 2372
rect 94608 2360 94636 2400
rect 95234 2388 95240 2440
rect 95292 2428 95298 2440
rect 95292 2400 99052 2428
rect 95292 2388 95298 2400
rect 97902 2360 97908 2372
rect 94608 2332 97908 2360
rect 97902 2320 97908 2332
rect 97960 2320 97966 2372
rect 54846 2252 54852 2304
rect 54904 2292 54910 2304
rect 56594 2292 56600 2304
rect 54904 2264 56600 2292
rect 54904 2252 54910 2264
rect 56594 2252 56600 2264
rect 56652 2252 56658 2304
rect 59446 2252 59452 2304
rect 59504 2292 59510 2304
rect 60829 2295 60887 2301
rect 60829 2292 60841 2295
rect 59504 2264 60841 2292
rect 59504 2252 59510 2264
rect 60829 2261 60841 2264
rect 60875 2261 60887 2295
rect 60829 2255 60887 2261
rect 63221 2295 63279 2301
rect 63221 2261 63233 2295
rect 63267 2292 63279 2295
rect 63310 2292 63316 2304
rect 63267 2264 63316 2292
rect 63267 2261 63279 2264
rect 63221 2255 63279 2261
rect 63310 2252 63316 2264
rect 63368 2252 63374 2304
rect 81066 2252 81072 2304
rect 81124 2292 81130 2304
rect 98270 2292 98276 2304
rect 81124 2264 98276 2292
rect 81124 2252 81130 2264
rect 98270 2252 98276 2264
rect 98328 2252 98334 2304
rect 99024 2292 99052 2400
rect 99098 2388 99104 2440
rect 99156 2428 99162 2440
rect 99469 2431 99527 2437
rect 99469 2428 99481 2431
rect 99156 2400 99481 2428
rect 99156 2388 99162 2400
rect 99469 2397 99481 2400
rect 99515 2397 99527 2431
rect 99469 2391 99527 2397
rect 101769 2431 101827 2437
rect 101769 2397 101781 2431
rect 101815 2428 101827 2431
rect 102594 2428 102600 2440
rect 101815 2400 102600 2428
rect 101815 2397 101827 2400
rect 101769 2391 101827 2397
rect 102594 2388 102600 2400
rect 102652 2388 102658 2440
rect 102704 2428 102732 2468
rect 103241 2465 103253 2499
rect 103287 2496 103299 2499
rect 103514 2496 103520 2508
rect 103287 2468 103520 2496
rect 103287 2465 103299 2468
rect 103241 2459 103299 2465
rect 103514 2456 103520 2468
rect 103572 2456 103578 2508
rect 105173 2499 105231 2505
rect 105173 2465 105185 2499
rect 105219 2465 105231 2499
rect 105173 2459 105231 2465
rect 104342 2428 104348 2440
rect 102704 2400 104348 2428
rect 104342 2388 104348 2400
rect 104400 2388 104406 2440
rect 105188 2428 105216 2459
rect 106458 2456 106464 2508
rect 106516 2496 106522 2508
rect 109604 2505 109632 2536
rect 111886 2524 111892 2536
rect 111944 2524 111950 2576
rect 113284 2564 113312 2604
rect 114186 2592 114192 2604
rect 114244 2592 114250 2644
rect 117225 2635 117283 2641
rect 117225 2632 117237 2635
rect 114296 2604 117237 2632
rect 114296 2564 114324 2604
rect 117225 2601 117237 2604
rect 117271 2601 117283 2635
rect 118234 2632 118240 2644
rect 118195 2604 118240 2632
rect 117225 2595 117283 2601
rect 118234 2592 118240 2604
rect 118292 2592 118298 2644
rect 118970 2592 118976 2644
rect 119028 2632 119034 2644
rect 122009 2635 122067 2641
rect 122009 2632 122021 2635
rect 119028 2604 122021 2632
rect 119028 2592 119034 2604
rect 122009 2601 122021 2604
rect 122055 2601 122067 2635
rect 122009 2595 122067 2601
rect 123662 2592 123668 2644
rect 123720 2632 123726 2644
rect 123757 2635 123815 2641
rect 123757 2632 123769 2635
rect 123720 2604 123769 2632
rect 123720 2592 123726 2604
rect 123757 2601 123769 2604
rect 123803 2601 123815 2635
rect 125594 2632 125600 2644
rect 123757 2595 123815 2601
rect 124508 2604 125600 2632
rect 115198 2564 115204 2576
rect 113284 2536 114324 2564
rect 115159 2536 115204 2564
rect 115198 2524 115204 2536
rect 115256 2524 115262 2576
rect 124306 2564 124312 2576
rect 117056 2536 117452 2564
rect 106553 2499 106611 2505
rect 106553 2496 106565 2499
rect 106516 2468 106565 2496
rect 106516 2456 106522 2468
rect 106553 2465 106565 2468
rect 106599 2465 106611 2499
rect 106553 2459 106611 2465
rect 109589 2499 109647 2505
rect 109589 2465 109601 2499
rect 109635 2465 109647 2499
rect 109589 2459 109647 2465
rect 110598 2456 110604 2508
rect 110656 2496 110662 2508
rect 110785 2499 110843 2505
rect 110785 2496 110797 2499
rect 110656 2468 110797 2496
rect 110656 2456 110662 2468
rect 110785 2465 110797 2468
rect 110831 2465 110843 2499
rect 110785 2459 110843 2465
rect 112257 2499 112315 2505
rect 112257 2465 112269 2499
rect 112303 2496 112315 2499
rect 114097 2499 114155 2505
rect 112303 2468 113128 2496
rect 112303 2465 112315 2468
rect 112257 2459 112315 2465
rect 107197 2431 107255 2437
rect 105188 2400 107148 2428
rect 105265 2363 105323 2369
rect 105265 2360 105277 2363
rect 99760 2332 105277 2360
rect 99760 2292 99788 2332
rect 105265 2329 105277 2332
rect 105311 2329 105323 2363
rect 107120 2360 107148 2400
rect 107197 2397 107209 2431
rect 107243 2428 107255 2431
rect 108666 2428 108672 2440
rect 107243 2400 108672 2428
rect 107243 2397 107255 2400
rect 107197 2391 107255 2397
rect 108666 2388 108672 2400
rect 108724 2388 108730 2440
rect 108850 2388 108856 2440
rect 108908 2428 108914 2440
rect 108908 2400 109172 2428
rect 108908 2388 108914 2400
rect 109034 2360 109040 2372
rect 107120 2332 109040 2360
rect 105265 2323 105323 2329
rect 109034 2320 109040 2332
rect 109092 2320 109098 2372
rect 109144 2360 109172 2400
rect 109218 2388 109224 2440
rect 109276 2428 109282 2440
rect 110046 2428 110052 2440
rect 109276 2400 110052 2428
rect 109276 2388 109282 2400
rect 110046 2388 110052 2400
rect 110104 2388 110110 2440
rect 112346 2428 112352 2440
rect 112307 2400 112352 2428
rect 112346 2388 112352 2400
rect 112404 2388 112410 2440
rect 113100 2428 113128 2468
rect 114097 2465 114109 2499
rect 114143 2465 114155 2499
rect 114097 2459 114155 2465
rect 115109 2499 115167 2505
rect 115109 2465 115121 2499
rect 115155 2496 115167 2499
rect 116854 2496 116860 2508
rect 115155 2468 116860 2496
rect 115155 2465 115167 2468
rect 115109 2459 115167 2465
rect 113818 2428 113824 2440
rect 113100 2400 113824 2428
rect 113818 2388 113824 2400
rect 113876 2388 113882 2440
rect 114112 2428 114140 2459
rect 116854 2456 116860 2468
rect 116912 2456 116918 2508
rect 117056 2428 117084 2536
rect 117130 2456 117136 2508
rect 117188 2496 117194 2508
rect 117424 2496 117452 2536
rect 123588 2536 124312 2564
rect 117866 2496 117872 2508
rect 117188 2468 117233 2496
rect 117424 2468 117872 2496
rect 117188 2456 117194 2468
rect 117866 2456 117872 2468
rect 117924 2456 117930 2508
rect 118142 2496 118148 2508
rect 118103 2468 118148 2496
rect 118142 2456 118148 2468
rect 118200 2456 118206 2508
rect 119157 2499 119215 2505
rect 119157 2465 119169 2499
rect 119203 2465 119215 2499
rect 120166 2496 120172 2508
rect 120127 2468 120172 2496
rect 119157 2459 119215 2465
rect 114112 2400 117084 2428
rect 119172 2428 119200 2459
rect 120166 2456 120172 2468
rect 120224 2496 120230 2508
rect 120261 2499 120319 2505
rect 120261 2496 120273 2499
rect 120224 2468 120273 2496
rect 120224 2456 120230 2468
rect 120261 2465 120273 2468
rect 120307 2465 120319 2499
rect 120261 2459 120319 2465
rect 121917 2499 121975 2505
rect 121917 2465 121929 2499
rect 121963 2496 121975 2499
rect 123588 2496 123616 2536
rect 124306 2524 124312 2536
rect 124364 2524 124370 2576
rect 121963 2468 123616 2496
rect 123665 2499 123723 2505
rect 121963 2465 121975 2468
rect 121917 2459 121975 2465
rect 123665 2465 123677 2499
rect 123711 2496 123723 2499
rect 124508 2496 124536 2604
rect 125594 2592 125600 2604
rect 125652 2592 125658 2644
rect 125778 2632 125784 2644
rect 125739 2604 125784 2632
rect 125778 2592 125784 2604
rect 125836 2592 125842 2644
rect 126974 2632 126980 2644
rect 125888 2604 126980 2632
rect 124769 2567 124827 2573
rect 124769 2533 124781 2567
rect 124815 2564 124827 2567
rect 125888 2564 125916 2604
rect 126974 2592 126980 2604
rect 127032 2592 127038 2644
rect 128633 2635 128691 2641
rect 128633 2601 128645 2635
rect 128679 2632 128691 2635
rect 129550 2632 129556 2644
rect 128679 2604 129556 2632
rect 128679 2601 128691 2604
rect 128633 2595 128691 2601
rect 129550 2592 129556 2604
rect 129608 2592 129614 2644
rect 129918 2592 129924 2644
rect 129976 2632 129982 2644
rect 131666 2632 131672 2644
rect 129976 2604 131672 2632
rect 129976 2592 129982 2604
rect 131666 2592 131672 2604
rect 131724 2592 131730 2644
rect 131945 2635 132003 2641
rect 131945 2601 131957 2635
rect 131991 2632 132003 2635
rect 132126 2632 132132 2644
rect 131991 2604 132132 2632
rect 131991 2601 132003 2604
rect 131945 2595 132003 2601
rect 132126 2592 132132 2604
rect 132184 2592 132190 2644
rect 132586 2592 132592 2644
rect 132644 2632 132650 2644
rect 133782 2632 133788 2644
rect 132644 2604 133788 2632
rect 132644 2592 132650 2604
rect 133782 2592 133788 2604
rect 133840 2592 133846 2644
rect 133884 2604 134748 2632
rect 124815 2536 125916 2564
rect 127636 2536 127940 2564
rect 124815 2533 124827 2536
rect 124769 2527 124827 2533
rect 123711 2468 124536 2496
rect 124585 2499 124643 2505
rect 123711 2465 123723 2468
rect 123665 2459 123723 2465
rect 124585 2465 124597 2499
rect 124631 2496 124643 2499
rect 124674 2496 124680 2508
rect 124631 2468 124680 2496
rect 124631 2465 124643 2468
rect 124585 2459 124643 2465
rect 124674 2456 124680 2468
rect 124732 2456 124738 2508
rect 125597 2499 125655 2505
rect 125597 2465 125609 2499
rect 125643 2496 125655 2499
rect 125686 2496 125692 2508
rect 125643 2468 125692 2496
rect 125643 2465 125655 2468
rect 125597 2459 125655 2465
rect 125686 2456 125692 2468
rect 125744 2456 125750 2508
rect 127529 2499 127587 2505
rect 127529 2465 127541 2499
rect 127575 2496 127587 2499
rect 127636 2496 127664 2536
rect 127575 2468 127664 2496
rect 127912 2496 127940 2536
rect 128170 2524 128176 2576
rect 128228 2564 128234 2576
rect 132218 2564 132224 2576
rect 128228 2536 132224 2564
rect 128228 2524 128234 2536
rect 132218 2524 132224 2536
rect 132276 2524 132282 2576
rect 132310 2524 132316 2576
rect 132368 2564 132374 2576
rect 133884 2564 133912 2604
rect 132368 2536 133912 2564
rect 134720 2564 134748 2604
rect 134794 2592 134800 2644
rect 134852 2632 134858 2644
rect 138658 2632 138664 2644
rect 134852 2604 138664 2632
rect 134852 2592 134858 2604
rect 138658 2592 138664 2604
rect 138716 2592 138722 2644
rect 138750 2592 138756 2644
rect 138808 2632 138814 2644
rect 138845 2635 138903 2641
rect 138845 2632 138857 2635
rect 138808 2604 138857 2632
rect 138808 2592 138814 2604
rect 138845 2601 138857 2604
rect 138891 2601 138903 2635
rect 139670 2632 139676 2644
rect 138845 2595 138903 2601
rect 138960 2604 139676 2632
rect 138960 2564 138988 2604
rect 139670 2592 139676 2604
rect 139728 2592 139734 2644
rect 139854 2632 139860 2644
rect 139815 2604 139860 2632
rect 139854 2592 139860 2604
rect 139912 2592 139918 2644
rect 139946 2592 139952 2644
rect 140004 2632 140010 2644
rect 144178 2632 144184 2644
rect 140004 2604 144184 2632
rect 140004 2592 140010 2604
rect 144178 2592 144184 2604
rect 144236 2592 144242 2644
rect 144546 2632 144552 2644
rect 144288 2604 144552 2632
rect 144288 2564 144316 2604
rect 144546 2592 144552 2604
rect 144604 2592 144610 2644
rect 144641 2635 144699 2641
rect 144641 2601 144653 2635
rect 144687 2632 144699 2635
rect 147950 2632 147956 2644
rect 144687 2604 147956 2632
rect 144687 2601 144699 2604
rect 144641 2595 144699 2601
rect 147950 2592 147956 2604
rect 148008 2592 148014 2644
rect 149256 2604 162164 2632
rect 134720 2536 138988 2564
rect 139044 2536 144316 2564
rect 144380 2536 145328 2564
rect 132368 2524 132374 2536
rect 128446 2496 128452 2508
rect 127912 2468 128452 2496
rect 127575 2465 127587 2468
rect 127529 2459 127587 2465
rect 128446 2456 128452 2468
rect 128504 2456 128510 2508
rect 128541 2499 128599 2505
rect 128541 2465 128553 2499
rect 128587 2496 128599 2499
rect 129366 2496 129372 2508
rect 128587 2468 129372 2496
rect 128587 2465 128599 2468
rect 128541 2459 128599 2465
rect 129366 2456 129372 2468
rect 129424 2456 129430 2508
rect 129550 2496 129556 2508
rect 129511 2468 129556 2496
rect 129550 2456 129556 2468
rect 129608 2456 129614 2508
rect 130841 2499 130899 2505
rect 130841 2465 130853 2499
rect 130887 2496 130899 2499
rect 130930 2496 130936 2508
rect 130887 2468 130936 2496
rect 130887 2465 130899 2468
rect 130841 2459 130899 2465
rect 130930 2456 130936 2468
rect 130988 2456 130994 2508
rect 131850 2496 131856 2508
rect 131811 2468 131856 2496
rect 131850 2456 131856 2468
rect 131908 2456 131914 2508
rect 133141 2499 133199 2505
rect 133141 2465 133153 2499
rect 133187 2496 133199 2499
rect 133506 2496 133512 2508
rect 133187 2468 133512 2496
rect 133187 2465 133199 2468
rect 133141 2459 133199 2465
rect 133506 2456 133512 2468
rect 133564 2456 133570 2508
rect 134058 2456 134064 2508
rect 134116 2496 134122 2508
rect 135806 2496 135812 2508
rect 134116 2468 135812 2496
rect 134116 2456 134122 2468
rect 135806 2456 135812 2468
rect 135864 2456 135870 2508
rect 135901 2499 135959 2505
rect 135901 2465 135913 2499
rect 135947 2465 135959 2499
rect 135901 2459 135959 2465
rect 119172 2400 127848 2428
rect 109144 2332 111380 2360
rect 99024 2264 99788 2292
rect 100110 2252 100116 2304
rect 100168 2292 100174 2304
rect 107286 2292 107292 2304
rect 100168 2264 107292 2292
rect 100168 2252 100174 2264
rect 107286 2252 107292 2264
rect 107344 2252 107350 2304
rect 107378 2252 107384 2304
rect 107436 2292 107442 2304
rect 109221 2295 109279 2301
rect 109221 2292 109233 2295
rect 107436 2264 109233 2292
rect 107436 2252 107442 2264
rect 109221 2261 109233 2264
rect 109267 2261 109279 2295
rect 109221 2255 109279 2261
rect 109310 2252 109316 2304
rect 109368 2292 109374 2304
rect 110414 2292 110420 2304
rect 109368 2264 110420 2292
rect 109368 2252 109374 2264
rect 110414 2252 110420 2264
rect 110472 2252 110478 2304
rect 111153 2295 111211 2301
rect 111153 2261 111165 2295
rect 111199 2292 111211 2295
rect 111242 2292 111248 2304
rect 111199 2264 111248 2292
rect 111199 2261 111211 2264
rect 111153 2255 111211 2261
rect 111242 2252 111248 2264
rect 111300 2252 111306 2304
rect 111352 2292 111380 2332
rect 111426 2320 111432 2372
rect 111484 2360 111490 2372
rect 119249 2363 119307 2369
rect 119249 2360 119261 2363
rect 111484 2332 119261 2360
rect 111484 2320 111490 2332
rect 119249 2329 119261 2332
rect 119295 2329 119307 2363
rect 119249 2323 119307 2329
rect 120000 2332 124904 2360
rect 116210 2292 116216 2304
rect 111352 2264 116216 2292
rect 116210 2252 116216 2264
rect 116268 2252 116274 2304
rect 116302 2252 116308 2304
rect 116360 2292 116366 2304
rect 118234 2292 118240 2304
rect 116360 2264 118240 2292
rect 116360 2252 116366 2264
rect 118234 2252 118240 2264
rect 118292 2252 118298 2304
rect 118326 2252 118332 2304
rect 118384 2292 118390 2304
rect 120000 2292 120028 2332
rect 118384 2264 120028 2292
rect 118384 2252 118390 2264
rect 120166 2252 120172 2304
rect 120224 2292 120230 2304
rect 120353 2295 120411 2301
rect 120353 2292 120365 2295
rect 120224 2264 120365 2292
rect 120224 2252 120230 2264
rect 120353 2261 120365 2264
rect 120399 2261 120411 2295
rect 124876 2292 124904 2332
rect 125134 2320 125140 2372
rect 125192 2360 125198 2372
rect 127342 2360 127348 2372
rect 125192 2332 127348 2360
rect 125192 2320 125198 2332
rect 127342 2320 127348 2332
rect 127400 2320 127406 2372
rect 127434 2320 127440 2372
rect 127492 2360 127498 2372
rect 127621 2363 127679 2369
rect 127621 2360 127633 2363
rect 127492 2332 127633 2360
rect 127492 2320 127498 2332
rect 127621 2329 127633 2332
rect 127667 2329 127679 2363
rect 127820 2360 127848 2400
rect 128078 2388 128084 2440
rect 128136 2428 128142 2440
rect 129645 2431 129703 2437
rect 129645 2428 129657 2431
rect 128136 2400 129657 2428
rect 128136 2388 128142 2400
rect 129645 2397 129657 2400
rect 129691 2397 129703 2431
rect 129645 2391 129703 2397
rect 130194 2388 130200 2440
rect 130252 2428 130258 2440
rect 133233 2431 133291 2437
rect 133233 2428 133245 2431
rect 130252 2400 133245 2428
rect 130252 2388 130258 2400
rect 133233 2397 133245 2400
rect 133279 2397 133291 2431
rect 133233 2391 133291 2397
rect 133414 2388 133420 2440
rect 133472 2428 133478 2440
rect 134521 2431 134579 2437
rect 134521 2428 134533 2431
rect 133472 2400 134533 2428
rect 133472 2388 133478 2400
rect 134521 2397 134533 2400
rect 134567 2397 134579 2431
rect 134521 2391 134579 2397
rect 134610 2388 134616 2440
rect 134668 2428 134674 2440
rect 135622 2428 135628 2440
rect 134668 2400 135628 2428
rect 134668 2388 134674 2400
rect 135622 2388 135628 2400
rect 135680 2388 135686 2440
rect 129274 2360 129280 2372
rect 127820 2332 129280 2360
rect 127621 2323 127679 2329
rect 129274 2320 129280 2332
rect 129332 2320 129338 2372
rect 130378 2360 130384 2372
rect 129384 2332 130384 2360
rect 129384 2292 129412 2332
rect 130378 2320 130384 2332
rect 130436 2320 130442 2372
rect 130933 2363 130991 2369
rect 130933 2329 130945 2363
rect 130979 2360 130991 2363
rect 135530 2360 135536 2372
rect 130979 2332 135536 2360
rect 130979 2329 130991 2332
rect 130933 2323 130991 2329
rect 135530 2320 135536 2332
rect 135588 2320 135594 2372
rect 135806 2360 135812 2372
rect 135767 2332 135812 2360
rect 135806 2320 135812 2332
rect 135864 2320 135870 2372
rect 135916 2360 135944 2459
rect 136174 2456 136180 2508
rect 136232 2496 136238 2508
rect 137649 2499 137707 2505
rect 136232 2468 137600 2496
rect 136232 2456 136238 2468
rect 137572 2428 137600 2468
rect 137649 2465 137661 2499
rect 137695 2496 137707 2499
rect 137830 2496 137836 2508
rect 137695 2468 137836 2496
rect 137695 2465 137707 2468
rect 137649 2459 137707 2465
rect 137830 2456 137836 2468
rect 137888 2456 137894 2508
rect 138014 2456 138020 2508
rect 138072 2496 138078 2508
rect 138382 2496 138388 2508
rect 138072 2468 138388 2496
rect 138072 2456 138078 2468
rect 138382 2456 138388 2468
rect 138440 2456 138446 2508
rect 138777 2499 138835 2505
rect 138777 2465 138789 2499
rect 138823 2496 138835 2499
rect 139044 2496 139072 2536
rect 138823 2468 139072 2496
rect 139765 2499 139823 2505
rect 138823 2465 138835 2468
rect 138777 2459 138835 2465
rect 139765 2465 139777 2499
rect 139811 2465 139823 2499
rect 139765 2459 139823 2465
rect 137738 2428 137744 2440
rect 136192 2400 137416 2428
rect 137572 2400 137744 2428
rect 136192 2360 136220 2400
rect 135916 2332 136220 2360
rect 136634 2320 136640 2372
rect 136692 2360 136698 2372
rect 137388 2360 137416 2400
rect 137738 2388 137744 2400
rect 137796 2388 137802 2440
rect 139780 2428 139808 2459
rect 140314 2456 140320 2508
rect 140372 2496 140378 2508
rect 144380 2496 144408 2536
rect 144546 2496 144552 2508
rect 140372 2468 144408 2496
rect 144507 2468 144552 2496
rect 140372 2456 140378 2468
rect 144546 2456 144552 2468
rect 144604 2456 144610 2508
rect 145300 2496 145328 2536
rect 145742 2524 145748 2576
rect 145800 2564 145806 2576
rect 149256 2564 149284 2604
rect 145800 2536 149284 2564
rect 145800 2524 145806 2536
rect 150250 2524 150256 2576
rect 150308 2564 150314 2576
rect 157886 2564 157892 2576
rect 150308 2536 157892 2564
rect 150308 2524 150314 2536
rect 157886 2524 157892 2536
rect 157944 2524 157950 2576
rect 157978 2524 157984 2576
rect 158036 2564 158042 2576
rect 162026 2564 162032 2576
rect 158036 2536 162032 2564
rect 158036 2524 158042 2536
rect 162026 2524 162032 2536
rect 162084 2524 162090 2576
rect 162136 2564 162164 2604
rect 162486 2592 162492 2644
rect 162544 2632 162550 2644
rect 164326 2632 164332 2644
rect 162544 2604 164332 2632
rect 162544 2592 162550 2604
rect 164326 2592 164332 2604
rect 164384 2592 164390 2644
rect 164789 2635 164847 2641
rect 164789 2601 164801 2635
rect 164835 2632 164847 2635
rect 165522 2632 165528 2644
rect 164835 2604 165528 2632
rect 164835 2601 164847 2604
rect 164789 2595 164847 2601
rect 165522 2592 165528 2604
rect 165580 2592 165586 2644
rect 169297 2635 169355 2641
rect 169297 2601 169309 2635
rect 169343 2632 169355 2635
rect 171134 2632 171140 2644
rect 169343 2604 171140 2632
rect 169343 2601 169355 2604
rect 169297 2595 169355 2601
rect 171134 2592 171140 2604
rect 171192 2592 171198 2644
rect 171229 2635 171287 2641
rect 171229 2601 171241 2635
rect 171275 2632 171287 2635
rect 171686 2632 171692 2644
rect 171275 2604 171692 2632
rect 171275 2601 171287 2604
rect 171229 2595 171287 2601
rect 171686 2592 171692 2604
rect 171744 2592 171750 2644
rect 175734 2632 175740 2644
rect 171796 2604 175740 2632
rect 163038 2564 163044 2576
rect 162136 2536 163044 2564
rect 163038 2524 163044 2536
rect 163096 2524 163102 2576
rect 167454 2564 167460 2576
rect 163608 2536 167460 2564
rect 145300 2468 146248 2496
rect 146110 2428 146116 2440
rect 137848 2400 139716 2428
rect 139780 2400 146116 2428
rect 137848 2360 137876 2400
rect 136692 2332 137324 2360
rect 137388 2332 137876 2360
rect 136692 2320 136698 2332
rect 124876 2264 129412 2292
rect 129461 2295 129519 2301
rect 120353 2255 120411 2261
rect 129461 2261 129473 2295
rect 129507 2292 129519 2295
rect 129550 2292 129556 2304
rect 129507 2264 129556 2292
rect 129507 2261 129519 2264
rect 129461 2255 129519 2261
rect 129550 2252 129556 2264
rect 129608 2292 129614 2304
rect 129734 2292 129740 2304
rect 129608 2264 129740 2292
rect 129608 2252 129614 2264
rect 129734 2252 129740 2264
rect 129792 2252 129798 2304
rect 129826 2252 129832 2304
rect 129884 2292 129890 2304
rect 130746 2292 130752 2304
rect 129884 2264 130752 2292
rect 129884 2252 129890 2264
rect 130746 2252 130752 2264
rect 130804 2252 130810 2304
rect 131022 2252 131028 2304
rect 131080 2292 131086 2304
rect 137186 2292 137192 2304
rect 131080 2264 137192 2292
rect 131080 2252 131086 2264
rect 137186 2252 137192 2264
rect 137244 2252 137250 2304
rect 137296 2292 137324 2332
rect 138198 2320 138204 2372
rect 138256 2360 138262 2372
rect 139688 2360 139716 2400
rect 146110 2388 146116 2400
rect 146168 2388 146174 2440
rect 146220 2428 146248 2468
rect 146662 2456 146668 2508
rect 146720 2496 146726 2508
rect 155310 2496 155316 2508
rect 146720 2468 155316 2496
rect 146720 2456 146726 2468
rect 155310 2456 155316 2468
rect 155368 2456 155374 2508
rect 155402 2456 155408 2508
rect 155460 2496 155466 2508
rect 156046 2496 156052 2508
rect 155460 2468 156052 2496
rect 155460 2456 155466 2468
rect 156046 2456 156052 2468
rect 156104 2456 156110 2508
rect 157058 2496 157064 2508
rect 157019 2468 157064 2496
rect 157058 2456 157064 2468
rect 157116 2456 157122 2508
rect 157150 2456 157156 2508
rect 157208 2496 157214 2508
rect 157518 2496 157524 2508
rect 157208 2468 157524 2496
rect 157208 2456 157214 2468
rect 157518 2456 157524 2468
rect 157576 2456 157582 2508
rect 157628 2468 158208 2496
rect 147398 2428 147404 2440
rect 146220 2400 147404 2428
rect 147398 2388 147404 2400
rect 147456 2388 147462 2440
rect 149054 2388 149060 2440
rect 149112 2428 149118 2440
rect 157628 2428 157656 2468
rect 149112 2400 157656 2428
rect 158073 2431 158131 2437
rect 149112 2388 149118 2400
rect 158073 2397 158085 2431
rect 158119 2397 158131 2431
rect 158180 2428 158208 2468
rect 158254 2456 158260 2508
rect 158312 2496 158318 2508
rect 161014 2496 161020 2508
rect 158312 2468 161020 2496
rect 158312 2456 158318 2468
rect 161014 2456 161020 2468
rect 161072 2456 161078 2508
rect 161193 2499 161251 2505
rect 161193 2465 161205 2499
rect 161239 2465 161251 2499
rect 161193 2459 161251 2465
rect 158806 2428 158812 2440
rect 158180 2400 158812 2428
rect 158073 2391 158131 2397
rect 144454 2360 144460 2372
rect 138256 2332 139624 2360
rect 139688 2332 144460 2360
rect 138256 2320 138262 2332
rect 137646 2292 137652 2304
rect 137296 2264 137652 2292
rect 137646 2252 137652 2264
rect 137704 2252 137710 2304
rect 137741 2295 137799 2301
rect 137741 2261 137753 2295
rect 137787 2292 137799 2295
rect 139486 2292 139492 2304
rect 137787 2264 139492 2292
rect 137787 2261 137799 2264
rect 137741 2255 137799 2261
rect 139486 2252 139492 2264
rect 139544 2252 139550 2304
rect 139596 2292 139624 2332
rect 144454 2320 144460 2332
rect 144512 2320 144518 2372
rect 144638 2320 144644 2372
rect 144696 2360 144702 2372
rect 145006 2360 145012 2372
rect 144696 2332 145012 2360
rect 144696 2320 144702 2332
rect 145006 2320 145012 2332
rect 145064 2320 145070 2372
rect 153654 2320 153660 2372
rect 153712 2360 153718 2372
rect 157978 2360 157984 2372
rect 153712 2332 157984 2360
rect 153712 2320 153718 2332
rect 157978 2320 157984 2332
rect 158036 2320 158042 2372
rect 158088 2360 158116 2391
rect 158806 2388 158812 2400
rect 158864 2388 158870 2440
rect 159082 2428 159088 2440
rect 159043 2400 159088 2428
rect 159082 2388 159088 2400
rect 159140 2388 159146 2440
rect 160097 2431 160155 2437
rect 160097 2397 160109 2431
rect 160143 2428 160155 2431
rect 161106 2428 161112 2440
rect 160143 2400 161112 2428
rect 160143 2397 160155 2400
rect 160097 2391 160155 2397
rect 161106 2388 161112 2400
rect 161164 2388 161170 2440
rect 161208 2428 161236 2459
rect 161290 2456 161296 2508
rect 161348 2496 161354 2508
rect 162394 2496 162400 2508
rect 161348 2468 162400 2496
rect 161348 2456 161354 2468
rect 162394 2456 162400 2468
rect 162452 2456 162458 2508
rect 162762 2456 162768 2508
rect 162820 2496 162826 2508
rect 163133 2499 163191 2505
rect 163133 2496 163145 2499
rect 162820 2468 163145 2496
rect 162820 2456 162826 2468
rect 163133 2465 163145 2468
rect 163179 2465 163191 2499
rect 163133 2459 163191 2465
rect 163222 2456 163228 2508
rect 163280 2496 163286 2508
rect 163608 2496 163636 2536
rect 167454 2524 167460 2536
rect 167512 2524 167518 2576
rect 169754 2564 169760 2576
rect 167564 2536 169760 2564
rect 163280 2468 163636 2496
rect 163280 2456 163286 2468
rect 163682 2456 163688 2508
rect 163740 2496 163746 2508
rect 164697 2499 164755 2505
rect 163740 2468 164648 2496
rect 163740 2456 163746 2468
rect 161474 2428 161480 2440
rect 161208 2400 161480 2428
rect 161474 2388 161480 2400
rect 161532 2388 161538 2440
rect 161566 2388 161572 2440
rect 161624 2428 161630 2440
rect 164418 2428 164424 2440
rect 161624 2400 164424 2428
rect 161624 2388 161630 2400
rect 164418 2388 164424 2400
rect 164476 2388 164482 2440
rect 164620 2428 164648 2468
rect 164697 2465 164709 2499
rect 164743 2496 164755 2499
rect 167270 2496 167276 2508
rect 164743 2468 167276 2496
rect 164743 2465 164755 2468
rect 164697 2459 164755 2465
rect 167270 2456 167276 2468
rect 167328 2456 167334 2508
rect 167564 2496 167592 2536
rect 169754 2524 169760 2536
rect 169812 2524 169818 2576
rect 171796 2564 171824 2604
rect 175734 2592 175740 2604
rect 175792 2592 175798 2644
rect 175918 2632 175924 2644
rect 175879 2604 175924 2632
rect 175918 2592 175924 2604
rect 175976 2592 175982 2644
rect 176856 2604 177160 2632
rect 176746 2564 176752 2576
rect 169864 2536 171824 2564
rect 174740 2536 176752 2564
rect 167380 2468 167592 2496
rect 167641 2499 167699 2505
rect 165430 2428 165436 2440
rect 164620 2400 165436 2428
rect 165430 2388 165436 2400
rect 165488 2388 165494 2440
rect 165709 2431 165767 2437
rect 165709 2397 165721 2431
rect 165755 2428 165767 2431
rect 167380 2428 167408 2468
rect 167641 2465 167653 2499
rect 167687 2496 167699 2499
rect 167730 2496 167736 2508
rect 167687 2468 167736 2496
rect 167687 2465 167699 2468
rect 167641 2459 167699 2465
rect 167730 2456 167736 2468
rect 167788 2456 167794 2508
rect 169110 2456 169116 2508
rect 169168 2496 169174 2508
rect 169205 2499 169263 2505
rect 169205 2496 169217 2499
rect 169168 2468 169217 2496
rect 169168 2456 169174 2468
rect 169205 2465 169217 2468
rect 169251 2465 169263 2499
rect 169205 2459 169263 2465
rect 169294 2456 169300 2508
rect 169352 2496 169358 2508
rect 169864 2496 169892 2536
rect 169352 2468 169892 2496
rect 171137 2499 171195 2505
rect 169352 2456 169358 2468
rect 171137 2465 171149 2499
rect 171183 2496 171195 2499
rect 173342 2496 173348 2508
rect 171183 2468 173348 2496
rect 171183 2465 171195 2468
rect 171137 2459 171195 2465
rect 173342 2456 173348 2468
rect 173400 2456 173406 2508
rect 173986 2496 173992 2508
rect 173947 2468 173992 2496
rect 173986 2456 173992 2468
rect 174044 2456 174050 2508
rect 165755 2400 167408 2428
rect 165755 2397 165767 2400
rect 165709 2391 165767 2397
rect 167546 2388 167552 2440
rect 167604 2428 167610 2440
rect 172425 2431 172483 2437
rect 172425 2428 172437 2431
rect 167604 2400 172437 2428
rect 167604 2388 167610 2400
rect 172425 2397 172437 2400
rect 172471 2397 172483 2431
rect 172425 2391 172483 2397
rect 173897 2431 173955 2437
rect 173897 2397 173909 2431
rect 173943 2428 173955 2431
rect 174740 2428 174768 2536
rect 176746 2524 176752 2536
rect 176804 2524 176810 2576
rect 174817 2499 174875 2505
rect 174817 2465 174829 2499
rect 174863 2465 174875 2499
rect 174817 2459 174875 2465
rect 173943 2400 174768 2428
rect 174832 2428 174860 2459
rect 174906 2456 174912 2508
rect 174964 2496 174970 2508
rect 175826 2496 175832 2508
rect 174964 2468 175009 2496
rect 175787 2468 175832 2496
rect 174964 2456 174970 2468
rect 175826 2456 175832 2468
rect 175884 2456 175890 2508
rect 176856 2496 176884 2604
rect 177132 2564 177160 2604
rect 178126 2592 178132 2644
rect 178184 2632 178190 2644
rect 184382 2632 184388 2644
rect 178184 2604 184388 2632
rect 178184 2592 178190 2604
rect 184382 2592 184388 2604
rect 184440 2592 184446 2644
rect 185118 2592 185124 2644
rect 185176 2632 185182 2644
rect 192665 2635 192723 2641
rect 185176 2604 191696 2632
rect 185176 2592 185182 2604
rect 177132 2536 178816 2564
rect 176396 2468 176884 2496
rect 176933 2499 176991 2505
rect 176286 2428 176292 2440
rect 174832 2400 176292 2428
rect 173943 2397 173955 2400
rect 173897 2391 173955 2397
rect 176286 2388 176292 2400
rect 176344 2388 176350 2440
rect 176396 2360 176424 2468
rect 176933 2465 176945 2499
rect 176979 2496 176991 2499
rect 177022 2496 177028 2508
rect 176979 2468 177028 2496
rect 176979 2465 176991 2468
rect 176933 2459 176991 2465
rect 177022 2456 177028 2468
rect 177080 2456 177086 2508
rect 178788 2505 178816 2536
rect 182744 2536 185164 2564
rect 178773 2499 178831 2505
rect 178773 2465 178785 2499
rect 178819 2465 178831 2499
rect 178773 2459 178831 2465
rect 180337 2499 180395 2505
rect 180337 2465 180349 2499
rect 180383 2496 180395 2499
rect 181070 2496 181076 2508
rect 180383 2468 181076 2496
rect 180383 2465 180395 2468
rect 180337 2459 180395 2465
rect 181070 2456 181076 2468
rect 181128 2456 181134 2508
rect 182744 2505 182772 2536
rect 182729 2499 182787 2505
rect 182729 2465 182741 2499
rect 182775 2465 182787 2499
rect 182729 2459 182787 2465
rect 183649 2499 183707 2505
rect 183649 2465 183661 2499
rect 183695 2496 183707 2499
rect 184566 2496 184572 2508
rect 183695 2468 184572 2496
rect 183695 2465 183707 2468
rect 183649 2459 183707 2465
rect 184566 2456 184572 2468
rect 184624 2456 184630 2508
rect 181160 2431 181218 2437
rect 181160 2397 181172 2431
rect 181206 2428 181218 2431
rect 184474 2428 184480 2440
rect 181206 2400 184480 2428
rect 181206 2397 181218 2400
rect 181160 2391 181218 2397
rect 184474 2388 184480 2400
rect 184532 2388 184538 2440
rect 185136 2428 185164 2536
rect 185670 2524 185676 2576
rect 185728 2564 185734 2576
rect 186866 2564 186872 2576
rect 185728 2536 186872 2564
rect 185728 2524 185734 2536
rect 186866 2524 186872 2536
rect 186924 2524 186930 2576
rect 189350 2564 189356 2576
rect 187620 2536 189212 2564
rect 189311 2536 189356 2564
rect 185213 2499 185271 2505
rect 185213 2465 185225 2499
rect 185259 2496 185271 2499
rect 185946 2496 185952 2508
rect 185259 2468 185952 2496
rect 185259 2465 185271 2468
rect 185213 2459 185271 2465
rect 185946 2456 185952 2468
rect 186004 2456 186010 2508
rect 187620 2505 187648 2536
rect 187605 2499 187663 2505
rect 187605 2465 187617 2499
rect 187651 2465 187663 2499
rect 187605 2459 187663 2465
rect 186038 2428 186044 2440
rect 185136 2400 185256 2428
rect 185999 2400 186044 2428
rect 158088 2332 176424 2360
rect 180245 2363 180303 2369
rect 180245 2329 180257 2363
rect 180291 2329 180303 2363
rect 180245 2323 180303 2329
rect 146386 2292 146392 2304
rect 139596 2264 146392 2292
rect 146386 2252 146392 2264
rect 146444 2252 146450 2304
rect 153010 2252 153016 2304
rect 153068 2292 153074 2304
rect 160922 2292 160928 2304
rect 153068 2264 160928 2292
rect 153068 2252 153074 2264
rect 160922 2252 160928 2264
rect 160980 2252 160986 2304
rect 161293 2295 161351 2301
rect 161293 2261 161305 2295
rect 161339 2292 161351 2295
rect 163130 2292 163136 2304
rect 161339 2264 163136 2292
rect 161339 2261 161351 2264
rect 161293 2255 161351 2261
rect 163130 2252 163136 2264
rect 163188 2252 163194 2304
rect 163225 2295 163283 2301
rect 163225 2261 163237 2295
rect 163271 2292 163283 2295
rect 163314 2292 163320 2304
rect 163271 2264 163320 2292
rect 163271 2261 163283 2264
rect 163225 2255 163283 2261
rect 163314 2252 163320 2264
rect 163372 2252 163378 2304
rect 164878 2252 164884 2304
rect 164936 2292 164942 2304
rect 167086 2292 167092 2304
rect 164936 2264 167092 2292
rect 164936 2252 164942 2264
rect 167086 2252 167092 2264
rect 167144 2252 167150 2304
rect 167178 2252 167184 2304
rect 167236 2292 167242 2304
rect 177025 2295 177083 2301
rect 177025 2292 177037 2295
rect 167236 2264 177037 2292
rect 167236 2252 167242 2264
rect 177025 2261 177037 2264
rect 177071 2261 177083 2295
rect 177025 2255 177083 2261
rect 177758 2252 177764 2304
rect 177816 2292 177822 2304
rect 179598 2292 179604 2304
rect 177816 2264 179604 2292
rect 177816 2252 177822 2264
rect 179598 2252 179604 2264
rect 179656 2252 179662 2304
rect 180260 2292 180288 2323
rect 181254 2320 181260 2372
rect 181312 2360 181318 2372
rect 182542 2360 182548 2372
rect 181312 2332 182548 2360
rect 181312 2320 181318 2332
rect 182542 2320 182548 2332
rect 182600 2320 182606 2372
rect 182637 2363 182695 2369
rect 182637 2329 182649 2363
rect 182683 2360 182695 2363
rect 184934 2360 184940 2372
rect 182683 2332 184940 2360
rect 182683 2329 182695 2332
rect 182637 2323 182695 2329
rect 184934 2320 184940 2332
rect 184992 2320 184998 2372
rect 185118 2360 185124 2372
rect 185079 2332 185124 2360
rect 185118 2320 185124 2332
rect 185176 2320 185182 2372
rect 185228 2360 185256 2400
rect 186038 2388 186044 2400
rect 186096 2388 186102 2440
rect 187418 2428 187424 2440
rect 187379 2400 187424 2428
rect 187418 2388 187424 2400
rect 187476 2388 187482 2440
rect 189184 2428 189212 2536
rect 189350 2524 189356 2536
rect 189408 2524 189414 2576
rect 190178 2524 190184 2576
rect 190236 2564 190242 2576
rect 191668 2564 191696 2604
rect 192665 2601 192677 2635
rect 192711 2632 192723 2635
rect 192754 2632 192760 2644
rect 192711 2604 192760 2632
rect 192711 2601 192723 2604
rect 192665 2595 192723 2601
rect 192754 2592 192760 2604
rect 192812 2592 192818 2644
rect 193858 2632 193864 2644
rect 193819 2604 193864 2632
rect 193858 2592 193864 2604
rect 193916 2592 193922 2644
rect 194042 2592 194048 2644
rect 194100 2592 194106 2644
rect 194962 2632 194968 2644
rect 194923 2604 194968 2632
rect 194962 2592 194968 2604
rect 195020 2592 195026 2644
rect 195054 2592 195060 2644
rect 195112 2632 195118 2644
rect 195977 2635 196035 2641
rect 195977 2632 195989 2635
rect 195112 2604 195989 2632
rect 195112 2592 195118 2604
rect 195977 2601 195989 2604
rect 196023 2601 196035 2635
rect 195977 2595 196035 2601
rect 196434 2592 196440 2644
rect 196492 2632 196498 2644
rect 196989 2635 197047 2641
rect 196989 2632 197001 2635
rect 196492 2604 197001 2632
rect 196492 2592 196498 2604
rect 196989 2601 197001 2604
rect 197035 2601 197047 2635
rect 196989 2595 197047 2601
rect 194060 2564 194088 2592
rect 190236 2536 191604 2564
rect 191668 2536 194088 2564
rect 190236 2524 190242 2536
rect 189261 2499 189319 2505
rect 189261 2465 189273 2499
rect 189307 2496 189319 2499
rect 189718 2496 189724 2508
rect 189307 2468 189724 2496
rect 189307 2465 189319 2468
rect 189261 2459 189319 2465
rect 189718 2456 189724 2468
rect 189776 2456 189782 2508
rect 190546 2496 190552 2508
rect 190507 2468 190552 2496
rect 190546 2456 190552 2468
rect 190604 2456 190610 2508
rect 190641 2499 190699 2505
rect 190641 2465 190653 2499
rect 190687 2496 190699 2499
rect 190730 2496 190736 2508
rect 190687 2468 190736 2496
rect 190687 2465 190699 2468
rect 190641 2459 190699 2465
rect 190730 2456 190736 2468
rect 190788 2456 190794 2508
rect 191576 2505 191604 2536
rect 191561 2499 191619 2505
rect 191561 2465 191573 2499
rect 191607 2465 191619 2499
rect 191561 2459 191619 2465
rect 192573 2499 192631 2505
rect 192573 2465 192585 2499
rect 192619 2465 192631 2499
rect 192573 2459 192631 2465
rect 191653 2431 191711 2437
rect 191653 2428 191665 2431
rect 189184 2400 191665 2428
rect 191653 2397 191665 2400
rect 191699 2397 191711 2431
rect 191653 2391 191711 2397
rect 186590 2360 186596 2372
rect 185228 2332 186596 2360
rect 186590 2320 186596 2332
rect 186648 2320 186654 2372
rect 191006 2320 191012 2372
rect 191064 2360 191070 2372
rect 192588 2360 192616 2459
rect 193214 2456 193220 2508
rect 193272 2496 193278 2508
rect 193769 2499 193827 2505
rect 193769 2496 193781 2499
rect 193272 2468 193781 2496
rect 193272 2456 193278 2468
rect 193769 2465 193781 2468
rect 193815 2465 193827 2499
rect 193769 2459 193827 2465
rect 194042 2456 194048 2508
rect 194100 2496 194106 2508
rect 194873 2499 194931 2505
rect 194873 2496 194885 2499
rect 194100 2468 194885 2496
rect 194100 2456 194106 2468
rect 194873 2465 194885 2468
rect 194919 2465 194931 2499
rect 194873 2459 194931 2465
rect 195885 2499 195943 2505
rect 195885 2465 195897 2499
rect 195931 2465 195943 2499
rect 196894 2496 196900 2508
rect 196855 2468 196900 2496
rect 195885 2459 195943 2465
rect 192754 2388 192760 2440
rect 192812 2428 192818 2440
rect 195900 2428 195928 2459
rect 196894 2456 196900 2468
rect 196952 2456 196958 2508
rect 192812 2400 195928 2428
rect 192812 2388 192818 2400
rect 191064 2332 192616 2360
rect 191064 2320 191070 2332
rect 192662 2320 192668 2372
rect 192720 2360 192726 2372
rect 193490 2360 193496 2372
rect 192720 2332 193496 2360
rect 192720 2320 192726 2332
rect 193490 2320 193496 2332
rect 193548 2320 193554 2372
rect 187326 2292 187332 2304
rect 180260 2264 187332 2292
rect 187326 2252 187332 2264
rect 187384 2252 187390 2304
rect 187510 2252 187516 2304
rect 187568 2292 187574 2304
rect 193306 2292 193312 2304
rect 187568 2264 193312 2292
rect 187568 2252 187574 2264
rect 193306 2252 193312 2264
rect 193364 2252 193370 2304
rect 1104 2202 198812 2224
rect 1104 2150 4078 2202
rect 4130 2150 44078 2202
rect 44130 2150 84078 2202
rect 84130 2150 124078 2202
rect 124130 2150 164078 2202
rect 164130 2150 198812 2202
rect 1104 2128 198812 2150
rect 5353 2091 5411 2097
rect 5353 2057 5365 2091
rect 5399 2088 5411 2091
rect 5718 2088 5724 2100
rect 5399 2060 5724 2088
rect 5399 2057 5411 2060
rect 5353 2051 5411 2057
rect 5718 2048 5724 2060
rect 5776 2048 5782 2100
rect 6362 2048 6368 2100
rect 6420 2088 6426 2100
rect 6917 2091 6975 2097
rect 6917 2088 6929 2091
rect 6420 2060 6929 2088
rect 6420 2048 6426 2060
rect 6917 2057 6929 2060
rect 6963 2057 6975 2091
rect 6917 2051 6975 2057
rect 7466 2048 7472 2100
rect 7524 2088 7530 2100
rect 7929 2091 7987 2097
rect 7929 2088 7941 2091
rect 7524 2060 7941 2088
rect 7524 2048 7530 2060
rect 7929 2057 7941 2060
rect 7975 2057 7987 2091
rect 8938 2088 8944 2100
rect 8899 2060 8944 2088
rect 7929 2051 7987 2057
rect 8938 2048 8944 2060
rect 8996 2048 9002 2100
rect 9950 2088 9956 2100
rect 9911 2060 9956 2088
rect 9950 2048 9956 2060
rect 10008 2048 10014 2100
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 11425 2091 11483 2097
rect 11425 2088 11437 2091
rect 11204 2060 11437 2088
rect 11204 2048 11210 2060
rect 11425 2057 11437 2060
rect 11471 2057 11483 2091
rect 11425 2051 11483 2057
rect 12805 2091 12863 2097
rect 12805 2057 12817 2091
rect 12851 2088 12863 2091
rect 13538 2088 13544 2100
rect 12851 2060 13544 2088
rect 12851 2057 12863 2060
rect 12805 2051 12863 2057
rect 13538 2048 13544 2060
rect 13596 2048 13602 2100
rect 13814 2088 13820 2100
rect 13775 2060 13820 2088
rect 13814 2048 13820 2060
rect 13872 2048 13878 2100
rect 16301 2091 16359 2097
rect 16301 2057 16313 2091
rect 16347 2088 16359 2091
rect 16666 2088 16672 2100
rect 16347 2060 16672 2088
rect 16347 2057 16359 2060
rect 16301 2051 16359 2057
rect 16666 2048 16672 2060
rect 16724 2048 16730 2100
rect 18141 2091 18199 2097
rect 18141 2057 18153 2091
rect 18187 2088 18199 2091
rect 19426 2088 19432 2100
rect 18187 2060 19432 2088
rect 18187 2057 18199 2060
rect 18141 2051 18199 2057
rect 19426 2048 19432 2060
rect 19484 2048 19490 2100
rect 20530 2088 20536 2100
rect 20491 2060 20536 2088
rect 20530 2048 20536 2060
rect 20588 2048 20594 2100
rect 21637 2091 21695 2097
rect 21637 2057 21649 2091
rect 21683 2088 21695 2091
rect 23566 2088 23572 2100
rect 21683 2060 23572 2088
rect 21683 2057 21695 2060
rect 21637 2051 21695 2057
rect 23566 2048 23572 2060
rect 23624 2048 23630 2100
rect 23753 2091 23811 2097
rect 23753 2057 23765 2091
rect 23799 2088 23811 2091
rect 25038 2088 25044 2100
rect 23799 2060 25044 2088
rect 23799 2057 23811 2060
rect 23753 2051 23811 2057
rect 25038 2048 25044 2060
rect 25096 2048 25102 2100
rect 26697 2091 26755 2097
rect 26697 2057 26709 2091
rect 26743 2088 26755 2091
rect 27890 2088 27896 2100
rect 26743 2060 27896 2088
rect 26743 2057 26755 2060
rect 26697 2051 26755 2057
rect 27890 2048 27896 2060
rect 27948 2048 27954 2100
rect 30285 2091 30343 2097
rect 30285 2057 30297 2091
rect 30331 2088 30343 2091
rect 30466 2088 30472 2100
rect 30331 2060 30472 2088
rect 30331 2057 30343 2060
rect 30285 2051 30343 2057
rect 30466 2048 30472 2060
rect 30524 2048 30530 2100
rect 32306 2088 32312 2100
rect 32267 2060 32312 2088
rect 32306 2048 32312 2060
rect 32364 2048 32370 2100
rect 32766 2048 32772 2100
rect 32824 2088 32830 2100
rect 33321 2091 33379 2097
rect 33321 2088 33333 2091
rect 32824 2060 33333 2088
rect 32824 2048 32830 2060
rect 33321 2057 33333 2060
rect 33367 2057 33379 2091
rect 34974 2088 34980 2100
rect 34935 2060 34980 2088
rect 33321 2051 33379 2057
rect 34974 2048 34980 2060
rect 35032 2048 35038 2100
rect 37829 2091 37887 2097
rect 37829 2057 37841 2091
rect 37875 2088 37887 2091
rect 37918 2088 37924 2100
rect 37875 2060 37924 2088
rect 37875 2057 37887 2060
rect 37829 2051 37887 2057
rect 37918 2048 37924 2060
rect 37976 2048 37982 2100
rect 39390 2088 39396 2100
rect 39351 2060 39396 2088
rect 39390 2048 39396 2060
rect 39448 2048 39454 2100
rect 41138 2088 41144 2100
rect 41099 2060 41144 2088
rect 41138 2048 41144 2060
rect 41196 2048 41202 2100
rect 42334 2088 42340 2100
rect 42295 2060 42340 2088
rect 42334 2048 42340 2060
rect 42392 2048 42398 2100
rect 43441 2091 43499 2097
rect 43441 2057 43453 2091
rect 43487 2088 43499 2091
rect 44266 2088 44272 2100
rect 43487 2060 44272 2088
rect 43487 2057 43499 2060
rect 43441 2051 43499 2057
rect 44266 2048 44272 2060
rect 44324 2048 44330 2100
rect 44450 2088 44456 2100
rect 44411 2060 44456 2088
rect 44450 2048 44456 2060
rect 44508 2048 44514 2100
rect 46198 2048 46204 2100
rect 46256 2088 46262 2100
rect 46293 2091 46351 2097
rect 46293 2088 46305 2091
rect 46256 2060 46305 2088
rect 46256 2048 46262 2060
rect 46293 2057 46305 2060
rect 46339 2057 46351 2091
rect 47302 2088 47308 2100
rect 47263 2060 47308 2088
rect 46293 2051 46351 2057
rect 47302 2048 47308 2060
rect 47360 2048 47366 2100
rect 48317 2091 48375 2097
rect 48317 2057 48329 2091
rect 48363 2088 48375 2091
rect 49694 2088 49700 2100
rect 48363 2060 49700 2088
rect 48363 2057 48375 2060
rect 48317 2051 48375 2057
rect 49694 2048 49700 2060
rect 49752 2048 49758 2100
rect 50709 2091 50767 2097
rect 50709 2057 50721 2091
rect 50755 2088 50767 2091
rect 54846 2088 54852 2100
rect 50755 2060 54852 2088
rect 50755 2057 50767 2060
rect 50709 2051 50767 2057
rect 54846 2048 54852 2060
rect 54904 2048 54910 2100
rect 57330 2088 57336 2100
rect 55508 2060 57336 2088
rect 22649 2023 22707 2029
rect 22649 1989 22661 2023
rect 22695 2020 22707 2023
rect 24762 2020 24768 2032
rect 22695 1992 24768 2020
rect 22695 1989 22707 1992
rect 22649 1983 22707 1989
rect 24762 1980 24768 1992
rect 24820 1980 24826 2032
rect 30190 1980 30196 2032
rect 30248 2020 30254 2032
rect 31297 2023 31355 2029
rect 31297 2020 31309 2023
rect 30248 1992 31309 2020
rect 30248 1980 30254 1992
rect 31297 1989 31309 1992
rect 31343 1989 31355 2023
rect 31297 1983 31355 1989
rect 33410 1980 33416 2032
rect 33468 2020 33474 2032
rect 36357 2023 36415 2029
rect 36357 2020 36369 2023
rect 33468 1992 36369 2020
rect 33468 1980 33474 1992
rect 36357 1989 36369 1992
rect 36403 1989 36415 2023
rect 55508 2020 55536 2060
rect 57330 2048 57336 2060
rect 57388 2048 57394 2100
rect 57425 2091 57483 2097
rect 57425 2057 57437 2091
rect 57471 2088 57483 2091
rect 59538 2088 59544 2100
rect 57471 2060 59544 2088
rect 57471 2057 57483 2060
rect 57425 2051 57483 2057
rect 59538 2048 59544 2060
rect 59596 2048 59602 2100
rect 64969 2091 65027 2097
rect 64969 2057 64981 2091
rect 65015 2088 65027 2091
rect 67726 2088 67732 2100
rect 65015 2060 67732 2088
rect 65015 2057 65027 2060
rect 64969 2051 65027 2057
rect 67726 2048 67732 2060
rect 67784 2048 67790 2100
rect 69658 2048 69664 2100
rect 69716 2088 69722 2100
rect 93210 2088 93216 2100
rect 69716 2060 93216 2088
rect 69716 2048 69722 2060
rect 93210 2048 93216 2060
rect 93268 2048 93274 2100
rect 94498 2048 94504 2100
rect 94556 2088 94562 2100
rect 100202 2088 100208 2100
rect 94556 2060 100064 2088
rect 100163 2060 100208 2088
rect 94556 2048 94562 2060
rect 58894 2020 58900 2032
rect 36357 1983 36415 1989
rect 53760 1992 55536 2020
rect 55600 1992 58900 2020
rect 15838 1912 15844 1964
rect 15896 1952 15902 1964
rect 15896 1924 20484 1952
rect 15896 1912 15902 1924
rect 4522 1844 4528 1896
rect 4580 1884 4586 1896
rect 5261 1887 5319 1893
rect 5261 1884 5273 1887
rect 4580 1856 5273 1884
rect 4580 1844 4586 1856
rect 5261 1853 5273 1856
rect 5307 1853 5319 1887
rect 5261 1847 5319 1853
rect 5350 1844 5356 1896
rect 5408 1884 5414 1896
rect 6825 1887 6883 1893
rect 6825 1884 6837 1887
rect 5408 1856 6837 1884
rect 5408 1844 5414 1856
rect 6825 1853 6837 1856
rect 6871 1853 6883 1887
rect 6825 1847 6883 1853
rect 7837 1887 7895 1893
rect 7837 1853 7849 1887
rect 7883 1853 7895 1887
rect 7837 1847 7895 1853
rect 8849 1887 8907 1893
rect 8849 1853 8861 1887
rect 8895 1884 8907 1887
rect 9306 1884 9312 1896
rect 8895 1856 9312 1884
rect 8895 1853 8907 1856
rect 8849 1847 8907 1853
rect 6270 1776 6276 1828
rect 6328 1816 6334 1828
rect 7852 1816 7880 1847
rect 9306 1844 9312 1856
rect 9364 1844 9370 1896
rect 9861 1887 9919 1893
rect 9861 1853 9873 1887
rect 9907 1884 9919 1887
rect 10134 1884 10140 1896
rect 9907 1856 10140 1884
rect 9907 1853 9919 1856
rect 9861 1847 9919 1853
rect 10134 1844 10140 1856
rect 10192 1844 10198 1896
rect 11054 1844 11060 1896
rect 11112 1884 11118 1896
rect 11333 1887 11391 1893
rect 11333 1884 11345 1887
rect 11112 1856 11345 1884
rect 11112 1844 11118 1856
rect 11333 1853 11345 1856
rect 11379 1853 11391 1887
rect 11333 1847 11391 1853
rect 12713 1887 12771 1893
rect 12713 1853 12725 1887
rect 12759 1884 12771 1887
rect 13262 1884 13268 1896
rect 12759 1856 13268 1884
rect 12759 1853 12771 1856
rect 12713 1847 12771 1853
rect 13262 1844 13268 1856
rect 13320 1844 13326 1896
rect 13725 1887 13783 1893
rect 13725 1853 13737 1887
rect 13771 1853 13783 1887
rect 13725 1847 13783 1853
rect 6328 1788 7880 1816
rect 6328 1776 6334 1788
rect 11882 1776 11888 1828
rect 11940 1816 11946 1828
rect 13740 1816 13768 1847
rect 15378 1844 15384 1896
rect 15436 1884 15442 1896
rect 16209 1887 16267 1893
rect 16209 1884 16221 1887
rect 15436 1856 16221 1884
rect 15436 1844 15442 1856
rect 16209 1853 16221 1856
rect 16255 1853 16267 1887
rect 16209 1847 16267 1853
rect 16666 1844 16672 1896
rect 16724 1884 16730 1896
rect 20456 1893 20484 1924
rect 21634 1912 21640 1964
rect 21692 1952 21698 1964
rect 21692 1924 23704 1952
rect 21692 1912 21698 1924
rect 23676 1893 23704 1924
rect 24578 1912 24584 1964
rect 24636 1952 24642 1964
rect 29730 1952 29736 1964
rect 24636 1924 26648 1952
rect 24636 1912 24642 1924
rect 26620 1893 26648 1924
rect 28000 1924 29736 1952
rect 18049 1887 18107 1893
rect 18049 1884 18061 1887
rect 16724 1856 18061 1884
rect 16724 1844 16730 1856
rect 18049 1853 18061 1856
rect 18095 1853 18107 1887
rect 18049 1847 18107 1853
rect 20441 1887 20499 1893
rect 20441 1853 20453 1887
rect 20487 1853 20499 1887
rect 21545 1887 21603 1893
rect 21545 1884 21557 1887
rect 20441 1847 20499 1853
rect 20548 1856 21557 1884
rect 11940 1788 13768 1816
rect 11940 1776 11946 1788
rect 17586 1776 17592 1828
rect 17644 1816 17650 1828
rect 20548 1816 20576 1856
rect 21545 1853 21557 1856
rect 21591 1853 21603 1887
rect 21545 1847 21603 1853
rect 22557 1887 22615 1893
rect 22557 1853 22569 1887
rect 22603 1853 22615 1887
rect 22557 1847 22615 1853
rect 23661 1887 23719 1893
rect 23661 1853 23673 1887
rect 23707 1853 23719 1887
rect 23661 1847 23719 1853
rect 25593 1887 25651 1893
rect 25593 1853 25605 1887
rect 25639 1853 25651 1887
rect 25593 1847 25651 1853
rect 26613 1887 26671 1893
rect 26613 1853 26625 1887
rect 26659 1853 26671 1887
rect 26613 1847 26671 1853
rect 17644 1788 20576 1816
rect 17644 1776 17650 1788
rect 21082 1776 21088 1828
rect 21140 1816 21146 1828
rect 22572 1816 22600 1847
rect 21140 1788 22600 1816
rect 21140 1776 21146 1788
rect 22830 1776 22836 1828
rect 22888 1816 22894 1828
rect 25608 1816 25636 1847
rect 22888 1788 25636 1816
rect 25685 1819 25743 1825
rect 22888 1776 22894 1788
rect 25685 1785 25697 1819
rect 25731 1816 25743 1819
rect 28000 1816 28028 1924
rect 29730 1912 29736 1924
rect 29788 1912 29794 1964
rect 30282 1912 30288 1964
rect 30340 1952 30346 1964
rect 30340 1924 31892 1952
rect 30340 1912 30346 1924
rect 28074 1844 28080 1896
rect 28132 1884 28138 1896
rect 30193 1887 30251 1893
rect 30193 1884 30205 1887
rect 28132 1856 30205 1884
rect 28132 1844 28138 1856
rect 30193 1853 30205 1856
rect 30239 1853 30251 1887
rect 30193 1847 30251 1853
rect 31205 1887 31263 1893
rect 31205 1853 31217 1887
rect 31251 1853 31263 1887
rect 31205 1847 31263 1853
rect 25731 1788 28028 1816
rect 25731 1785 25743 1788
rect 25685 1779 25743 1785
rect 28902 1776 28908 1828
rect 28960 1816 28966 1828
rect 31220 1816 31248 1847
rect 28960 1788 31248 1816
rect 31864 1816 31892 1924
rect 31938 1912 31944 1964
rect 31996 1952 32002 1964
rect 31996 1924 34928 1952
rect 31996 1912 32002 1924
rect 34900 1893 34928 1924
rect 41414 1912 41420 1964
rect 41472 1952 41478 1964
rect 41472 1924 43392 1952
rect 41472 1912 41478 1924
rect 32225 1887 32283 1893
rect 32225 1853 32237 1887
rect 32271 1853 32283 1887
rect 33229 1887 33287 1893
rect 33229 1884 33241 1887
rect 32225 1847 32283 1853
rect 32508 1856 33241 1884
rect 32232 1816 32260 1847
rect 31864 1788 32260 1816
rect 28960 1776 28966 1788
rect 21450 1708 21456 1760
rect 21508 1748 21514 1760
rect 23750 1748 23756 1760
rect 21508 1720 23756 1748
rect 21508 1708 21514 1720
rect 23750 1708 23756 1720
rect 23808 1708 23814 1760
rect 27614 1708 27620 1760
rect 27672 1748 27678 1760
rect 32508 1748 32536 1856
rect 33229 1853 33241 1856
rect 33275 1853 33287 1887
rect 33229 1847 33287 1853
rect 34885 1887 34943 1893
rect 34885 1853 34897 1887
rect 34931 1853 34943 1887
rect 36265 1887 36323 1893
rect 36265 1884 36277 1887
rect 34885 1847 34943 1853
rect 34992 1856 36277 1884
rect 32858 1776 32864 1828
rect 32916 1816 32922 1828
rect 34992 1816 35020 1856
rect 36265 1853 36277 1856
rect 36311 1853 36323 1887
rect 37734 1884 37740 1896
rect 37695 1856 37740 1884
rect 36265 1847 36323 1853
rect 37734 1844 37740 1856
rect 37792 1844 37798 1896
rect 39301 1887 39359 1893
rect 39301 1853 39313 1887
rect 39347 1853 39359 1887
rect 39301 1847 39359 1853
rect 41049 1887 41107 1893
rect 41049 1853 41061 1887
rect 41095 1853 41107 1887
rect 41049 1847 41107 1853
rect 42245 1887 42303 1893
rect 42245 1853 42257 1887
rect 42291 1884 42303 1887
rect 42886 1884 42892 1896
rect 42291 1856 42892 1884
rect 42291 1853 42303 1856
rect 42245 1847 42303 1853
rect 32916 1788 35020 1816
rect 32916 1776 32922 1788
rect 35894 1776 35900 1828
rect 35952 1816 35958 1828
rect 39316 1816 39344 1847
rect 35952 1788 39344 1816
rect 35952 1776 35958 1788
rect 27672 1720 32536 1748
rect 27672 1708 27678 1720
rect 36722 1708 36728 1760
rect 36780 1748 36786 1760
rect 41064 1748 41092 1847
rect 42886 1844 42892 1856
rect 42944 1844 42950 1896
rect 43364 1893 43392 1924
rect 43349 1887 43407 1893
rect 43349 1853 43361 1887
rect 43395 1853 43407 1887
rect 43349 1847 43407 1853
rect 43438 1844 43444 1896
rect 43496 1884 43502 1896
rect 44361 1887 44419 1893
rect 44361 1884 44373 1887
rect 43496 1856 44373 1884
rect 43496 1844 43502 1856
rect 44361 1853 44373 1856
rect 44407 1853 44419 1887
rect 44361 1847 44419 1853
rect 46201 1887 46259 1893
rect 46201 1853 46213 1887
rect 46247 1853 46259 1887
rect 46201 1847 46259 1853
rect 41506 1776 41512 1828
rect 41564 1816 41570 1828
rect 46216 1816 46244 1847
rect 46382 1844 46388 1896
rect 46440 1884 46446 1896
rect 47213 1887 47271 1893
rect 47213 1884 47225 1887
rect 46440 1856 47225 1884
rect 46440 1844 46446 1856
rect 47213 1853 47225 1856
rect 47259 1853 47271 1887
rect 47213 1847 47271 1853
rect 47670 1844 47676 1896
rect 47728 1884 47734 1896
rect 48225 1887 48283 1893
rect 48225 1884 48237 1887
rect 47728 1856 48237 1884
rect 47728 1844 47734 1856
rect 48225 1853 48237 1856
rect 48271 1853 48283 1887
rect 48225 1847 48283 1853
rect 50617 1887 50675 1893
rect 50617 1853 50629 1887
rect 50663 1884 50675 1887
rect 50706 1884 50712 1896
rect 50663 1856 50712 1884
rect 50663 1853 50675 1856
rect 50617 1847 50675 1853
rect 50706 1844 50712 1856
rect 50764 1844 50770 1896
rect 52365 1887 52423 1893
rect 52365 1853 52377 1887
rect 52411 1853 52423 1887
rect 52365 1847 52423 1853
rect 52457 1887 52515 1893
rect 52457 1853 52469 1887
rect 52503 1884 52515 1887
rect 53558 1884 53564 1896
rect 52503 1856 53564 1884
rect 52503 1853 52515 1856
rect 52457 1847 52515 1853
rect 41564 1788 46244 1816
rect 52380 1816 52408 1847
rect 53558 1844 53564 1856
rect 53616 1844 53622 1896
rect 53760 1893 53788 1992
rect 55600 1952 55628 1992
rect 58894 1980 58900 1992
rect 58952 1980 58958 2032
rect 62298 2020 62304 2032
rect 59280 1992 62304 2020
rect 53852 1924 55628 1952
rect 55677 1955 55735 1961
rect 53745 1887 53803 1893
rect 53745 1853 53757 1887
rect 53791 1853 53803 1887
rect 53745 1847 53803 1853
rect 53852 1816 53880 1924
rect 55677 1921 55689 1955
rect 55723 1952 55735 1955
rect 57698 1952 57704 1964
rect 55723 1924 57704 1952
rect 55723 1921 55735 1924
rect 55677 1915 55735 1921
rect 57698 1912 57704 1924
rect 57756 1912 57762 1964
rect 54018 1884 54024 1896
rect 53979 1856 54024 1884
rect 54018 1844 54024 1856
rect 54076 1844 54082 1896
rect 55122 1884 55128 1896
rect 55083 1856 55128 1884
rect 55122 1844 55128 1856
rect 55180 1844 55186 1896
rect 59280 1893 59308 1992
rect 62298 1980 62304 1992
rect 62356 1980 62362 2032
rect 65978 2020 65984 2032
rect 63696 1992 65984 2020
rect 59541 1955 59599 1961
rect 59541 1921 59553 1955
rect 59587 1952 59599 1955
rect 62022 1952 62028 1964
rect 59587 1924 62028 1952
rect 59587 1921 59599 1924
rect 59541 1915 59599 1921
rect 62022 1912 62028 1924
rect 62080 1912 62086 1964
rect 63696 1961 63724 1992
rect 65978 1980 65984 1992
rect 66036 1980 66042 2032
rect 71866 2020 71872 2032
rect 66088 1992 71872 2020
rect 63681 1955 63739 1961
rect 63681 1921 63693 1955
rect 63727 1921 63739 1955
rect 63681 1915 63739 1921
rect 57333 1887 57391 1893
rect 57333 1853 57345 1887
rect 57379 1853 57391 1887
rect 57333 1847 57391 1853
rect 59265 1887 59323 1893
rect 59265 1853 59277 1887
rect 59311 1853 59323 1887
rect 59265 1847 59323 1853
rect 61013 1887 61071 1893
rect 61013 1853 61025 1887
rect 61059 1884 61071 1887
rect 62114 1884 62120 1896
rect 61059 1856 62120 1884
rect 61059 1853 61071 1856
rect 61013 1847 61071 1853
rect 52380 1788 53880 1816
rect 41564 1776 41570 1788
rect 54662 1776 54668 1828
rect 54720 1816 54726 1828
rect 57348 1816 57376 1847
rect 62114 1844 62120 1856
rect 62172 1844 62178 1896
rect 63405 1887 63463 1893
rect 63405 1853 63417 1887
rect 63451 1853 63463 1887
rect 63405 1847 63463 1853
rect 65153 1887 65211 1893
rect 65153 1853 65165 1887
rect 65199 1884 65211 1887
rect 66088 1884 66116 1992
rect 71866 1980 71872 1992
rect 71924 1980 71930 2032
rect 81434 1980 81440 2032
rect 81492 2020 81498 2032
rect 81986 2020 81992 2032
rect 81492 1992 81992 2020
rect 81492 1980 81498 1992
rect 81986 1980 81992 1992
rect 82044 1980 82050 2032
rect 82998 1980 83004 2032
rect 83056 1980 83062 2032
rect 83274 1980 83280 2032
rect 83332 2020 83338 2032
rect 89714 2020 89720 2032
rect 83332 1992 89720 2020
rect 83332 1980 83338 1992
rect 89714 1980 89720 1992
rect 89772 1980 89778 2032
rect 100036 2020 100064 2060
rect 100202 2048 100208 2060
rect 100260 2048 100266 2100
rect 105262 2048 105268 2100
rect 105320 2088 105326 2100
rect 108390 2088 108396 2100
rect 105320 2060 108396 2088
rect 105320 2048 105326 2060
rect 108390 2048 108396 2060
rect 108448 2048 108454 2100
rect 108758 2048 108764 2100
rect 108816 2048 108822 2100
rect 108942 2048 108948 2100
rect 109000 2088 109006 2100
rect 109310 2088 109316 2100
rect 109000 2060 109316 2088
rect 109000 2048 109006 2060
rect 109310 2048 109316 2060
rect 109368 2048 109374 2100
rect 109402 2048 109408 2100
rect 109460 2088 109466 2100
rect 113910 2088 113916 2100
rect 109460 2060 113916 2088
rect 109460 2048 109466 2060
rect 113910 2048 113916 2060
rect 113968 2048 113974 2100
rect 114002 2048 114008 2100
rect 114060 2088 114066 2100
rect 115201 2091 115259 2097
rect 115201 2088 115213 2091
rect 114060 2060 115213 2088
rect 114060 2048 114066 2060
rect 115201 2057 115213 2060
rect 115247 2057 115259 2091
rect 116210 2088 116216 2100
rect 116171 2060 116216 2088
rect 115201 2051 115259 2057
rect 116210 2048 116216 2060
rect 116268 2048 116274 2100
rect 117409 2091 117467 2097
rect 117409 2057 117421 2091
rect 117455 2088 117467 2091
rect 117590 2088 117596 2100
rect 117455 2060 117596 2088
rect 117455 2057 117467 2060
rect 117409 2051 117467 2057
rect 117590 2048 117596 2060
rect 117648 2048 117654 2100
rect 118602 2048 118608 2100
rect 118660 2088 118666 2100
rect 118660 2060 120212 2088
rect 118660 2048 118666 2060
rect 101217 2023 101275 2029
rect 101217 2020 101229 2023
rect 95528 1992 99972 2020
rect 100036 1992 101229 2020
rect 69842 1912 69848 1964
rect 69900 1952 69906 1964
rect 74169 1955 74227 1961
rect 74169 1952 74181 1955
rect 69900 1924 74181 1952
rect 69900 1912 69906 1924
rect 74169 1921 74181 1924
rect 74215 1921 74227 1955
rect 81710 1952 81716 1964
rect 74169 1915 74227 1921
rect 76668 1924 81716 1952
rect 66254 1884 66260 1896
rect 65199 1856 66116 1884
rect 66215 1856 66260 1884
rect 65199 1853 65211 1856
rect 65153 1847 65211 1853
rect 54720 1788 57376 1816
rect 61105 1819 61163 1825
rect 54720 1776 54726 1788
rect 61105 1785 61117 1819
rect 61151 1816 61163 1819
rect 62942 1816 62948 1828
rect 61151 1788 62948 1816
rect 61151 1785 61163 1788
rect 61105 1779 61163 1785
rect 62942 1776 62948 1788
rect 63000 1776 63006 1828
rect 36780 1720 41092 1748
rect 36780 1708 36786 1720
rect 43530 1708 43536 1760
rect 43588 1748 43594 1760
rect 47026 1748 47032 1760
rect 43588 1720 47032 1748
rect 43588 1708 43594 1720
rect 47026 1708 47032 1720
rect 47084 1708 47090 1760
rect 63420 1748 63448 1847
rect 66254 1844 66260 1856
rect 66312 1844 66318 1896
rect 68922 1884 68928 1896
rect 68883 1856 68928 1884
rect 68922 1844 68928 1856
rect 68980 1844 68986 1896
rect 70578 1884 70584 1896
rect 70539 1856 70584 1884
rect 70578 1844 70584 1856
rect 70636 1844 70642 1896
rect 72418 1884 72424 1896
rect 72379 1856 72424 1884
rect 72418 1844 72424 1856
rect 72476 1844 72482 1896
rect 73522 1844 73528 1896
rect 73580 1884 73586 1896
rect 76668 1893 76696 1924
rect 81710 1912 81716 1924
rect 81768 1912 81774 1964
rect 83016 1952 83044 1980
rect 93026 1952 93032 1964
rect 82004 1924 83044 1952
rect 83108 1924 93032 1952
rect 74261 1887 74319 1893
rect 74261 1884 74273 1887
rect 73580 1856 74273 1884
rect 73580 1844 73586 1856
rect 74261 1853 74273 1856
rect 74307 1853 74319 1887
rect 74261 1847 74319 1853
rect 76653 1887 76711 1893
rect 76653 1853 76665 1887
rect 76699 1853 76711 1887
rect 78214 1884 78220 1896
rect 78175 1856 78220 1884
rect 76653 1847 76711 1853
rect 78214 1844 78220 1856
rect 78272 1844 78278 1896
rect 80146 1884 80152 1896
rect 80107 1856 80152 1884
rect 80146 1844 80152 1856
rect 80204 1844 80210 1896
rect 82004 1893 82032 1924
rect 81989 1887 82047 1893
rect 81989 1853 82001 1887
rect 82035 1853 82047 1887
rect 81989 1847 82047 1853
rect 82170 1844 82176 1896
rect 82228 1884 82234 1896
rect 83108 1884 83136 1924
rect 93026 1912 93032 1924
rect 93084 1912 93090 1964
rect 95528 1961 95556 1992
rect 95513 1955 95571 1961
rect 95513 1921 95525 1955
rect 95559 1921 95571 1955
rect 96246 1952 96252 1964
rect 95513 1915 95571 1921
rect 95620 1924 96252 1952
rect 82228 1856 83136 1884
rect 83553 1887 83611 1893
rect 82228 1844 82234 1856
rect 83553 1853 83565 1887
rect 83599 1884 83611 1887
rect 84654 1884 84660 1896
rect 83599 1856 84660 1884
rect 83599 1853 83611 1856
rect 83553 1847 83611 1853
rect 84654 1844 84660 1856
rect 84712 1844 84718 1896
rect 85850 1884 85856 1896
rect 85811 1856 85856 1884
rect 85850 1844 85856 1856
rect 85908 1844 85914 1896
rect 87785 1887 87843 1893
rect 87785 1853 87797 1887
rect 87831 1884 87843 1887
rect 88426 1884 88432 1896
rect 87831 1856 88432 1884
rect 87831 1853 87843 1856
rect 87785 1847 87843 1853
rect 88426 1844 88432 1856
rect 88484 1844 88490 1896
rect 88794 1884 88800 1896
rect 88755 1856 88800 1884
rect 88794 1844 88800 1856
rect 88852 1844 88858 1896
rect 91370 1884 91376 1896
rect 91331 1856 91376 1884
rect 91370 1844 91376 1856
rect 91428 1844 91434 1896
rect 92842 1884 92848 1896
rect 92803 1856 92848 1884
rect 92842 1844 92848 1856
rect 92900 1844 92906 1896
rect 95421 1887 95479 1893
rect 95421 1853 95433 1887
rect 95467 1884 95479 1887
rect 95620 1884 95648 1924
rect 96246 1912 96252 1924
rect 96304 1912 96310 1964
rect 99193 1955 99251 1961
rect 99193 1921 99205 1955
rect 99239 1952 99251 1955
rect 99944 1952 99972 1992
rect 101217 1989 101229 1992
rect 101263 1989 101275 2023
rect 101217 1983 101275 1989
rect 105446 1980 105452 2032
rect 105504 2020 105510 2032
rect 108114 2020 108120 2032
rect 105504 1992 108120 2020
rect 105504 1980 105510 1992
rect 108114 1980 108120 1992
rect 108172 1980 108178 2032
rect 108776 2020 108804 2048
rect 110874 2020 110880 2032
rect 108776 1992 110880 2020
rect 110874 1980 110880 1992
rect 110932 1980 110938 2032
rect 110966 1980 110972 2032
rect 111024 2020 111030 2032
rect 113358 2020 113364 2032
rect 111024 1992 113364 2020
rect 111024 1980 111030 1992
rect 113358 1980 113364 1992
rect 113416 1980 113422 2032
rect 119982 2020 119988 2032
rect 113468 1992 119988 2020
rect 100846 1952 100852 1964
rect 99239 1924 99880 1952
rect 99944 1924 100852 1952
rect 99239 1921 99251 1924
rect 99193 1915 99251 1921
rect 95467 1856 95648 1884
rect 95467 1853 95479 1856
rect 95421 1847 95479 1853
rect 95970 1844 95976 1896
rect 96028 1884 96034 1896
rect 96709 1887 96767 1893
rect 96709 1884 96721 1887
rect 96028 1856 96721 1884
rect 96028 1844 96034 1856
rect 96709 1853 96721 1856
rect 96755 1853 96767 1887
rect 96709 1847 96767 1853
rect 97074 1844 97080 1896
rect 97132 1884 97138 1896
rect 98549 1887 98607 1893
rect 98549 1884 98561 1887
rect 97132 1856 98561 1884
rect 97132 1844 97138 1856
rect 98549 1853 98561 1856
rect 98595 1853 98607 1887
rect 98549 1847 98607 1853
rect 63770 1776 63776 1828
rect 63828 1816 63834 1828
rect 66073 1819 66131 1825
rect 66073 1816 66085 1819
rect 63828 1788 66085 1816
rect 63828 1776 63834 1788
rect 66073 1785 66085 1788
rect 66119 1785 66131 1819
rect 66073 1779 66131 1785
rect 66162 1776 66168 1828
rect 66220 1816 66226 1828
rect 68557 1819 68615 1825
rect 68557 1816 68569 1819
rect 66220 1788 68569 1816
rect 66220 1776 66226 1788
rect 68557 1785 68569 1788
rect 68603 1785 68615 1819
rect 68557 1779 68615 1785
rect 69566 1776 69572 1828
rect 69624 1816 69630 1828
rect 70489 1819 70547 1825
rect 70489 1816 70501 1819
rect 69624 1788 70501 1816
rect 69624 1776 69630 1788
rect 70489 1785 70501 1788
rect 70535 1785 70547 1819
rect 70489 1779 70547 1785
rect 70762 1776 70768 1828
rect 70820 1816 70826 1828
rect 72053 1819 72111 1825
rect 72053 1816 72065 1819
rect 70820 1788 72065 1816
rect 70820 1776 70826 1788
rect 72053 1785 72065 1788
rect 72099 1785 72111 1819
rect 72053 1779 72111 1785
rect 76745 1819 76803 1825
rect 76745 1785 76757 1819
rect 76791 1816 76803 1819
rect 77754 1816 77760 1828
rect 76791 1788 77760 1816
rect 76791 1785 76803 1788
rect 76745 1779 76803 1785
rect 77754 1776 77760 1788
rect 77812 1776 77818 1828
rect 89441 1819 89499 1825
rect 89441 1785 89453 1819
rect 89487 1816 89499 1819
rect 89898 1816 89904 1828
rect 89487 1788 89904 1816
rect 89487 1785 89499 1788
rect 89441 1779 89499 1785
rect 89898 1776 89904 1788
rect 89956 1776 89962 1828
rect 91741 1819 91799 1825
rect 91741 1785 91753 1819
rect 91787 1816 91799 1819
rect 92934 1816 92940 1828
rect 91787 1788 92940 1816
rect 91787 1785 91799 1788
rect 91741 1779 91799 1785
rect 92934 1776 92940 1788
rect 92992 1776 92998 1828
rect 93305 1819 93363 1825
rect 93305 1785 93317 1819
rect 93351 1816 93363 1819
rect 96430 1816 96436 1828
rect 93351 1788 96436 1816
rect 93351 1785 93363 1788
rect 93305 1779 93363 1785
rect 96430 1776 96436 1788
rect 96488 1776 96494 1828
rect 97353 1819 97411 1825
rect 97353 1785 97365 1819
rect 97399 1816 97411 1819
rect 98178 1816 98184 1828
rect 97399 1788 98184 1816
rect 97399 1785 97411 1788
rect 97353 1779 97411 1785
rect 98178 1776 98184 1788
rect 98236 1776 98242 1828
rect 98270 1776 98276 1828
rect 98328 1816 98334 1828
rect 99852 1816 99880 1924
rect 100846 1912 100852 1924
rect 100904 1912 100910 1964
rect 105357 1955 105415 1961
rect 105357 1921 105369 1955
rect 105403 1952 105415 1955
rect 106642 1952 106648 1964
rect 105403 1924 106648 1952
rect 105403 1921 105415 1924
rect 105357 1915 105415 1921
rect 106642 1912 106648 1924
rect 106700 1912 106706 1964
rect 107746 1912 107752 1964
rect 107804 1952 107810 1964
rect 108577 1955 108635 1961
rect 107804 1924 108344 1952
rect 107804 1912 107810 1924
rect 100113 1887 100171 1893
rect 100113 1853 100125 1887
rect 100159 1884 100171 1887
rect 100159 1856 101076 1884
rect 100159 1853 100171 1856
rect 100113 1847 100171 1853
rect 100662 1816 100668 1828
rect 98328 1788 99788 1816
rect 99852 1788 100668 1816
rect 98328 1776 98334 1788
rect 66898 1748 66904 1760
rect 63420 1720 66904 1748
rect 66898 1708 66904 1720
rect 66956 1708 66962 1760
rect 78033 1751 78091 1757
rect 78033 1717 78045 1751
rect 78079 1748 78091 1751
rect 78122 1748 78128 1760
rect 78079 1720 78128 1748
rect 78079 1717 78091 1720
rect 78033 1711 78091 1717
rect 78122 1708 78128 1720
rect 78180 1708 78186 1760
rect 79870 1708 79876 1760
rect 79928 1748 79934 1760
rect 80057 1751 80115 1757
rect 80057 1748 80069 1751
rect 79928 1720 80069 1748
rect 79928 1708 79934 1720
rect 80057 1717 80069 1720
rect 80103 1717 80115 1751
rect 81618 1748 81624 1760
rect 81579 1720 81624 1748
rect 80057 1711 80115 1717
rect 81618 1708 81624 1720
rect 81676 1708 81682 1760
rect 83366 1748 83372 1760
rect 83327 1720 83372 1748
rect 83366 1708 83372 1720
rect 83424 1708 83430 1760
rect 85574 1708 85580 1760
rect 85632 1748 85638 1760
rect 85669 1751 85727 1757
rect 85669 1748 85681 1751
rect 85632 1720 85681 1748
rect 85632 1708 85638 1720
rect 85669 1717 85681 1720
rect 85715 1717 85727 1751
rect 85669 1711 85727 1717
rect 87322 1708 87328 1760
rect 87380 1748 87386 1760
rect 87417 1751 87475 1757
rect 87417 1748 87429 1751
rect 87380 1720 87429 1748
rect 87380 1708 87386 1720
rect 87417 1717 87429 1720
rect 87463 1717 87475 1751
rect 87417 1711 87475 1717
rect 93210 1708 93216 1760
rect 93268 1748 93274 1760
rect 96982 1748 96988 1760
rect 93268 1720 96988 1748
rect 93268 1708 93274 1720
rect 96982 1708 96988 1720
rect 97040 1708 97046 1760
rect 99760 1748 99788 1788
rect 100662 1776 100668 1788
rect 100720 1776 100726 1828
rect 101048 1816 101076 1856
rect 101122 1844 101128 1896
rect 101180 1884 101186 1896
rect 102778 1884 102784 1896
rect 101180 1856 101225 1884
rect 102739 1856 102784 1884
rect 101180 1844 101186 1856
rect 102778 1844 102784 1856
rect 102836 1844 102842 1896
rect 102888 1856 105216 1884
rect 102888 1816 102916 1856
rect 101048 1788 102916 1816
rect 102965 1819 103023 1825
rect 102965 1785 102977 1819
rect 103011 1816 103023 1819
rect 104250 1816 104256 1828
rect 103011 1788 104256 1816
rect 103011 1785 103023 1788
rect 102965 1779 103023 1785
rect 104250 1776 104256 1788
rect 104308 1776 104314 1828
rect 105188 1816 105216 1856
rect 105262 1844 105268 1896
rect 105320 1884 105326 1896
rect 106829 1887 106887 1893
rect 105320 1856 105365 1884
rect 105320 1844 105326 1856
rect 106829 1853 106841 1887
rect 106875 1884 106887 1887
rect 107838 1884 107844 1896
rect 106875 1856 107844 1884
rect 106875 1853 106887 1856
rect 106829 1847 106887 1853
rect 107838 1844 107844 1856
rect 107896 1844 107902 1896
rect 106734 1816 106740 1828
rect 105188 1788 106740 1816
rect 106734 1776 106740 1788
rect 106792 1776 106798 1828
rect 106921 1819 106979 1825
rect 106921 1785 106933 1819
rect 106967 1816 106979 1819
rect 108206 1816 108212 1828
rect 106967 1788 108212 1816
rect 106967 1785 106979 1788
rect 106921 1779 106979 1785
rect 108206 1776 108212 1788
rect 108264 1776 108270 1828
rect 108316 1816 108344 1924
rect 108577 1921 108589 1955
rect 108623 1952 108635 1955
rect 108623 1924 108988 1952
rect 108623 1921 108635 1924
rect 108577 1915 108635 1921
rect 108482 1884 108488 1896
rect 108443 1856 108488 1884
rect 108482 1844 108488 1856
rect 108540 1844 108546 1896
rect 108960 1884 108988 1924
rect 109954 1884 109960 1896
rect 108960 1856 109960 1884
rect 109954 1844 109960 1856
rect 110012 1844 110018 1896
rect 110325 1887 110383 1893
rect 110325 1853 110337 1887
rect 110371 1884 110383 1887
rect 110782 1884 110788 1896
rect 110371 1856 110788 1884
rect 110371 1853 110383 1856
rect 110325 1847 110383 1853
rect 110782 1844 110788 1856
rect 110840 1844 110846 1896
rect 111981 1887 112039 1893
rect 111981 1853 111993 1887
rect 112027 1853 112039 1887
rect 111981 1847 112039 1853
rect 109773 1819 109831 1825
rect 109773 1816 109785 1819
rect 108316 1788 109785 1816
rect 109773 1785 109785 1788
rect 109819 1785 109831 1819
rect 109773 1779 109831 1785
rect 110414 1776 110420 1828
rect 110472 1816 110478 1828
rect 111702 1816 111708 1828
rect 110472 1788 111708 1816
rect 110472 1776 110478 1788
rect 111702 1776 111708 1788
rect 111760 1776 111766 1828
rect 111996 1816 112024 1847
rect 112070 1844 112076 1896
rect 112128 1884 112134 1896
rect 113468 1893 113496 1992
rect 119982 1980 119988 1992
rect 120040 1980 120046 2032
rect 120184 2020 120212 2060
rect 120258 2048 120264 2100
rect 120316 2088 120322 2100
rect 123573 2091 123631 2097
rect 120316 2060 120361 2088
rect 120316 2048 120322 2060
rect 123573 2057 123585 2091
rect 123619 2088 123631 2091
rect 124490 2088 124496 2100
rect 123619 2060 124496 2088
rect 123619 2057 123631 2060
rect 123573 2051 123631 2057
rect 124490 2048 124496 2060
rect 124548 2048 124554 2100
rect 124769 2091 124827 2097
rect 124769 2057 124781 2091
rect 124815 2088 124827 2091
rect 124858 2088 124864 2100
rect 124815 2060 124864 2088
rect 124815 2057 124827 2060
rect 124769 2051 124827 2057
rect 124858 2048 124864 2060
rect 124916 2048 124922 2100
rect 125318 2048 125324 2100
rect 125376 2088 125382 2100
rect 126514 2088 126520 2100
rect 125376 2060 126520 2088
rect 125376 2048 125382 2060
rect 126514 2048 126520 2060
rect 126572 2048 126578 2100
rect 126701 2091 126759 2097
rect 126701 2057 126713 2091
rect 126747 2088 126759 2091
rect 126790 2088 126796 2100
rect 126747 2060 126796 2088
rect 126747 2057 126759 2060
rect 126701 2051 126759 2057
rect 126790 2048 126796 2060
rect 126848 2048 126854 2100
rect 127802 2048 127808 2100
rect 127860 2088 127866 2100
rect 129093 2091 129151 2097
rect 129093 2088 129105 2091
rect 127860 2060 129105 2088
rect 127860 2048 127866 2060
rect 129093 2057 129105 2060
rect 129139 2057 129151 2091
rect 132862 2088 132868 2100
rect 129093 2051 129151 2057
rect 131224 2060 132724 2088
rect 132823 2060 132868 2088
rect 122561 2023 122619 2029
rect 122561 2020 122573 2023
rect 120184 1992 122573 2020
rect 122561 1989 122573 1992
rect 122607 1989 122619 2023
rect 122561 1983 122619 1989
rect 122834 1980 122840 2032
rect 122892 2020 122898 2032
rect 125873 2023 125931 2029
rect 125873 2020 125885 2023
rect 122892 1992 125885 2020
rect 122892 1980 122898 1992
rect 125873 1989 125885 1992
rect 125919 1989 125931 2023
rect 131022 2020 131028 2032
rect 125873 1983 125931 1989
rect 128924 1992 131028 2020
rect 113542 1912 113548 1964
rect 113600 1952 113606 1964
rect 113600 1924 113645 1952
rect 113600 1912 113606 1924
rect 113818 1912 113824 1964
rect 113876 1952 113882 1964
rect 117130 1952 117136 1964
rect 113876 1924 117136 1952
rect 113876 1912 113882 1924
rect 117130 1912 117136 1924
rect 117188 1912 117194 1964
rect 117225 1955 117283 1961
rect 117225 1921 117237 1955
rect 117271 1952 117283 1955
rect 118326 1952 118332 1964
rect 117271 1924 118332 1952
rect 117271 1921 117283 1924
rect 117225 1915 117283 1921
rect 113453 1887 113511 1893
rect 112128 1856 112173 1884
rect 112128 1844 112134 1856
rect 113453 1853 113465 1887
rect 113499 1853 113511 1887
rect 113453 1847 113511 1853
rect 113634 1844 113640 1896
rect 113692 1884 113698 1896
rect 114462 1884 114468 1896
rect 113692 1856 114468 1884
rect 113692 1844 113698 1856
rect 114462 1844 114468 1856
rect 114520 1844 114526 1896
rect 115106 1884 115112 1896
rect 115067 1856 115112 1884
rect 115106 1844 115112 1856
rect 115164 1844 115170 1896
rect 115198 1844 115204 1896
rect 115256 1844 115262 1896
rect 117332 1893 117360 1924
rect 118326 1912 118332 1924
rect 118384 1912 118390 1964
rect 128170 1952 128176 1964
rect 118436 1924 128176 1952
rect 116121 1887 116179 1893
rect 116121 1853 116133 1887
rect 116167 1884 116179 1887
rect 117317 1887 117375 1893
rect 116167 1856 117268 1884
rect 116167 1853 116179 1856
rect 116121 1847 116179 1853
rect 115216 1816 115244 1844
rect 111996 1788 115244 1816
rect 117240 1816 117268 1856
rect 117317 1853 117329 1887
rect 117363 1884 117375 1887
rect 117363 1856 117397 1884
rect 117363 1853 117375 1856
rect 117317 1847 117375 1853
rect 118050 1844 118056 1896
rect 118108 1884 118114 1896
rect 118436 1884 118464 1924
rect 128170 1912 128176 1924
rect 128228 1912 128234 1964
rect 118602 1884 118608 1896
rect 118108 1856 118464 1884
rect 118528 1856 118608 1884
rect 118108 1844 118114 1856
rect 118528 1816 118556 1856
rect 118602 1844 118608 1856
rect 118660 1844 118666 1896
rect 119065 1887 119123 1893
rect 119065 1853 119077 1887
rect 119111 1884 119123 1887
rect 119890 1884 119896 1896
rect 119111 1856 119896 1884
rect 119111 1853 119123 1856
rect 119065 1847 119123 1853
rect 119890 1844 119896 1856
rect 119948 1844 119954 1896
rect 120169 1887 120227 1893
rect 120169 1853 120181 1887
rect 120215 1853 120227 1887
rect 120169 1847 120227 1853
rect 121181 1887 121239 1893
rect 121181 1853 121193 1887
rect 121227 1853 121239 1887
rect 121181 1847 121239 1853
rect 122469 1887 122527 1893
rect 122469 1853 122481 1887
rect 122515 1884 122527 1887
rect 123481 1887 123539 1893
rect 122515 1856 123432 1884
rect 122515 1853 122527 1856
rect 122469 1847 122527 1853
rect 119154 1816 119160 1828
rect 117240 1788 118556 1816
rect 119115 1788 119160 1816
rect 119154 1776 119160 1788
rect 119212 1776 119218 1828
rect 120074 1816 120080 1828
rect 120035 1788 120080 1816
rect 120074 1776 120080 1788
rect 120132 1816 120138 1828
rect 120184 1816 120212 1847
rect 120132 1788 120212 1816
rect 121196 1816 121224 1847
rect 123018 1816 123024 1828
rect 121196 1788 123024 1816
rect 120132 1776 120138 1788
rect 123018 1776 123024 1788
rect 123076 1776 123082 1828
rect 123404 1816 123432 1856
rect 123481 1853 123493 1887
rect 123527 1884 123539 1887
rect 123938 1884 123944 1896
rect 123527 1856 123944 1884
rect 123527 1853 123539 1856
rect 123481 1847 123539 1853
rect 123938 1844 123944 1856
rect 123996 1844 124002 1896
rect 124677 1887 124735 1893
rect 124677 1853 124689 1887
rect 124723 1884 124735 1887
rect 125689 1887 125747 1893
rect 124723 1856 125088 1884
rect 124723 1853 124735 1856
rect 124677 1847 124735 1853
rect 124950 1816 124956 1828
rect 123404 1788 124956 1816
rect 124950 1776 124956 1788
rect 125008 1776 125014 1828
rect 125060 1760 125088 1856
rect 125689 1853 125701 1887
rect 125735 1884 125747 1887
rect 125778 1884 125784 1896
rect 125735 1856 125784 1884
rect 125735 1853 125747 1856
rect 125689 1847 125747 1853
rect 125778 1844 125784 1856
rect 125836 1844 125842 1896
rect 126790 1884 126796 1896
rect 126751 1856 126796 1884
rect 126790 1844 126796 1856
rect 126848 1844 126854 1896
rect 126882 1844 126888 1896
rect 126940 1884 126946 1896
rect 127989 1887 128047 1893
rect 126940 1856 126985 1884
rect 126940 1844 126946 1856
rect 127989 1853 128001 1887
rect 128035 1884 128047 1887
rect 128924 1884 128952 1992
rect 131022 1980 131028 1992
rect 131080 1980 131086 2032
rect 131224 1952 131252 2060
rect 131298 1980 131304 2032
rect 131356 2020 131362 2032
rect 131758 2020 131764 2032
rect 131356 1992 131764 2020
rect 131356 1980 131362 1992
rect 131758 1980 131764 1992
rect 131816 1980 131822 2032
rect 132696 2020 132724 2060
rect 132862 2048 132868 2060
rect 132920 2048 132926 2100
rect 133877 2091 133935 2097
rect 133877 2057 133889 2091
rect 133923 2088 133935 2091
rect 133966 2088 133972 2100
rect 133923 2060 133972 2088
rect 133923 2057 133935 2060
rect 133877 2051 133935 2057
rect 133966 2048 133972 2060
rect 134024 2048 134030 2100
rect 134058 2048 134064 2100
rect 134116 2088 134122 2100
rect 136726 2088 136732 2100
rect 134116 2060 136732 2088
rect 134116 2048 134122 2060
rect 136726 2048 136732 2060
rect 136784 2048 136790 2100
rect 137465 2091 137523 2097
rect 137465 2057 137477 2091
rect 137511 2088 137523 2091
rect 137554 2088 137560 2100
rect 137511 2060 137560 2088
rect 137511 2057 137523 2060
rect 137465 2051 137523 2057
rect 137554 2048 137560 2060
rect 137612 2048 137618 2100
rect 137646 2048 137652 2100
rect 137704 2088 137710 2100
rect 138477 2091 138535 2097
rect 138477 2088 138489 2091
rect 137704 2060 138489 2088
rect 137704 2048 137710 2060
rect 138477 2057 138489 2060
rect 138523 2057 138535 2091
rect 138477 2051 138535 2057
rect 138566 2048 138572 2100
rect 138624 2088 138630 2100
rect 139489 2091 139547 2097
rect 139489 2088 139501 2091
rect 138624 2060 139501 2088
rect 138624 2048 138630 2060
rect 139489 2057 139501 2060
rect 139535 2057 139547 2091
rect 139489 2051 139547 2057
rect 139578 2048 139584 2100
rect 139636 2088 139642 2100
rect 140501 2091 140559 2097
rect 140501 2088 140513 2091
rect 139636 2060 140513 2088
rect 139636 2048 139642 2060
rect 140501 2057 140513 2060
rect 140547 2057 140559 2091
rect 140501 2051 140559 2057
rect 143350 2048 143356 2100
rect 143408 2088 143414 2100
rect 145009 2091 145067 2097
rect 145009 2088 145021 2091
rect 143408 2060 145021 2088
rect 143408 2048 143414 2060
rect 145009 2057 145021 2060
rect 145055 2057 145067 2091
rect 146113 2091 146171 2097
rect 146113 2088 146125 2091
rect 145009 2051 145067 2057
rect 145116 2060 146125 2088
rect 137738 2020 137744 2032
rect 132696 1992 137744 2020
rect 137738 1980 137744 1992
rect 137796 1980 137802 2032
rect 137830 1980 137836 2032
rect 137888 2020 137894 2032
rect 143997 2023 144055 2029
rect 143997 2020 144009 2023
rect 137888 1992 144009 2020
rect 137888 1980 137894 1992
rect 143997 1989 144009 1992
rect 144043 1989 144055 2023
rect 143997 1983 144055 1989
rect 144178 1980 144184 2032
rect 144236 2020 144242 2032
rect 144236 1992 144408 2020
rect 144236 1980 144242 1992
rect 138198 1952 138204 1964
rect 129016 1924 131252 1952
rect 131316 1924 138204 1952
rect 129016 1893 129044 1924
rect 128035 1856 128952 1884
rect 129001 1887 129059 1893
rect 128035 1853 128047 1856
rect 127989 1847 128047 1853
rect 129001 1853 129013 1887
rect 129047 1853 129059 1887
rect 130286 1884 130292 1896
rect 130247 1856 130292 1884
rect 129001 1847 129059 1853
rect 130286 1844 130292 1856
rect 130344 1844 130350 1896
rect 131206 1884 131212 1896
rect 130396 1856 131212 1884
rect 125318 1776 125324 1828
rect 125376 1816 125382 1828
rect 125376 1788 127020 1816
rect 125376 1776 125382 1788
rect 104526 1748 104532 1760
rect 99760 1720 104532 1748
rect 104526 1708 104532 1720
rect 104584 1708 104590 1760
rect 104618 1708 104624 1760
rect 104676 1748 104682 1760
rect 108758 1748 108764 1760
rect 104676 1720 108764 1748
rect 104676 1708 104682 1720
rect 108758 1708 108764 1720
rect 108816 1708 108822 1760
rect 110598 1708 110604 1760
rect 110656 1748 110662 1760
rect 114278 1748 114284 1760
rect 110656 1720 114284 1748
rect 110656 1708 110662 1720
rect 114278 1708 114284 1720
rect 114336 1708 114342 1760
rect 114370 1708 114376 1760
rect 114428 1748 114434 1760
rect 116026 1748 116032 1760
rect 114428 1720 116032 1748
rect 114428 1708 114434 1720
rect 116026 1708 116032 1720
rect 116084 1708 116090 1760
rect 116118 1708 116124 1760
rect 116176 1748 116182 1760
rect 121273 1751 121331 1757
rect 121273 1748 121285 1751
rect 116176 1720 121285 1748
rect 116176 1708 116182 1720
rect 121273 1717 121285 1720
rect 121319 1717 121331 1751
rect 121273 1711 121331 1717
rect 121914 1708 121920 1760
rect 121972 1748 121978 1760
rect 124674 1748 124680 1760
rect 121972 1720 124680 1748
rect 121972 1708 121978 1720
rect 124674 1708 124680 1720
rect 124732 1708 124738 1760
rect 125042 1748 125048 1760
rect 125003 1720 125048 1748
rect 125042 1708 125048 1720
rect 125100 1708 125106 1760
rect 126992 1748 127020 1788
rect 129182 1776 129188 1828
rect 129240 1816 129246 1828
rect 130396 1816 130424 1856
rect 131206 1844 131212 1856
rect 131264 1844 131270 1896
rect 131316 1893 131344 1924
rect 138198 1912 138204 1924
rect 138256 1912 138262 1964
rect 140038 1952 140044 1964
rect 138400 1924 140044 1952
rect 131301 1887 131359 1893
rect 131301 1853 131313 1887
rect 131347 1853 131359 1887
rect 131301 1847 131359 1853
rect 132773 1887 132831 1893
rect 132773 1853 132785 1887
rect 132819 1884 132831 1887
rect 133690 1884 133696 1896
rect 132819 1856 133696 1884
rect 132819 1853 132831 1856
rect 132773 1847 132831 1853
rect 133690 1844 133696 1856
rect 133748 1844 133754 1896
rect 133785 1887 133843 1893
rect 133785 1853 133797 1887
rect 133831 1884 133843 1887
rect 133874 1884 133880 1896
rect 133831 1856 133880 1884
rect 133831 1853 133843 1856
rect 133785 1847 133843 1853
rect 133874 1844 133880 1856
rect 133932 1844 133938 1896
rect 134610 1884 134616 1896
rect 133984 1856 134616 1884
rect 129240 1788 130424 1816
rect 129240 1776 129246 1788
rect 130746 1776 130752 1828
rect 130804 1816 130810 1828
rect 131393 1819 131451 1825
rect 131393 1816 131405 1819
rect 130804 1788 131405 1816
rect 130804 1776 130810 1788
rect 131393 1785 131405 1788
rect 131439 1785 131451 1819
rect 131393 1779 131451 1785
rect 131666 1776 131672 1828
rect 131724 1816 131730 1828
rect 133984 1816 134012 1856
rect 134610 1844 134616 1856
rect 134668 1844 134674 1896
rect 134794 1884 134800 1896
rect 134755 1856 134800 1884
rect 134794 1844 134800 1856
rect 134852 1844 134858 1896
rect 135346 1844 135352 1896
rect 135404 1884 135410 1896
rect 135806 1884 135812 1896
rect 135404 1856 135812 1884
rect 135404 1844 135410 1856
rect 135806 1844 135812 1856
rect 135864 1844 135870 1896
rect 135901 1887 135959 1893
rect 135901 1853 135913 1887
rect 135947 1853 135959 1887
rect 135901 1847 135959 1853
rect 131724 1788 134012 1816
rect 131724 1776 131730 1788
rect 134242 1776 134248 1828
rect 134300 1816 134306 1828
rect 135916 1816 135944 1847
rect 135990 1844 135996 1896
rect 136048 1884 136054 1896
rect 137278 1884 137284 1896
rect 136048 1856 137284 1884
rect 136048 1844 136054 1856
rect 137278 1844 137284 1856
rect 137336 1844 137342 1896
rect 138400 1893 138428 1924
rect 140038 1912 140044 1924
rect 140096 1912 140102 1964
rect 140130 1912 140136 1964
rect 140188 1952 140194 1964
rect 144270 1952 144276 1964
rect 140188 1924 144276 1952
rect 140188 1912 140194 1924
rect 144270 1912 144276 1924
rect 144328 1912 144334 1964
rect 144380 1952 144408 1992
rect 144454 1980 144460 2032
rect 144512 2020 144518 2032
rect 145116 2020 145144 2060
rect 146113 2057 146125 2060
rect 146159 2057 146171 2091
rect 146113 2051 146171 2057
rect 147122 2048 147128 2100
rect 147180 2088 147186 2100
rect 147217 2091 147275 2097
rect 147217 2088 147229 2091
rect 147180 2060 147229 2088
rect 147180 2048 147186 2060
rect 147217 2057 147229 2060
rect 147263 2057 147275 2091
rect 147217 2051 147275 2057
rect 147306 2048 147312 2100
rect 147364 2088 147370 2100
rect 148229 2091 148287 2097
rect 148229 2088 148241 2091
rect 147364 2060 148241 2088
rect 147364 2048 147370 2060
rect 148229 2057 148241 2060
rect 148275 2057 148287 2091
rect 148229 2051 148287 2057
rect 148870 2048 148876 2100
rect 148928 2088 148934 2100
rect 153197 2091 153255 2097
rect 148928 2060 150204 2088
rect 148928 2048 148934 2060
rect 146938 2020 146944 2032
rect 144512 1992 145144 2020
rect 145852 1992 146944 2020
rect 144512 1980 144518 1992
rect 145852 1952 145880 1992
rect 146938 1980 146944 1992
rect 146996 1980 147002 2032
rect 147398 1980 147404 2032
rect 147456 2020 147462 2032
rect 150066 2020 150072 2032
rect 147456 1992 150072 2020
rect 147456 1980 147462 1992
rect 150066 1980 150072 1992
rect 150124 1980 150130 2032
rect 150176 2020 150204 2060
rect 153197 2057 153209 2091
rect 153243 2088 153255 2091
rect 153470 2088 153476 2100
rect 153243 2060 153476 2088
rect 153243 2057 153255 2060
rect 153197 2051 153255 2057
rect 153470 2048 153476 2060
rect 153528 2048 153534 2100
rect 159358 2088 159364 2100
rect 153580 2060 159364 2088
rect 153580 2020 153608 2060
rect 159358 2048 159364 2060
rect 159416 2048 159422 2100
rect 159450 2048 159456 2100
rect 159508 2088 159514 2100
rect 160830 2088 160836 2100
rect 159508 2060 159680 2088
rect 160791 2060 160836 2088
rect 159508 2048 159514 2060
rect 150176 1992 153608 2020
rect 153838 1980 153844 2032
rect 153896 2020 153902 2032
rect 155678 2020 155684 2032
rect 153896 1992 155684 2020
rect 153896 1980 153902 1992
rect 155678 1980 155684 1992
rect 155736 1980 155742 2032
rect 159542 2020 159548 2032
rect 155788 1992 159548 2020
rect 150894 1952 150900 1964
rect 144380 1924 145880 1952
rect 146220 1924 147260 1952
rect 137373 1887 137431 1893
rect 137373 1853 137385 1887
rect 137419 1884 137431 1887
rect 138385 1887 138443 1893
rect 137419 1856 138336 1884
rect 137419 1853 137431 1856
rect 137373 1847 137431 1853
rect 138014 1816 138020 1828
rect 134300 1788 135024 1816
rect 135916 1788 138020 1816
rect 134300 1776 134306 1788
rect 128081 1751 128139 1757
rect 128081 1748 128093 1751
rect 126992 1720 128093 1748
rect 128081 1717 128093 1720
rect 128127 1717 128139 1751
rect 128081 1711 128139 1717
rect 128170 1708 128176 1760
rect 128228 1748 128234 1760
rect 129550 1748 129556 1760
rect 128228 1720 129556 1748
rect 128228 1708 128234 1720
rect 129550 1708 129556 1720
rect 129608 1708 129614 1760
rect 130381 1751 130439 1757
rect 130381 1717 130393 1751
rect 130427 1748 130439 1751
rect 134150 1748 134156 1760
rect 130427 1720 134156 1748
rect 130427 1717 130439 1720
rect 130381 1711 130439 1717
rect 134150 1708 134156 1720
rect 134208 1708 134214 1760
rect 134610 1708 134616 1760
rect 134668 1748 134674 1760
rect 134889 1751 134947 1757
rect 134889 1748 134901 1751
rect 134668 1720 134901 1748
rect 134668 1708 134674 1720
rect 134889 1717 134901 1720
rect 134935 1717 134947 1751
rect 134996 1748 135024 1788
rect 138014 1776 138020 1788
rect 138072 1776 138078 1828
rect 138308 1816 138336 1856
rect 138385 1853 138397 1887
rect 138431 1853 138443 1887
rect 139210 1884 139216 1896
rect 138385 1847 138443 1853
rect 138676 1856 139216 1884
rect 138676 1816 138704 1856
rect 139210 1844 139216 1856
rect 139268 1844 139274 1896
rect 139397 1887 139455 1893
rect 139397 1853 139409 1887
rect 139443 1884 139455 1887
rect 140409 1887 140467 1893
rect 139443 1856 140360 1884
rect 139443 1853 139455 1856
rect 139397 1847 139455 1853
rect 138308 1788 138704 1816
rect 138842 1776 138848 1828
rect 138900 1816 138906 1828
rect 139670 1816 139676 1828
rect 138900 1788 139676 1816
rect 138900 1776 138906 1788
rect 139670 1776 139676 1788
rect 139728 1776 139734 1828
rect 140332 1816 140360 1856
rect 140409 1853 140421 1887
rect 140455 1884 140467 1887
rect 143905 1887 143963 1893
rect 140455 1856 143856 1884
rect 140455 1853 140467 1856
rect 140409 1847 140467 1853
rect 140866 1816 140872 1828
rect 140332 1788 140872 1816
rect 140866 1776 140872 1788
rect 140924 1776 140930 1828
rect 143828 1816 143856 1856
rect 143905 1853 143917 1887
rect 143951 1884 143963 1887
rect 144730 1884 144736 1896
rect 143951 1856 144736 1884
rect 143951 1853 143963 1856
rect 143905 1847 143963 1853
rect 144730 1844 144736 1856
rect 144788 1844 144794 1896
rect 144917 1887 144975 1893
rect 144917 1853 144929 1887
rect 144963 1884 144975 1887
rect 145466 1884 145472 1896
rect 144963 1856 145472 1884
rect 144963 1853 144975 1856
rect 144917 1847 144975 1853
rect 145466 1844 145472 1856
rect 145524 1844 145530 1896
rect 145558 1844 145564 1896
rect 145616 1884 145622 1896
rect 146021 1887 146079 1893
rect 145616 1856 145880 1884
rect 145616 1844 145622 1856
rect 145282 1816 145288 1828
rect 143828 1788 145288 1816
rect 145282 1776 145288 1788
rect 145340 1776 145346 1828
rect 145852 1816 145880 1856
rect 146021 1853 146033 1887
rect 146067 1884 146079 1887
rect 146220 1884 146248 1924
rect 146067 1856 146248 1884
rect 147125 1887 147183 1893
rect 146067 1853 146079 1856
rect 146021 1847 146079 1853
rect 147125 1853 147137 1887
rect 147171 1853 147183 1887
rect 147232 1884 147260 1924
rect 148060 1924 150900 1952
rect 148060 1884 148088 1924
rect 150894 1912 150900 1924
rect 150952 1912 150958 1964
rect 155218 1952 155224 1964
rect 153120 1924 155224 1952
rect 153120 1893 153148 1924
rect 155218 1912 155224 1924
rect 155276 1912 155282 1964
rect 155788 1893 155816 1992
rect 159542 1980 159548 1992
rect 159600 1980 159606 2032
rect 159652 2020 159680 2060
rect 160830 2048 160836 2060
rect 160888 2048 160894 2100
rect 160922 2048 160928 2100
rect 160980 2088 160986 2100
rect 162394 2088 162400 2100
rect 160980 2060 162400 2088
rect 160980 2048 160986 2060
rect 162394 2048 162400 2060
rect 162452 2048 162458 2100
rect 162504 2060 164464 2088
rect 162504 2020 162532 2060
rect 159652 1992 162532 2020
rect 163222 1980 163228 2032
rect 163280 2020 163286 2032
rect 164326 2020 164332 2032
rect 163280 1992 164332 2020
rect 163280 1980 163286 1992
rect 164326 1980 164332 1992
rect 164384 1980 164390 2032
rect 164436 2020 164464 2060
rect 164510 2048 164516 2100
rect 164568 2088 164574 2100
rect 164568 2060 165936 2088
rect 164568 2048 164574 2060
rect 164436 1992 164924 2020
rect 155865 1955 155923 1961
rect 155865 1921 155877 1955
rect 155911 1952 155923 1955
rect 155954 1952 155960 1964
rect 155911 1924 155960 1952
rect 155911 1921 155923 1924
rect 155865 1915 155923 1921
rect 155954 1912 155960 1924
rect 156012 1912 156018 1964
rect 158714 1952 158720 1964
rect 158675 1924 158720 1952
rect 158714 1912 158720 1924
rect 158772 1912 158778 1964
rect 159726 1952 159732 1964
rect 159687 1924 159732 1952
rect 159726 1912 159732 1924
rect 159784 1912 159790 1964
rect 159818 1912 159824 1964
rect 159876 1952 159882 1964
rect 162210 1952 162216 1964
rect 159876 1924 162216 1952
rect 159876 1912 159882 1924
rect 162210 1912 162216 1924
rect 162268 1912 162274 1964
rect 163777 1955 163835 1961
rect 162688 1924 163728 1952
rect 147232 1856 148088 1884
rect 148137 1887 148195 1893
rect 147125 1847 147183 1853
rect 148137 1853 148149 1887
rect 148183 1884 148195 1887
rect 152461 1887 152519 1893
rect 152461 1884 152473 1887
rect 148183 1856 152473 1884
rect 148183 1853 148195 1856
rect 148137 1847 148195 1853
rect 152461 1853 152473 1856
rect 152507 1853 152519 1887
rect 152461 1847 152519 1853
rect 153105 1887 153163 1893
rect 153105 1853 153117 1887
rect 153151 1853 153163 1887
rect 153105 1847 153163 1853
rect 155773 1887 155831 1893
rect 155773 1853 155785 1887
rect 155819 1853 155831 1887
rect 155773 1847 155831 1853
rect 157245 1887 157303 1893
rect 157245 1853 157257 1887
rect 157291 1884 157303 1887
rect 160554 1884 160560 1896
rect 157291 1856 160560 1884
rect 157291 1853 157303 1856
rect 157245 1847 157303 1853
rect 146846 1816 146852 1828
rect 145852 1788 146852 1816
rect 146846 1776 146852 1788
rect 146904 1776 146910 1828
rect 147140 1816 147168 1847
rect 160554 1844 160560 1856
rect 160612 1844 160618 1896
rect 160738 1884 160744 1896
rect 160699 1856 160744 1884
rect 160738 1844 160744 1856
rect 160796 1844 160802 1896
rect 161106 1844 161112 1896
rect 161164 1884 161170 1896
rect 161566 1884 161572 1896
rect 161164 1856 161572 1884
rect 161164 1844 161170 1856
rect 161566 1844 161572 1856
rect 161624 1844 161630 1896
rect 161750 1884 161756 1896
rect 161711 1856 161756 1884
rect 161750 1844 161756 1856
rect 161808 1844 161814 1896
rect 161845 1887 161903 1893
rect 161845 1853 161857 1887
rect 161891 1884 161903 1887
rect 162688 1884 162716 1924
rect 161891 1856 162716 1884
rect 162765 1887 162823 1893
rect 161891 1853 161903 1856
rect 161845 1847 161903 1853
rect 162765 1853 162777 1887
rect 162811 1853 162823 1887
rect 162765 1847 162823 1853
rect 162857 1887 162915 1893
rect 162857 1853 162869 1887
rect 162903 1884 162915 1887
rect 163038 1884 163044 1896
rect 162903 1856 163044 1884
rect 162903 1853 162915 1856
rect 162857 1847 162915 1853
rect 149606 1816 149612 1828
rect 147140 1788 149612 1816
rect 149606 1776 149612 1788
rect 149664 1776 149670 1828
rect 149716 1788 158392 1816
rect 135993 1751 136051 1757
rect 135993 1748 136005 1751
rect 134996 1720 136005 1748
rect 134889 1711 134947 1717
rect 135993 1717 136005 1720
rect 136039 1717 136051 1751
rect 135993 1711 136051 1717
rect 136174 1708 136180 1760
rect 136232 1748 136238 1760
rect 136634 1748 136640 1760
rect 136232 1720 136640 1748
rect 136232 1708 136238 1720
rect 136634 1708 136640 1720
rect 136692 1708 136698 1760
rect 137094 1708 137100 1760
rect 137152 1748 137158 1760
rect 138106 1748 138112 1760
rect 137152 1720 138112 1748
rect 137152 1708 137158 1720
rect 138106 1708 138112 1720
rect 138164 1708 138170 1760
rect 138290 1708 138296 1760
rect 138348 1748 138354 1760
rect 140130 1748 140136 1760
rect 138348 1720 140136 1748
rect 138348 1708 138354 1720
rect 140130 1708 140136 1720
rect 140188 1708 140194 1760
rect 140222 1708 140228 1760
rect 140280 1748 140286 1760
rect 145098 1748 145104 1760
rect 140280 1720 145104 1748
rect 140280 1708 140286 1720
rect 145098 1708 145104 1720
rect 145156 1708 145162 1760
rect 145190 1708 145196 1760
rect 145248 1748 145254 1760
rect 149716 1748 149744 1788
rect 145248 1720 149744 1748
rect 152461 1751 152519 1757
rect 145248 1708 145254 1720
rect 152461 1717 152473 1751
rect 152507 1748 152519 1751
rect 155954 1748 155960 1760
rect 152507 1720 155960 1748
rect 152507 1717 152519 1720
rect 152461 1711 152519 1717
rect 155954 1708 155960 1720
rect 156012 1708 156018 1760
rect 156046 1708 156052 1760
rect 156104 1748 156110 1760
rect 157337 1751 157395 1757
rect 157337 1748 157349 1751
rect 156104 1720 157349 1748
rect 156104 1708 156110 1720
rect 157337 1717 157349 1720
rect 157383 1717 157395 1751
rect 158364 1748 158392 1788
rect 159358 1776 159364 1828
rect 159416 1816 159422 1828
rect 161474 1816 161480 1828
rect 159416 1788 161480 1816
rect 159416 1776 159422 1788
rect 161474 1776 161480 1788
rect 161532 1776 161538 1828
rect 162780 1816 162808 1847
rect 163038 1844 163044 1856
rect 163096 1844 163102 1896
rect 163700 1884 163728 1924
rect 163777 1921 163789 1955
rect 163823 1952 163835 1955
rect 163823 1924 164556 1952
rect 163823 1921 163835 1924
rect 163777 1915 163835 1921
rect 164234 1884 164240 1896
rect 163700 1856 164240 1884
rect 164234 1844 164240 1856
rect 164292 1844 164298 1896
rect 163590 1816 163596 1828
rect 162780 1788 163596 1816
rect 163590 1776 163596 1788
rect 163648 1776 163654 1828
rect 163682 1776 163688 1828
rect 163740 1816 163746 1828
rect 164528 1816 164556 1924
rect 164694 1912 164700 1964
rect 164752 1952 164758 1964
rect 164896 1952 164924 1992
rect 165246 1980 165252 2032
rect 165304 2020 165310 2032
rect 165614 2020 165620 2032
rect 165304 1992 165620 2020
rect 165304 1980 165310 1992
rect 165614 1980 165620 1992
rect 165672 1980 165678 2032
rect 165706 1980 165712 2032
rect 165764 2020 165770 2032
rect 165908 2020 165936 2060
rect 167086 2048 167092 2100
rect 167144 2088 167150 2100
rect 168558 2088 168564 2100
rect 167144 2060 167684 2088
rect 168519 2060 168564 2088
rect 167144 2048 167150 2060
rect 167178 2020 167184 2032
rect 165764 1992 165809 2020
rect 165908 1992 167184 2020
rect 165764 1980 165770 1992
rect 167178 1980 167184 1992
rect 167236 1980 167242 2032
rect 167546 2020 167552 2032
rect 167380 1992 167552 2020
rect 166994 1952 167000 1964
rect 164752 1924 164797 1952
rect 164896 1924 167000 1952
rect 164752 1912 164758 1924
rect 166994 1912 167000 1924
rect 167052 1912 167058 1964
rect 167380 1952 167408 1992
rect 167546 1980 167552 1992
rect 167604 1980 167610 2032
rect 167457 1955 167515 1961
rect 167457 1952 167469 1955
rect 167380 1924 167469 1952
rect 167457 1921 167469 1924
rect 167503 1921 167515 1955
rect 167656 1952 167684 2060
rect 168558 2048 168564 2060
rect 168616 2048 168622 2100
rect 168650 2048 168656 2100
rect 168708 2088 168714 2100
rect 173897 2091 173955 2097
rect 173897 2088 173909 2091
rect 168708 2060 173909 2088
rect 168708 2048 168714 2060
rect 173897 2057 173909 2060
rect 173943 2057 173955 2091
rect 173897 2051 173955 2057
rect 173986 2048 173992 2100
rect 174044 2088 174050 2100
rect 175277 2091 175335 2097
rect 175277 2088 175289 2091
rect 174044 2060 175289 2088
rect 174044 2048 174050 2060
rect 175277 2057 175289 2060
rect 175323 2057 175335 2091
rect 175277 2051 175335 2057
rect 175734 2048 175740 2100
rect 175792 2088 175798 2100
rect 177758 2088 177764 2100
rect 175792 2060 177764 2088
rect 175792 2048 175798 2060
rect 177758 2048 177764 2060
rect 177816 2048 177822 2100
rect 177850 2048 177856 2100
rect 177908 2088 177914 2100
rect 179509 2091 179567 2097
rect 179509 2088 179521 2091
rect 177908 2060 179521 2088
rect 177908 2048 177914 2060
rect 179509 2057 179521 2060
rect 179555 2057 179567 2091
rect 179509 2051 179567 2057
rect 179598 2048 179604 2100
rect 179656 2088 179662 2100
rect 181990 2088 181996 2100
rect 179656 2060 180472 2088
rect 181951 2060 181996 2088
rect 179656 2048 179662 2060
rect 171226 1980 171232 2032
rect 171284 2020 171290 2032
rect 176470 2020 176476 2032
rect 171284 1992 176476 2020
rect 171284 1980 171290 1992
rect 176470 1980 176476 1992
rect 176528 1980 176534 2032
rect 178218 1980 178224 2032
rect 178276 2020 178282 2032
rect 180334 2020 180340 2032
rect 178276 1992 180340 2020
rect 178276 1980 178282 1992
rect 180334 1980 180340 1992
rect 180392 1980 180398 2032
rect 180444 2020 180472 2060
rect 181990 2048 181996 2060
rect 182048 2048 182054 2100
rect 183741 2091 183799 2097
rect 183741 2057 183753 2091
rect 183787 2088 183799 2091
rect 184842 2088 184848 2100
rect 183787 2060 184848 2088
rect 183787 2057 183799 2060
rect 183741 2051 183799 2057
rect 184842 2048 184848 2060
rect 184900 2048 184906 2100
rect 185394 2088 185400 2100
rect 185355 2060 185400 2088
rect 185394 2048 185400 2060
rect 185452 2048 185458 2100
rect 186314 2088 186320 2100
rect 185504 2060 186320 2088
rect 185504 2020 185532 2060
rect 186314 2048 186320 2060
rect 186372 2048 186378 2100
rect 186406 2048 186412 2100
rect 186464 2088 186470 2100
rect 189258 2088 189264 2100
rect 186464 2060 189264 2088
rect 186464 2048 186470 2060
rect 189258 2048 189264 2060
rect 189316 2048 189322 2100
rect 192938 2088 192944 2100
rect 192899 2060 192944 2088
rect 192938 2048 192944 2060
rect 192996 2048 193002 2100
rect 195054 2048 195060 2100
rect 195112 2088 195118 2100
rect 195882 2088 195888 2100
rect 195112 2060 195888 2088
rect 195112 2048 195118 2060
rect 195882 2048 195888 2060
rect 195940 2048 195946 2100
rect 180444 1992 185532 2020
rect 186222 1980 186228 2032
rect 186280 2020 186286 2032
rect 186501 2023 186559 2029
rect 186501 2020 186513 2023
rect 186280 1992 186513 2020
rect 186280 1980 186286 1992
rect 186501 1989 186513 1992
rect 186547 1989 186559 2023
rect 186501 1983 186559 1989
rect 186590 1980 186596 2032
rect 186648 2020 186654 2032
rect 187973 2023 188031 2029
rect 187973 2020 187985 2023
rect 186648 1992 187985 2020
rect 186648 1980 186654 1992
rect 187973 1989 187985 1992
rect 188019 1989 188031 2023
rect 187973 1983 188031 1989
rect 189442 1980 189448 2032
rect 189500 2020 189506 2032
rect 195793 2023 195851 2029
rect 195793 2020 195805 2023
rect 189500 1992 195805 2020
rect 189500 1980 189506 1992
rect 195793 1989 195805 1992
rect 195839 1989 195851 2023
rect 195793 1983 195851 1989
rect 171413 1955 171471 1961
rect 171413 1952 171425 1955
rect 167656 1924 171425 1952
rect 167457 1915 167515 1921
rect 171413 1921 171425 1924
rect 171459 1921 171471 1955
rect 171413 1915 171471 1921
rect 172885 1955 172943 1961
rect 172885 1921 172897 1955
rect 172931 1952 172943 1955
rect 176838 1952 176844 1964
rect 172931 1924 176844 1952
rect 172931 1921 172943 1924
rect 172885 1915 172943 1921
rect 176838 1912 176844 1924
rect 176896 1912 176902 1964
rect 177209 1955 177267 1961
rect 177209 1952 177221 1955
rect 176948 1924 177221 1952
rect 164605 1887 164663 1893
rect 164605 1853 164617 1887
rect 164651 1884 164663 1887
rect 165430 1884 165436 1896
rect 164651 1856 165436 1884
rect 164651 1853 164663 1856
rect 164605 1847 164663 1853
rect 165430 1844 165436 1856
rect 165488 1844 165494 1896
rect 165617 1887 165675 1893
rect 165617 1853 165629 1887
rect 165663 1884 165675 1887
rect 168374 1884 168380 1896
rect 165663 1856 168380 1884
rect 165663 1853 165675 1856
rect 165617 1847 165675 1853
rect 168374 1844 168380 1856
rect 168432 1844 168438 1896
rect 168469 1887 168527 1893
rect 168469 1853 168481 1887
rect 168515 1884 168527 1887
rect 169478 1884 169484 1896
rect 168515 1856 169484 1884
rect 168515 1853 168527 1856
rect 168469 1847 168527 1853
rect 169478 1844 169484 1856
rect 169536 1844 169542 1896
rect 169573 1887 169631 1893
rect 169573 1853 169585 1887
rect 169619 1884 169631 1887
rect 169662 1884 169668 1896
rect 169619 1856 169668 1884
rect 169619 1853 169631 1856
rect 169573 1847 169631 1853
rect 169662 1844 169668 1856
rect 169720 1844 169726 1896
rect 169938 1844 169944 1896
rect 169996 1884 170002 1896
rect 171870 1884 171876 1896
rect 169996 1856 171876 1884
rect 169996 1844 170002 1856
rect 171870 1844 171876 1856
rect 171928 1844 171934 1896
rect 172974 1884 172980 1896
rect 172935 1856 172980 1884
rect 172974 1844 172980 1856
rect 173032 1844 173038 1896
rect 173066 1844 173072 1896
rect 173124 1884 173130 1896
rect 173618 1884 173624 1896
rect 173124 1856 173624 1884
rect 173124 1844 173130 1856
rect 173618 1844 173624 1856
rect 173676 1844 173682 1896
rect 173802 1884 173808 1896
rect 173763 1856 173808 1884
rect 173802 1844 173808 1856
rect 173860 1844 173866 1896
rect 175185 1887 175243 1893
rect 175185 1853 175197 1887
rect 175231 1884 175243 1887
rect 176194 1884 176200 1896
rect 175231 1856 176200 1884
rect 175231 1853 175243 1856
rect 175185 1847 175243 1853
rect 176194 1844 176200 1856
rect 176252 1844 176258 1896
rect 176286 1844 176292 1896
rect 176344 1884 176350 1896
rect 176948 1884 176976 1924
rect 177209 1921 177221 1924
rect 177255 1921 177267 1955
rect 180981 1955 181039 1961
rect 180981 1952 180993 1955
rect 177209 1915 177267 1921
rect 178328 1924 180993 1952
rect 176344 1856 176976 1884
rect 177117 1887 177175 1893
rect 176344 1844 176350 1856
rect 177117 1853 177129 1887
rect 177163 1884 177175 1887
rect 178218 1884 178224 1896
rect 177163 1856 178224 1884
rect 177163 1853 177175 1856
rect 177117 1847 177175 1853
rect 178218 1844 178224 1856
rect 178276 1844 178282 1896
rect 178328 1816 178356 1924
rect 180981 1921 180993 1924
rect 181027 1921 181039 1955
rect 180981 1915 181039 1921
rect 181070 1912 181076 1964
rect 181128 1952 181134 1964
rect 186038 1952 186044 1964
rect 181128 1924 186044 1952
rect 181128 1912 181134 1924
rect 186038 1912 186044 1924
rect 186096 1912 186102 1964
rect 187694 1952 187700 1964
rect 186424 1924 187700 1952
rect 178405 1887 178463 1893
rect 178405 1853 178417 1887
rect 178451 1884 178463 1887
rect 179322 1884 179328 1896
rect 178451 1856 179328 1884
rect 178451 1853 178463 1856
rect 178405 1847 178463 1853
rect 179322 1844 179328 1856
rect 179380 1844 179386 1896
rect 179417 1887 179475 1893
rect 179417 1853 179429 1887
rect 179463 1853 179475 1887
rect 179417 1847 179475 1853
rect 178497 1819 178555 1825
rect 178497 1816 178509 1819
rect 163740 1788 164372 1816
rect 164528 1788 178356 1816
rect 178420 1788 178509 1816
rect 163740 1776 163746 1788
rect 161934 1748 161940 1760
rect 158364 1720 161940 1748
rect 157337 1711 157395 1717
rect 161934 1708 161940 1720
rect 161992 1708 161998 1760
rect 162026 1708 162032 1760
rect 162084 1748 162090 1760
rect 163777 1751 163835 1757
rect 163777 1748 163789 1751
rect 162084 1720 163789 1748
rect 162084 1708 162090 1720
rect 163777 1717 163789 1720
rect 163823 1717 163835 1751
rect 164344 1748 164372 1788
rect 169665 1751 169723 1757
rect 169665 1748 169677 1751
rect 164344 1720 169677 1748
rect 163777 1711 163835 1717
rect 169665 1717 169677 1720
rect 169711 1717 169723 1751
rect 169665 1711 169723 1717
rect 169754 1708 169760 1760
rect 169812 1748 169818 1760
rect 172422 1748 172428 1760
rect 169812 1720 172428 1748
rect 169812 1708 169818 1720
rect 172422 1708 172428 1720
rect 172480 1708 172486 1760
rect 172974 1708 172980 1760
rect 173032 1748 173038 1760
rect 176010 1748 176016 1760
rect 173032 1720 176016 1748
rect 173032 1708 173038 1720
rect 176010 1708 176016 1720
rect 176068 1708 176074 1760
rect 176102 1708 176108 1760
rect 176160 1748 176166 1760
rect 178420 1748 178448 1788
rect 178497 1785 178509 1788
rect 178543 1785 178555 1819
rect 179432 1816 179460 1847
rect 179506 1844 179512 1896
rect 179564 1884 179570 1896
rect 180702 1884 180708 1896
rect 179564 1856 180708 1884
rect 179564 1844 179570 1856
rect 180702 1844 180708 1856
rect 180760 1844 180766 1896
rect 180889 1887 180947 1893
rect 180889 1853 180901 1887
rect 180935 1884 180947 1887
rect 181901 1887 181959 1893
rect 180935 1856 181760 1884
rect 180935 1853 180947 1856
rect 180889 1847 180947 1853
rect 181622 1816 181628 1828
rect 179432 1788 181628 1816
rect 178497 1779 178555 1785
rect 181622 1776 181628 1788
rect 181680 1776 181686 1828
rect 176160 1720 178448 1748
rect 181732 1748 181760 1856
rect 181901 1853 181913 1887
rect 181947 1884 181959 1887
rect 183649 1887 183707 1893
rect 181947 1856 183600 1884
rect 181947 1853 181959 1856
rect 181901 1847 181959 1853
rect 183462 1748 183468 1760
rect 181732 1720 183468 1748
rect 176160 1708 176166 1720
rect 183462 1708 183468 1720
rect 183520 1708 183526 1760
rect 183572 1748 183600 1856
rect 183649 1853 183661 1887
rect 183695 1853 183707 1887
rect 183649 1847 183707 1853
rect 183664 1816 183692 1847
rect 183738 1844 183744 1896
rect 183796 1884 183802 1896
rect 184934 1884 184940 1896
rect 183796 1856 184940 1884
rect 183796 1844 183802 1856
rect 184934 1844 184940 1856
rect 184992 1844 184998 1896
rect 186424 1893 186452 1924
rect 187694 1912 187700 1924
rect 187752 1912 187758 1964
rect 191466 1952 191472 1964
rect 189460 1924 191472 1952
rect 185305 1887 185363 1893
rect 185305 1853 185317 1887
rect 185351 1884 185363 1887
rect 186409 1887 186467 1893
rect 185351 1856 186360 1884
rect 185351 1853 185363 1856
rect 185305 1847 185363 1853
rect 186332 1828 186360 1856
rect 186409 1853 186421 1887
rect 186455 1853 186467 1887
rect 186409 1847 186467 1853
rect 187881 1887 187939 1893
rect 187881 1853 187893 1887
rect 187927 1884 187939 1887
rect 189460 1884 189488 1924
rect 191466 1912 191472 1924
rect 191524 1912 191530 1964
rect 191926 1912 191932 1964
rect 191984 1952 191990 1964
rect 194686 1952 194692 1964
rect 191984 1924 193996 1952
rect 194647 1924 194692 1952
rect 191984 1912 191990 1924
rect 187927 1856 189488 1884
rect 189537 1887 189595 1893
rect 187927 1853 187939 1856
rect 187881 1847 187939 1853
rect 189537 1853 189549 1887
rect 189583 1884 189595 1887
rect 190454 1884 190460 1896
rect 189583 1856 190460 1884
rect 189583 1853 189595 1856
rect 189537 1847 189595 1853
rect 190454 1844 190460 1856
rect 190512 1844 190518 1896
rect 190549 1887 190607 1893
rect 190549 1853 190561 1887
rect 190595 1853 190607 1887
rect 190549 1847 190607 1853
rect 185762 1816 185768 1828
rect 183664 1788 185768 1816
rect 185762 1776 185768 1788
rect 185820 1776 185826 1828
rect 186314 1776 186320 1828
rect 186372 1776 186378 1828
rect 189258 1776 189264 1828
rect 189316 1816 189322 1828
rect 190564 1816 190592 1847
rect 190638 1844 190644 1896
rect 190696 1884 190702 1896
rect 192849 1887 192907 1893
rect 190696 1856 190741 1884
rect 190696 1844 190702 1856
rect 192849 1853 192861 1887
rect 192895 1853 192907 1887
rect 192849 1847 192907 1853
rect 189316 1788 190592 1816
rect 192864 1816 192892 1847
rect 193306 1844 193312 1896
rect 193364 1884 193370 1896
rect 193861 1887 193919 1893
rect 193861 1884 193873 1887
rect 193364 1856 193873 1884
rect 193364 1844 193370 1856
rect 193861 1853 193873 1856
rect 193907 1853 193919 1887
rect 193968 1884 193996 1924
rect 194686 1912 194692 1924
rect 194744 1912 194750 1964
rect 195701 1887 195759 1893
rect 195701 1884 195713 1887
rect 193968 1856 195713 1884
rect 193861 1847 193919 1853
rect 195701 1853 195713 1856
rect 195747 1853 195759 1887
rect 195701 1847 195759 1853
rect 197262 1816 197268 1828
rect 192864 1788 197268 1816
rect 189316 1776 189322 1788
rect 197262 1776 197268 1788
rect 197320 1776 197326 1828
rect 185302 1748 185308 1760
rect 183572 1720 185308 1748
rect 185302 1708 185308 1720
rect 185360 1708 185366 1760
rect 185946 1708 185952 1760
rect 186004 1748 186010 1760
rect 189629 1751 189687 1757
rect 189629 1748 189641 1751
rect 186004 1720 189641 1748
rect 186004 1708 186010 1720
rect 189629 1717 189641 1720
rect 189675 1717 189687 1751
rect 189629 1711 189687 1717
rect 189810 1708 189816 1760
rect 189868 1748 189874 1760
rect 195146 1748 195152 1760
rect 189868 1720 195152 1748
rect 189868 1708 189874 1720
rect 195146 1708 195152 1720
rect 195204 1708 195210 1760
rect 1104 1658 198812 1680
rect 1104 1606 24078 1658
rect 24130 1606 64078 1658
rect 64130 1606 104078 1658
rect 104130 1606 144078 1658
rect 144130 1606 184078 1658
rect 184130 1606 198812 1658
rect 1104 1584 198812 1606
rect 5353 1547 5411 1553
rect 5353 1513 5365 1547
rect 5399 1544 5411 1547
rect 5902 1544 5908 1556
rect 5399 1516 5908 1544
rect 5399 1513 5411 1516
rect 5353 1507 5411 1513
rect 5902 1504 5908 1516
rect 5960 1504 5966 1556
rect 7009 1547 7067 1553
rect 7009 1513 7021 1547
rect 7055 1544 7067 1547
rect 7190 1544 7196 1556
rect 7055 1516 7196 1544
rect 7055 1513 7067 1516
rect 7009 1507 7067 1513
rect 7190 1504 7196 1516
rect 7248 1504 7254 1556
rect 7926 1504 7932 1556
rect 7984 1544 7990 1556
rect 8021 1547 8079 1553
rect 8021 1544 8033 1547
rect 7984 1516 8033 1544
rect 7984 1504 7990 1516
rect 8021 1513 8033 1516
rect 8067 1513 8079 1547
rect 8021 1507 8079 1513
rect 15841 1547 15899 1553
rect 15841 1513 15853 1547
rect 15887 1544 15899 1547
rect 16574 1544 16580 1556
rect 15887 1516 16580 1544
rect 15887 1513 15899 1516
rect 15841 1507 15899 1513
rect 16574 1504 16580 1516
rect 16632 1504 16638 1556
rect 16850 1544 16856 1556
rect 16811 1516 16856 1544
rect 16850 1504 16856 1516
rect 16908 1504 16914 1556
rect 20165 1547 20223 1553
rect 20165 1513 20177 1547
rect 20211 1544 20223 1547
rect 21910 1544 21916 1556
rect 20211 1516 21916 1544
rect 20211 1513 20223 1516
rect 20165 1507 20223 1513
rect 21910 1504 21916 1516
rect 21968 1504 21974 1556
rect 22002 1504 22008 1556
rect 22060 1544 22066 1556
rect 22465 1547 22523 1553
rect 22465 1544 22477 1547
rect 22060 1516 22477 1544
rect 22060 1504 22066 1516
rect 22465 1513 22477 1516
rect 22511 1513 22523 1547
rect 22465 1507 22523 1513
rect 24213 1547 24271 1553
rect 24213 1513 24225 1547
rect 24259 1544 24271 1547
rect 24946 1544 24952 1556
rect 24259 1516 24952 1544
rect 24259 1513 24271 1516
rect 24213 1507 24271 1513
rect 24946 1504 24952 1516
rect 25004 1504 25010 1556
rect 25225 1547 25283 1553
rect 25225 1513 25237 1547
rect 25271 1544 25283 1547
rect 25314 1544 25320 1556
rect 25271 1516 25320 1544
rect 25271 1513 25283 1516
rect 25225 1507 25283 1513
rect 25314 1504 25320 1516
rect 25372 1504 25378 1556
rect 28534 1544 28540 1556
rect 28495 1516 28540 1544
rect 28534 1504 28540 1516
rect 28592 1504 28598 1556
rect 32950 1544 32956 1556
rect 32911 1516 32956 1544
rect 32950 1504 32956 1516
rect 33008 1504 33014 1556
rect 33870 1504 33876 1556
rect 33928 1544 33934 1556
rect 33965 1547 34023 1553
rect 33965 1544 33977 1547
rect 33928 1516 33977 1544
rect 33928 1504 33934 1516
rect 33965 1513 33977 1516
rect 34011 1513 34023 1547
rect 33965 1507 34023 1513
rect 35529 1547 35587 1553
rect 35529 1513 35541 1547
rect 35575 1544 35587 1547
rect 35986 1544 35992 1556
rect 35575 1516 35992 1544
rect 35575 1513 35587 1516
rect 35529 1507 35587 1513
rect 35986 1504 35992 1516
rect 36044 1504 36050 1556
rect 39114 1544 39120 1556
rect 39075 1516 39120 1544
rect 39114 1504 39120 1516
rect 39172 1504 39178 1556
rect 42981 1547 43039 1553
rect 42981 1513 42993 1547
rect 43027 1544 43039 1547
rect 43530 1544 43536 1556
rect 43027 1516 43536 1544
rect 43027 1513 43039 1516
rect 42981 1507 43039 1513
rect 43530 1504 43536 1516
rect 43588 1504 43594 1556
rect 43622 1504 43628 1556
rect 43680 1544 43686 1556
rect 44453 1547 44511 1553
rect 44453 1544 44465 1547
rect 43680 1516 44465 1544
rect 43680 1504 43686 1516
rect 44453 1513 44465 1516
rect 44499 1513 44511 1547
rect 44453 1507 44511 1513
rect 45370 1504 45376 1556
rect 45428 1544 45434 1556
rect 45465 1547 45523 1553
rect 45465 1544 45477 1547
rect 45428 1516 45477 1544
rect 45428 1504 45434 1516
rect 45465 1513 45477 1516
rect 45511 1513 45523 1547
rect 45465 1507 45523 1513
rect 49789 1547 49847 1553
rect 49789 1513 49801 1547
rect 49835 1544 49847 1547
rect 50338 1544 50344 1556
rect 49835 1516 50344 1544
rect 49835 1513 49847 1516
rect 49789 1507 49847 1513
rect 50338 1504 50344 1516
rect 50396 1504 50402 1556
rect 50801 1547 50859 1553
rect 50801 1513 50813 1547
rect 50847 1544 50859 1547
rect 52546 1544 52552 1556
rect 50847 1516 52552 1544
rect 50847 1513 50859 1516
rect 50801 1507 50859 1513
rect 52546 1504 52552 1516
rect 52604 1504 52610 1556
rect 52641 1547 52699 1553
rect 52641 1513 52653 1547
rect 52687 1544 52699 1547
rect 53834 1544 53840 1556
rect 52687 1516 53840 1544
rect 52687 1513 52699 1516
rect 52641 1507 52699 1513
rect 53834 1504 53840 1516
rect 53892 1504 53898 1556
rect 54110 1544 54116 1556
rect 54071 1516 54116 1544
rect 54110 1504 54116 1516
rect 54168 1504 54174 1556
rect 59541 1547 59599 1553
rect 59541 1513 59553 1547
rect 59587 1544 59599 1547
rect 62482 1544 62488 1556
rect 59587 1516 62488 1544
rect 59587 1513 59599 1516
rect 59541 1507 59599 1513
rect 62482 1504 62488 1516
rect 62540 1504 62546 1556
rect 74077 1547 74135 1553
rect 74077 1513 74089 1547
rect 74123 1544 74135 1547
rect 75362 1544 75368 1556
rect 74123 1516 75368 1544
rect 74123 1513 74135 1516
rect 74077 1507 74135 1513
rect 75362 1504 75368 1516
rect 75420 1504 75426 1556
rect 79962 1544 79968 1556
rect 79923 1516 79968 1544
rect 79962 1504 79968 1516
rect 80020 1504 80026 1556
rect 81434 1544 81440 1556
rect 80072 1516 81440 1544
rect 14090 1436 14096 1488
rect 14148 1476 14154 1488
rect 14148 1448 16804 1476
rect 14148 1436 14154 1448
rect 3970 1368 3976 1420
rect 4028 1408 4034 1420
rect 5261 1411 5319 1417
rect 5261 1408 5273 1411
rect 4028 1380 5273 1408
rect 4028 1368 4034 1380
rect 5261 1377 5273 1380
rect 5307 1377 5319 1411
rect 6917 1411 6975 1417
rect 6917 1408 6929 1411
rect 5261 1371 5319 1377
rect 5368 1380 6929 1408
rect 4982 1300 4988 1352
rect 5040 1340 5046 1352
rect 5368 1340 5396 1380
rect 6917 1377 6929 1380
rect 6963 1377 6975 1411
rect 6917 1371 6975 1377
rect 7558 1368 7564 1420
rect 7616 1408 7622 1420
rect 7929 1411 7987 1417
rect 7929 1408 7941 1411
rect 7616 1380 7941 1408
rect 7616 1368 7622 1380
rect 7929 1377 7941 1380
rect 7975 1377 7987 1411
rect 7929 1371 7987 1377
rect 15749 1411 15807 1417
rect 15749 1377 15761 1411
rect 15795 1408 15807 1411
rect 16298 1408 16304 1420
rect 15795 1380 16304 1408
rect 15795 1377 15807 1380
rect 15749 1371 15807 1377
rect 16298 1368 16304 1380
rect 16356 1368 16362 1420
rect 16776 1417 16804 1448
rect 20622 1436 20628 1488
rect 20680 1476 20686 1488
rect 20680 1448 22416 1476
rect 20680 1436 20686 1448
rect 16753 1411 16811 1417
rect 16753 1377 16765 1411
rect 16799 1377 16811 1411
rect 16753 1371 16811 1377
rect 18874 1368 18880 1420
rect 18932 1408 18938 1420
rect 20073 1411 20131 1417
rect 20073 1408 20085 1411
rect 18932 1380 20085 1408
rect 18932 1368 18938 1380
rect 20073 1377 20085 1380
rect 20119 1377 20131 1411
rect 21361 1411 21419 1417
rect 21361 1408 21373 1411
rect 20073 1371 20131 1377
rect 20180 1380 21373 1408
rect 5040 1312 5396 1340
rect 5040 1300 5046 1312
rect 19794 1300 19800 1352
rect 19852 1340 19858 1352
rect 20180 1340 20208 1380
rect 21361 1377 21373 1380
rect 21407 1377 21419 1411
rect 21361 1371 21419 1377
rect 21450 1368 21456 1420
rect 21508 1408 21514 1420
rect 22388 1417 22416 1448
rect 32398 1436 32404 1488
rect 32456 1476 32462 1488
rect 32456 1448 35480 1476
rect 32456 1436 32462 1448
rect 22373 1411 22431 1417
rect 21508 1380 21553 1408
rect 21508 1368 21514 1380
rect 22373 1377 22385 1411
rect 22419 1377 22431 1411
rect 24121 1411 24179 1417
rect 24121 1408 24133 1411
rect 22373 1371 22431 1377
rect 22480 1380 24133 1408
rect 19852 1312 20208 1340
rect 19852 1300 19858 1312
rect 21910 1300 21916 1352
rect 21968 1340 21974 1352
rect 22480 1340 22508 1380
rect 24121 1377 24133 1380
rect 24167 1377 24179 1411
rect 25133 1411 25191 1417
rect 25133 1408 25145 1411
rect 24121 1371 24179 1377
rect 24228 1380 25145 1408
rect 21968 1312 22508 1340
rect 21968 1300 21974 1312
rect 22554 1300 22560 1352
rect 22612 1340 22618 1352
rect 24228 1340 24256 1380
rect 25133 1377 25145 1380
rect 25179 1377 25191 1411
rect 28445 1411 28503 1417
rect 28445 1408 28457 1411
rect 25133 1371 25191 1377
rect 25240 1380 28457 1408
rect 22612 1312 24256 1340
rect 22612 1300 22618 1312
rect 23658 1232 23664 1284
rect 23716 1272 23722 1284
rect 25240 1272 25268 1380
rect 28445 1377 28457 1380
rect 28491 1377 28503 1411
rect 28445 1371 28503 1377
rect 30650 1368 30656 1420
rect 30708 1408 30714 1420
rect 32861 1411 32919 1417
rect 32861 1408 32873 1411
rect 30708 1380 32873 1408
rect 30708 1368 30714 1380
rect 32861 1377 32873 1380
rect 32907 1377 32919 1411
rect 32861 1371 32919 1377
rect 33042 1368 33048 1420
rect 33100 1408 33106 1420
rect 35452 1417 35480 1448
rect 38102 1436 38108 1488
rect 38160 1476 38166 1488
rect 38160 1448 42932 1476
rect 38160 1436 38166 1448
rect 33873 1411 33931 1417
rect 33873 1408 33885 1411
rect 33100 1380 33885 1408
rect 33100 1368 33106 1380
rect 33873 1377 33885 1380
rect 33919 1377 33931 1411
rect 33873 1371 33931 1377
rect 35437 1411 35495 1417
rect 35437 1377 35449 1411
rect 35483 1377 35495 1411
rect 39025 1411 39083 1417
rect 39025 1408 39037 1411
rect 35437 1371 35495 1377
rect 35820 1380 39037 1408
rect 34974 1300 34980 1352
rect 35032 1340 35038 1352
rect 35820 1340 35848 1380
rect 39025 1377 39037 1380
rect 39071 1377 39083 1411
rect 39025 1371 39083 1377
rect 41598 1368 41604 1420
rect 41656 1408 41662 1420
rect 42904 1417 42932 1448
rect 43070 1436 43076 1488
rect 43128 1476 43134 1488
rect 43128 1448 45416 1476
rect 43128 1436 43134 1448
rect 45388 1417 45416 1448
rect 51166 1436 51172 1488
rect 51224 1476 51230 1488
rect 63494 1476 63500 1488
rect 51224 1448 54064 1476
rect 51224 1436 51230 1448
rect 42889 1411 42947 1417
rect 41656 1380 42840 1408
rect 41656 1368 41662 1380
rect 35032 1312 35848 1340
rect 42812 1340 42840 1380
rect 42889 1377 42901 1411
rect 42935 1377 42947 1411
rect 44361 1411 44419 1417
rect 44361 1408 44373 1411
rect 42889 1371 42947 1377
rect 42996 1380 44373 1408
rect 42996 1340 43024 1380
rect 44361 1377 44373 1380
rect 44407 1377 44419 1411
rect 44361 1371 44419 1377
rect 45373 1411 45431 1417
rect 45373 1377 45385 1411
rect 45419 1377 45431 1411
rect 45373 1371 45431 1377
rect 47486 1368 47492 1420
rect 47544 1408 47550 1420
rect 49697 1411 49755 1417
rect 49697 1408 49709 1411
rect 47544 1380 49709 1408
rect 47544 1368 47550 1380
rect 49697 1377 49709 1380
rect 49743 1377 49755 1411
rect 49697 1371 49755 1377
rect 49878 1368 49884 1420
rect 49936 1408 49942 1420
rect 50709 1411 50767 1417
rect 50709 1408 50721 1411
rect 49936 1380 50721 1408
rect 49936 1368 49942 1380
rect 50709 1377 50721 1380
rect 50755 1377 50767 1411
rect 50709 1371 50767 1377
rect 52549 1411 52607 1417
rect 52549 1377 52561 1411
rect 52595 1408 52607 1411
rect 52914 1408 52920 1420
rect 52595 1380 52920 1408
rect 52595 1377 52607 1380
rect 52549 1371 52607 1377
rect 52914 1368 52920 1380
rect 52972 1368 52978 1420
rect 54036 1417 54064 1448
rect 59740 1448 63500 1476
rect 54021 1411 54079 1417
rect 54021 1377 54033 1411
rect 54067 1377 54079 1411
rect 54021 1371 54079 1377
rect 56873 1411 56931 1417
rect 56873 1377 56885 1411
rect 56919 1408 56931 1411
rect 58618 1408 58624 1420
rect 56919 1380 58624 1408
rect 56919 1377 56931 1380
rect 56873 1371 56931 1377
rect 58618 1368 58624 1380
rect 58676 1368 58682 1420
rect 59740 1417 59768 1448
rect 63494 1436 63500 1448
rect 63552 1436 63558 1488
rect 65058 1436 65064 1488
rect 65116 1476 65122 1488
rect 69661 1479 69719 1485
rect 69661 1476 69673 1479
rect 65116 1448 69673 1476
rect 65116 1436 65122 1448
rect 69661 1445 69673 1448
rect 69707 1445 69719 1479
rect 69661 1439 69719 1445
rect 78953 1479 79011 1485
rect 78953 1445 78965 1479
rect 78999 1476 79011 1479
rect 79042 1476 79048 1488
rect 78999 1448 79048 1476
rect 78999 1445 79011 1448
rect 78953 1439 79011 1445
rect 79042 1436 79048 1448
rect 79100 1436 79106 1488
rect 59725 1411 59783 1417
rect 59725 1377 59737 1411
rect 59771 1377 59783 1411
rect 59725 1371 59783 1377
rect 59814 1368 59820 1420
rect 59872 1408 59878 1420
rect 61105 1411 61163 1417
rect 61105 1408 61117 1411
rect 59872 1380 61117 1408
rect 59872 1368 59878 1380
rect 61105 1377 61117 1380
rect 61151 1377 61163 1411
rect 61470 1408 61476 1420
rect 61431 1380 61476 1408
rect 61105 1371 61163 1377
rect 61470 1368 61476 1380
rect 61528 1368 61534 1420
rect 64230 1368 64236 1420
rect 64288 1408 64294 1420
rect 66162 1408 66168 1420
rect 64288 1380 66168 1408
rect 64288 1368 64294 1380
rect 66162 1368 66168 1380
rect 66220 1368 66226 1420
rect 69474 1368 69480 1420
rect 69532 1408 69538 1420
rect 69753 1411 69811 1417
rect 69753 1408 69765 1411
rect 69532 1380 69765 1408
rect 69532 1368 69538 1380
rect 69753 1377 69765 1380
rect 69799 1377 69811 1411
rect 69753 1371 69811 1377
rect 70302 1368 70308 1420
rect 70360 1408 70366 1420
rect 72602 1408 72608 1420
rect 70360 1380 72464 1408
rect 72563 1380 72608 1408
rect 70360 1368 70366 1380
rect 42812 1312 43024 1340
rect 35032 1300 35038 1312
rect 55950 1300 55956 1352
rect 56008 1340 56014 1352
rect 56229 1343 56287 1349
rect 56229 1340 56241 1343
rect 56008 1312 56241 1340
rect 56008 1300 56014 1312
rect 56229 1309 56241 1312
rect 56275 1309 56287 1343
rect 72436 1340 72464 1380
rect 72602 1368 72608 1380
rect 72660 1368 72666 1420
rect 75454 1408 75460 1420
rect 75415 1380 75460 1408
rect 75454 1368 75460 1380
rect 75512 1368 75518 1420
rect 76101 1411 76159 1417
rect 76101 1377 76113 1411
rect 76147 1408 76159 1411
rect 76374 1408 76380 1420
rect 76147 1380 76380 1408
rect 76147 1377 76159 1380
rect 76101 1371 76159 1377
rect 76374 1368 76380 1380
rect 76432 1368 76438 1420
rect 77113 1411 77171 1417
rect 77113 1377 77125 1411
rect 77159 1408 77171 1411
rect 78861 1411 78919 1417
rect 77159 1380 78812 1408
rect 77159 1377 77171 1380
rect 77113 1371 77171 1377
rect 72513 1343 72571 1349
rect 72513 1340 72525 1343
rect 72436 1312 72525 1340
rect 56229 1303 56287 1309
rect 72513 1309 72525 1312
rect 72559 1309 72571 1343
rect 78784 1340 78812 1380
rect 78861 1377 78873 1411
rect 78907 1408 78919 1411
rect 80072 1408 80100 1516
rect 81434 1504 81440 1516
rect 81492 1504 81498 1556
rect 81805 1547 81863 1553
rect 81805 1513 81817 1547
rect 81851 1544 81863 1547
rect 82170 1544 82176 1556
rect 81851 1516 82176 1544
rect 81851 1513 81863 1516
rect 81805 1507 81863 1513
rect 82170 1504 82176 1516
rect 82228 1504 82234 1556
rect 82817 1547 82875 1553
rect 82817 1513 82829 1547
rect 82863 1544 82875 1547
rect 83274 1544 83280 1556
rect 82863 1516 83280 1544
rect 82863 1513 82875 1516
rect 82817 1507 82875 1513
rect 83274 1504 83280 1516
rect 83332 1504 83338 1556
rect 85577 1547 85635 1553
rect 85577 1513 85589 1547
rect 85623 1544 85635 1547
rect 86310 1544 86316 1556
rect 85623 1516 86316 1544
rect 85623 1513 85635 1516
rect 85577 1507 85635 1513
rect 86310 1504 86316 1516
rect 86368 1504 86374 1556
rect 91186 1544 91192 1556
rect 86420 1516 91048 1544
rect 91147 1516 91192 1544
rect 84473 1411 84531 1417
rect 78907 1380 80100 1408
rect 80164 1380 84424 1408
rect 78907 1377 78919 1380
rect 78861 1371 78919 1377
rect 80164 1340 80192 1380
rect 78784 1312 80192 1340
rect 72513 1303 72571 1309
rect 23716 1244 25268 1272
rect 84396 1272 84424 1380
rect 84473 1377 84485 1411
rect 84519 1377 84531 1411
rect 84654 1408 84660 1420
rect 84615 1380 84660 1408
rect 84473 1371 84531 1377
rect 84488 1340 84516 1371
rect 84654 1368 84660 1380
rect 84712 1368 84718 1420
rect 85666 1408 85672 1420
rect 84764 1380 85672 1408
rect 84764 1340 84792 1380
rect 85666 1368 85672 1380
rect 85724 1368 85730 1420
rect 86420 1408 86448 1516
rect 91020 1476 91048 1516
rect 91186 1504 91192 1516
rect 91244 1504 91250 1556
rect 94041 1547 94099 1553
rect 94041 1513 94053 1547
rect 94087 1544 94099 1547
rect 95510 1544 95516 1556
rect 94087 1516 95516 1544
rect 94087 1513 94099 1516
rect 94041 1507 94099 1513
rect 95510 1504 95516 1516
rect 95568 1504 95574 1556
rect 96982 1544 96988 1556
rect 96943 1516 96988 1544
rect 96982 1504 96988 1516
rect 97040 1504 97046 1556
rect 104618 1544 104624 1556
rect 99208 1516 104624 1544
rect 92750 1476 92756 1488
rect 91020 1448 92756 1476
rect 92750 1436 92756 1448
rect 92808 1436 92814 1488
rect 93026 1436 93032 1488
rect 93084 1476 93090 1488
rect 93084 1448 95096 1476
rect 93084 1436 93090 1448
rect 87414 1408 87420 1420
rect 85776 1380 86448 1408
rect 87375 1380 87420 1408
rect 84488 1312 84792 1340
rect 85776 1272 85804 1380
rect 87414 1368 87420 1380
rect 87472 1368 87478 1420
rect 88521 1411 88579 1417
rect 88521 1377 88533 1411
rect 88567 1408 88579 1411
rect 89622 1408 89628 1420
rect 88567 1380 89628 1408
rect 88567 1377 88579 1380
rect 88521 1371 88579 1377
rect 89622 1368 89628 1380
rect 89680 1368 89686 1420
rect 90174 1408 90180 1420
rect 90135 1380 90180 1408
rect 90174 1368 90180 1380
rect 90232 1368 90238 1420
rect 90358 1408 90364 1420
rect 90319 1380 90364 1408
rect 90358 1368 90364 1380
rect 90416 1368 90422 1420
rect 92106 1368 92112 1420
rect 92164 1408 92170 1420
rect 92477 1411 92535 1417
rect 92477 1408 92489 1411
rect 92164 1380 92489 1408
rect 92164 1368 92170 1380
rect 92477 1377 92489 1380
rect 92523 1377 92535 1411
rect 93118 1408 93124 1420
rect 93079 1380 93124 1408
rect 92477 1371 92535 1377
rect 93118 1368 93124 1380
rect 93176 1368 93182 1420
rect 86402 1300 86408 1352
rect 86460 1340 86466 1352
rect 86773 1343 86831 1349
rect 86773 1340 86785 1343
rect 86460 1312 86785 1340
rect 86460 1300 86466 1312
rect 86773 1309 86785 1312
rect 86819 1309 86831 1343
rect 95068 1340 95096 1448
rect 95234 1436 95240 1488
rect 95292 1476 95298 1488
rect 95329 1479 95387 1485
rect 95329 1476 95341 1479
rect 95292 1448 95341 1476
rect 95292 1436 95298 1448
rect 95329 1445 95341 1448
rect 95375 1445 95387 1479
rect 98914 1476 98920 1488
rect 95329 1439 95387 1445
rect 95528 1448 98920 1476
rect 95142 1368 95148 1420
rect 95200 1408 95206 1420
rect 95421 1411 95479 1417
rect 95421 1408 95433 1411
rect 95200 1380 95433 1408
rect 95200 1368 95206 1380
rect 95421 1377 95433 1380
rect 95467 1377 95479 1411
rect 95421 1371 95479 1377
rect 95528 1340 95556 1448
rect 98914 1436 98920 1448
rect 98972 1436 98978 1488
rect 96893 1411 96951 1417
rect 96893 1377 96905 1411
rect 96939 1408 96951 1411
rect 99101 1411 99159 1417
rect 96939 1380 99052 1408
rect 96939 1377 96951 1380
rect 96893 1371 96951 1377
rect 95068 1312 95556 1340
rect 86773 1303 86831 1309
rect 84396 1244 85804 1272
rect 99024 1272 99052 1380
rect 99101 1377 99113 1411
rect 99147 1377 99159 1411
rect 99101 1371 99159 1377
rect 99116 1340 99144 1371
rect 99208 1340 99236 1516
rect 104618 1504 104624 1516
rect 104676 1504 104682 1556
rect 105722 1544 105728 1556
rect 105683 1516 105728 1544
rect 105722 1504 105728 1516
rect 105780 1504 105786 1556
rect 109034 1544 109040 1556
rect 107304 1516 109040 1544
rect 99282 1436 99288 1488
rect 99340 1476 99346 1488
rect 102137 1479 102195 1485
rect 99340 1448 101996 1476
rect 99340 1436 99346 1448
rect 99116 1312 99236 1340
rect 101968 1340 101996 1448
rect 102137 1445 102149 1479
rect 102183 1476 102195 1479
rect 104710 1476 104716 1488
rect 102183 1448 104716 1476
rect 102183 1445 102195 1448
rect 102137 1439 102195 1445
rect 104710 1436 104716 1448
rect 104768 1436 104774 1488
rect 107304 1476 107332 1516
rect 109034 1504 109040 1516
rect 109092 1504 109098 1556
rect 109494 1544 109500 1556
rect 109144 1516 109500 1544
rect 105648 1448 107332 1476
rect 107473 1479 107531 1485
rect 102045 1411 102103 1417
rect 102045 1377 102057 1411
rect 102091 1408 102103 1411
rect 102226 1408 102232 1420
rect 102091 1380 102232 1408
rect 102091 1377 102103 1380
rect 102045 1371 102103 1377
rect 102226 1368 102232 1380
rect 102284 1368 102290 1420
rect 104621 1411 104679 1417
rect 102336 1380 104480 1408
rect 102336 1340 102364 1380
rect 101968 1312 102364 1340
rect 99282 1272 99288 1284
rect 99024 1244 99288 1272
rect 23716 1232 23722 1244
rect 99282 1232 99288 1244
rect 99340 1232 99346 1284
rect 104452 1272 104480 1380
rect 104621 1377 104633 1411
rect 104667 1408 104679 1411
rect 105538 1408 105544 1420
rect 104667 1380 105544 1408
rect 104667 1377 104679 1380
rect 104621 1371 104679 1377
rect 105538 1368 105544 1380
rect 105596 1368 105602 1420
rect 105648 1417 105676 1448
rect 107473 1445 107485 1479
rect 107519 1476 107531 1479
rect 109144 1476 109172 1516
rect 109494 1504 109500 1516
rect 109552 1504 109558 1556
rect 109678 1544 109684 1556
rect 109639 1516 109684 1544
rect 109678 1504 109684 1516
rect 109736 1504 109742 1556
rect 109770 1504 109776 1556
rect 109828 1544 109834 1556
rect 114370 1544 114376 1556
rect 109828 1516 114376 1544
rect 109828 1504 109834 1516
rect 114370 1504 114376 1516
rect 114428 1504 114434 1556
rect 115750 1504 115756 1556
rect 115808 1544 115814 1556
rect 116397 1547 116455 1553
rect 116397 1544 116409 1547
rect 115808 1516 116409 1544
rect 115808 1504 115814 1516
rect 116397 1513 116409 1516
rect 116443 1513 116455 1547
rect 116397 1507 116455 1513
rect 117682 1504 117688 1556
rect 117740 1544 117746 1556
rect 118237 1547 118295 1553
rect 118237 1544 118249 1547
rect 117740 1516 118249 1544
rect 117740 1504 117746 1516
rect 118237 1513 118249 1516
rect 118283 1513 118295 1547
rect 118237 1507 118295 1513
rect 119154 1504 119160 1556
rect 119212 1544 119218 1556
rect 120442 1544 120448 1556
rect 119212 1516 120448 1544
rect 119212 1504 119218 1516
rect 120442 1504 120448 1516
rect 120500 1504 120506 1556
rect 121086 1504 121092 1556
rect 121144 1544 121150 1556
rect 121457 1547 121515 1553
rect 121457 1544 121469 1547
rect 121144 1516 121469 1544
rect 121144 1504 121150 1516
rect 121457 1513 121469 1516
rect 121503 1513 121515 1547
rect 121457 1507 121515 1513
rect 121822 1504 121828 1556
rect 121880 1544 121886 1556
rect 122837 1547 122895 1553
rect 122837 1544 122849 1547
rect 121880 1516 122849 1544
rect 121880 1504 121886 1516
rect 122837 1513 122849 1516
rect 122883 1513 122895 1547
rect 122837 1507 122895 1513
rect 123754 1504 123760 1556
rect 123812 1544 123818 1556
rect 127894 1544 127900 1556
rect 123812 1516 127900 1544
rect 123812 1504 123818 1516
rect 127894 1504 127900 1516
rect 127952 1504 127958 1556
rect 128078 1504 128084 1556
rect 128136 1544 128142 1556
rect 140314 1544 140320 1556
rect 128136 1516 140320 1544
rect 128136 1504 128142 1516
rect 140314 1504 140320 1516
rect 140372 1504 140378 1556
rect 141234 1544 141240 1556
rect 141195 1516 141240 1544
rect 141234 1504 141240 1516
rect 141292 1504 141298 1556
rect 141694 1504 141700 1556
rect 141752 1544 141758 1556
rect 143074 1544 143080 1556
rect 141752 1516 143080 1544
rect 141752 1504 141758 1516
rect 143074 1504 143080 1516
rect 143132 1504 143138 1556
rect 146202 1504 146208 1556
rect 146260 1544 146266 1556
rect 146757 1547 146815 1553
rect 146757 1544 146769 1547
rect 146260 1516 146769 1544
rect 146260 1504 146266 1516
rect 146757 1513 146769 1516
rect 146803 1513 146815 1547
rect 146757 1507 146815 1513
rect 146846 1504 146852 1556
rect 146904 1544 146910 1556
rect 147398 1544 147404 1556
rect 146904 1516 147404 1544
rect 146904 1504 146910 1516
rect 147398 1504 147404 1516
rect 147456 1504 147462 1556
rect 150342 1544 150348 1556
rect 150303 1516 150348 1544
rect 150342 1504 150348 1516
rect 150400 1504 150406 1556
rect 152458 1544 152464 1556
rect 152419 1516 152464 1544
rect 152458 1504 152464 1516
rect 152516 1504 152522 1556
rect 154022 1504 154028 1556
rect 154080 1544 154086 1556
rect 154209 1547 154267 1553
rect 154209 1544 154221 1547
rect 154080 1516 154221 1544
rect 154080 1504 154086 1516
rect 154209 1513 154221 1516
rect 154255 1513 154267 1547
rect 154209 1507 154267 1513
rect 155236 1516 155448 1544
rect 114281 1479 114339 1485
rect 114281 1476 114293 1479
rect 107519 1448 109172 1476
rect 109512 1448 114293 1476
rect 107519 1445 107531 1448
rect 107473 1439 107531 1445
rect 105633 1411 105691 1417
rect 105633 1377 105645 1411
rect 105679 1377 105691 1411
rect 105633 1371 105691 1377
rect 105814 1368 105820 1420
rect 105872 1408 105878 1420
rect 106826 1408 106832 1420
rect 105872 1380 106688 1408
rect 106787 1380 106832 1408
rect 105872 1368 105878 1380
rect 104526 1300 104532 1352
rect 104584 1340 104590 1352
rect 104713 1343 104771 1349
rect 104713 1340 104725 1343
rect 104584 1312 104725 1340
rect 104584 1300 104590 1312
rect 104713 1309 104725 1312
rect 104759 1309 104771 1343
rect 106660 1340 106688 1380
rect 106826 1368 106832 1380
rect 106884 1368 106890 1420
rect 108485 1411 108543 1417
rect 106936 1380 108436 1408
rect 106936 1340 106964 1380
rect 106660 1312 106964 1340
rect 108408 1340 108436 1380
rect 108485 1377 108497 1411
rect 108531 1408 108543 1411
rect 109402 1408 109408 1420
rect 108531 1380 109408 1408
rect 108531 1377 108543 1380
rect 108485 1371 108543 1377
rect 109402 1368 109408 1380
rect 109460 1368 109466 1420
rect 108577 1343 108635 1349
rect 108577 1340 108589 1343
rect 108408 1312 108589 1340
rect 104713 1303 104771 1309
rect 108577 1309 108589 1312
rect 108623 1309 108635 1343
rect 108577 1303 108635 1309
rect 108298 1272 108304 1284
rect 104452 1244 108304 1272
rect 108298 1232 108304 1244
rect 108356 1232 108362 1284
rect 99190 1204 99196 1216
rect 99151 1176 99196 1204
rect 99190 1164 99196 1176
rect 99248 1164 99254 1216
rect 108574 1164 108580 1216
rect 108632 1204 108638 1216
rect 109512 1204 109540 1448
rect 114281 1445 114293 1448
rect 114327 1445 114339 1479
rect 118878 1476 118884 1488
rect 114281 1439 114339 1445
rect 115216 1448 118884 1476
rect 109589 1411 109647 1417
rect 109589 1377 109601 1411
rect 109635 1408 109647 1411
rect 110598 1408 110604 1420
rect 109635 1380 110460 1408
rect 110559 1380 110604 1408
rect 109635 1377 109647 1380
rect 109589 1371 109647 1377
rect 110432 1340 110460 1380
rect 110598 1368 110604 1380
rect 110656 1368 110662 1420
rect 110690 1368 110696 1420
rect 110748 1408 110754 1420
rect 112346 1408 112352 1420
rect 110748 1380 110793 1408
rect 110892 1380 112352 1408
rect 110748 1368 110754 1380
rect 110892 1340 110920 1380
rect 112346 1368 112352 1380
rect 112404 1368 112410 1420
rect 112441 1411 112499 1417
rect 112441 1377 112453 1411
rect 112487 1408 112499 1411
rect 114189 1411 114247 1417
rect 112487 1380 114140 1408
rect 112487 1377 112499 1380
rect 112441 1371 112499 1377
rect 112530 1340 112536 1352
rect 110432 1312 110920 1340
rect 112491 1312 112536 1340
rect 112530 1300 112536 1312
rect 112588 1300 112594 1352
rect 114112 1340 114140 1380
rect 114189 1377 114201 1411
rect 114235 1408 114247 1411
rect 115216 1408 115244 1448
rect 118878 1436 118884 1448
rect 118936 1436 118942 1488
rect 122190 1476 122196 1488
rect 119172 1448 122196 1476
rect 114235 1380 115244 1408
rect 114235 1377 114247 1380
rect 114189 1371 114247 1377
rect 115290 1368 115296 1420
rect 115348 1408 115354 1420
rect 116305 1411 116363 1417
rect 115348 1380 115393 1408
rect 115348 1368 115354 1380
rect 116305 1377 116317 1411
rect 116351 1408 116363 1411
rect 118050 1408 118056 1420
rect 116351 1380 118056 1408
rect 116351 1377 116363 1380
rect 116305 1371 116363 1377
rect 118050 1368 118056 1380
rect 118108 1368 118114 1420
rect 118145 1411 118203 1417
rect 118145 1377 118157 1411
rect 118191 1408 118203 1411
rect 118786 1408 118792 1420
rect 118191 1380 118792 1408
rect 118191 1377 118203 1380
rect 118145 1371 118203 1377
rect 118786 1368 118792 1380
rect 118844 1368 118850 1420
rect 119172 1417 119200 1448
rect 122190 1436 122196 1448
rect 122248 1436 122254 1488
rect 122282 1436 122288 1488
rect 122340 1476 122346 1488
rect 123941 1479 123999 1485
rect 123941 1476 123953 1479
rect 122340 1448 123953 1476
rect 122340 1436 122346 1448
rect 123941 1445 123953 1448
rect 123987 1445 123999 1479
rect 123941 1439 123999 1445
rect 124674 1436 124680 1488
rect 124732 1476 124738 1488
rect 124953 1479 125011 1485
rect 124953 1476 124965 1479
rect 124732 1448 124965 1476
rect 124732 1436 124738 1448
rect 124953 1445 124965 1448
rect 124999 1445 125011 1479
rect 124953 1439 125011 1445
rect 125226 1436 125232 1488
rect 125284 1476 125290 1488
rect 127529 1479 127587 1485
rect 127529 1476 127541 1479
rect 125284 1448 127541 1476
rect 125284 1436 125290 1448
rect 127529 1445 127541 1448
rect 127575 1445 127587 1479
rect 127529 1439 127587 1445
rect 128541 1479 128599 1485
rect 128541 1445 128553 1479
rect 128587 1476 128599 1479
rect 129182 1476 129188 1488
rect 128587 1448 129188 1476
rect 128587 1445 128599 1448
rect 128541 1439 128599 1445
rect 129182 1436 129188 1448
rect 129240 1436 129246 1488
rect 129458 1436 129464 1488
rect 129516 1476 129522 1488
rect 135349 1479 135407 1485
rect 129516 1448 130516 1476
rect 129516 1436 129522 1448
rect 119157 1411 119215 1417
rect 119157 1377 119169 1411
rect 119203 1377 119215 1411
rect 121362 1408 121368 1420
rect 121323 1380 121368 1408
rect 119157 1371 119215 1377
rect 121362 1368 121368 1380
rect 121420 1368 121426 1420
rect 122745 1411 122803 1417
rect 122745 1377 122757 1411
rect 122791 1408 122803 1411
rect 123754 1408 123760 1420
rect 122791 1380 123760 1408
rect 122791 1377 122803 1380
rect 122745 1371 122803 1377
rect 123754 1368 123760 1380
rect 123812 1368 123818 1420
rect 123849 1411 123907 1417
rect 123849 1377 123861 1411
rect 123895 1408 123907 1411
rect 124858 1408 124864 1420
rect 123895 1380 124720 1408
rect 124819 1380 124864 1408
rect 123895 1377 123907 1380
rect 123849 1371 123907 1377
rect 116486 1340 116492 1352
rect 114112 1312 116492 1340
rect 116486 1300 116492 1312
rect 116544 1300 116550 1352
rect 119338 1300 119344 1352
rect 119396 1340 119402 1352
rect 123386 1340 123392 1352
rect 119396 1312 123392 1340
rect 119396 1300 119402 1312
rect 123386 1300 123392 1312
rect 123444 1300 123450 1352
rect 124692 1340 124720 1380
rect 124858 1368 124864 1380
rect 124916 1368 124922 1420
rect 125042 1368 125048 1420
rect 125100 1408 125106 1420
rect 127437 1411 127495 1417
rect 125100 1380 127388 1408
rect 125100 1368 125106 1380
rect 125134 1340 125140 1352
rect 124692 1312 125140 1340
rect 125134 1300 125140 1312
rect 125192 1300 125198 1352
rect 127360 1340 127388 1380
rect 127437 1377 127449 1411
rect 127483 1408 127495 1411
rect 128078 1408 128084 1420
rect 127483 1380 128084 1408
rect 127483 1377 127495 1380
rect 127437 1371 127495 1377
rect 128078 1368 128084 1380
rect 128136 1368 128142 1420
rect 128446 1408 128452 1420
rect 128407 1380 128452 1408
rect 128446 1368 128452 1380
rect 128504 1368 128510 1420
rect 129553 1411 129611 1417
rect 129553 1377 129565 1411
rect 129599 1408 129611 1411
rect 129642 1408 129648 1420
rect 129599 1380 129648 1408
rect 129599 1377 129611 1380
rect 129553 1371 129611 1377
rect 129642 1368 129648 1380
rect 129700 1368 129706 1420
rect 127802 1340 127808 1352
rect 127360 1312 127808 1340
rect 127802 1300 127808 1312
rect 127860 1300 127866 1352
rect 130488 1340 130516 1448
rect 130580 1448 135116 1476
rect 130580 1417 130608 1448
rect 130565 1411 130623 1417
rect 130565 1377 130577 1411
rect 130611 1377 130623 1411
rect 130565 1371 130623 1377
rect 130657 1411 130715 1417
rect 130657 1377 130669 1411
rect 130703 1377 130715 1411
rect 132402 1408 132408 1420
rect 132363 1380 132408 1408
rect 130657 1371 130715 1377
rect 130672 1340 130700 1371
rect 132402 1368 132408 1380
rect 132460 1368 132466 1420
rect 132497 1411 132555 1417
rect 132497 1377 132509 1411
rect 132543 1408 132555 1411
rect 133230 1408 133236 1420
rect 132543 1380 133236 1408
rect 132543 1377 132555 1380
rect 132497 1371 132555 1377
rect 133230 1368 133236 1380
rect 133288 1368 133294 1420
rect 133414 1408 133420 1420
rect 133375 1380 133420 1408
rect 133414 1368 133420 1380
rect 133472 1368 133478 1420
rect 133509 1411 133567 1417
rect 133509 1377 133521 1411
rect 133555 1408 133567 1411
rect 134058 1408 134064 1420
rect 133555 1380 134064 1408
rect 133555 1377 133567 1380
rect 133509 1371 133567 1377
rect 134058 1368 134064 1380
rect 134116 1368 134122 1420
rect 134978 1340 134984 1352
rect 130488 1312 130700 1340
rect 131684 1312 134984 1340
rect 112162 1232 112168 1284
rect 112220 1272 112226 1284
rect 115385 1275 115443 1281
rect 115385 1272 115397 1275
rect 112220 1244 115397 1272
rect 112220 1232 112226 1244
rect 115385 1241 115397 1244
rect 115431 1241 115443 1275
rect 115385 1235 115443 1241
rect 118142 1232 118148 1284
rect 118200 1272 118206 1284
rect 127526 1272 127532 1284
rect 118200 1244 127532 1272
rect 118200 1232 118206 1244
rect 127526 1232 127532 1244
rect 127584 1232 127590 1284
rect 127894 1232 127900 1284
rect 127952 1272 127958 1284
rect 129090 1272 129096 1284
rect 127952 1244 129096 1272
rect 127952 1232 127958 1244
rect 129090 1232 129096 1244
rect 129148 1232 129154 1284
rect 129274 1232 129280 1284
rect 129332 1272 129338 1284
rect 129645 1275 129703 1281
rect 129645 1272 129657 1275
rect 129332 1244 129657 1272
rect 129332 1232 129338 1244
rect 129645 1241 129657 1244
rect 129691 1241 129703 1275
rect 129645 1235 129703 1241
rect 108632 1176 109540 1204
rect 108632 1164 108638 1176
rect 117038 1164 117044 1216
rect 117096 1204 117102 1216
rect 119249 1207 119307 1213
rect 119249 1204 119261 1207
rect 117096 1176 119261 1204
rect 117096 1164 117102 1176
rect 119249 1173 119261 1176
rect 119295 1173 119307 1207
rect 119249 1167 119307 1173
rect 120534 1164 120540 1216
rect 120592 1204 120598 1216
rect 125226 1204 125232 1216
rect 120592 1176 125232 1204
rect 120592 1164 120598 1176
rect 125226 1164 125232 1176
rect 125284 1164 125290 1216
rect 125962 1164 125968 1216
rect 126020 1204 126026 1216
rect 127434 1204 127440 1216
rect 126020 1176 127440 1204
rect 126020 1164 126026 1176
rect 127434 1164 127440 1176
rect 127492 1164 127498 1216
rect 127618 1164 127624 1216
rect 127676 1204 127682 1216
rect 131684 1204 131712 1312
rect 134978 1300 134984 1312
rect 135036 1300 135042 1352
rect 135088 1340 135116 1448
rect 135349 1445 135361 1479
rect 135395 1476 135407 1479
rect 135438 1476 135444 1488
rect 135395 1448 135444 1476
rect 135395 1445 135407 1448
rect 135349 1439 135407 1445
rect 135438 1436 135444 1448
rect 135496 1436 135502 1488
rect 135622 1436 135628 1488
rect 135680 1476 135686 1488
rect 136174 1476 136180 1488
rect 135680 1448 136180 1476
rect 135680 1436 135686 1448
rect 136174 1436 136180 1448
rect 136232 1436 136238 1488
rect 136358 1476 136364 1488
rect 136319 1448 136364 1476
rect 136358 1436 136364 1448
rect 136416 1436 136422 1488
rect 136818 1436 136824 1488
rect 136876 1476 136882 1488
rect 137830 1476 137836 1488
rect 136876 1448 137836 1476
rect 136876 1436 136882 1448
rect 137830 1436 137836 1448
rect 137888 1436 137894 1488
rect 137922 1436 137928 1488
rect 137980 1476 137986 1488
rect 138842 1476 138848 1488
rect 137980 1448 138848 1476
rect 137980 1436 137986 1448
rect 138842 1436 138848 1448
rect 138900 1436 138906 1488
rect 142982 1476 142988 1488
rect 141068 1448 142988 1476
rect 135254 1408 135260 1420
rect 135215 1380 135260 1408
rect 135254 1368 135260 1380
rect 135312 1368 135318 1420
rect 136269 1411 136327 1417
rect 136269 1377 136281 1411
rect 136315 1408 136327 1411
rect 137002 1408 137008 1420
rect 136315 1380 137008 1408
rect 136315 1377 136327 1380
rect 136269 1371 136327 1377
rect 137002 1368 137008 1380
rect 137060 1368 137066 1420
rect 137186 1368 137192 1420
rect 137244 1408 137250 1420
rect 138566 1408 138572 1420
rect 137244 1380 138572 1408
rect 137244 1368 137250 1380
rect 138566 1368 138572 1380
rect 138624 1368 138630 1420
rect 138934 1408 138940 1420
rect 138895 1380 138940 1408
rect 138934 1368 138940 1380
rect 138992 1368 138998 1420
rect 139026 1368 139032 1420
rect 139084 1408 139090 1420
rect 139084 1380 139129 1408
rect 139084 1368 139090 1380
rect 139670 1368 139676 1420
rect 139728 1408 139734 1420
rect 141068 1408 141096 1448
rect 142982 1436 142988 1448
rect 143040 1436 143046 1488
rect 144914 1476 144920 1488
rect 144012 1448 144920 1476
rect 139728 1380 141096 1408
rect 139728 1368 139734 1380
rect 141142 1368 141148 1420
rect 141200 1408 141206 1420
rect 141200 1380 141245 1408
rect 141200 1368 141206 1380
rect 141510 1368 141516 1420
rect 141568 1408 141574 1420
rect 143810 1408 143816 1420
rect 141568 1380 143816 1408
rect 141568 1368 141574 1380
rect 143810 1368 143816 1380
rect 143868 1368 143874 1420
rect 144012 1417 144040 1448
rect 144914 1436 144920 1448
rect 144972 1436 144978 1488
rect 145098 1436 145104 1488
rect 145156 1476 145162 1488
rect 145156 1448 145201 1476
rect 145392 1448 146892 1476
rect 145156 1436 145162 1448
rect 143997 1411 144055 1417
rect 143997 1377 144009 1411
rect 144043 1377 144055 1411
rect 143997 1371 144055 1377
rect 144089 1411 144147 1417
rect 144089 1377 144101 1411
rect 144135 1408 144147 1411
rect 144638 1408 144644 1420
rect 144135 1380 144644 1408
rect 144135 1377 144147 1380
rect 144089 1371 144147 1377
rect 144638 1368 144644 1380
rect 144696 1368 144702 1420
rect 145009 1411 145067 1417
rect 145009 1377 145021 1411
rect 145055 1377 145067 1411
rect 145009 1371 145067 1377
rect 137094 1340 137100 1352
rect 135088 1312 137100 1340
rect 137094 1300 137100 1312
rect 137152 1300 137158 1352
rect 137278 1300 137284 1352
rect 137336 1340 137342 1352
rect 140961 1343 141019 1349
rect 140961 1340 140973 1343
rect 137336 1312 140973 1340
rect 137336 1300 137342 1312
rect 140961 1309 140973 1312
rect 141007 1309 141019 1343
rect 145024 1340 145052 1371
rect 145392 1340 145420 1448
rect 145466 1368 145472 1420
rect 145524 1408 145530 1420
rect 146662 1408 146668 1420
rect 145524 1380 145696 1408
rect 146623 1380 146668 1408
rect 145524 1368 145530 1380
rect 145024 1312 145420 1340
rect 140961 1303 141019 1309
rect 133325 1275 133383 1281
rect 133325 1241 133337 1275
rect 133371 1272 133383 1275
rect 133414 1272 133420 1284
rect 133371 1244 133420 1272
rect 133371 1241 133383 1244
rect 133325 1235 133383 1241
rect 133414 1232 133420 1244
rect 133472 1272 133478 1284
rect 141510 1272 141516 1284
rect 133472 1244 141516 1272
rect 133472 1232 133478 1244
rect 141510 1232 141516 1244
rect 141568 1232 141574 1284
rect 144638 1272 144644 1284
rect 141804 1244 144644 1272
rect 127676 1176 131712 1204
rect 127676 1164 127682 1176
rect 133690 1164 133696 1216
rect 133748 1204 133754 1216
rect 138842 1204 138848 1216
rect 133748 1176 138848 1204
rect 133748 1164 133754 1176
rect 138842 1164 138848 1176
rect 138900 1164 138906 1216
rect 139118 1164 139124 1216
rect 139176 1204 139182 1216
rect 140682 1204 140688 1216
rect 139176 1176 140688 1204
rect 139176 1164 139182 1176
rect 140682 1164 140688 1176
rect 140740 1164 140746 1216
rect 140961 1207 141019 1213
rect 140961 1173 140973 1207
rect 141007 1204 141019 1207
rect 141804 1204 141832 1244
rect 144638 1232 144644 1244
rect 144696 1232 144702 1284
rect 141007 1176 141832 1204
rect 141007 1173 141019 1176
rect 140961 1167 141019 1173
rect 142890 1164 142896 1216
rect 142948 1204 142954 1216
rect 145006 1204 145012 1216
rect 142948 1176 145012 1204
rect 142948 1164 142954 1176
rect 145006 1164 145012 1176
rect 145064 1164 145070 1216
rect 145668 1204 145696 1380
rect 146662 1368 146668 1380
rect 146720 1368 146726 1420
rect 146864 1408 146892 1448
rect 146938 1436 146944 1488
rect 146996 1476 147002 1488
rect 148778 1476 148784 1488
rect 146996 1448 148784 1476
rect 146996 1436 147002 1448
rect 148778 1436 148784 1448
rect 148836 1436 148842 1488
rect 155236 1476 155264 1516
rect 154132 1448 155264 1476
rect 155420 1476 155448 1516
rect 155678 1504 155684 1556
rect 155736 1544 155742 1556
rect 161014 1544 161020 1556
rect 155736 1516 159956 1544
rect 160975 1516 161020 1544
rect 155736 1504 155742 1516
rect 159818 1476 159824 1488
rect 155420 1448 159680 1476
rect 159779 1448 159824 1476
rect 149054 1408 149060 1420
rect 146864 1380 149060 1408
rect 149054 1368 149060 1380
rect 149112 1368 149118 1420
rect 150250 1408 150256 1420
rect 150211 1380 150256 1408
rect 150250 1368 150256 1380
rect 150308 1368 150314 1420
rect 152369 1411 152427 1417
rect 152369 1377 152381 1411
rect 152415 1408 152427 1411
rect 153838 1408 153844 1420
rect 152415 1380 153844 1408
rect 152415 1377 152427 1380
rect 152369 1371 152427 1377
rect 153838 1368 153844 1380
rect 153896 1368 153902 1420
rect 154132 1417 154160 1448
rect 154117 1411 154175 1417
rect 154117 1377 154129 1411
rect 154163 1377 154175 1411
rect 155213 1411 155271 1417
rect 155213 1408 155225 1411
rect 154117 1371 154175 1377
rect 155144 1380 155225 1408
rect 155034 1300 155040 1352
rect 155092 1340 155098 1352
rect 155144 1340 155172 1380
rect 155213 1377 155225 1380
rect 155259 1377 155271 1411
rect 156322 1408 156328 1420
rect 155213 1371 155271 1377
rect 155420 1380 156328 1408
rect 155092 1312 155172 1340
rect 155313 1343 155371 1349
rect 155092 1300 155098 1312
rect 155313 1309 155325 1343
rect 155359 1340 155371 1343
rect 155420 1340 155448 1380
rect 156322 1368 156328 1380
rect 156380 1368 156386 1420
rect 157242 1368 157248 1420
rect 157300 1408 157306 1420
rect 158993 1411 159051 1417
rect 158993 1408 159005 1411
rect 157300 1380 159005 1408
rect 157300 1368 157306 1380
rect 158993 1377 159005 1380
rect 159039 1377 159051 1411
rect 159652 1408 159680 1448
rect 159818 1436 159824 1448
rect 159876 1436 159882 1488
rect 159928 1476 159956 1516
rect 161014 1504 161020 1516
rect 161072 1504 161078 1556
rect 161198 1504 161204 1556
rect 161256 1544 161262 1556
rect 162486 1544 162492 1556
rect 161256 1516 162492 1544
rect 161256 1504 161262 1516
rect 162486 1504 162492 1516
rect 162544 1504 162550 1556
rect 163682 1544 163688 1556
rect 162596 1516 163688 1544
rect 162118 1476 162124 1488
rect 159928 1448 162124 1476
rect 162118 1436 162124 1448
rect 162176 1436 162182 1488
rect 160646 1408 160652 1420
rect 159652 1380 160652 1408
rect 158993 1371 159051 1377
rect 160646 1368 160652 1380
rect 160704 1368 160710 1420
rect 160925 1411 160983 1417
rect 160925 1377 160937 1411
rect 160971 1408 160983 1411
rect 162596 1408 162624 1516
rect 163682 1504 163688 1516
rect 163740 1504 163746 1556
rect 164344 1516 164924 1544
rect 164344 1476 164372 1516
rect 164510 1476 164516 1488
rect 162688 1448 164372 1476
rect 164471 1448 164516 1476
rect 162688 1417 162716 1448
rect 164510 1436 164516 1448
rect 164568 1436 164574 1488
rect 164896 1476 164924 1516
rect 164970 1504 164976 1556
rect 165028 1544 165034 1556
rect 168377 1547 168435 1553
rect 165028 1516 168052 1544
rect 165028 1504 165034 1516
rect 165246 1476 165252 1488
rect 164896 1448 165252 1476
rect 165246 1436 165252 1448
rect 165304 1436 165310 1488
rect 165522 1436 165528 1488
rect 165580 1476 165586 1488
rect 165580 1448 165625 1476
rect 165580 1436 165586 1448
rect 160971 1380 162624 1408
rect 162673 1411 162731 1417
rect 160971 1377 160983 1380
rect 160925 1371 160983 1377
rect 162673 1377 162685 1411
rect 162719 1377 162731 1411
rect 162673 1371 162731 1377
rect 162762 1368 162768 1420
rect 162820 1408 162826 1420
rect 162820 1380 162865 1408
rect 162820 1368 162826 1380
rect 163590 1368 163596 1420
rect 163648 1408 163654 1420
rect 164970 1408 164976 1420
rect 163648 1380 164976 1408
rect 163648 1368 163654 1380
rect 164970 1368 164976 1380
rect 165028 1368 165034 1420
rect 165062 1368 165068 1420
rect 165120 1408 165126 1420
rect 167914 1408 167920 1420
rect 165120 1380 167920 1408
rect 165120 1368 165126 1380
rect 167914 1368 167920 1380
rect 167972 1368 167978 1420
rect 168024 1408 168052 1516
rect 168377 1513 168389 1547
rect 168423 1544 168435 1547
rect 169294 1544 169300 1556
rect 168423 1516 169300 1544
rect 168423 1513 168435 1516
rect 168377 1507 168435 1513
rect 169294 1504 169300 1516
rect 169352 1504 169358 1556
rect 169849 1547 169907 1553
rect 169849 1513 169861 1547
rect 169895 1544 169907 1547
rect 170030 1544 170036 1556
rect 169895 1516 170036 1544
rect 169895 1513 169907 1516
rect 169849 1507 169907 1513
rect 170030 1504 170036 1516
rect 170088 1504 170094 1556
rect 174906 1544 174912 1556
rect 171060 1516 174912 1544
rect 168098 1436 168104 1488
rect 168156 1476 168162 1488
rect 169938 1476 169944 1488
rect 168156 1448 169944 1476
rect 168156 1436 168162 1448
rect 169938 1436 169944 1448
rect 169996 1436 170002 1488
rect 169386 1408 169392 1420
rect 168024 1380 169392 1408
rect 169386 1368 169392 1380
rect 169444 1368 169450 1420
rect 169757 1411 169815 1417
rect 169757 1377 169769 1411
rect 169803 1408 169815 1411
rect 171060 1408 171088 1516
rect 174906 1504 174912 1516
rect 174964 1504 174970 1556
rect 175734 1544 175740 1556
rect 175016 1516 175740 1544
rect 171318 1476 171324 1488
rect 171279 1448 171324 1476
rect 171318 1436 171324 1448
rect 171376 1436 171382 1488
rect 173066 1476 173072 1488
rect 172348 1448 173072 1476
rect 171226 1408 171232 1420
rect 169803 1380 171088 1408
rect 171187 1380 171232 1408
rect 169803 1377 169815 1380
rect 169757 1371 169815 1377
rect 171226 1368 171232 1380
rect 171284 1368 171290 1420
rect 172348 1417 172376 1448
rect 173066 1436 173072 1448
rect 173124 1436 173130 1488
rect 173437 1479 173495 1485
rect 173437 1476 173449 1479
rect 173268 1448 173449 1476
rect 173268 1420 173296 1448
rect 173437 1445 173449 1448
rect 173483 1445 173495 1479
rect 173437 1439 173495 1445
rect 173618 1436 173624 1488
rect 173676 1476 173682 1488
rect 174446 1476 174452 1488
rect 173676 1448 174452 1476
rect 173676 1436 173682 1448
rect 174446 1436 174452 1448
rect 174504 1436 174510 1488
rect 172333 1411 172391 1417
rect 172333 1377 172345 1411
rect 172379 1377 172391 1411
rect 172333 1371 172391 1377
rect 172422 1368 172428 1420
rect 172480 1408 172486 1420
rect 172480 1380 172525 1408
rect 172480 1368 172486 1380
rect 173250 1368 173256 1420
rect 173308 1368 173314 1420
rect 173342 1368 173348 1420
rect 173400 1408 173406 1420
rect 173400 1380 173445 1408
rect 173400 1368 173406 1380
rect 173526 1368 173532 1420
rect 173584 1408 173590 1420
rect 175016 1408 175044 1516
rect 175734 1504 175740 1516
rect 175792 1504 175798 1556
rect 176562 1504 176568 1556
rect 176620 1544 176626 1556
rect 178221 1547 178279 1553
rect 178221 1544 178233 1547
rect 176620 1516 178233 1544
rect 176620 1504 176626 1516
rect 178221 1513 178233 1516
rect 178267 1513 178279 1547
rect 178221 1507 178279 1513
rect 178310 1504 178316 1556
rect 178368 1544 178374 1556
rect 179233 1547 179291 1553
rect 179233 1544 179245 1547
rect 178368 1516 179245 1544
rect 178368 1504 178374 1516
rect 179233 1513 179245 1516
rect 179279 1513 179291 1547
rect 179233 1507 179291 1513
rect 179322 1504 179328 1556
rect 179380 1544 179386 1556
rect 182266 1544 182272 1556
rect 179380 1516 182272 1544
rect 179380 1504 179386 1516
rect 182266 1504 182272 1516
rect 182324 1504 182330 1556
rect 182361 1547 182419 1553
rect 182361 1513 182373 1547
rect 182407 1544 182419 1547
rect 183554 1544 183560 1556
rect 182407 1516 183560 1544
rect 182407 1513 182419 1516
rect 182361 1507 182419 1513
rect 183554 1504 183560 1516
rect 183612 1504 183618 1556
rect 184661 1547 184719 1553
rect 184661 1513 184673 1547
rect 184707 1544 184719 1547
rect 184750 1544 184756 1556
rect 184707 1516 184756 1544
rect 184707 1513 184719 1516
rect 184661 1507 184719 1513
rect 184750 1504 184756 1516
rect 184808 1504 184814 1556
rect 185486 1504 185492 1556
rect 185544 1544 185550 1556
rect 187329 1547 187387 1553
rect 187329 1544 187341 1547
rect 185544 1516 187341 1544
rect 185544 1504 185550 1516
rect 187329 1513 187341 1516
rect 187375 1513 187387 1547
rect 187329 1507 187387 1513
rect 187878 1504 187884 1556
rect 187936 1544 187942 1556
rect 188341 1547 188399 1553
rect 188341 1544 188353 1547
rect 187936 1516 188353 1544
rect 187936 1504 187942 1516
rect 188341 1513 188353 1516
rect 188387 1513 188399 1547
rect 188341 1507 188399 1513
rect 188982 1504 188988 1556
rect 189040 1544 189046 1556
rect 189537 1547 189595 1553
rect 189537 1544 189549 1547
rect 189040 1516 189549 1544
rect 189040 1504 189046 1516
rect 189537 1513 189549 1516
rect 189583 1513 189595 1547
rect 191285 1547 191343 1553
rect 191285 1544 191297 1547
rect 189537 1507 189595 1513
rect 191116 1516 191297 1544
rect 175200 1448 176792 1476
rect 175200 1417 175228 1448
rect 173584 1380 175044 1408
rect 175185 1411 175243 1417
rect 173584 1368 173590 1380
rect 175185 1377 175197 1411
rect 175231 1377 175243 1411
rect 176102 1408 176108 1420
rect 175185 1371 175243 1377
rect 175292 1380 176108 1408
rect 155359 1312 155448 1340
rect 155359 1309 155371 1312
rect 155313 1303 155371 1309
rect 155494 1300 155500 1352
rect 155552 1340 155558 1352
rect 156046 1340 156052 1352
rect 155552 1312 156052 1340
rect 155552 1300 155558 1312
rect 156046 1300 156052 1312
rect 156104 1300 156110 1352
rect 159082 1300 159088 1352
rect 159140 1340 159146 1352
rect 162026 1340 162032 1352
rect 159140 1312 162032 1340
rect 159140 1300 159146 1312
rect 162026 1300 162032 1312
rect 162084 1300 162090 1352
rect 162394 1300 162400 1352
rect 162452 1340 162458 1352
rect 164326 1340 164332 1352
rect 162452 1312 164332 1340
rect 162452 1300 162458 1312
rect 164326 1300 164332 1312
rect 164384 1300 164390 1352
rect 164878 1300 164884 1352
rect 164936 1340 164942 1352
rect 166902 1340 166908 1352
rect 164936 1312 166908 1340
rect 164936 1300 164942 1312
rect 166902 1300 166908 1312
rect 166960 1300 166966 1352
rect 167362 1340 167368 1352
rect 167323 1312 167368 1340
rect 167362 1300 167368 1312
rect 167420 1300 167426 1352
rect 167454 1300 167460 1352
rect 167512 1340 167518 1352
rect 175292 1340 175320 1380
rect 176102 1368 176108 1380
rect 176160 1368 176166 1420
rect 176197 1411 176255 1417
rect 176197 1377 176209 1411
rect 176243 1408 176255 1411
rect 176764 1408 176792 1448
rect 176838 1436 176844 1488
rect 176896 1476 176902 1488
rect 186130 1476 186136 1488
rect 176896 1448 186136 1476
rect 176896 1436 176902 1448
rect 186130 1436 186136 1448
rect 186188 1436 186194 1488
rect 186314 1436 186320 1488
rect 186372 1476 186378 1488
rect 188798 1476 188804 1488
rect 186372 1448 188804 1476
rect 186372 1436 186378 1448
rect 188798 1436 188804 1448
rect 188856 1436 188862 1488
rect 188890 1436 188896 1488
rect 188948 1476 188954 1488
rect 191116 1476 191144 1516
rect 191285 1513 191297 1516
rect 191331 1513 191343 1547
rect 191285 1507 191343 1513
rect 191374 1504 191380 1556
rect 191432 1544 191438 1556
rect 194962 1544 194968 1556
rect 191432 1516 194968 1544
rect 191432 1504 191438 1516
rect 194962 1504 194968 1516
rect 195020 1504 195026 1556
rect 193125 1479 193183 1485
rect 193125 1476 193137 1479
rect 188948 1448 191144 1476
rect 191208 1448 193137 1476
rect 188948 1436 188954 1448
rect 177482 1408 177488 1420
rect 176243 1380 176700 1408
rect 176764 1380 177488 1408
rect 176243 1377 176255 1380
rect 176197 1371 176255 1377
rect 167512 1312 175320 1340
rect 167512 1300 167518 1312
rect 175366 1300 175372 1352
rect 175424 1300 175430 1352
rect 176672 1340 176700 1380
rect 177482 1368 177488 1380
rect 177540 1368 177546 1420
rect 178126 1408 178132 1420
rect 178087 1380 178132 1408
rect 178126 1368 178132 1380
rect 178184 1368 178190 1420
rect 179141 1411 179199 1417
rect 178236 1380 179092 1408
rect 178236 1340 178264 1380
rect 176672 1312 178264 1340
rect 179064 1340 179092 1380
rect 179141 1377 179153 1411
rect 179187 1408 179199 1411
rect 181254 1408 181260 1420
rect 179187 1380 181116 1408
rect 181215 1380 181260 1408
rect 179187 1377 179199 1380
rect 179141 1371 179199 1377
rect 180518 1340 180524 1352
rect 179064 1312 180524 1340
rect 180518 1300 180524 1312
rect 180576 1300 180582 1352
rect 181088 1340 181116 1380
rect 181254 1368 181260 1380
rect 181312 1368 181318 1420
rect 182269 1411 182327 1417
rect 181364 1380 182220 1408
rect 181364 1340 181392 1380
rect 181088 1312 181392 1340
rect 182192 1340 182220 1380
rect 182269 1377 182281 1411
rect 182315 1408 182327 1411
rect 184569 1411 184627 1417
rect 182315 1380 184520 1408
rect 182315 1377 182327 1380
rect 182269 1371 182327 1377
rect 183186 1340 183192 1352
rect 182192 1312 183192 1340
rect 183186 1300 183192 1312
rect 183244 1300 183250 1352
rect 184492 1340 184520 1380
rect 184569 1377 184581 1411
rect 184615 1408 184627 1411
rect 186682 1408 186688 1420
rect 184615 1380 186688 1408
rect 184615 1377 184627 1380
rect 184569 1371 184627 1377
rect 186682 1368 186688 1380
rect 186740 1368 186746 1420
rect 186866 1368 186872 1420
rect 186924 1408 186930 1420
rect 187142 1408 187148 1420
rect 186924 1380 187148 1408
rect 186924 1368 186930 1380
rect 187142 1368 187148 1380
rect 187200 1368 187206 1420
rect 187237 1411 187295 1417
rect 187237 1377 187249 1411
rect 187283 1408 187295 1411
rect 188249 1411 188307 1417
rect 187283 1380 188200 1408
rect 187283 1377 187295 1380
rect 187237 1371 187295 1377
rect 186222 1340 186228 1352
rect 184492 1312 186228 1340
rect 186222 1300 186228 1312
rect 186280 1300 186286 1352
rect 145742 1232 145748 1284
rect 145800 1272 145806 1284
rect 175182 1272 175188 1284
rect 145800 1244 175188 1272
rect 145800 1232 145806 1244
rect 175182 1232 175188 1244
rect 175240 1232 175246 1284
rect 175277 1275 175335 1281
rect 175277 1241 175289 1275
rect 175323 1272 175335 1275
rect 175384 1272 175412 1300
rect 175323 1244 175412 1272
rect 175323 1241 175335 1244
rect 175277 1235 175335 1241
rect 175458 1232 175464 1284
rect 175516 1272 175522 1284
rect 176289 1275 176347 1281
rect 176289 1272 176301 1275
rect 175516 1244 176301 1272
rect 175516 1232 175522 1244
rect 176289 1241 176301 1244
rect 176335 1241 176347 1275
rect 186590 1272 186596 1284
rect 176289 1235 176347 1241
rect 176396 1244 186596 1272
rect 147858 1204 147864 1216
rect 145668 1176 147864 1204
rect 147858 1164 147864 1176
rect 147916 1164 147922 1216
rect 148226 1164 148232 1216
rect 148284 1204 148290 1216
rect 160094 1204 160100 1216
rect 148284 1176 160100 1204
rect 148284 1164 148290 1176
rect 160094 1164 160100 1176
rect 160152 1164 160158 1216
rect 162302 1164 162308 1216
rect 162360 1204 162366 1216
rect 162762 1204 162768 1216
rect 162360 1176 162768 1204
rect 162360 1164 162366 1176
rect 162762 1164 162768 1176
rect 162820 1164 162826 1216
rect 162854 1164 162860 1216
rect 162912 1204 162918 1216
rect 176396 1204 176424 1244
rect 186590 1232 186596 1244
rect 186648 1232 186654 1284
rect 188172 1272 188200 1380
rect 188249 1377 188261 1411
rect 188295 1377 188307 1411
rect 188249 1371 188307 1377
rect 188264 1340 188292 1371
rect 188430 1368 188436 1420
rect 188488 1408 188494 1420
rect 191208 1417 191236 1448
rect 193125 1445 193137 1448
rect 193171 1445 193183 1479
rect 193125 1439 193183 1445
rect 189445 1411 189503 1417
rect 189445 1408 189457 1411
rect 188488 1380 189457 1408
rect 188488 1368 188494 1380
rect 189445 1377 189457 1380
rect 189491 1377 189503 1411
rect 189445 1371 189503 1377
rect 191201 1411 191259 1417
rect 191201 1377 191213 1411
rect 191247 1377 191259 1411
rect 193306 1408 193312 1420
rect 193267 1380 193312 1408
rect 191201 1371 191259 1377
rect 193306 1368 193312 1380
rect 193364 1368 193370 1420
rect 194045 1411 194103 1417
rect 194045 1377 194057 1411
rect 194091 1408 194103 1411
rect 195054 1408 195060 1420
rect 194091 1380 195060 1408
rect 194091 1377 194103 1380
rect 194045 1371 194103 1377
rect 195054 1368 195060 1380
rect 195112 1368 195118 1420
rect 195146 1368 195152 1420
rect 195204 1408 195210 1420
rect 195977 1411 196035 1417
rect 195204 1380 195249 1408
rect 195204 1368 195210 1380
rect 195977 1377 195989 1411
rect 196023 1408 196035 1411
rect 198458 1408 198464 1420
rect 196023 1380 198464 1408
rect 196023 1377 196035 1380
rect 195977 1371 196035 1377
rect 198458 1368 198464 1380
rect 198516 1368 198522 1420
rect 191374 1340 191380 1352
rect 188264 1312 191380 1340
rect 191374 1300 191380 1312
rect 191432 1300 191438 1352
rect 193125 1343 193183 1349
rect 193125 1309 193137 1343
rect 193171 1340 193183 1343
rect 196710 1340 196716 1352
rect 193171 1312 196716 1340
rect 193171 1309 193183 1312
rect 193125 1303 193183 1309
rect 196710 1300 196716 1312
rect 196768 1300 196774 1352
rect 195790 1272 195796 1284
rect 188172 1244 195796 1272
rect 195790 1232 195796 1244
rect 195848 1232 195854 1284
rect 162912 1176 176424 1204
rect 162912 1164 162918 1176
rect 176470 1164 176476 1216
rect 176528 1204 176534 1216
rect 178770 1204 178776 1216
rect 176528 1176 178776 1204
rect 176528 1164 176534 1176
rect 178770 1164 178776 1176
rect 178828 1164 178834 1216
rect 181346 1204 181352 1216
rect 181307 1176 181352 1204
rect 181346 1164 181352 1176
rect 181404 1164 181410 1216
rect 181622 1164 181628 1216
rect 181680 1204 181686 1216
rect 182266 1204 182272 1216
rect 181680 1176 182272 1204
rect 181680 1164 181686 1176
rect 182266 1164 182272 1176
rect 182324 1164 182330 1216
rect 1104 1114 198812 1136
rect 1104 1062 4078 1114
rect 4130 1062 44078 1114
rect 44130 1062 84078 1114
rect 84130 1062 124078 1114
rect 124130 1062 164078 1114
rect 164130 1062 198812 1114
rect 1104 1040 198812 1062
rect 108114 960 108120 1012
rect 108172 1000 108178 1012
rect 112162 1000 112168 1012
rect 108172 972 112168 1000
rect 108172 960 108178 972
rect 112162 960 112168 972
rect 112220 960 112226 1012
rect 117774 960 117780 1012
rect 117832 1000 117838 1012
rect 117832 972 133184 1000
rect 117832 960 117838 972
rect 108022 892 108028 944
rect 108080 932 108086 944
rect 113450 932 113456 944
rect 108080 904 113456 932
rect 108080 892 108086 904
rect 113450 892 113456 904
rect 113508 892 113514 944
rect 115658 932 115664 944
rect 113560 904 115664 932
rect 106734 824 106740 876
rect 106792 864 106798 876
rect 113560 864 113588 904
rect 115658 892 115664 904
rect 115716 892 115722 944
rect 118878 892 118884 944
rect 118936 932 118942 944
rect 123938 932 123944 944
rect 118936 904 123944 932
rect 118936 892 118942 904
rect 123938 892 123944 904
rect 123996 892 124002 944
rect 126238 892 126244 944
rect 126296 932 126302 944
rect 130010 932 130016 944
rect 126296 904 130016 932
rect 126296 892 126302 904
rect 130010 892 130016 904
rect 130068 892 130074 944
rect 130102 892 130108 944
rect 130160 932 130166 944
rect 133046 932 133052 944
rect 130160 904 133052 932
rect 130160 892 130166 904
rect 133046 892 133052 904
rect 133104 892 133110 944
rect 106792 836 113588 864
rect 106792 824 106798 836
rect 115106 824 115112 876
rect 115164 864 115170 876
rect 127618 864 127624 876
rect 115164 836 127624 864
rect 115164 824 115170 836
rect 127618 824 127624 836
rect 127676 824 127682 876
rect 127986 824 127992 876
rect 128044 864 128050 876
rect 132494 864 132500 876
rect 128044 836 132500 864
rect 128044 824 128050 836
rect 132494 824 132500 836
rect 132552 824 132558 876
rect 133156 864 133184 972
rect 133782 960 133788 1012
rect 133840 1000 133846 1012
rect 134794 1000 134800 1012
rect 133840 972 134800 1000
rect 133840 960 133846 972
rect 134794 960 134800 972
rect 134852 960 134858 1012
rect 134886 960 134892 1012
rect 134944 1000 134950 1012
rect 137278 1000 137284 1012
rect 134944 972 137284 1000
rect 134944 960 134950 972
rect 137278 960 137284 972
rect 137336 960 137342 1012
rect 137557 1003 137615 1009
rect 137557 969 137569 1003
rect 137603 1000 137615 1003
rect 144917 1003 144975 1009
rect 144917 1000 144929 1003
rect 137603 972 144929 1000
rect 137603 969 137615 972
rect 137557 963 137615 969
rect 144917 969 144929 972
rect 144963 969 144975 1003
rect 144917 963 144975 969
rect 145009 1003 145067 1009
rect 145009 969 145021 1003
rect 145055 1000 145067 1003
rect 149698 1000 149704 1012
rect 145055 972 149704 1000
rect 145055 969 145067 972
rect 145009 963 145067 969
rect 149698 960 149704 972
rect 149756 960 149762 1012
rect 152918 960 152924 1012
rect 152976 1000 152982 1012
rect 162854 1000 162860 1012
rect 152976 972 162860 1000
rect 152976 960 152982 972
rect 162854 960 162860 972
rect 162912 960 162918 1012
rect 162946 960 162952 1012
rect 163004 1000 163010 1012
rect 165985 1003 166043 1009
rect 165985 1000 165997 1003
rect 163004 972 165997 1000
rect 163004 960 163010 972
rect 165985 969 165997 972
rect 166031 969 166043 1003
rect 165985 963 166043 969
rect 166074 960 166080 1012
rect 166132 1000 166138 1012
rect 166132 972 168420 1000
rect 166132 960 166138 972
rect 133233 935 133291 941
rect 133233 901 133245 935
rect 133279 932 133291 935
rect 140498 932 140504 944
rect 133279 904 140504 932
rect 133279 901 133291 904
rect 133233 895 133291 901
rect 140498 892 140504 904
rect 140556 892 140562 944
rect 140682 892 140688 944
rect 140740 932 140746 944
rect 143721 935 143779 941
rect 143721 932 143733 935
rect 140740 904 143733 932
rect 140740 892 140746 904
rect 143721 901 143733 904
rect 143767 901 143779 935
rect 143721 895 143779 901
rect 144546 892 144552 944
rect 144604 932 144610 944
rect 149793 935 149851 941
rect 149793 932 149805 935
rect 144604 904 149805 932
rect 144604 892 144610 904
rect 149793 901 149805 904
rect 149839 901 149851 935
rect 149793 895 149851 901
rect 156874 892 156880 944
rect 156932 932 156938 944
rect 160462 932 160468 944
rect 156932 904 160468 932
rect 156932 892 156938 904
rect 160462 892 160468 904
rect 160520 892 160526 944
rect 160554 892 160560 944
rect 160612 932 160618 944
rect 161937 935 161995 941
rect 161937 932 161949 935
rect 160612 904 161949 932
rect 160612 892 160618 904
rect 161937 901 161949 904
rect 161983 901 161995 935
rect 161937 895 161995 901
rect 162026 892 162032 944
rect 162084 932 162090 944
rect 168282 932 168288 944
rect 162084 904 168288 932
rect 162084 892 162090 904
rect 168282 892 168288 904
rect 168340 892 168346 944
rect 168392 932 168420 972
rect 169110 960 169116 1012
rect 169168 1000 169174 1012
rect 169168 972 172836 1000
rect 169168 960 169174 972
rect 172698 932 172704 944
rect 168392 904 172704 932
rect 172698 892 172704 904
rect 172756 892 172762 944
rect 172808 932 172836 972
rect 182100 972 182220 1000
rect 181438 932 181444 944
rect 172808 904 181444 932
rect 181438 892 181444 904
rect 181496 892 181502 944
rect 181530 892 181536 944
rect 181588 932 181594 944
rect 182100 932 182128 972
rect 182192 941 182220 972
rect 181588 904 182128 932
rect 182177 935 182235 941
rect 181588 892 181594 904
rect 182177 901 182189 935
rect 182223 901 182235 935
rect 182177 895 182235 901
rect 141881 867 141939 873
rect 141881 864 141893 867
rect 133156 836 141893 864
rect 141881 833 141893 836
rect 141927 833 141939 867
rect 141881 827 141939 833
rect 143810 824 143816 876
rect 143868 864 143874 876
rect 148226 864 148232 876
rect 143868 836 148232 864
rect 143868 824 143874 836
rect 148226 824 148232 836
rect 148284 824 148290 876
rect 152734 864 152740 876
rect 148796 836 152740 864
rect 119706 756 119712 808
rect 119764 796 119770 808
rect 129829 799 129887 805
rect 129829 796 129841 799
rect 119764 768 129841 796
rect 119764 756 119770 768
rect 129829 765 129841 768
rect 129875 765 129887 799
rect 129829 759 129887 765
rect 132402 756 132408 808
rect 132460 796 132466 808
rect 132460 768 135208 796
rect 132460 756 132466 768
rect 121362 688 121368 740
rect 121420 728 121426 740
rect 135073 731 135131 737
rect 135073 728 135085 731
rect 121420 700 135085 728
rect 121420 688 121426 700
rect 135073 697 135085 700
rect 135119 697 135131 731
rect 135073 691 135131 697
rect 133233 663 133291 669
rect 133233 660 133245 663
rect 129752 632 133245 660
rect 115290 552 115296 604
rect 115348 592 115354 604
rect 129752 592 129780 632
rect 133233 629 133245 632
rect 133279 629 133291 663
rect 135180 660 135208 768
rect 137094 756 137100 808
rect 137152 796 137158 808
rect 142890 796 142896 808
rect 137152 768 142896 796
rect 137152 756 137158 768
rect 142890 756 142896 768
rect 142948 756 142954 808
rect 142982 756 142988 808
rect 143040 796 143046 808
rect 145009 799 145067 805
rect 145009 796 145021 799
rect 143040 768 145021 796
rect 143040 756 143046 768
rect 145009 765 145021 768
rect 145055 765 145067 799
rect 145009 759 145067 765
rect 146021 799 146079 805
rect 146021 765 146033 799
rect 146067 796 146079 799
rect 148796 796 148824 836
rect 152734 824 152740 836
rect 152792 824 152798 876
rect 155954 824 155960 876
rect 156012 864 156018 876
rect 166994 864 167000 876
rect 156012 836 167000 864
rect 156012 824 156018 836
rect 166994 824 167000 836
rect 167052 824 167058 876
rect 169018 824 169024 876
rect 169076 864 169082 876
rect 175274 864 175280 876
rect 169076 836 175280 864
rect 169076 824 169082 836
rect 175274 824 175280 836
rect 175332 824 175338 876
rect 175826 824 175832 876
rect 175884 864 175890 876
rect 181806 864 181812 876
rect 175884 836 181812 864
rect 175884 824 175890 836
rect 181806 824 181812 836
rect 181864 824 181870 876
rect 163406 796 163412 808
rect 146067 768 148824 796
rect 148888 768 163412 796
rect 146067 765 146079 768
rect 146021 759 146079 765
rect 135257 731 135315 737
rect 135257 697 135269 731
rect 135303 728 135315 731
rect 142522 728 142528 740
rect 135303 700 142528 728
rect 135303 697 135315 700
rect 135257 691 135315 697
rect 142522 688 142528 700
rect 142580 688 142586 740
rect 143718 688 143724 740
rect 143776 728 143782 740
rect 144638 728 144644 740
rect 143776 700 144644 728
rect 143776 688 143782 700
rect 144638 688 144644 700
rect 144696 688 144702 740
rect 144914 688 144920 740
rect 144972 728 144978 740
rect 148888 728 148916 768
rect 163406 756 163412 768
rect 163464 756 163470 808
rect 163774 756 163780 808
rect 163832 796 163838 808
rect 171134 796 171140 808
rect 163832 768 171140 796
rect 163832 756 163838 768
rect 171134 756 171140 768
rect 171192 756 171198 808
rect 182177 799 182235 805
rect 182177 765 182189 799
rect 182223 796 182235 799
rect 188062 796 188068 808
rect 182223 768 188068 796
rect 182223 765 182235 768
rect 182177 759 182235 765
rect 188062 756 188068 768
rect 188120 756 188126 808
rect 144972 700 148916 728
rect 149793 731 149851 737
rect 144972 688 144978 700
rect 149793 697 149805 731
rect 149839 728 149851 731
rect 164786 728 164792 740
rect 149839 700 164792 728
rect 149839 697 149851 700
rect 149793 691 149851 697
rect 164786 688 164792 700
rect 164844 688 164850 740
rect 165985 731 166043 737
rect 165985 697 165997 731
rect 166031 728 166043 731
rect 169570 728 169576 740
rect 166031 700 169576 728
rect 166031 697 166043 700
rect 165985 691 166043 697
rect 169570 688 169576 700
rect 169628 688 169634 740
rect 155586 660 155592 672
rect 135180 632 155592 660
rect 133233 623 133291 629
rect 155586 620 155592 632
rect 155644 620 155650 672
rect 156046 620 156052 672
rect 156104 660 156110 672
rect 165614 660 165620 672
rect 156104 632 165620 660
rect 156104 620 156110 632
rect 165614 620 165620 632
rect 165672 620 165678 672
rect 166258 620 166264 672
rect 166316 660 166322 672
rect 173894 660 173900 672
rect 166316 632 173900 660
rect 166316 620 166322 632
rect 173894 620 173900 632
rect 173952 620 173958 672
rect 115348 564 129780 592
rect 129829 595 129887 601
rect 115348 552 115354 564
rect 129829 561 129841 595
rect 129875 592 129887 595
rect 140590 592 140596 604
rect 129875 564 140596 592
rect 129875 561 129887 564
rect 129829 555 129887 561
rect 140590 552 140596 564
rect 140648 552 140654 604
rect 140777 595 140835 601
rect 140777 561 140789 595
rect 140823 592 140835 595
rect 143626 592 143632 604
rect 140823 564 143632 592
rect 140823 561 140835 564
rect 140777 555 140835 561
rect 143626 552 143632 564
rect 143684 552 143690 604
rect 143721 595 143779 601
rect 143721 561 143733 595
rect 143767 592 143779 595
rect 149238 592 149244 604
rect 143767 564 149244 592
rect 143767 561 143779 564
rect 143721 555 143779 561
rect 149238 552 149244 564
rect 149296 552 149302 604
rect 151446 552 151452 604
rect 151504 592 151510 604
rect 171318 592 171324 604
rect 151504 564 171324 592
rect 151504 552 151510 564
rect 171318 552 171324 564
rect 171376 552 171382 604
rect 130930 484 130936 536
rect 130988 524 130994 536
rect 156966 524 156972 536
rect 130988 496 156972 524
rect 130988 484 130994 496
rect 156966 484 156972 496
rect 157024 484 157030 536
rect 160646 484 160652 536
rect 160704 524 160710 536
rect 166534 524 166540 536
rect 160704 496 166540 524
rect 160704 484 160710 496
rect 166534 484 166540 496
rect 166592 484 166598 536
rect 166813 527 166871 533
rect 166813 493 166825 527
rect 166859 524 166871 527
rect 167362 524 167368 536
rect 166859 496 167368 524
rect 166859 493 166871 496
rect 166813 487 166871 493
rect 167362 484 167368 496
rect 167420 484 167426 536
rect 128446 416 128452 468
rect 128504 456 128510 468
rect 155402 456 155408 468
rect 128504 428 155408 456
rect 128504 416 128510 428
rect 155402 416 155408 428
rect 155460 416 155466 468
rect 156230 416 156236 468
rect 156288 456 156294 468
rect 161750 456 161756 468
rect 156288 428 161756 456
rect 156288 416 156294 428
rect 161750 416 161756 428
rect 161808 416 161814 468
rect 161845 459 161903 465
rect 161845 425 161857 459
rect 161891 456 161903 459
rect 173526 456 173532 468
rect 161891 428 173532 456
rect 161891 425 161903 428
rect 161845 419 161903 425
rect 173526 416 173532 428
rect 173584 416 173590 468
rect 119890 348 119896 400
rect 119948 388 119954 400
rect 140777 391 140835 397
rect 140777 388 140789 391
rect 119948 360 140789 388
rect 119948 348 119954 360
rect 140777 357 140789 360
rect 140823 357 140835 391
rect 140777 351 140835 357
rect 141881 391 141939 397
rect 141881 357 141893 391
rect 141927 388 141939 391
rect 150802 388 150808 400
rect 141927 360 150808 388
rect 141927 357 141939 360
rect 141881 351 141939 357
rect 150802 348 150808 360
rect 150860 348 150866 400
rect 155034 348 155040 400
rect 155092 388 155098 400
rect 177850 388 177856 400
rect 155092 360 177856 388
rect 155092 348 155098 360
rect 177850 348 177856 360
rect 177908 348 177914 400
rect 129366 280 129372 332
rect 129424 320 129430 332
rect 137557 323 137615 329
rect 137557 320 137569 323
rect 129424 292 137569 320
rect 129424 280 129430 292
rect 137557 289 137569 292
rect 137603 289 137615 323
rect 137557 283 137615 289
rect 137646 280 137652 332
rect 137704 320 137710 332
rect 156506 320 156512 332
rect 137704 292 156512 320
rect 137704 280 137710 292
rect 156506 280 156512 292
rect 156564 280 156570 332
rect 157518 280 157524 332
rect 157576 320 157582 332
rect 157576 292 159220 320
rect 157576 280 157582 292
rect 129642 212 129648 264
rect 129700 252 129706 264
rect 157794 252 157800 264
rect 129700 224 157800 252
rect 129700 212 129706 224
rect 157794 212 157800 224
rect 157852 212 157858 264
rect 130286 144 130292 196
rect 130344 184 130350 196
rect 159082 184 159088 196
rect 130344 156 159088 184
rect 130344 144 130350 156
rect 159082 144 159088 156
rect 159140 144 159146 196
rect 159192 184 159220 292
rect 159266 280 159272 332
rect 159324 320 159330 332
rect 161845 323 161903 329
rect 161845 320 161857 323
rect 159324 292 161857 320
rect 159324 280 159330 292
rect 161845 289 161857 292
rect 161891 289 161903 323
rect 161845 283 161903 289
rect 161937 323 161995 329
rect 161937 289 161949 323
rect 161983 320 161995 323
rect 178310 320 178316 332
rect 161983 292 178316 320
rect 161983 289 161995 292
rect 161937 283 161995 289
rect 178310 280 178316 292
rect 178368 280 178374 332
rect 159542 212 159548 264
rect 159600 252 159606 264
rect 166813 255 166871 261
rect 166813 252 166825 255
rect 159600 224 166825 252
rect 159600 212 159606 224
rect 166813 221 166825 224
rect 166859 221 166871 255
rect 166813 215 166871 221
rect 166902 212 166908 264
rect 166960 252 166966 264
rect 170030 252 170036 264
rect 166960 224 170036 252
rect 166960 212 166966 224
rect 170030 212 170036 224
rect 170088 212 170094 264
rect 160646 184 160652 196
rect 159192 156 160652 184
rect 160646 144 160652 156
rect 160704 144 160710 196
rect 160738 144 160744 196
rect 160796 184 160802 196
rect 179598 184 179604 196
rect 160796 156 179604 184
rect 160796 144 160802 156
rect 179598 144 179604 156
rect 179656 144 179662 196
rect 128998 76 129004 128
rect 129056 116 129062 128
rect 132862 116 132868 128
rect 129056 88 132868 116
rect 129056 76 129062 88
rect 132862 76 132868 88
rect 132920 76 132926 128
rect 133138 76 133144 128
rect 133196 116 133202 128
rect 163038 116 163044 128
rect 133196 88 163044 116
rect 133196 76 133202 88
rect 163038 76 163044 88
rect 163096 76 163102 128
rect 163222 76 163228 128
rect 163280 116 163286 128
rect 168466 116 168472 128
rect 163280 88 168472 116
rect 163280 76 163286 88
rect 168466 76 168472 88
rect 168524 76 168530 128
rect 131114 8 131120 60
rect 131172 48 131178 60
rect 162578 48 162584 60
rect 131172 20 162584 48
rect 131172 8 131178 20
rect 162578 8 162584 20
rect 162636 8 162642 60
rect 162762 8 162768 60
rect 162820 48 162826 60
rect 172146 48 172152 60
rect 162820 20 172152 48
rect 162820 8 162826 20
rect 172146 8 172152 20
rect 172204 8 172210 60
<< via1 >>
rect 147312 10548 147364 10600
rect 124404 10480 124456 10532
rect 133604 10480 133656 10532
rect 82176 10412 82228 10464
rect 132960 10412 133012 10464
rect 119804 10344 119856 10396
rect 128912 10344 128964 10396
rect 97816 10276 97868 10328
rect 145564 10276 145616 10328
rect 119712 10208 119764 10260
rect 128544 10208 128596 10260
rect 130384 10208 130436 10260
rect 140964 10208 141016 10260
rect 145840 10208 145892 10260
rect 169576 10208 169628 10260
rect 75184 10140 75236 10192
rect 142988 10140 143040 10192
rect 159088 10140 159140 10192
rect 169944 10140 169996 10192
rect 171324 10140 171376 10192
rect 185676 10140 185728 10192
rect 95700 10072 95752 10124
rect 121276 10072 121328 10124
rect 129004 10072 129056 10124
rect 144368 10072 144420 10124
rect 149704 10072 149756 10124
rect 195152 10072 195204 10124
rect 97540 10004 97592 10056
rect 105636 10004 105688 10056
rect 106096 10004 106148 10056
rect 121184 10004 121236 10056
rect 125140 10004 125192 10056
rect 136916 10004 136968 10056
rect 104440 9936 104492 9988
rect 131764 9936 131816 9988
rect 135444 9936 135496 9988
rect 141792 10004 141844 10056
rect 151268 10004 151320 10056
rect 181260 10004 181312 10056
rect 182088 10004 182140 10056
rect 187056 10004 187108 10056
rect 140412 9936 140464 9988
rect 77852 9868 77904 9920
rect 86040 9868 86092 9920
rect 94320 9911 94372 9920
rect 94320 9877 94329 9911
rect 94329 9877 94363 9911
rect 94363 9877 94372 9911
rect 94320 9868 94372 9877
rect 96068 9868 96120 9920
rect 99932 9868 99984 9920
rect 107936 9868 107988 9920
rect 140780 9868 140832 9920
rect 156052 9936 156104 9988
rect 159180 9936 159232 9988
rect 165252 9936 165304 9988
rect 177028 9936 177080 9988
rect 166172 9868 166224 9920
rect 166264 9868 166316 9920
rect 181536 9936 181588 9988
rect 182732 9936 182784 9988
rect 198832 9936 198884 9988
rect 179512 9868 179564 9920
rect 183192 9868 183244 9920
rect 191104 9868 191156 9920
rect 198004 9868 198056 9920
rect 4078 9766 4130 9818
rect 44078 9766 44130 9818
rect 84078 9766 84130 9818
rect 124078 9766 124130 9818
rect 164078 9766 164130 9818
rect 1032 9664 1084 9716
rect 85856 9664 85908 9716
rect 134800 9664 134852 9716
rect 136180 9664 136232 9716
rect 139124 9664 139176 9716
rect 152096 9664 152148 9716
rect 204 9528 256 9580
rect 1492 9460 1544 9512
rect 3332 9460 3384 9512
rect 5540 9503 5592 9512
rect 5540 9469 5549 9503
rect 5549 9469 5583 9503
rect 5583 9469 5592 9503
rect 5540 9460 5592 9469
rect 11336 9528 11388 9580
rect 43720 9528 43772 9580
rect 73160 9596 73212 9648
rect 75368 9596 75420 9648
rect 83832 9596 83884 9648
rect 85948 9596 86000 9648
rect 110328 9596 110380 9648
rect 111708 9596 111760 9648
rect 86132 9528 86184 9580
rect 94320 9571 94372 9580
rect 94320 9537 94329 9571
rect 94329 9537 94363 9571
rect 94363 9537 94372 9571
rect 94320 9528 94372 9537
rect 6920 9503 6972 9512
rect 6920 9469 6929 9503
rect 6929 9469 6963 9503
rect 6963 9469 6972 9503
rect 6920 9460 6972 9469
rect 7104 9460 7156 9512
rect 15292 9460 15344 9512
rect 17040 9503 17092 9512
rect 17040 9469 17049 9503
rect 17049 9469 17083 9503
rect 17083 9469 17092 9503
rect 17040 9460 17092 9469
rect 40960 9460 41012 9512
rect 61292 9503 61344 9512
rect 43628 9392 43680 9444
rect 61292 9469 61301 9503
rect 61301 9469 61335 9503
rect 61335 9469 61344 9503
rect 61292 9460 61344 9469
rect 61476 9503 61528 9512
rect 61476 9469 61485 9503
rect 61485 9469 61519 9503
rect 61519 9469 61528 9503
rect 61476 9460 61528 9469
rect 61568 9460 61620 9512
rect 71412 9460 71464 9512
rect 71596 9392 71648 9444
rect 73436 9392 73488 9444
rect 89444 9460 89496 9512
rect 95424 9460 95476 9512
rect 108212 9528 108264 9580
rect 111248 9528 111300 9580
rect 113916 9571 113968 9580
rect 96068 9503 96120 9512
rect 87236 9392 87288 9444
rect 96068 9469 96077 9503
rect 96077 9469 96111 9503
rect 96111 9469 96120 9503
rect 96068 9460 96120 9469
rect 98000 9460 98052 9512
rect 98644 9460 98696 9512
rect 99380 9460 99432 9512
rect 111524 9503 111576 9512
rect 111524 9469 111533 9503
rect 111533 9469 111567 9503
rect 111567 9469 111576 9503
rect 111524 9460 111576 9469
rect 95976 9392 96028 9444
rect 97908 9392 97960 9444
rect 105636 9392 105688 9444
rect 113916 9537 113925 9571
rect 113925 9537 113959 9571
rect 113959 9537 113968 9571
rect 113916 9528 113968 9537
rect 119436 9528 119488 9580
rect 119620 9571 119672 9580
rect 119620 9537 119629 9571
rect 119629 9537 119663 9571
rect 119663 9537 119672 9571
rect 119620 9528 119672 9537
rect 124680 9528 124732 9580
rect 125508 9571 125560 9580
rect 125508 9537 125517 9571
rect 125517 9537 125551 9571
rect 125551 9537 125560 9571
rect 125508 9528 125560 9537
rect 129280 9528 129332 9580
rect 130384 9528 130436 9580
rect 130568 9571 130620 9580
rect 130568 9537 130577 9571
rect 130577 9537 130611 9571
rect 130611 9537 130620 9571
rect 130568 9528 130620 9537
rect 115204 9460 115256 9512
rect 119804 9460 119856 9512
rect 124496 9460 124548 9512
rect 129464 9460 129516 9512
rect 132316 9460 132368 9512
rect 136272 9596 136324 9648
rect 142620 9596 142672 9648
rect 156696 9639 156748 9648
rect 156696 9605 156705 9639
rect 156705 9605 156739 9639
rect 156739 9605 156748 9639
rect 156696 9596 156748 9605
rect 158076 9596 158128 9648
rect 164148 9596 164200 9648
rect 165252 9639 165304 9648
rect 165252 9605 165261 9639
rect 165261 9605 165295 9639
rect 165295 9605 165304 9639
rect 165252 9596 165304 9605
rect 165344 9596 165396 9648
rect 168380 9596 168432 9648
rect 171324 9639 171376 9648
rect 171324 9605 171333 9639
rect 171333 9605 171367 9639
rect 171367 9605 171376 9639
rect 171324 9596 171376 9605
rect 134524 9528 134576 9580
rect 151268 9571 151320 9580
rect 151268 9537 151277 9571
rect 151277 9537 151311 9571
rect 151311 9537 151320 9571
rect 151268 9528 151320 9537
rect 153844 9571 153896 9580
rect 153844 9537 153853 9571
rect 153853 9537 153887 9571
rect 153887 9537 153896 9571
rect 153844 9528 153896 9537
rect 159088 9528 159140 9580
rect 150624 9460 150676 9512
rect 153476 9503 153528 9512
rect 153476 9469 153485 9503
rect 153485 9469 153519 9503
rect 153519 9469 153528 9503
rect 153476 9460 153528 9469
rect 156328 9503 156380 9512
rect 11244 9324 11296 9376
rect 27896 9324 27948 9376
rect 40868 9324 40920 9376
rect 46112 9324 46164 9376
rect 46940 9324 46992 9376
rect 59360 9324 59412 9376
rect 62672 9367 62724 9376
rect 62672 9333 62681 9367
rect 62681 9333 62715 9367
rect 62715 9333 62724 9367
rect 62672 9324 62724 9333
rect 64696 9367 64748 9376
rect 64696 9333 64705 9367
rect 64705 9333 64739 9367
rect 64739 9333 64748 9367
rect 64696 9324 64748 9333
rect 65708 9367 65760 9376
rect 65708 9333 65717 9367
rect 65717 9333 65751 9367
rect 65751 9333 65760 9367
rect 65708 9324 65760 9333
rect 70492 9324 70544 9376
rect 73712 9324 73764 9376
rect 73988 9324 74040 9376
rect 76380 9367 76432 9376
rect 76380 9333 76389 9367
rect 76389 9333 76423 9367
rect 76423 9333 76432 9367
rect 76380 9324 76432 9333
rect 78220 9367 78272 9376
rect 78220 9333 78229 9367
rect 78229 9333 78263 9367
rect 78263 9333 78272 9367
rect 78220 9324 78272 9333
rect 80704 9324 80756 9376
rect 82636 9367 82688 9376
rect 82636 9333 82645 9367
rect 82645 9333 82679 9367
rect 82679 9333 82688 9367
rect 82636 9324 82688 9333
rect 82728 9324 82780 9376
rect 85580 9324 85632 9376
rect 85672 9324 85724 9376
rect 96896 9367 96948 9376
rect 96896 9333 96905 9367
rect 96905 9333 96939 9367
rect 96939 9333 96948 9367
rect 96896 9324 96948 9333
rect 96988 9324 97040 9376
rect 99196 9367 99248 9376
rect 99196 9333 99205 9367
rect 99205 9333 99239 9367
rect 99239 9333 99248 9367
rect 99196 9324 99248 9333
rect 99564 9324 99616 9376
rect 110420 9324 110472 9376
rect 114652 9324 114704 9376
rect 116584 9324 116636 9376
rect 128360 9324 128412 9376
rect 128452 9324 128504 9376
rect 136364 9392 136416 9444
rect 140964 9435 141016 9444
rect 133420 9367 133472 9376
rect 133420 9333 133429 9367
rect 133429 9333 133463 9367
rect 133463 9333 133472 9367
rect 133420 9324 133472 9333
rect 133604 9324 133656 9376
rect 135720 9324 135772 9376
rect 139124 9367 139176 9376
rect 139124 9333 139133 9367
rect 139133 9333 139167 9367
rect 139167 9333 139176 9367
rect 139124 9324 139176 9333
rect 140964 9401 140973 9435
rect 140973 9401 141007 9435
rect 141007 9401 141016 9435
rect 140964 9392 141016 9401
rect 146116 9392 146168 9444
rect 151636 9392 151688 9444
rect 156328 9469 156337 9503
rect 156337 9469 156371 9503
rect 156371 9469 156380 9503
rect 156328 9460 156380 9469
rect 160100 9460 160152 9512
rect 164884 9503 164936 9512
rect 164884 9469 164893 9503
rect 164893 9469 164927 9503
rect 164927 9469 164936 9503
rect 164884 9460 164936 9469
rect 165068 9528 165120 9580
rect 166264 9528 166316 9580
rect 172152 9528 172204 9580
rect 167736 9503 167788 9512
rect 167736 9469 167745 9503
rect 167745 9469 167779 9503
rect 167779 9469 167788 9503
rect 167736 9460 167788 9469
rect 169760 9460 169812 9512
rect 171416 9503 171468 9512
rect 171416 9469 171425 9503
rect 171425 9469 171459 9503
rect 171459 9469 171468 9503
rect 171416 9460 171468 9469
rect 172336 9503 172388 9512
rect 172336 9469 172345 9503
rect 172345 9469 172379 9503
rect 172379 9469 172388 9503
rect 172336 9460 172388 9469
rect 173716 9503 173768 9512
rect 173716 9469 173725 9503
rect 173725 9469 173759 9503
rect 173759 9469 173768 9503
rect 173716 9460 173768 9469
rect 175464 9503 175516 9512
rect 175464 9469 175473 9503
rect 175473 9469 175507 9503
rect 175507 9469 175516 9503
rect 175464 9460 175516 9469
rect 179236 9596 179288 9648
rect 181260 9571 181312 9580
rect 155592 9392 155644 9444
rect 157432 9392 157484 9444
rect 142068 9324 142120 9376
rect 144920 9324 144972 9376
rect 147680 9367 147732 9376
rect 147680 9333 147689 9367
rect 147689 9333 147723 9367
rect 147723 9333 147732 9367
rect 147680 9324 147732 9333
rect 148416 9324 148468 9376
rect 155500 9324 155552 9376
rect 156604 9324 156656 9376
rect 157340 9324 157392 9376
rect 162216 9392 162268 9444
rect 175924 9392 175976 9444
rect 181260 9537 181269 9571
rect 181269 9537 181303 9571
rect 181303 9537 181312 9571
rect 181260 9528 181312 9537
rect 181536 9664 181588 9716
rect 183928 9664 183980 9716
rect 187424 9664 187476 9716
rect 191932 9664 191984 9716
rect 181628 9596 181680 9648
rect 182548 9596 182600 9648
rect 182732 9639 182784 9648
rect 182732 9605 182741 9639
rect 182741 9605 182775 9639
rect 182775 9605 182784 9639
rect 182732 9596 182784 9605
rect 191104 9596 191156 9648
rect 196256 9596 196308 9648
rect 199752 9596 199804 9648
rect 190184 9528 190236 9580
rect 194508 9528 194560 9580
rect 195152 9571 195204 9580
rect 195152 9537 195161 9571
rect 195161 9537 195195 9571
rect 195195 9537 195204 9571
rect 195152 9528 195204 9537
rect 177856 9460 177908 9512
rect 182640 9460 182692 9512
rect 182824 9503 182876 9512
rect 182824 9469 182833 9503
rect 182833 9469 182867 9503
rect 182867 9469 182876 9503
rect 182824 9460 182876 9469
rect 183744 9460 183796 9512
rect 184020 9392 184072 9444
rect 188988 9460 189040 9512
rect 189448 9503 189500 9512
rect 189448 9469 189457 9503
rect 189457 9469 189491 9503
rect 189491 9469 189500 9503
rect 189448 9460 189500 9469
rect 192668 9503 192720 9512
rect 191196 9392 191248 9444
rect 192668 9469 192677 9503
rect 192677 9469 192711 9503
rect 192711 9469 192720 9503
rect 192668 9460 192720 9469
rect 194232 9503 194284 9512
rect 194232 9469 194241 9503
rect 194241 9469 194275 9503
rect 194275 9469 194284 9503
rect 194232 9460 194284 9469
rect 197360 9460 197412 9512
rect 195060 9392 195112 9444
rect 164332 9324 164384 9376
rect 169116 9324 169168 9376
rect 174912 9324 174964 9376
rect 191932 9324 191984 9376
rect 24078 9222 24130 9274
rect 64078 9222 64130 9274
rect 104078 9222 104130 9274
rect 144078 9222 144130 9274
rect 184078 9222 184130 9274
rect 6920 9120 6972 9172
rect 7104 9163 7156 9172
rect 7104 9129 7113 9163
rect 7113 9129 7147 9163
rect 7147 9129 7156 9163
rect 7104 9120 7156 9129
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 61292 9120 61344 9172
rect 64696 9120 64748 9172
rect 74448 9120 74500 9172
rect 4068 9052 4120 9104
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 27068 9052 27120 9104
rect 11244 9027 11296 9036
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 11612 8984 11664 9036
rect 15200 8984 15252 9036
rect 27896 9027 27948 9036
rect 27896 8993 27905 9027
rect 27905 8993 27939 9027
rect 27939 8993 27948 9027
rect 27896 8984 27948 8993
rect 41328 9052 41380 9104
rect 38292 8984 38344 9036
rect 40868 9027 40920 9036
rect 40868 8993 40877 9027
rect 40877 8993 40911 9027
rect 40911 8993 40920 9027
rect 40868 8984 40920 8993
rect 43444 8984 43496 9036
rect 43812 9052 43864 9104
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6828 8916 6880 8968
rect 4528 8848 4580 8900
rect 14372 8916 14424 8968
rect 16764 8916 16816 8968
rect 20444 8916 20496 8968
rect 29276 8916 29328 8968
rect 31116 8916 31168 8968
rect 32128 8959 32180 8968
rect 32128 8925 32137 8959
rect 32137 8925 32171 8959
rect 32171 8925 32180 8959
rect 32128 8916 32180 8925
rect 32220 8916 32272 8968
rect 39120 8916 39172 8968
rect 39396 8916 39448 8968
rect 42708 8916 42760 8968
rect 43720 8959 43772 8968
rect 43720 8925 43729 8959
rect 43729 8925 43763 8959
rect 43763 8925 43772 8959
rect 43720 8916 43772 8925
rect 44180 8916 44232 8968
rect 46940 8916 46992 8968
rect 49056 8984 49108 9036
rect 47584 8916 47636 8968
rect 55864 8916 55916 8968
rect 60464 9027 60516 9036
rect 40224 8848 40276 8900
rect 53104 8848 53156 8900
rect 60464 8993 60473 9027
rect 60473 8993 60507 9027
rect 60507 8993 60516 9027
rect 60464 8984 60516 8993
rect 61200 8984 61252 9036
rect 65708 8984 65760 9036
rect 77208 9052 77260 9104
rect 73712 9027 73764 9036
rect 73712 8993 73721 9027
rect 73721 8993 73755 9027
rect 73755 8993 73764 9027
rect 73712 8984 73764 8993
rect 75276 9027 75328 9036
rect 75276 8993 75285 9027
rect 75285 8993 75319 9027
rect 75319 8993 75328 9027
rect 75276 8984 75328 8993
rect 75460 8984 75512 9036
rect 77852 8984 77904 9036
rect 86960 9120 87012 9172
rect 99288 9120 99340 9172
rect 105636 9163 105688 9172
rect 105636 9129 105645 9163
rect 105645 9129 105679 9163
rect 105679 9129 105688 9163
rect 105636 9120 105688 9129
rect 105728 9120 105780 9172
rect 110788 9120 110840 9172
rect 85488 9052 85540 9104
rect 85948 9027 86000 9036
rect 59544 8916 59596 8968
rect 60556 8959 60608 8968
rect 60556 8925 60565 8959
rect 60565 8925 60599 8959
rect 60599 8925 60608 8959
rect 60556 8916 60608 8925
rect 61108 8916 61160 8968
rect 62580 8916 62632 8968
rect 66076 8916 66128 8968
rect 67824 8916 67876 8968
rect 69940 8916 69992 8968
rect 70308 8959 70360 8968
rect 70308 8925 70317 8959
rect 70317 8925 70351 8959
rect 70351 8925 70360 8959
rect 70308 8916 70360 8925
rect 72240 8916 72292 8968
rect 75184 8959 75236 8968
rect 75184 8925 75193 8959
rect 75193 8925 75227 8959
rect 75227 8925 75236 8959
rect 75184 8916 75236 8925
rect 77392 8959 77444 8968
rect 77392 8925 77401 8959
rect 77401 8925 77435 8959
rect 77435 8925 77444 8959
rect 77392 8916 77444 8925
rect 70952 8848 71004 8900
rect 76840 8848 76892 8900
rect 81532 8916 81584 8968
rect 12256 8780 12308 8832
rect 82820 8780 82872 8832
rect 85948 8993 85957 9027
rect 85957 8993 85991 9027
rect 85991 8993 86000 9027
rect 85948 8984 86000 8993
rect 99196 9052 99248 9104
rect 106924 9052 106976 9104
rect 95148 8984 95200 9036
rect 97080 8984 97132 9036
rect 97908 9027 97960 9036
rect 97908 8993 97917 9027
rect 97917 8993 97951 9027
rect 97951 8993 97960 9027
rect 97908 8984 97960 8993
rect 100852 8984 100904 9036
rect 107936 9027 107988 9036
rect 107936 8993 107945 9027
rect 107945 8993 107979 9027
rect 107979 8993 107988 9027
rect 107936 8984 107988 8993
rect 142068 9120 142120 9172
rect 148324 9120 148376 9172
rect 152096 9163 152148 9172
rect 152096 9129 152105 9163
rect 152105 9129 152139 9163
rect 152139 9129 152148 9163
rect 152096 9120 152148 9129
rect 155776 9120 155828 9172
rect 158812 9120 158864 9172
rect 160100 9163 160152 9172
rect 160100 9129 160109 9163
rect 160109 9129 160143 9163
rect 160143 9129 160152 9163
rect 160100 9120 160152 9129
rect 160284 9120 160336 9172
rect 166632 9120 166684 9172
rect 111248 9027 111300 9036
rect 111248 8993 111257 9027
rect 111257 8993 111291 9027
rect 111291 8993 111300 9027
rect 111248 8984 111300 8993
rect 83556 8916 83608 8968
rect 85856 8959 85908 8968
rect 85856 8925 85865 8959
rect 85865 8925 85899 8959
rect 85899 8925 85908 8959
rect 85856 8916 85908 8925
rect 89260 8959 89312 8968
rect 89260 8925 89269 8959
rect 89269 8925 89303 8959
rect 89303 8925 89312 8959
rect 89260 8916 89312 8925
rect 90364 8959 90416 8968
rect 90364 8925 90373 8959
rect 90373 8925 90407 8959
rect 90407 8925 90416 8959
rect 90364 8916 90416 8925
rect 91836 8959 91888 8968
rect 91836 8925 91845 8959
rect 91845 8925 91879 8959
rect 91879 8925 91888 8959
rect 91836 8916 91888 8925
rect 95424 8916 95476 8968
rect 97816 8916 97868 8968
rect 98092 8959 98144 8968
rect 98092 8925 98101 8959
rect 98101 8925 98135 8959
rect 98135 8925 98144 8959
rect 98092 8916 98144 8925
rect 99104 8916 99156 8968
rect 99932 8916 99984 8968
rect 102048 8959 102100 8968
rect 102048 8925 102057 8959
rect 102057 8925 102091 8959
rect 102091 8925 102100 8959
rect 102048 8916 102100 8925
rect 103060 8959 103112 8968
rect 103060 8925 103069 8959
rect 103069 8925 103103 8959
rect 103103 8925 103112 8959
rect 103060 8916 103112 8925
rect 109224 8916 109276 8968
rect 119712 9027 119764 9036
rect 119712 8993 119721 9027
rect 119721 8993 119755 9027
rect 119755 8993 119764 9027
rect 119712 8984 119764 8993
rect 122196 8984 122248 9036
rect 124404 9027 124456 9036
rect 124404 8993 124413 9027
rect 124413 8993 124447 9027
rect 124447 8993 124456 9027
rect 124404 8984 124456 8993
rect 128084 8984 128136 9036
rect 128452 9027 128504 9036
rect 128452 8993 128461 9027
rect 128461 8993 128495 9027
rect 128495 8993 128504 9027
rect 128452 8984 128504 8993
rect 129556 9027 129608 9036
rect 129556 8993 129565 9027
rect 129565 8993 129599 9027
rect 129599 8993 129608 9027
rect 129556 8984 129608 8993
rect 130384 8984 130436 9036
rect 134524 9027 134576 9036
rect 120356 8916 120408 8968
rect 117228 8848 117280 8900
rect 119712 8848 119764 8900
rect 130476 8916 130528 8968
rect 130844 8959 130896 8968
rect 130844 8925 130853 8959
rect 130853 8925 130887 8959
rect 130887 8925 130896 8959
rect 130844 8916 130896 8925
rect 125876 8891 125928 8900
rect 125876 8857 125885 8891
rect 125885 8857 125919 8891
rect 125919 8857 125928 8891
rect 125876 8848 125928 8857
rect 129372 8848 129424 8900
rect 88616 8780 88668 8832
rect 97448 8780 97500 8832
rect 102600 8780 102652 8832
rect 107292 8780 107344 8832
rect 111156 8780 111208 8832
rect 118424 8780 118476 8832
rect 125232 8780 125284 8832
rect 127808 8780 127860 8832
rect 133328 8916 133380 8968
rect 134524 8993 134533 9027
rect 134533 8993 134567 9027
rect 134567 8993 134576 9027
rect 134524 8984 134576 8993
rect 135076 8984 135128 9036
rect 136916 9027 136968 9036
rect 136916 8993 136925 9027
rect 136925 8993 136959 9027
rect 136959 8993 136968 9027
rect 136916 8984 136968 8993
rect 138388 8984 138440 9036
rect 147680 9052 147732 9104
rect 150716 9052 150768 9104
rect 162124 9052 162176 9104
rect 137836 8916 137888 8968
rect 145472 9027 145524 9036
rect 145472 8993 145481 9027
rect 145481 8993 145515 9027
rect 145515 8993 145524 9027
rect 145472 8984 145524 8993
rect 141148 8959 141200 8968
rect 141148 8925 141157 8959
rect 141157 8925 141191 8959
rect 141191 8925 141200 8959
rect 141148 8916 141200 8925
rect 142160 8959 142212 8968
rect 142160 8925 142169 8959
rect 142169 8925 142203 8959
rect 142203 8925 142212 8959
rect 142160 8916 142212 8925
rect 144736 8916 144788 8968
rect 150440 8984 150492 9036
rect 156696 9027 156748 9036
rect 156696 8993 156705 9027
rect 156705 8993 156739 9027
rect 156739 8993 156748 9027
rect 156696 8984 156748 8993
rect 156880 8984 156932 9036
rect 160192 8984 160244 9036
rect 165620 9052 165672 9104
rect 166448 9052 166500 9104
rect 170956 9052 171008 9104
rect 164332 8984 164384 9036
rect 169024 9027 169076 9036
rect 169024 8993 169033 9027
rect 169033 8993 169067 9027
rect 169067 8993 169076 9027
rect 169024 8984 169076 8993
rect 169944 9027 169996 9036
rect 169944 8993 169953 9027
rect 169953 8993 169987 9027
rect 169987 8993 169996 9027
rect 169944 8984 169996 8993
rect 171232 9027 171284 9036
rect 171232 8993 171241 9027
rect 171241 8993 171275 9027
rect 171275 8993 171284 9027
rect 171232 8984 171284 8993
rect 145840 8959 145892 8968
rect 145840 8925 145849 8959
rect 145849 8925 145883 8959
rect 145883 8925 145892 8959
rect 145840 8916 145892 8925
rect 151084 8959 151136 8968
rect 151084 8925 151093 8959
rect 151093 8925 151127 8959
rect 151127 8925 151136 8959
rect 151084 8916 151136 8925
rect 152832 8916 152884 8968
rect 154488 8959 154540 8968
rect 154488 8925 154497 8959
rect 154497 8925 154531 8959
rect 154531 8925 154540 8959
rect 154488 8916 154540 8925
rect 156236 8916 156288 8968
rect 157984 8959 158036 8968
rect 157984 8925 157993 8959
rect 157993 8925 158027 8959
rect 158027 8925 158036 8959
rect 157984 8916 158036 8925
rect 160008 8916 160060 8968
rect 161940 8959 161992 8968
rect 161940 8925 161949 8959
rect 161949 8925 161983 8959
rect 161983 8925 161992 8959
rect 161940 8916 161992 8925
rect 140228 8891 140280 8900
rect 132224 8780 132276 8832
rect 139124 8780 139176 8832
rect 140228 8857 140237 8891
rect 140237 8857 140271 8891
rect 140271 8857 140280 8891
rect 140228 8848 140280 8857
rect 148232 8891 148284 8900
rect 148232 8857 148241 8891
rect 148241 8857 148275 8891
rect 148275 8857 148284 8891
rect 148232 8848 148284 8857
rect 164424 8891 164476 8900
rect 141240 8780 141292 8832
rect 157156 8780 157208 8832
rect 160468 8780 160520 8832
rect 164424 8857 164433 8891
rect 164433 8857 164467 8891
rect 164467 8857 164476 8891
rect 164424 8848 164476 8857
rect 164792 8848 164844 8900
rect 169208 8916 169260 8968
rect 179512 9120 179564 9172
rect 184480 9120 184532 9172
rect 171508 9052 171560 9104
rect 192116 9120 192168 9172
rect 197360 9163 197412 9172
rect 197360 9129 197369 9163
rect 197369 9129 197403 9163
rect 197403 9129 197412 9163
rect 197360 9120 197412 9129
rect 187884 9052 187936 9104
rect 198464 9052 198516 9104
rect 174912 9027 174964 9036
rect 174912 8993 174921 9027
rect 174921 8993 174955 9027
rect 174955 8993 174964 9027
rect 174912 8984 174964 8993
rect 173716 8916 173768 8968
rect 178040 8959 178092 8968
rect 178040 8925 178049 8959
rect 178049 8925 178083 8959
rect 178083 8925 178092 8959
rect 178040 8916 178092 8925
rect 172520 8848 172572 8900
rect 181628 8984 181680 9036
rect 181996 9027 182048 9036
rect 181996 8993 182005 9027
rect 182005 8993 182039 9027
rect 182039 8993 182048 9027
rect 181996 8984 182048 8993
rect 182640 8984 182692 9036
rect 184572 8984 184624 9036
rect 186228 9027 186280 9036
rect 186228 8993 186237 9027
rect 186237 8993 186271 9027
rect 186271 8993 186280 9027
rect 186228 8984 186280 8993
rect 189356 8984 189408 9036
rect 191932 9027 191984 9036
rect 191932 8993 191941 9027
rect 191941 8993 191975 9027
rect 191975 8993 191984 9027
rect 191932 8984 191984 8993
rect 196440 9027 196492 9036
rect 184848 8959 184900 8968
rect 184848 8925 184857 8959
rect 184857 8925 184891 8959
rect 184891 8925 184900 8959
rect 184848 8916 184900 8925
rect 184940 8916 184992 8968
rect 187516 8916 187568 8968
rect 191472 8916 191524 8968
rect 192300 8916 192352 8968
rect 182088 8891 182140 8900
rect 182088 8857 182097 8891
rect 182097 8857 182131 8891
rect 182131 8857 182140 8891
rect 182088 8848 182140 8857
rect 173164 8780 173216 8832
rect 174268 8780 174320 8832
rect 176752 8780 176804 8832
rect 176844 8780 176896 8832
rect 183560 8848 183612 8900
rect 189724 8848 189776 8900
rect 190736 8848 190788 8900
rect 196440 8993 196449 9027
rect 196449 8993 196483 9027
rect 196483 8993 196492 9027
rect 196440 8984 196492 8993
rect 197268 9027 197320 9036
rect 197268 8993 197277 9027
rect 197277 8993 197311 9027
rect 197311 8993 197320 9027
rect 197268 8984 197320 8993
rect 194876 8959 194928 8968
rect 194876 8925 194885 8959
rect 194885 8925 194919 8959
rect 194919 8925 194928 8959
rect 194876 8916 194928 8925
rect 195336 8916 195388 8968
rect 182824 8780 182876 8832
rect 197360 8780 197412 8832
rect 4078 8678 4130 8730
rect 44078 8678 44130 8730
rect 84078 8678 84130 8730
rect 124078 8678 124130 8730
rect 164078 8678 164130 8730
rect 48504 8576 48556 8628
rect 11520 8508 11572 8560
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 4988 8440 5040 8492
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 19800 8508 19852 8560
rect 16764 8483 16816 8492
rect 16764 8449 16773 8483
rect 16773 8449 16807 8483
rect 16807 8449 16816 8483
rect 16764 8440 16816 8449
rect 20444 8483 20496 8492
rect 20444 8449 20453 8483
rect 20453 8449 20487 8483
rect 20487 8449 20496 8483
rect 20444 8440 20496 8449
rect 28080 8508 28132 8560
rect 31576 8508 31628 8560
rect 46388 8508 46440 8560
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 32220 8440 32272 8492
rect 33232 8483 33284 8492
rect 33232 8449 33241 8483
rect 33241 8449 33275 8483
rect 33275 8449 33284 8483
rect 33232 8440 33284 8449
rect 34152 8440 34204 8492
rect 39120 8483 39172 8492
rect 39120 8449 39129 8483
rect 39129 8449 39163 8483
rect 39163 8449 39172 8483
rect 39120 8440 39172 8449
rect 40960 8483 41012 8492
rect 40960 8449 40969 8483
rect 40969 8449 41003 8483
rect 41003 8449 41012 8483
rect 40960 8440 41012 8449
rect 41420 8440 41472 8492
rect 43720 8440 43772 8492
rect 47584 8483 47636 8492
rect 47584 8449 47593 8483
rect 47593 8449 47627 8483
rect 47627 8449 47636 8483
rect 47584 8440 47636 8449
rect 77392 8576 77444 8628
rect 82268 8576 82320 8628
rect 82820 8576 82872 8628
rect 83924 8576 83976 8628
rect 91100 8576 91152 8628
rect 96712 8576 96764 8628
rect 99564 8576 99616 8628
rect 60464 8508 60516 8560
rect 59544 8483 59596 8492
rect 59544 8449 59553 8483
rect 59553 8449 59587 8483
rect 59587 8449 59596 8483
rect 59544 8440 59596 8449
rect 60832 8483 60884 8492
rect 60832 8449 60841 8483
rect 60841 8449 60875 8483
rect 60875 8449 60884 8483
rect 60832 8440 60884 8449
rect 66076 8483 66128 8492
rect 66076 8449 66085 8483
rect 66085 8449 66119 8483
rect 66119 8449 66128 8483
rect 66076 8440 66128 8449
rect 67088 8483 67140 8492
rect 67088 8449 67097 8483
rect 67097 8449 67131 8483
rect 67131 8449 67140 8483
rect 67088 8440 67140 8449
rect 75828 8508 75880 8560
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 5724 8372 5776 8424
rect 11428 8372 11480 8424
rect 18972 8372 19024 8424
rect 24952 8415 25004 8424
rect 24952 8381 24961 8415
rect 24961 8381 24995 8415
rect 24995 8381 25004 8415
rect 24952 8372 25004 8381
rect 26056 8415 26108 8424
rect 26056 8381 26065 8415
rect 26065 8381 26099 8415
rect 26099 8381 26108 8415
rect 26056 8372 26108 8381
rect 29092 8372 29144 8424
rect 33048 8415 33100 8424
rect 33048 8381 33057 8415
rect 33057 8381 33091 8415
rect 33091 8381 33100 8415
rect 33048 8372 33100 8381
rect 37556 8372 37608 8424
rect 41972 8415 42024 8424
rect 7380 8304 7432 8356
rect 11520 8304 11572 8356
rect 35992 8304 36044 8356
rect 41972 8381 41981 8415
rect 41981 8381 42015 8415
rect 42015 8381 42024 8415
rect 41972 8372 42024 8381
rect 43536 8415 43588 8424
rect 43536 8381 43545 8415
rect 43545 8381 43579 8415
rect 43579 8381 43588 8415
rect 43536 8372 43588 8381
rect 46480 8372 46532 8424
rect 52092 8372 52144 8424
rect 54668 8415 54720 8424
rect 48964 8304 49016 8356
rect 54116 8304 54168 8356
rect 54668 8381 54677 8415
rect 54677 8381 54711 8415
rect 54711 8381 54720 8415
rect 54668 8372 54720 8381
rect 59636 8372 59688 8424
rect 63684 8372 63736 8424
rect 70952 8415 71004 8424
rect 70952 8381 70961 8415
rect 70961 8381 70995 8415
rect 70995 8381 71004 8415
rect 70952 8372 71004 8381
rect 71320 8415 71372 8424
rect 71320 8381 71329 8415
rect 71329 8381 71363 8415
rect 71363 8381 71372 8415
rect 71320 8372 71372 8381
rect 71596 8372 71648 8424
rect 73068 8372 73120 8424
rect 75092 8440 75144 8492
rect 80244 8508 80296 8560
rect 82176 8551 82228 8560
rect 82176 8517 82185 8551
rect 82185 8517 82219 8551
rect 82219 8517 82228 8551
rect 82176 8508 82228 8517
rect 80704 8483 80756 8492
rect 80704 8449 80713 8483
rect 80713 8449 80747 8483
rect 80747 8449 80756 8483
rect 80704 8440 80756 8449
rect 74448 8415 74500 8424
rect 74448 8381 74457 8415
rect 74457 8381 74491 8415
rect 74491 8381 74500 8415
rect 74448 8372 74500 8381
rect 69020 8347 69072 8356
rect 69020 8313 69029 8347
rect 69029 8313 69063 8347
rect 69063 8313 69072 8347
rect 69020 8304 69072 8313
rect 75368 8372 75420 8424
rect 76840 8415 76892 8424
rect 76840 8381 76849 8415
rect 76849 8381 76883 8415
rect 76883 8381 76892 8415
rect 76840 8372 76892 8381
rect 82912 8440 82964 8492
rect 83556 8483 83608 8492
rect 83556 8449 83565 8483
rect 83565 8449 83599 8483
rect 83599 8449 83608 8483
rect 83556 8440 83608 8449
rect 86960 8440 87012 8492
rect 85672 8415 85724 8424
rect 85672 8381 85681 8415
rect 85681 8381 85715 8415
rect 85715 8381 85724 8415
rect 85672 8372 85724 8381
rect 85948 8372 86000 8424
rect 87236 8415 87288 8424
rect 11152 8236 11204 8288
rect 27344 8279 27396 8288
rect 27344 8245 27353 8279
rect 27353 8245 27387 8279
rect 27387 8245 27396 8279
rect 27344 8236 27396 8245
rect 34888 8279 34940 8288
rect 34888 8245 34897 8279
rect 34897 8245 34931 8279
rect 34931 8245 34940 8279
rect 34888 8236 34940 8245
rect 44364 8279 44416 8288
rect 44364 8245 44373 8279
rect 44373 8245 44407 8279
rect 44407 8245 44416 8279
rect 44364 8236 44416 8245
rect 58532 8279 58584 8288
rect 58532 8245 58541 8279
rect 58541 8245 58575 8279
rect 58575 8245 58584 8279
rect 58532 8236 58584 8245
rect 63960 8279 64012 8288
rect 63960 8245 63969 8279
rect 63969 8245 64003 8279
rect 64003 8245 64012 8279
rect 63960 8236 64012 8245
rect 64972 8279 65024 8288
rect 64972 8245 64981 8279
rect 64981 8245 65015 8279
rect 65015 8245 65024 8279
rect 64972 8236 65024 8245
rect 78404 8304 78456 8356
rect 84384 8304 84436 8356
rect 87236 8381 87245 8415
rect 87245 8381 87279 8415
rect 87279 8381 87288 8415
rect 87236 8372 87288 8381
rect 92388 8508 92440 8560
rect 88340 8372 88392 8424
rect 88892 8415 88944 8424
rect 88892 8381 88901 8415
rect 88901 8381 88935 8415
rect 88935 8381 88944 8415
rect 88892 8372 88944 8381
rect 93400 8440 93452 8492
rect 93676 8483 93728 8492
rect 93676 8449 93685 8483
rect 93685 8449 93719 8483
rect 93719 8449 93728 8483
rect 93676 8440 93728 8449
rect 98552 8508 98604 8560
rect 103520 8576 103572 8628
rect 108856 8576 108908 8628
rect 105268 8508 105320 8560
rect 109132 8508 109184 8560
rect 93768 8415 93820 8424
rect 93768 8381 93777 8415
rect 93777 8381 93811 8415
rect 93811 8381 93820 8415
rect 93768 8372 93820 8381
rect 97264 8440 97316 8492
rect 102048 8440 102100 8492
rect 96620 8415 96672 8424
rect 90824 8304 90876 8356
rect 96620 8381 96629 8415
rect 96629 8381 96663 8415
rect 96663 8381 96672 8415
rect 96620 8372 96672 8381
rect 97080 8372 97132 8424
rect 97540 8372 97592 8424
rect 99104 8415 99156 8424
rect 99104 8381 99113 8415
rect 99113 8381 99147 8415
rect 99147 8381 99156 8415
rect 99104 8372 99156 8381
rect 104532 8372 104584 8424
rect 105728 8372 105780 8424
rect 106096 8415 106148 8424
rect 106096 8381 106105 8415
rect 106105 8381 106139 8415
rect 106139 8381 106148 8415
rect 106096 8372 106148 8381
rect 98000 8304 98052 8356
rect 80980 8236 81032 8288
rect 84660 8236 84712 8288
rect 85672 8236 85724 8288
rect 90272 8236 90324 8288
rect 91376 8236 91428 8288
rect 99472 8304 99524 8356
rect 99288 8236 99340 8288
rect 102232 8279 102284 8288
rect 102232 8245 102241 8279
rect 102241 8245 102275 8279
rect 102275 8245 102284 8279
rect 102232 8236 102284 8245
rect 108764 8440 108816 8492
rect 109224 8440 109276 8492
rect 109960 8440 110012 8492
rect 110144 8415 110196 8424
rect 109684 8304 109736 8356
rect 110144 8381 110153 8415
rect 110153 8381 110187 8415
rect 110187 8381 110196 8415
rect 110144 8372 110196 8381
rect 111708 8415 111760 8424
rect 111708 8381 111717 8415
rect 111717 8381 111751 8415
rect 111751 8381 111760 8415
rect 111708 8372 111760 8381
rect 111892 8372 111944 8424
rect 129004 8508 129056 8560
rect 114652 8483 114704 8492
rect 114652 8449 114661 8483
rect 114661 8449 114695 8483
rect 114695 8449 114704 8483
rect 114652 8440 114704 8449
rect 121092 8440 121144 8492
rect 124588 8440 124640 8492
rect 125140 8483 125192 8492
rect 125140 8449 125149 8483
rect 125149 8449 125183 8483
rect 125183 8449 125192 8483
rect 125140 8440 125192 8449
rect 126612 8483 126664 8492
rect 126612 8449 126621 8483
rect 126621 8449 126655 8483
rect 126655 8449 126664 8483
rect 126612 8440 126664 8449
rect 127808 8483 127860 8492
rect 127808 8449 127817 8483
rect 127817 8449 127851 8483
rect 127851 8449 127860 8483
rect 127808 8440 127860 8449
rect 136364 8576 136416 8628
rect 138204 8576 138256 8628
rect 144828 8576 144880 8628
rect 151084 8576 151136 8628
rect 159824 8576 159876 8628
rect 159916 8576 159968 8628
rect 164332 8576 164384 8628
rect 164424 8576 164476 8628
rect 175740 8576 175792 8628
rect 176200 8576 176252 8628
rect 178960 8576 179012 8628
rect 131304 8508 131356 8560
rect 132224 8440 132276 8492
rect 132408 8483 132460 8492
rect 132408 8449 132417 8483
rect 132417 8449 132451 8483
rect 132451 8449 132460 8483
rect 132408 8440 132460 8449
rect 135720 8508 135772 8560
rect 135168 8440 135220 8492
rect 135536 8440 135588 8492
rect 136088 8440 136140 8492
rect 137928 8483 137980 8492
rect 137928 8449 137937 8483
rect 137937 8449 137971 8483
rect 137971 8449 137980 8483
rect 137928 8440 137980 8449
rect 121460 8372 121512 8424
rect 126704 8415 126756 8424
rect 126704 8381 126713 8415
rect 126713 8381 126747 8415
rect 126747 8381 126756 8415
rect 126704 8372 126756 8381
rect 129648 8372 129700 8424
rect 132132 8415 132184 8424
rect 132132 8381 132141 8415
rect 132141 8381 132175 8415
rect 132175 8381 132184 8415
rect 132132 8372 132184 8381
rect 132960 8372 133012 8424
rect 135996 8372 136048 8424
rect 142160 8508 142212 8560
rect 146116 8551 146168 8560
rect 146116 8517 146125 8551
rect 146125 8517 146159 8551
rect 146159 8517 146168 8551
rect 146116 8508 146168 8517
rect 159548 8508 159600 8560
rect 140412 8483 140464 8492
rect 139124 8372 139176 8424
rect 140412 8449 140421 8483
rect 140421 8449 140455 8483
rect 140455 8449 140464 8483
rect 140412 8440 140464 8449
rect 140780 8440 140832 8492
rect 144920 8440 144972 8492
rect 148416 8440 148468 8492
rect 148692 8483 148744 8492
rect 148692 8449 148701 8483
rect 148701 8449 148735 8483
rect 148735 8449 148744 8483
rect 148692 8440 148744 8449
rect 149704 8440 149756 8492
rect 150716 8440 150768 8492
rect 151636 8483 151688 8492
rect 151636 8449 151645 8483
rect 151645 8449 151679 8483
rect 151679 8449 151688 8483
rect 151636 8440 151688 8449
rect 152832 8483 152884 8492
rect 152832 8449 152841 8483
rect 152841 8449 152875 8483
rect 152875 8449 152884 8483
rect 152832 8440 152884 8449
rect 156236 8483 156288 8492
rect 156236 8449 156245 8483
rect 156245 8449 156279 8483
rect 156279 8449 156288 8483
rect 156236 8440 156288 8449
rect 146208 8415 146260 8424
rect 146208 8381 146217 8415
rect 146217 8381 146251 8415
rect 146251 8381 146260 8415
rect 146208 8372 146260 8381
rect 153844 8415 153896 8424
rect 112168 8304 112220 8356
rect 118700 8304 118752 8356
rect 120264 8347 120316 8356
rect 120264 8313 120273 8347
rect 120273 8313 120307 8347
rect 120307 8313 120316 8347
rect 120264 8304 120316 8313
rect 123300 8304 123352 8356
rect 126152 8304 126204 8356
rect 127900 8304 127952 8356
rect 130844 8304 130896 8356
rect 112812 8236 112864 8288
rect 113456 8279 113508 8288
rect 113456 8245 113465 8279
rect 113465 8245 113499 8279
rect 113499 8245 113508 8279
rect 113456 8236 113508 8245
rect 119988 8236 120040 8288
rect 133788 8236 133840 8288
rect 133880 8236 133932 8288
rect 140780 8236 140832 8288
rect 145564 8304 145616 8356
rect 153844 8381 153853 8415
rect 153853 8381 153887 8415
rect 153887 8381 153896 8415
rect 153844 8372 153896 8381
rect 155408 8415 155460 8424
rect 155408 8381 155417 8415
rect 155417 8381 155451 8415
rect 155451 8381 155460 8415
rect 155408 8372 155460 8381
rect 156144 8372 156196 8424
rect 159916 8440 159968 8492
rect 160008 8440 160060 8492
rect 170036 8508 170088 8560
rect 165344 8440 165396 8492
rect 166816 8440 166868 8492
rect 162584 8415 162636 8424
rect 154028 8304 154080 8356
rect 162584 8381 162593 8415
rect 162593 8381 162627 8415
rect 162627 8381 162636 8415
rect 162584 8372 162636 8381
rect 164240 8372 164292 8424
rect 168472 8483 168524 8492
rect 167184 8372 167236 8424
rect 159548 8304 159600 8356
rect 166540 8304 166592 8356
rect 168472 8449 168481 8483
rect 168481 8449 168515 8483
rect 168515 8449 168524 8483
rect 168472 8440 168524 8449
rect 171508 8508 171560 8560
rect 176844 8508 176896 8560
rect 170772 8372 170824 8424
rect 171784 8415 171836 8424
rect 171784 8381 171793 8415
rect 171793 8381 171827 8415
rect 171827 8381 171836 8415
rect 171784 8372 171836 8381
rect 176384 8415 176436 8424
rect 176384 8381 176393 8415
rect 176393 8381 176427 8415
rect 176427 8381 176436 8415
rect 176384 8372 176436 8381
rect 176568 8372 176620 8424
rect 171048 8304 171100 8356
rect 159640 8236 159692 8288
rect 160652 8236 160704 8288
rect 163964 8236 164016 8288
rect 164516 8279 164568 8288
rect 164516 8245 164525 8279
rect 164525 8245 164559 8279
rect 164559 8245 164568 8279
rect 164516 8236 164568 8245
rect 164608 8236 164660 8288
rect 167092 8236 167144 8288
rect 171140 8236 171192 8288
rect 176476 8304 176528 8356
rect 184664 8576 184716 8628
rect 184940 8508 184992 8560
rect 187884 8551 187936 8560
rect 187884 8517 187893 8551
rect 187893 8517 187927 8551
rect 187927 8517 187936 8551
rect 187884 8508 187936 8517
rect 181444 8415 181496 8424
rect 181444 8381 181453 8415
rect 181453 8381 181487 8415
rect 181487 8381 181496 8415
rect 181444 8372 181496 8381
rect 180984 8304 181036 8356
rect 183836 8440 183888 8492
rect 183928 8483 183980 8492
rect 183928 8449 183937 8483
rect 183937 8449 183971 8483
rect 183971 8449 183980 8483
rect 183928 8440 183980 8449
rect 184112 8440 184164 8492
rect 184756 8440 184808 8492
rect 183008 8372 183060 8424
rect 185492 8415 185544 8424
rect 185492 8381 185501 8415
rect 185501 8381 185535 8415
rect 185535 8381 185544 8415
rect 185492 8372 185544 8381
rect 188436 8440 188488 8492
rect 188068 8372 188120 8424
rect 188896 8304 188948 8356
rect 191196 8576 191248 8628
rect 194232 8576 194284 8628
rect 191012 8508 191064 8560
rect 190644 8372 190696 8424
rect 196256 8508 196308 8560
rect 192116 8440 192168 8492
rect 194968 8483 195020 8492
rect 194968 8449 194977 8483
rect 194977 8449 195011 8483
rect 195011 8449 195020 8483
rect 194968 8440 195020 8449
rect 193864 8372 193916 8424
rect 197544 8440 197596 8492
rect 173900 8236 173952 8288
rect 177488 8236 177540 8288
rect 179512 8236 179564 8288
rect 190552 8236 190604 8288
rect 194508 8236 194560 8288
rect 24078 8134 24130 8186
rect 64078 8134 64130 8186
rect 104078 8134 104130 8186
rect 144078 8134 144130 8186
rect 184078 8134 184130 8186
rect 7380 8075 7432 8084
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 24952 8032 25004 8084
rect 37556 8032 37608 8084
rect 41972 8032 42024 8084
rect 54668 8032 54720 8084
rect 55864 8075 55916 8084
rect 55864 8041 55873 8075
rect 55873 8041 55907 8075
rect 55907 8041 55916 8075
rect 55864 8032 55916 8041
rect 75276 8032 75328 8084
rect 81256 8032 81308 8084
rect 83096 8032 83148 8084
rect 29552 7964 29604 8016
rect 6092 7939 6144 7948
rect 6092 7905 6101 7939
rect 6101 7905 6135 7939
rect 6135 7905 6144 7939
rect 6092 7896 6144 7905
rect 11520 7896 11572 7948
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 16856 7896 16908 7948
rect 27344 7896 27396 7948
rect 32128 7939 32180 7948
rect 4344 7828 4396 7880
rect 3332 7760 3384 7812
rect 5356 7828 5408 7880
rect 7472 7828 7524 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 7288 7760 7340 7812
rect 12440 7828 12492 7880
rect 14832 7828 14884 7880
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 16948 7871 17000 7880
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 15844 7760 15896 7812
rect 20444 7828 20496 7880
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 23572 7828 23624 7880
rect 24860 7871 24912 7880
rect 24860 7837 24869 7871
rect 24869 7837 24903 7871
rect 24903 7837 24912 7871
rect 24860 7828 24912 7837
rect 25872 7828 25924 7880
rect 25136 7760 25188 7812
rect 32128 7905 32137 7939
rect 32137 7905 32171 7939
rect 32171 7905 32180 7939
rect 32128 7896 32180 7905
rect 32588 7964 32640 8016
rect 34888 7896 34940 7948
rect 47308 7964 47360 8016
rect 44364 7896 44416 7948
rect 44456 7896 44508 7948
rect 47400 7939 47452 7948
rect 47400 7905 47409 7939
rect 47409 7905 47443 7939
rect 47443 7905 47452 7939
rect 47400 7896 47452 7905
rect 58532 7939 58584 7948
rect 58532 7905 58541 7939
rect 58541 7905 58575 7939
rect 58575 7905 58584 7939
rect 58532 7896 58584 7905
rect 60740 7964 60792 8016
rect 61108 7896 61160 7948
rect 61292 7939 61344 7948
rect 61292 7905 61301 7939
rect 61301 7905 61335 7939
rect 61335 7905 61344 7939
rect 61292 7896 61344 7905
rect 63960 7964 64012 8016
rect 64972 7964 65024 8016
rect 67272 7964 67324 8016
rect 67824 7939 67876 7948
rect 29460 7828 29512 7880
rect 31852 7828 31904 7880
rect 30288 7760 30340 7812
rect 34980 7828 35032 7880
rect 41880 7828 41932 7880
rect 38936 7760 38988 7812
rect 41512 7692 41564 7744
rect 49240 7828 49292 7880
rect 51724 7871 51776 7880
rect 51724 7837 51733 7871
rect 51733 7837 51767 7871
rect 51767 7837 51776 7871
rect 51724 7828 51776 7837
rect 52552 7828 52604 7880
rect 51172 7760 51224 7812
rect 63040 7828 63092 7880
rect 62120 7760 62172 7812
rect 64512 7871 64564 7880
rect 64512 7837 64521 7871
rect 64521 7837 64555 7871
rect 64555 7837 64564 7871
rect 64512 7828 64564 7837
rect 63500 7760 63552 7812
rect 67824 7905 67833 7939
rect 67833 7905 67867 7939
rect 67867 7905 67876 7939
rect 67824 7896 67876 7905
rect 71780 7964 71832 8016
rect 71412 7939 71464 7948
rect 71412 7905 71421 7939
rect 71421 7905 71455 7939
rect 71455 7905 71464 7939
rect 71412 7896 71464 7905
rect 73436 7939 73488 7948
rect 64788 7828 64840 7880
rect 67916 7871 67968 7880
rect 67916 7837 67925 7871
rect 67925 7837 67959 7871
rect 67959 7837 67968 7871
rect 67916 7828 67968 7837
rect 68836 7828 68888 7880
rect 70124 7871 70176 7880
rect 70124 7837 70133 7871
rect 70133 7837 70167 7871
rect 70167 7837 70176 7871
rect 70124 7828 70176 7837
rect 71964 7828 72016 7880
rect 73436 7905 73445 7939
rect 73445 7905 73479 7939
rect 73479 7905 73488 7939
rect 73436 7896 73488 7905
rect 75276 7939 75328 7948
rect 75276 7905 75285 7939
rect 75285 7905 75319 7939
rect 75319 7905 75328 7939
rect 75276 7896 75328 7905
rect 78220 7939 78272 7948
rect 73528 7871 73580 7880
rect 73528 7837 73537 7871
rect 73537 7837 73571 7871
rect 73571 7837 73580 7871
rect 73528 7828 73580 7837
rect 75828 7828 75880 7880
rect 77024 7871 77076 7880
rect 77024 7837 77033 7871
rect 77033 7837 77067 7871
rect 77067 7837 77076 7871
rect 77024 7828 77076 7837
rect 75552 7760 75604 7812
rect 58256 7692 58308 7744
rect 78220 7905 78229 7939
rect 78229 7905 78263 7939
rect 78263 7905 78272 7939
rect 78220 7896 78272 7905
rect 80336 7964 80388 8016
rect 82728 7964 82780 8016
rect 80980 7939 81032 7948
rect 80980 7905 80989 7939
rect 80989 7905 81023 7939
rect 81023 7905 81032 7939
rect 80980 7896 81032 7905
rect 85488 7964 85540 8016
rect 83004 7939 83056 7948
rect 83004 7905 83013 7939
rect 83013 7905 83047 7939
rect 83047 7905 83056 7939
rect 83004 7896 83056 7905
rect 78496 7828 78548 7880
rect 80612 7871 80664 7880
rect 80612 7837 80621 7871
rect 80621 7837 80655 7871
rect 80655 7837 80664 7871
rect 80612 7828 80664 7837
rect 79508 7760 79560 7812
rect 81900 7760 81952 7812
rect 83280 7896 83332 7948
rect 85672 7939 85724 7948
rect 85672 7905 85681 7939
rect 85681 7905 85715 7939
rect 85715 7905 85724 7939
rect 85672 7896 85724 7905
rect 91652 8032 91704 8084
rect 94596 8032 94648 8084
rect 97908 8032 97960 8084
rect 98000 8032 98052 8084
rect 90916 7939 90968 7948
rect 85304 7871 85356 7880
rect 85304 7837 85313 7871
rect 85313 7837 85347 7871
rect 85347 7837 85356 7871
rect 85304 7828 85356 7837
rect 86316 7828 86368 7880
rect 89352 7828 89404 7880
rect 86960 7760 87012 7812
rect 85764 7692 85816 7744
rect 88800 7760 88852 7812
rect 90916 7905 90925 7939
rect 90925 7905 90959 7939
rect 90959 7905 90968 7939
rect 90916 7896 90968 7905
rect 91376 7939 91428 7948
rect 91376 7905 91385 7939
rect 91385 7905 91419 7939
rect 91419 7905 91428 7939
rect 91376 7896 91428 7905
rect 99932 7964 99984 8016
rect 94596 7939 94648 7948
rect 91008 7871 91060 7880
rect 91008 7837 91017 7871
rect 91017 7837 91051 7871
rect 91051 7837 91060 7871
rect 91008 7828 91060 7837
rect 92572 7871 92624 7880
rect 92572 7837 92581 7871
rect 92581 7837 92615 7871
rect 92615 7837 92624 7871
rect 92572 7828 92624 7837
rect 92848 7760 92900 7812
rect 94596 7905 94605 7939
rect 94605 7905 94639 7939
rect 94639 7905 94648 7939
rect 94596 7896 94648 7905
rect 95516 7939 95568 7948
rect 95516 7905 95525 7939
rect 95525 7905 95559 7939
rect 95559 7905 95568 7939
rect 95516 7896 95568 7905
rect 96068 7896 96120 7948
rect 96988 7939 97040 7948
rect 96988 7905 96997 7939
rect 96997 7905 97031 7939
rect 97031 7905 97040 7939
rect 96988 7896 97040 7905
rect 98460 7896 98512 7948
rect 98368 7871 98420 7880
rect 95608 7760 95660 7812
rect 94596 7692 94648 7744
rect 98368 7837 98377 7871
rect 98377 7837 98411 7871
rect 98411 7837 98420 7871
rect 98368 7828 98420 7837
rect 95792 7760 95844 7812
rect 98644 7760 98696 7812
rect 98828 7896 98880 7948
rect 102140 7896 102192 7948
rect 102232 7896 102284 7948
rect 104072 7896 104124 7948
rect 105360 7939 105412 7948
rect 105360 7905 105369 7939
rect 105369 7905 105403 7939
rect 105403 7905 105412 7939
rect 105360 7896 105412 7905
rect 110972 8032 111024 8084
rect 111064 8032 111116 8084
rect 124772 8032 124824 8084
rect 107752 7964 107804 8016
rect 107568 7939 107620 7948
rect 107568 7905 107577 7939
rect 107577 7905 107611 7939
rect 107611 7905 107620 7939
rect 107568 7896 107620 7905
rect 107660 7896 107712 7948
rect 109224 7939 109276 7948
rect 109224 7905 109233 7939
rect 109233 7905 109267 7939
rect 109267 7905 109276 7939
rect 109224 7896 109276 7905
rect 110420 7896 110472 7948
rect 122288 7964 122340 8016
rect 123208 7964 123260 8016
rect 115848 7896 115900 7948
rect 118700 7939 118752 7948
rect 118700 7905 118709 7939
rect 118709 7905 118743 7939
rect 118743 7905 118752 7939
rect 118700 7896 118752 7905
rect 123300 7939 123352 7948
rect 99472 7871 99524 7880
rect 99472 7837 99481 7871
rect 99481 7837 99515 7871
rect 99515 7837 99524 7871
rect 99472 7828 99524 7837
rect 99564 7828 99616 7880
rect 103428 7828 103480 7880
rect 106740 7828 106792 7880
rect 107752 7871 107804 7880
rect 107752 7837 107761 7871
rect 107761 7837 107795 7871
rect 107795 7837 107804 7871
rect 107752 7828 107804 7837
rect 112076 7828 112128 7880
rect 116308 7871 116360 7880
rect 116308 7837 116317 7871
rect 116317 7837 116351 7871
rect 116351 7837 116360 7871
rect 116308 7828 116360 7837
rect 119068 7828 119120 7880
rect 122656 7828 122708 7880
rect 103888 7803 103940 7812
rect 100944 7692 100996 7744
rect 103888 7769 103897 7803
rect 103897 7769 103931 7803
rect 103931 7769 103940 7803
rect 103888 7760 103940 7769
rect 106280 7760 106332 7812
rect 104808 7692 104860 7744
rect 109040 7735 109092 7744
rect 109040 7701 109049 7735
rect 109049 7701 109083 7735
rect 109083 7701 109092 7735
rect 109040 7692 109092 7701
rect 110788 7692 110840 7744
rect 111984 7692 112036 7744
rect 114192 7760 114244 7812
rect 119988 7760 120040 7812
rect 120172 7803 120224 7812
rect 120172 7769 120181 7803
rect 120181 7769 120215 7803
rect 120215 7769 120224 7803
rect 120172 7760 120224 7769
rect 118240 7692 118292 7744
rect 123300 7905 123309 7939
rect 123309 7905 123343 7939
rect 123343 7905 123352 7939
rect 123300 7896 123352 7905
rect 124864 7939 124916 7948
rect 124864 7905 124873 7939
rect 124873 7905 124907 7939
rect 124907 7905 124916 7939
rect 124864 7896 124916 7905
rect 124404 7760 124456 7812
rect 141148 8032 141200 8084
rect 141240 8032 141292 8084
rect 137836 7964 137888 8016
rect 125692 7871 125744 7880
rect 125692 7837 125701 7871
rect 125701 7837 125735 7871
rect 125735 7837 125744 7871
rect 125692 7828 125744 7837
rect 128360 7828 128412 7880
rect 131396 7896 131448 7948
rect 133236 7896 133288 7948
rect 134340 7896 134392 7948
rect 139492 7896 139544 7948
rect 139952 7896 140004 7948
rect 140504 7896 140556 7948
rect 141976 7964 142028 8016
rect 147220 7964 147272 8016
rect 145012 7896 145064 7948
rect 130844 7828 130896 7880
rect 140780 7828 140832 7880
rect 141148 7871 141200 7880
rect 141148 7837 141157 7871
rect 141157 7837 141191 7871
rect 141191 7837 141200 7871
rect 141148 7828 141200 7837
rect 142252 7828 142304 7880
rect 145932 7828 145984 7880
rect 160652 7964 160704 8016
rect 164240 8032 164292 8084
rect 164332 8032 164384 8084
rect 165068 8032 165120 8084
rect 167276 8032 167328 8084
rect 171140 8032 171192 8084
rect 172336 8032 172388 8084
rect 172704 8032 172756 8084
rect 181352 8032 181404 8084
rect 181536 8032 181588 8084
rect 183744 8032 183796 8084
rect 184848 8032 184900 8084
rect 184940 8032 184992 8084
rect 189448 8032 189500 8084
rect 190552 8032 190604 8084
rect 195336 8032 195388 8084
rect 197360 8075 197412 8084
rect 197360 8041 197369 8075
rect 197369 8041 197403 8075
rect 197403 8041 197412 8075
rect 197360 8032 197412 8041
rect 164608 7964 164660 8016
rect 168472 7964 168524 8016
rect 154120 7896 154172 7948
rect 147772 7828 147824 7880
rect 150072 7871 150124 7880
rect 150072 7837 150081 7871
rect 150081 7837 150115 7871
rect 150115 7837 150124 7871
rect 150072 7828 150124 7837
rect 151084 7871 151136 7880
rect 151084 7837 151093 7871
rect 151093 7837 151127 7871
rect 151127 7837 151136 7871
rect 151084 7828 151136 7837
rect 129832 7692 129884 7744
rect 133512 7760 133564 7812
rect 133604 7760 133656 7812
rect 134432 7760 134484 7812
rect 134616 7803 134668 7812
rect 134616 7769 134625 7803
rect 134625 7769 134659 7803
rect 134659 7769 134668 7803
rect 134616 7760 134668 7769
rect 134708 7760 134760 7812
rect 139952 7760 140004 7812
rect 140228 7803 140280 7812
rect 140228 7769 140237 7803
rect 140237 7769 140271 7803
rect 140271 7769 140280 7803
rect 140228 7760 140280 7769
rect 140320 7760 140372 7812
rect 153016 7828 153068 7880
rect 153292 7828 153344 7880
rect 152464 7760 152516 7812
rect 154304 7896 154356 7948
rect 155868 7896 155920 7948
rect 156788 7896 156840 7948
rect 156604 7828 156656 7880
rect 157708 7828 157760 7880
rect 157984 7896 158036 7948
rect 159916 7939 159968 7948
rect 159916 7905 159925 7939
rect 159925 7905 159959 7939
rect 159959 7905 159968 7939
rect 159916 7896 159968 7905
rect 164240 7896 164292 7948
rect 164516 7896 164568 7948
rect 158352 7828 158404 7880
rect 155960 7760 156012 7812
rect 161204 7828 161256 7880
rect 162308 7871 162360 7880
rect 162308 7837 162317 7871
rect 162317 7837 162351 7871
rect 162351 7837 162360 7871
rect 162308 7828 162360 7837
rect 167276 7828 167328 7880
rect 167000 7760 167052 7812
rect 173532 7939 173584 7948
rect 167736 7871 167788 7880
rect 167736 7837 167745 7871
rect 167745 7837 167779 7871
rect 167779 7837 167788 7871
rect 167736 7828 167788 7837
rect 173532 7905 173541 7939
rect 173541 7905 173575 7939
rect 173575 7905 173584 7939
rect 173532 7896 173584 7905
rect 173716 7896 173768 7948
rect 176476 7939 176528 7948
rect 176476 7905 176485 7939
rect 176485 7905 176519 7939
rect 176519 7905 176528 7939
rect 176476 7896 176528 7905
rect 178040 7939 178092 7948
rect 178040 7905 178049 7939
rect 178049 7905 178083 7939
rect 178083 7905 178092 7939
rect 178040 7896 178092 7905
rect 182088 7896 182140 7948
rect 182456 7939 182508 7948
rect 182456 7905 182465 7939
rect 182465 7905 182499 7939
rect 182499 7905 182508 7939
rect 182456 7896 182508 7905
rect 183560 7896 183612 7948
rect 179512 7871 179564 7880
rect 166448 7692 166500 7744
rect 172704 7760 172756 7812
rect 173900 7803 173952 7812
rect 173900 7769 173909 7803
rect 173909 7769 173943 7803
rect 173943 7769 173952 7803
rect 173900 7760 173952 7769
rect 176200 7803 176252 7812
rect 176200 7769 176209 7803
rect 176209 7769 176243 7803
rect 176243 7769 176252 7803
rect 176200 7760 176252 7769
rect 176384 7760 176436 7812
rect 178408 7760 178460 7812
rect 179512 7837 179521 7871
rect 179521 7837 179555 7871
rect 179555 7837 179564 7871
rect 179512 7828 179564 7837
rect 181168 7871 181220 7880
rect 181168 7837 181177 7871
rect 181177 7837 181211 7871
rect 181211 7837 181220 7871
rect 181168 7828 181220 7837
rect 182548 7871 182600 7880
rect 182548 7837 182557 7871
rect 182557 7837 182591 7871
rect 182591 7837 182600 7871
rect 182548 7828 182600 7837
rect 182824 7828 182876 7880
rect 187884 7896 187936 7948
rect 190552 7896 190604 7948
rect 191656 7939 191708 7948
rect 183560 7760 183612 7812
rect 184664 7760 184716 7812
rect 184848 7760 184900 7812
rect 189172 7760 189224 7812
rect 170036 7692 170088 7744
rect 171048 7692 171100 7744
rect 176568 7692 176620 7744
rect 176660 7692 176712 7744
rect 181812 7692 181864 7744
rect 182640 7692 182692 7744
rect 191656 7905 191665 7939
rect 191665 7905 191699 7939
rect 191699 7905 191708 7939
rect 191656 7896 191708 7905
rect 192760 7939 192812 7948
rect 192760 7905 192769 7939
rect 192769 7905 192803 7939
rect 192803 7905 192812 7939
rect 192760 7896 192812 7905
rect 194968 7896 195020 7948
rect 197084 7896 197136 7948
rect 192852 7871 192904 7880
rect 192852 7837 192861 7871
rect 192861 7837 192895 7871
rect 192895 7837 192904 7871
rect 192852 7828 192904 7837
rect 195796 7828 195848 7880
rect 192944 7760 192996 7812
rect 199292 7692 199344 7744
rect 4078 7590 4130 7642
rect 44078 7590 44130 7642
rect 84078 7590 84130 7642
rect 124078 7590 124130 7642
rect 164078 7590 164130 7642
rect 17592 7488 17644 7540
rect 7012 7420 7064 7472
rect 11060 7420 11112 7472
rect 22376 7420 22428 7472
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 7472 7352 7524 7404
rect 11152 7352 11204 7404
rect 6368 7284 6420 7336
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 6920 7216 6972 7268
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 13452 7395 13504 7404
rect 12440 7352 12492 7361
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 12992 7284 13044 7336
rect 13728 7284 13780 7336
rect 16672 7352 16724 7404
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 24860 7395 24912 7404
rect 24860 7361 24869 7395
rect 24869 7361 24903 7395
rect 24903 7361 24912 7395
rect 24860 7352 24912 7361
rect 83004 7488 83056 7540
rect 83832 7488 83884 7540
rect 25412 7420 25464 7472
rect 29460 7395 29512 7404
rect 29460 7361 29469 7395
rect 29469 7361 29503 7395
rect 29503 7361 29512 7395
rect 29460 7352 29512 7361
rect 18052 7327 18104 7336
rect 14188 7216 14240 7268
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 22008 7327 22060 7336
rect 17224 7216 17276 7268
rect 22008 7293 22017 7327
rect 22017 7293 22051 7327
rect 22051 7293 22060 7327
rect 22008 7284 22060 7293
rect 20536 7216 20588 7268
rect 24216 7216 24268 7268
rect 31852 7395 31904 7404
rect 31852 7361 31861 7395
rect 31861 7361 31895 7395
rect 31895 7361 31904 7395
rect 31852 7352 31904 7361
rect 41144 7420 41196 7472
rect 51540 7420 51592 7472
rect 33324 7352 33376 7404
rect 41880 7395 41932 7404
rect 41880 7361 41889 7395
rect 41889 7361 41923 7395
rect 41923 7361 41932 7395
rect 41880 7352 41932 7361
rect 30564 7327 30616 7336
rect 30564 7293 30573 7327
rect 30573 7293 30607 7327
rect 30607 7293 30616 7327
rect 30564 7284 30616 7293
rect 23664 7191 23716 7200
rect 23664 7157 23673 7191
rect 23673 7157 23707 7191
rect 23707 7157 23716 7191
rect 23664 7148 23716 7157
rect 27252 7191 27304 7200
rect 27252 7157 27261 7191
rect 27261 7157 27295 7191
rect 27295 7157 27304 7191
rect 27252 7148 27304 7157
rect 28540 7148 28592 7200
rect 37740 7284 37792 7336
rect 37924 7327 37976 7336
rect 37924 7293 37933 7327
rect 37933 7293 37967 7327
rect 37967 7293 37976 7327
rect 37924 7284 37976 7293
rect 39948 7284 40000 7336
rect 49240 7395 49292 7404
rect 49240 7361 49249 7395
rect 49249 7361 49283 7395
rect 49283 7361 49292 7395
rect 49240 7352 49292 7361
rect 49332 7352 49384 7404
rect 51724 7395 51776 7404
rect 51724 7361 51733 7395
rect 51733 7361 51767 7395
rect 51767 7361 51776 7395
rect 51724 7352 51776 7361
rect 55220 7420 55272 7472
rect 55680 7420 55732 7472
rect 63408 7420 63460 7472
rect 68468 7420 68520 7472
rect 80704 7420 80756 7472
rect 54116 7395 54168 7404
rect 54116 7361 54125 7395
rect 54125 7361 54159 7395
rect 54159 7361 54168 7395
rect 54116 7352 54168 7361
rect 42892 7327 42944 7336
rect 42892 7293 42901 7327
rect 42901 7293 42935 7327
rect 42935 7293 42944 7327
rect 42892 7284 42944 7293
rect 45376 7284 45428 7336
rect 46112 7327 46164 7336
rect 46112 7293 46121 7327
rect 46121 7293 46155 7327
rect 46155 7293 46164 7327
rect 46112 7284 46164 7293
rect 50344 7327 50396 7336
rect 43076 7216 43128 7268
rect 50344 7293 50353 7327
rect 50353 7293 50387 7327
rect 50387 7293 50396 7327
rect 50344 7284 50396 7293
rect 51816 7284 51868 7336
rect 55588 7327 55640 7336
rect 55588 7293 55597 7327
rect 55597 7293 55631 7327
rect 55631 7293 55640 7327
rect 55588 7284 55640 7293
rect 59360 7352 59412 7404
rect 59452 7352 59504 7404
rect 58440 7327 58492 7336
rect 58440 7293 58449 7327
rect 58449 7293 58483 7327
rect 58483 7293 58492 7327
rect 62672 7352 62724 7404
rect 62948 7352 63000 7404
rect 58440 7284 58492 7293
rect 61568 7327 61620 7336
rect 61568 7293 61577 7327
rect 61577 7293 61611 7327
rect 61611 7293 61620 7327
rect 61568 7284 61620 7293
rect 62488 7284 62540 7336
rect 63316 7327 63368 7336
rect 63316 7293 63325 7327
rect 63325 7293 63359 7327
rect 63359 7293 63368 7327
rect 63316 7284 63368 7293
rect 68560 7352 68612 7404
rect 64788 7327 64840 7336
rect 64788 7293 64797 7327
rect 64797 7293 64831 7327
rect 64831 7293 64840 7327
rect 64788 7284 64840 7293
rect 65064 7327 65116 7336
rect 65064 7293 65073 7327
rect 65073 7293 65107 7327
rect 65107 7293 65116 7327
rect 65064 7284 65116 7293
rect 68836 7327 68888 7336
rect 68836 7293 68845 7327
rect 68845 7293 68879 7327
rect 68879 7293 68888 7327
rect 68836 7284 68888 7293
rect 68928 7327 68980 7336
rect 68928 7293 68937 7327
rect 68937 7293 68971 7327
rect 68971 7293 68980 7327
rect 68928 7284 68980 7293
rect 60280 7148 60332 7200
rect 66260 7216 66312 7268
rect 70492 7284 70544 7336
rect 73988 7352 74040 7404
rect 72976 7284 73028 7336
rect 74632 7284 74684 7336
rect 76380 7352 76432 7404
rect 81164 7352 81216 7404
rect 74908 7327 74960 7336
rect 74908 7293 74917 7327
rect 74917 7293 74951 7327
rect 74951 7293 74960 7327
rect 74908 7284 74960 7293
rect 76748 7284 76800 7336
rect 77944 7327 77996 7336
rect 77944 7293 77953 7327
rect 77953 7293 77987 7327
rect 77987 7293 77996 7327
rect 77944 7284 77996 7293
rect 78588 7284 78640 7336
rect 81532 7327 81584 7336
rect 81532 7293 81541 7327
rect 81541 7293 81575 7327
rect 81575 7293 81584 7327
rect 81532 7284 81584 7293
rect 83188 7327 83240 7336
rect 81348 7216 81400 7268
rect 83188 7293 83197 7327
rect 83197 7293 83231 7327
rect 83231 7293 83240 7327
rect 83188 7284 83240 7293
rect 87788 7488 87840 7540
rect 85580 7327 85632 7336
rect 85580 7293 85589 7327
rect 85589 7293 85623 7327
rect 85623 7293 85632 7327
rect 85580 7284 85632 7293
rect 85856 7284 85908 7336
rect 87328 7420 87380 7472
rect 89260 7352 89312 7404
rect 87328 7327 87380 7336
rect 87328 7293 87337 7327
rect 87337 7293 87371 7327
rect 87371 7293 87380 7327
rect 87328 7284 87380 7293
rect 99472 7488 99524 7540
rect 112168 7488 112220 7540
rect 94504 7420 94556 7472
rect 90088 7352 90140 7404
rect 94228 7352 94280 7404
rect 91192 7216 91244 7268
rect 64696 7148 64748 7200
rect 66352 7148 66404 7200
rect 74540 7148 74592 7200
rect 91468 7284 91520 7336
rect 91744 7327 91796 7336
rect 91744 7293 91753 7327
rect 91753 7293 91787 7327
rect 91787 7293 91796 7327
rect 91744 7284 91796 7293
rect 92848 7284 92900 7336
rect 93308 7327 93360 7336
rect 93308 7293 93317 7327
rect 93317 7293 93351 7327
rect 93351 7293 93360 7327
rect 93308 7284 93360 7293
rect 98276 7420 98328 7472
rect 98460 7463 98512 7472
rect 98460 7429 98469 7463
rect 98469 7429 98503 7463
rect 98503 7429 98512 7463
rect 98460 7420 98512 7429
rect 102784 7420 102836 7472
rect 96896 7352 96948 7404
rect 95792 7284 95844 7336
rect 96160 7284 96212 7336
rect 98184 7284 98236 7336
rect 99656 7352 99708 7404
rect 100760 7352 100812 7404
rect 100944 7395 100996 7404
rect 100944 7361 100953 7395
rect 100953 7361 100987 7395
rect 100987 7361 100996 7395
rect 100944 7352 100996 7361
rect 99380 7327 99432 7336
rect 99380 7293 99389 7327
rect 99389 7293 99423 7327
rect 99423 7293 99432 7327
rect 99380 7284 99432 7293
rect 100392 7284 100444 7336
rect 101496 7284 101548 7336
rect 106004 7420 106056 7472
rect 107844 7420 107896 7472
rect 108028 7420 108080 7472
rect 111064 7420 111116 7472
rect 104072 7352 104124 7404
rect 109408 7352 109460 7404
rect 109684 7395 109736 7404
rect 109684 7361 109693 7395
rect 109693 7361 109727 7395
rect 109727 7361 109736 7395
rect 109684 7352 109736 7361
rect 112076 7395 112128 7404
rect 103612 7284 103664 7336
rect 105912 7327 105964 7336
rect 99472 7148 99524 7200
rect 102232 7148 102284 7200
rect 105912 7293 105921 7327
rect 105921 7293 105955 7327
rect 105955 7293 105964 7327
rect 105912 7284 105964 7293
rect 106372 7284 106424 7336
rect 108120 7327 108172 7336
rect 106464 7216 106516 7268
rect 108120 7293 108129 7327
rect 108129 7293 108163 7327
rect 108163 7293 108172 7327
rect 108120 7284 108172 7293
rect 109868 7284 109920 7336
rect 110512 7216 110564 7268
rect 112076 7361 112085 7395
rect 112085 7361 112119 7395
rect 112119 7361 112128 7395
rect 112076 7352 112128 7361
rect 113456 7352 113508 7404
rect 113916 7352 113968 7404
rect 114376 7352 114428 7404
rect 123208 7488 123260 7540
rect 132592 7488 132644 7540
rect 133972 7488 134024 7540
rect 116584 7395 116636 7404
rect 116584 7361 116593 7395
rect 116593 7361 116627 7395
rect 116627 7361 116636 7395
rect 116584 7352 116636 7361
rect 111708 7284 111760 7336
rect 115296 7327 115348 7336
rect 115296 7293 115305 7327
rect 115305 7293 115339 7327
rect 115339 7293 115348 7327
rect 115296 7284 115348 7293
rect 124772 7420 124824 7472
rect 126060 7420 126112 7472
rect 118056 7395 118108 7404
rect 118056 7361 118065 7395
rect 118065 7361 118099 7395
rect 118099 7361 118108 7395
rect 118056 7352 118108 7361
rect 127716 7395 127768 7404
rect 127716 7361 127725 7395
rect 127725 7361 127759 7395
rect 127759 7361 127768 7395
rect 127716 7352 127768 7361
rect 121552 7284 121604 7336
rect 126152 7284 126204 7336
rect 127808 7327 127860 7336
rect 127808 7293 127817 7327
rect 127817 7293 127851 7327
rect 127851 7293 127860 7327
rect 127808 7284 127860 7293
rect 134708 7420 134760 7472
rect 121000 7216 121052 7268
rect 124220 7216 124272 7268
rect 133052 7284 133104 7336
rect 133144 7284 133196 7336
rect 134616 7284 134668 7336
rect 135168 7420 135220 7472
rect 137192 7420 137244 7472
rect 137376 7463 137428 7472
rect 137376 7429 137385 7463
rect 137385 7429 137419 7463
rect 137419 7429 137428 7463
rect 137376 7420 137428 7429
rect 137468 7420 137520 7472
rect 140320 7420 140372 7472
rect 140504 7463 140556 7472
rect 140504 7429 140513 7463
rect 140513 7429 140547 7463
rect 140547 7429 140556 7463
rect 140504 7420 140556 7429
rect 142528 7488 142580 7540
rect 156788 7488 156840 7540
rect 136732 7352 136784 7404
rect 142252 7395 142304 7404
rect 142252 7361 142261 7395
rect 142261 7361 142295 7395
rect 142295 7361 142304 7395
rect 142252 7352 142304 7361
rect 142528 7352 142580 7404
rect 143448 7395 143500 7404
rect 143448 7361 143457 7395
rect 143457 7361 143491 7395
rect 143491 7361 143500 7395
rect 143448 7352 143500 7361
rect 145932 7395 145984 7404
rect 145932 7361 145941 7395
rect 145941 7361 145975 7395
rect 145975 7361 145984 7395
rect 145932 7352 145984 7361
rect 148968 7395 149020 7404
rect 148968 7361 148977 7395
rect 148977 7361 149011 7395
rect 149011 7361 149020 7395
rect 148968 7352 149020 7361
rect 150072 7420 150124 7472
rect 151728 7395 151780 7404
rect 135812 7284 135864 7336
rect 137008 7327 137060 7336
rect 104808 7148 104860 7200
rect 109316 7148 109368 7200
rect 109408 7148 109460 7200
rect 111340 7148 111392 7200
rect 120080 7148 120132 7200
rect 120816 7148 120868 7200
rect 125048 7148 125100 7200
rect 125232 7191 125284 7200
rect 125232 7157 125241 7191
rect 125241 7157 125275 7191
rect 125275 7157 125284 7191
rect 125232 7148 125284 7157
rect 126152 7148 126204 7200
rect 127440 7148 127492 7200
rect 128636 7191 128688 7200
rect 128636 7157 128645 7191
rect 128645 7157 128679 7191
rect 128679 7157 128688 7191
rect 128636 7148 128688 7157
rect 130292 7191 130344 7200
rect 130292 7157 130301 7191
rect 130301 7157 130335 7191
rect 130335 7157 130344 7191
rect 130292 7148 130344 7157
rect 133880 7216 133932 7268
rect 135352 7216 135404 7268
rect 137008 7293 137017 7327
rect 137017 7293 137051 7327
rect 137051 7293 137060 7327
rect 137008 7284 137060 7293
rect 137100 7284 137152 7336
rect 138756 7284 138808 7336
rect 140504 7284 140556 7336
rect 141976 7284 142028 7336
rect 139768 7216 139820 7268
rect 141240 7216 141292 7268
rect 147680 7327 147732 7336
rect 147680 7293 147689 7327
rect 147689 7293 147723 7327
rect 147723 7293 147732 7327
rect 148876 7327 148928 7336
rect 147680 7284 147732 7293
rect 148876 7293 148885 7327
rect 148885 7293 148919 7327
rect 148919 7293 148928 7327
rect 148876 7284 148928 7293
rect 150716 7284 150768 7336
rect 151728 7361 151737 7395
rect 151737 7361 151771 7395
rect 151771 7361 151780 7395
rect 151728 7352 151780 7361
rect 153844 7352 153896 7404
rect 157340 7420 157392 7472
rect 157708 7420 157760 7472
rect 158904 7488 158956 7540
rect 160284 7420 160336 7472
rect 162308 7420 162360 7472
rect 180892 7420 180944 7472
rect 181352 7488 181404 7540
rect 187976 7488 188028 7540
rect 184940 7420 184992 7472
rect 161848 7352 161900 7404
rect 161940 7352 161992 7404
rect 181536 7352 181588 7404
rect 181812 7352 181864 7404
rect 182640 7352 182692 7404
rect 182732 7352 182784 7404
rect 188804 7420 188856 7472
rect 142712 7216 142764 7268
rect 144276 7216 144328 7268
rect 150348 7216 150400 7268
rect 156052 7284 156104 7336
rect 157064 7284 157116 7336
rect 189172 7420 189224 7472
rect 196716 7420 196768 7472
rect 196992 7352 197044 7404
rect 133144 7148 133196 7200
rect 133696 7191 133748 7200
rect 133696 7157 133705 7191
rect 133705 7157 133739 7191
rect 133739 7157 133748 7191
rect 133696 7148 133748 7157
rect 133788 7148 133840 7200
rect 24078 7046 24130 7098
rect 64078 7046 64130 7098
rect 104078 7046 104130 7098
rect 144078 7046 144130 7098
rect 16948 6944 17000 6996
rect 18052 6944 18104 6996
rect 25320 6944 25372 6996
rect 30564 6944 30616 6996
rect 91744 6944 91796 6996
rect 95884 6944 95936 6996
rect 96528 6944 96580 6996
rect 99380 6944 99432 6996
rect 99472 6987 99524 6996
rect 99472 6953 99481 6987
rect 99481 6953 99515 6987
rect 99515 6953 99524 6987
rect 99472 6944 99524 6953
rect 105636 6944 105688 6996
rect 108028 6944 108080 6996
rect 120172 6944 120224 6996
rect 137468 6944 137520 6996
rect 137928 6944 137980 6996
rect 139584 6944 139636 6996
rect 139768 6987 139820 6996
rect 139768 6953 139777 6987
rect 139777 6953 139811 6987
rect 139811 6953 139820 6987
rect 139768 6944 139820 6953
rect 140320 6944 140372 6996
rect 144000 6944 144052 6996
rect 42432 6876 42484 6928
rect 49332 6876 49384 6928
rect 52460 6876 52512 6928
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 5724 6808 5776 6860
rect 7196 6808 7248 6860
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 9680 6808 9732 6860
rect 11704 6851 11756 6860
rect 11704 6817 11713 6851
rect 11713 6817 11747 6851
rect 11747 6817 11756 6851
rect 11704 6808 11756 6817
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 21732 6808 21784 6860
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 23572 6808 23624 6860
rect 24952 6851 25004 6860
rect 24952 6817 24961 6851
rect 24961 6817 24995 6851
rect 24995 6817 25004 6851
rect 24952 6808 25004 6817
rect 27252 6808 27304 6860
rect 27712 6851 27764 6860
rect 27712 6817 27721 6851
rect 27721 6817 27755 6851
rect 27755 6817 27764 6851
rect 27712 6808 27764 6817
rect 28448 6808 28500 6860
rect 30288 6808 30340 6860
rect 33324 6851 33376 6860
rect 33324 6817 33333 6851
rect 33333 6817 33367 6851
rect 33367 6817 33376 6851
rect 33324 6808 33376 6817
rect 33968 6808 34020 6860
rect 35900 6808 35952 6860
rect 37740 6808 37792 6860
rect 38200 6808 38252 6860
rect 39948 6808 40000 6860
rect 42892 6808 42944 6860
rect 45560 6851 45612 6860
rect 45560 6817 45569 6851
rect 45569 6817 45603 6851
rect 45603 6817 45612 6851
rect 45560 6808 45612 6817
rect 47308 6808 47360 6860
rect 47584 6851 47636 6860
rect 47584 6817 47593 6851
rect 47593 6817 47627 6851
rect 47627 6817 47636 6851
rect 47584 6808 47636 6817
rect 48964 6851 49016 6860
rect 48964 6817 48973 6851
rect 48973 6817 49007 6851
rect 49007 6817 49016 6851
rect 48964 6808 49016 6817
rect 49148 6808 49200 6860
rect 52552 6808 52604 6860
rect 52644 6808 52696 6860
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 6736 6740 6788 6792
rect 8484 6740 8536 6792
rect 9772 6740 9824 6792
rect 12348 6740 12400 6792
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 17960 6740 18012 6792
rect 21916 6740 21968 6792
rect 23756 6740 23808 6792
rect 26700 6740 26752 6792
rect 28632 6740 28684 6792
rect 29644 6740 29696 6792
rect 37832 6740 37884 6792
rect 40684 6740 40736 6792
rect 572 6672 624 6724
rect 2320 6604 2372 6656
rect 3792 6604 3844 6656
rect 3976 6672 4028 6724
rect 11336 6672 11388 6724
rect 30196 6672 30248 6724
rect 37188 6672 37240 6724
rect 41420 6672 41472 6724
rect 42616 6740 42668 6792
rect 45928 6740 45980 6792
rect 47676 6740 47728 6792
rect 7840 6604 7892 6656
rect 28908 6604 28960 6656
rect 33232 6604 33284 6656
rect 50436 6604 50488 6656
rect 53012 6740 53064 6792
rect 56600 6808 56652 6860
rect 58624 6808 58676 6860
rect 58808 6851 58860 6860
rect 58808 6817 58817 6851
rect 58817 6817 58851 6851
rect 58851 6817 58860 6851
rect 58808 6808 58860 6817
rect 57336 6740 57388 6792
rect 57704 6740 57756 6792
rect 62580 6808 62632 6860
rect 63776 6808 63828 6860
rect 64052 6851 64104 6860
rect 64052 6817 64061 6851
rect 64061 6817 64095 6851
rect 64095 6817 64104 6851
rect 64052 6808 64104 6817
rect 64236 6808 64288 6860
rect 66352 6808 66404 6860
rect 61660 6740 61712 6792
rect 65524 6740 65576 6792
rect 67180 6808 67232 6860
rect 66812 6740 66864 6792
rect 66444 6672 66496 6724
rect 69020 6808 69072 6860
rect 70308 6808 70360 6860
rect 69480 6783 69532 6792
rect 69480 6749 69489 6783
rect 69489 6749 69523 6783
rect 69523 6749 69532 6783
rect 69480 6740 69532 6749
rect 69848 6740 69900 6792
rect 70216 6672 70268 6724
rect 74264 6808 74316 6860
rect 73252 6672 73304 6724
rect 74540 6740 74592 6792
rect 76472 6808 76524 6860
rect 82636 6851 82688 6860
rect 81532 6740 81584 6792
rect 82636 6817 82645 6851
rect 82645 6817 82679 6851
rect 82679 6817 82688 6851
rect 82636 6808 82688 6817
rect 83372 6851 83424 6860
rect 83004 6783 83056 6792
rect 83004 6749 83013 6783
rect 83013 6749 83047 6783
rect 83047 6749 83056 6783
rect 83004 6740 83056 6749
rect 83372 6817 83381 6851
rect 83381 6817 83415 6851
rect 83415 6817 83424 6851
rect 83372 6808 83424 6817
rect 85120 6808 85172 6860
rect 86960 6876 87012 6928
rect 84292 6740 84344 6792
rect 89904 6808 89956 6860
rect 90364 6851 90416 6860
rect 90364 6817 90373 6851
rect 90373 6817 90407 6851
rect 90407 6817 90416 6851
rect 90364 6808 90416 6817
rect 92112 6808 92164 6860
rect 95148 6851 95200 6860
rect 95148 6817 95157 6851
rect 95157 6817 95191 6851
rect 95191 6817 95200 6851
rect 95148 6808 95200 6817
rect 97908 6876 97960 6928
rect 105912 6876 105964 6928
rect 96344 6808 96396 6860
rect 96712 6808 96764 6860
rect 97448 6808 97500 6860
rect 96252 6740 96304 6792
rect 99564 6808 99616 6860
rect 99748 6808 99800 6860
rect 103060 6808 103112 6860
rect 106556 6876 106608 6928
rect 99288 6740 99340 6792
rect 104440 6740 104492 6792
rect 105084 6740 105136 6792
rect 58624 6647 58676 6656
rect 58624 6613 58633 6647
rect 58633 6613 58667 6647
rect 58667 6613 58676 6647
rect 58624 6604 58676 6613
rect 58900 6604 58952 6656
rect 62304 6647 62356 6656
rect 62304 6613 62313 6647
rect 62313 6613 62347 6647
rect 62347 6613 62356 6647
rect 62304 6604 62356 6613
rect 63500 6604 63552 6656
rect 66260 6604 66312 6656
rect 67640 6647 67692 6656
rect 67640 6613 67649 6647
rect 67649 6613 67683 6647
rect 67683 6613 67692 6647
rect 67640 6604 67692 6613
rect 67732 6604 67784 6656
rect 68836 6604 68888 6656
rect 69020 6604 69072 6656
rect 70124 6604 70176 6656
rect 71504 6647 71556 6656
rect 71504 6613 71513 6647
rect 71513 6613 71547 6647
rect 71547 6613 71556 6647
rect 71504 6604 71556 6613
rect 72792 6604 72844 6656
rect 76196 6604 76248 6656
rect 80796 6604 80848 6656
rect 83464 6604 83516 6656
rect 84660 6604 84712 6656
rect 90180 6647 90232 6656
rect 90180 6613 90189 6647
rect 90189 6613 90223 6647
rect 90223 6613 90232 6647
rect 90180 6604 90232 6613
rect 91652 6604 91704 6656
rect 93584 6604 93636 6656
rect 97632 6604 97684 6656
rect 97816 6647 97868 6656
rect 97816 6613 97825 6647
rect 97825 6613 97859 6647
rect 97859 6613 97868 6647
rect 97816 6604 97868 6613
rect 98000 6672 98052 6724
rect 101680 6672 101732 6724
rect 102692 6672 102744 6724
rect 106096 6672 106148 6724
rect 111064 6808 111116 6860
rect 115112 6851 115164 6860
rect 106280 6740 106332 6792
rect 108856 6783 108908 6792
rect 108856 6749 108865 6783
rect 108865 6749 108899 6783
rect 108899 6749 108908 6783
rect 108856 6740 108908 6749
rect 109500 6740 109552 6792
rect 115112 6817 115121 6851
rect 115121 6817 115155 6851
rect 115155 6817 115164 6851
rect 115112 6808 115164 6817
rect 127716 6876 127768 6928
rect 115664 6808 115716 6860
rect 116308 6851 116360 6860
rect 116308 6817 116317 6851
rect 116317 6817 116351 6851
rect 116351 6817 116360 6851
rect 116308 6808 116360 6817
rect 119804 6808 119856 6860
rect 120172 6851 120224 6860
rect 120172 6817 120181 6851
rect 120181 6817 120215 6851
rect 120215 6817 120224 6851
rect 120172 6808 120224 6817
rect 120264 6808 120316 6860
rect 123668 6808 123720 6860
rect 124588 6851 124640 6860
rect 124588 6817 124597 6851
rect 124597 6817 124631 6851
rect 124631 6817 124640 6851
rect 124588 6808 124640 6817
rect 125508 6808 125560 6860
rect 125968 6808 126020 6860
rect 129096 6808 129148 6860
rect 129280 6851 129332 6860
rect 129280 6817 129289 6851
rect 129289 6817 129323 6851
rect 129323 6817 129332 6851
rect 129280 6808 129332 6817
rect 114468 6740 114520 6792
rect 114836 6740 114888 6792
rect 106648 6672 106700 6724
rect 99196 6604 99248 6656
rect 106832 6672 106884 6724
rect 115756 6672 115808 6724
rect 118148 6740 118200 6792
rect 118700 6783 118752 6792
rect 118700 6749 118709 6783
rect 118709 6749 118743 6783
rect 118743 6749 118752 6783
rect 118700 6740 118752 6749
rect 118884 6740 118936 6792
rect 122104 6740 122156 6792
rect 124220 6740 124272 6792
rect 124312 6740 124364 6792
rect 124956 6740 125008 6792
rect 127624 6740 127676 6792
rect 127900 6783 127952 6792
rect 127900 6749 127909 6783
rect 127909 6749 127943 6783
rect 127943 6749 127952 6783
rect 127900 6740 127952 6749
rect 131304 6808 131356 6860
rect 131488 6851 131540 6860
rect 131488 6817 131497 6851
rect 131497 6817 131531 6851
rect 131531 6817 131540 6851
rect 131488 6808 131540 6817
rect 134064 6808 134116 6860
rect 134340 6808 134392 6860
rect 134432 6808 134484 6860
rect 135536 6808 135588 6860
rect 135720 6851 135772 6860
rect 135720 6817 135729 6851
rect 135729 6817 135763 6851
rect 135763 6817 135772 6851
rect 135720 6808 135772 6817
rect 131764 6783 131816 6792
rect 131764 6749 131773 6783
rect 131773 6749 131807 6783
rect 131807 6749 131816 6783
rect 131764 6740 131816 6749
rect 132500 6740 132552 6792
rect 133328 6740 133380 6792
rect 135260 6740 135312 6792
rect 135628 6783 135680 6792
rect 135628 6749 135637 6783
rect 135637 6749 135671 6783
rect 135671 6749 135680 6783
rect 135628 6740 135680 6749
rect 110604 6604 110656 6656
rect 110788 6647 110840 6656
rect 110788 6613 110797 6647
rect 110797 6613 110831 6647
rect 110831 6613 110840 6647
rect 110788 6604 110840 6613
rect 112260 6604 112312 6656
rect 118332 6604 118384 6656
rect 128820 6672 128872 6724
rect 131212 6672 131264 6724
rect 132040 6672 132092 6724
rect 132592 6672 132644 6724
rect 140688 6876 140740 6928
rect 147864 6876 147916 6928
rect 141056 6808 141108 6860
rect 141148 6808 141200 6860
rect 136640 6740 136692 6792
rect 137652 6740 137704 6792
rect 138480 6672 138532 6724
rect 139032 6740 139084 6792
rect 143632 6808 143684 6860
rect 147772 6808 147824 6860
rect 147956 6851 148008 6860
rect 147956 6817 147965 6851
rect 147965 6817 147999 6851
rect 147999 6817 148008 6851
rect 147956 6808 148008 6817
rect 150716 6851 150768 6860
rect 150716 6817 150725 6851
rect 150725 6817 150759 6851
rect 150759 6817 150768 6851
rect 150716 6808 150768 6817
rect 151084 6808 151136 6860
rect 153016 6851 153068 6860
rect 153016 6817 153025 6851
rect 153025 6817 153059 6851
rect 153059 6817 153068 6851
rect 153016 6808 153068 6817
rect 144920 6740 144972 6792
rect 141148 6672 141200 6724
rect 152556 6740 152608 6792
rect 153108 6783 153160 6792
rect 153108 6749 153117 6783
rect 153117 6749 153151 6783
rect 153151 6749 153160 6783
rect 153108 6740 153160 6749
rect 125784 6604 125836 6656
rect 125968 6604 126020 6656
rect 130200 6604 130252 6656
rect 130476 6604 130528 6656
rect 154856 6604 154908 6656
rect 4078 6502 4130 6554
rect 44078 6502 44130 6554
rect 84078 6502 84130 6554
rect 124078 6502 124130 6554
rect 3792 6400 3844 6452
rect 7288 6400 7340 6452
rect 27160 6400 27212 6452
rect 1860 6332 1912 6384
rect 6920 6332 6972 6384
rect 4620 6264 4672 6316
rect 8760 6332 8812 6384
rect 15016 6332 15068 6384
rect 17132 6332 17184 6384
rect 19340 6332 19392 6384
rect 20904 6332 20956 6384
rect 26884 6332 26936 6384
rect 27620 6332 27672 6384
rect 29368 6332 29420 6384
rect 1952 6196 2004 6248
rect 6736 6196 6788 6248
rect 6920 6196 6972 6248
rect 7564 6196 7616 6248
rect 7840 6128 7892 6180
rect 8392 6264 8444 6316
rect 15568 6307 15620 6316
rect 15568 6273 15577 6307
rect 15577 6273 15611 6307
rect 15611 6273 15620 6307
rect 15568 6264 15620 6273
rect 18420 6264 18472 6316
rect 20628 6264 20680 6316
rect 23664 6307 23716 6316
rect 23664 6273 23673 6307
rect 23673 6273 23707 6307
rect 23707 6273 23716 6307
rect 23664 6264 23716 6273
rect 25044 6307 25096 6316
rect 25044 6273 25053 6307
rect 25053 6273 25087 6307
rect 25087 6273 25096 6307
rect 25044 6264 25096 6273
rect 26332 6264 26384 6316
rect 29644 6307 29696 6316
rect 29644 6273 29653 6307
rect 29653 6273 29687 6307
rect 29687 6273 29696 6307
rect 29644 6264 29696 6273
rect 36360 6400 36412 6452
rect 35440 6332 35492 6384
rect 37648 6332 37700 6384
rect 50712 6400 50764 6452
rect 60832 6400 60884 6452
rect 37832 6307 37884 6316
rect 37832 6273 37841 6307
rect 37841 6273 37875 6307
rect 37875 6273 37884 6307
rect 37832 6264 37884 6273
rect 42616 6307 42668 6316
rect 42616 6273 42625 6307
rect 42625 6273 42659 6307
rect 42659 6273 42668 6307
rect 42616 6264 42668 6273
rect 43720 6332 43772 6384
rect 44640 6332 44692 6384
rect 52920 6332 52972 6384
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 19432 6239 19484 6248
rect 19432 6205 19441 6239
rect 19441 6205 19475 6239
rect 19475 6205 19484 6239
rect 19432 6196 19484 6205
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 24860 6239 24912 6248
rect 24860 6205 24869 6239
rect 24869 6205 24903 6239
rect 24903 6205 24912 6239
rect 24860 6196 24912 6205
rect 27620 6196 27672 6248
rect 27896 6239 27948 6248
rect 27896 6205 27905 6239
rect 27905 6205 27939 6239
rect 27939 6205 27948 6239
rect 27896 6196 27948 6205
rect 13728 6128 13780 6180
rect 21916 6128 21968 6180
rect 32404 6196 32456 6248
rect 33876 6196 33928 6248
rect 36084 6196 36136 6248
rect 36544 6239 36596 6248
rect 36544 6205 36553 6239
rect 36553 6205 36587 6239
rect 36587 6205 36596 6239
rect 36544 6196 36596 6205
rect 39396 6239 39448 6248
rect 39396 6205 39405 6239
rect 39405 6205 39439 6239
rect 39439 6205 39448 6239
rect 39396 6196 39448 6205
rect 43996 6196 44048 6248
rect 44272 6196 44324 6248
rect 46112 6239 46164 6248
rect 46112 6205 46121 6239
rect 46121 6205 46155 6239
rect 46155 6205 46164 6239
rect 46112 6196 46164 6205
rect 47032 6196 47084 6248
rect 32772 6128 32824 6180
rect 39856 6128 39908 6180
rect 49424 6264 49476 6316
rect 53012 6307 53064 6316
rect 53012 6273 53021 6307
rect 53021 6273 53055 6307
rect 53055 6273 53064 6307
rect 53012 6264 53064 6273
rect 57244 6332 57296 6384
rect 57336 6307 57388 6316
rect 57336 6273 57345 6307
rect 57345 6273 57379 6307
rect 57379 6273 57388 6307
rect 57336 6264 57388 6273
rect 62120 6332 62172 6384
rect 66996 6332 67048 6384
rect 73712 6400 73764 6452
rect 106832 6400 106884 6452
rect 108396 6400 108448 6452
rect 110604 6400 110656 6452
rect 68836 6332 68888 6384
rect 64052 6264 64104 6316
rect 67180 6307 67232 6316
rect 67180 6273 67189 6307
rect 67189 6273 67223 6307
rect 67223 6273 67232 6307
rect 67180 6264 67232 6273
rect 48504 6239 48556 6248
rect 48504 6205 48513 6239
rect 48513 6205 48547 6239
rect 48547 6205 48556 6239
rect 48504 6196 48556 6205
rect 49700 6239 49752 6248
rect 49700 6205 49709 6239
rect 49709 6205 49743 6239
rect 49743 6205 49752 6239
rect 49700 6196 49752 6205
rect 54116 6239 54168 6248
rect 54116 6205 54125 6239
rect 54125 6205 54159 6239
rect 54159 6205 54168 6239
rect 54116 6196 54168 6205
rect 59452 6196 59504 6248
rect 63868 6239 63920 6248
rect 63868 6205 63877 6239
rect 63877 6205 63911 6239
rect 63911 6205 63920 6239
rect 63868 6196 63920 6205
rect 64604 6196 64656 6248
rect 64696 6196 64748 6248
rect 66904 6196 66956 6248
rect 70952 6332 71004 6384
rect 72056 6332 72108 6384
rect 72700 6332 72752 6384
rect 78220 6375 78272 6384
rect 78220 6341 78229 6375
rect 78229 6341 78263 6375
rect 78263 6341 78272 6375
rect 78220 6332 78272 6341
rect 79324 6332 79376 6384
rect 69020 6196 69072 6248
rect 69572 6264 69624 6316
rect 70400 6239 70452 6248
rect 70400 6205 70409 6239
rect 70409 6205 70443 6239
rect 70443 6205 70452 6239
rect 70676 6239 70728 6248
rect 70400 6196 70452 6205
rect 70676 6205 70685 6239
rect 70685 6205 70719 6239
rect 70719 6205 70728 6239
rect 70676 6196 70728 6205
rect 71780 6239 71832 6248
rect 71780 6205 71789 6239
rect 71789 6205 71823 6239
rect 71823 6205 71832 6239
rect 71780 6196 71832 6205
rect 71872 6196 71924 6248
rect 73344 6264 73396 6316
rect 77300 6264 77352 6316
rect 79048 6264 79100 6316
rect 76656 6239 76708 6248
rect 76656 6205 76665 6239
rect 76665 6205 76699 6239
rect 76699 6205 76708 6239
rect 76656 6196 76708 6205
rect 77760 6196 77812 6248
rect 78404 6239 78456 6248
rect 78404 6205 78413 6239
rect 78413 6205 78447 6239
rect 78447 6205 78456 6239
rect 78404 6196 78456 6205
rect 79876 6196 79928 6248
rect 80060 6239 80112 6248
rect 80060 6205 80069 6239
rect 80069 6205 80103 6239
rect 80103 6205 80112 6239
rect 81992 6332 82044 6384
rect 88432 6332 88484 6384
rect 89260 6332 89312 6384
rect 80060 6196 80112 6205
rect 81440 6239 81492 6248
rect 81440 6205 81449 6239
rect 81449 6205 81483 6239
rect 81483 6205 81492 6239
rect 81440 6196 81492 6205
rect 81716 6239 81768 6248
rect 81716 6205 81725 6239
rect 81725 6205 81759 6239
rect 81759 6205 81768 6239
rect 81716 6196 81768 6205
rect 81900 6239 81952 6248
rect 81900 6205 81909 6239
rect 81909 6205 81943 6239
rect 81943 6205 81952 6239
rect 81900 6196 81952 6205
rect 82912 6239 82964 6248
rect 82912 6205 82921 6239
rect 82921 6205 82955 6239
rect 82955 6205 82964 6239
rect 82912 6196 82964 6205
rect 83464 6239 83516 6248
rect 83464 6205 83473 6239
rect 83473 6205 83507 6239
rect 83507 6205 83516 6239
rect 83464 6196 83516 6205
rect 85212 6196 85264 6248
rect 85764 6239 85816 6248
rect 85764 6205 85773 6239
rect 85773 6205 85807 6239
rect 85807 6205 85816 6239
rect 85764 6196 85816 6205
rect 86868 6196 86920 6248
rect 87144 6239 87196 6248
rect 87144 6205 87153 6239
rect 87153 6205 87187 6239
rect 87187 6205 87196 6239
rect 87144 6196 87196 6205
rect 87420 6196 87472 6248
rect 88156 6196 88208 6248
rect 89812 6264 89864 6316
rect 89168 6196 89220 6248
rect 61844 6128 61896 6180
rect 81808 6128 81860 6180
rect 82176 6128 82228 6180
rect 91744 6332 91796 6384
rect 95148 6332 95200 6384
rect 97540 6264 97592 6316
rect 99288 6332 99340 6384
rect 99932 6264 99984 6316
rect 100116 6332 100168 6384
rect 100576 6264 100628 6316
rect 91560 6196 91612 6248
rect 92940 6239 92992 6248
rect 92940 6205 92949 6239
rect 92949 6205 92983 6239
rect 92983 6205 92992 6239
rect 92940 6196 92992 6205
rect 93124 6196 93176 6248
rect 93860 6196 93912 6248
rect 94964 6239 95016 6248
rect 94964 6205 94973 6239
rect 94973 6205 95007 6239
rect 95007 6205 95016 6239
rect 94964 6196 95016 6205
rect 95148 6239 95200 6248
rect 95148 6205 95157 6239
rect 95157 6205 95191 6239
rect 95191 6205 95200 6239
rect 95148 6196 95200 6205
rect 96804 6196 96856 6248
rect 91744 6128 91796 6180
rect 96896 6128 96948 6180
rect 3240 6060 3292 6112
rect 6828 6060 6880 6112
rect 6920 6060 6972 6112
rect 9680 6060 9732 6112
rect 21548 6060 21600 6112
rect 22468 6060 22520 6112
rect 29828 6060 29880 6112
rect 30380 6060 30432 6112
rect 45468 6060 45520 6112
rect 50436 6060 50488 6112
rect 50528 6060 50580 6112
rect 54576 6060 54628 6112
rect 56784 6060 56836 6112
rect 59176 6060 59228 6112
rect 59820 6060 59872 6112
rect 61936 6060 61988 6112
rect 67732 6060 67784 6112
rect 69112 6060 69164 6112
rect 77024 6060 77076 6112
rect 91560 6060 91612 6112
rect 96988 6060 97040 6112
rect 97356 6196 97408 6248
rect 98000 6196 98052 6248
rect 98644 6239 98696 6248
rect 98644 6205 98653 6239
rect 98653 6205 98687 6239
rect 98687 6205 98696 6239
rect 98644 6196 98696 6205
rect 98828 6239 98880 6248
rect 98828 6205 98837 6239
rect 98837 6205 98871 6239
rect 98871 6205 98880 6239
rect 98828 6196 98880 6205
rect 99472 6196 99524 6248
rect 104716 6264 104768 6316
rect 106280 6307 106332 6316
rect 103888 6239 103940 6248
rect 99012 6060 99064 6112
rect 99288 6060 99340 6112
rect 100024 6060 100076 6112
rect 101220 6060 101272 6112
rect 103888 6205 103897 6239
rect 103897 6205 103931 6239
rect 103931 6205 103940 6239
rect 103888 6196 103940 6205
rect 106280 6273 106289 6307
rect 106289 6273 106323 6307
rect 106323 6273 106332 6307
rect 106280 6264 106332 6273
rect 106556 6332 106608 6384
rect 108580 6332 108632 6384
rect 108672 6332 108724 6384
rect 109868 6264 109920 6316
rect 105360 6239 105412 6248
rect 105360 6205 105369 6239
rect 105369 6205 105403 6239
rect 105403 6205 105412 6239
rect 105360 6196 105412 6205
rect 105544 6196 105596 6248
rect 108028 6239 108080 6248
rect 108028 6205 108037 6239
rect 108037 6205 108071 6239
rect 108071 6205 108080 6239
rect 108028 6196 108080 6205
rect 108212 6239 108264 6248
rect 108212 6205 108221 6239
rect 108221 6205 108255 6239
rect 108255 6205 108264 6239
rect 108212 6196 108264 6205
rect 108396 6239 108448 6248
rect 108396 6205 108405 6239
rect 108405 6205 108439 6239
rect 108439 6205 108448 6239
rect 108396 6196 108448 6205
rect 109592 6239 109644 6248
rect 109592 6205 109601 6239
rect 109601 6205 109635 6239
rect 109635 6205 109644 6239
rect 109592 6196 109644 6205
rect 109776 6239 109828 6248
rect 109776 6205 109785 6239
rect 109785 6205 109819 6239
rect 109819 6205 109828 6239
rect 109776 6196 109828 6205
rect 110052 6332 110104 6384
rect 111248 6332 111300 6384
rect 116032 6332 116084 6384
rect 111432 6196 111484 6248
rect 112536 6196 112588 6248
rect 116400 6239 116452 6248
rect 116400 6205 116409 6239
rect 116409 6205 116443 6239
rect 116443 6205 116452 6239
rect 116400 6196 116452 6205
rect 106556 6060 106608 6112
rect 106648 6060 106700 6112
rect 107568 6060 107620 6112
rect 107660 6060 107712 6112
rect 117504 6128 117556 6180
rect 118700 6264 118752 6316
rect 119068 6307 119120 6316
rect 119068 6273 119077 6307
rect 119077 6273 119111 6307
rect 119111 6273 119120 6307
rect 119068 6264 119120 6273
rect 119804 6400 119856 6452
rect 122012 6400 122064 6452
rect 122104 6400 122156 6452
rect 122748 6400 122800 6452
rect 123116 6400 123168 6452
rect 126060 6400 126112 6452
rect 124404 6332 124456 6384
rect 120540 6307 120592 6316
rect 120540 6273 120549 6307
rect 120549 6273 120583 6307
rect 120583 6273 120592 6307
rect 120540 6264 120592 6273
rect 121460 6307 121512 6316
rect 121460 6273 121469 6307
rect 121469 6273 121503 6307
rect 121503 6273 121512 6307
rect 121460 6264 121512 6273
rect 125968 6264 126020 6316
rect 128268 6264 128320 6316
rect 131764 6332 131816 6384
rect 131948 6400 132000 6452
rect 138296 6400 138348 6452
rect 149980 6400 150032 6452
rect 120080 6128 120132 6180
rect 120632 6239 120684 6248
rect 120632 6205 120641 6239
rect 120641 6205 120675 6239
rect 120675 6205 120684 6239
rect 120632 6196 120684 6205
rect 120816 6196 120868 6248
rect 122840 6239 122892 6248
rect 122840 6205 122849 6239
rect 122849 6205 122883 6239
rect 122883 6205 122892 6239
rect 122840 6196 122892 6205
rect 123760 6196 123812 6248
rect 124404 6196 124456 6248
rect 124680 6239 124732 6248
rect 124680 6205 124689 6239
rect 124689 6205 124723 6239
rect 124723 6205 124732 6239
rect 124680 6196 124732 6205
rect 125784 6239 125836 6248
rect 125784 6205 125793 6239
rect 125793 6205 125827 6239
rect 125827 6205 125836 6239
rect 125784 6196 125836 6205
rect 130936 6196 130988 6248
rect 132592 6264 132644 6316
rect 132776 6307 132828 6316
rect 132776 6273 132785 6307
rect 132785 6273 132819 6307
rect 132819 6273 132828 6307
rect 132776 6264 132828 6273
rect 132224 6196 132276 6248
rect 113548 6060 113600 6112
rect 118608 6060 118660 6112
rect 120816 6060 120868 6112
rect 125508 6060 125560 6112
rect 125692 6060 125744 6112
rect 127624 6060 127676 6112
rect 130200 6128 130252 6180
rect 129188 6060 129240 6112
rect 131120 6060 131172 6112
rect 131580 6128 131632 6180
rect 133604 6264 133656 6316
rect 133972 6264 134024 6316
rect 135904 6264 135956 6316
rect 137560 6307 137612 6316
rect 133512 6196 133564 6248
rect 134432 6196 134484 6248
rect 133604 6060 133656 6112
rect 133972 6128 134024 6180
rect 134984 6196 135036 6248
rect 136548 6196 136600 6248
rect 136732 6196 136784 6248
rect 137560 6273 137569 6307
rect 137569 6273 137603 6307
rect 137603 6273 137612 6307
rect 137560 6264 137612 6273
rect 155316 6332 155368 6384
rect 138480 6239 138532 6248
rect 138480 6205 138489 6239
rect 138489 6205 138523 6239
rect 138523 6205 138532 6239
rect 138480 6196 138532 6205
rect 139584 6239 139636 6248
rect 139584 6205 139593 6239
rect 139593 6205 139627 6239
rect 139627 6205 139636 6239
rect 139584 6196 139636 6205
rect 140504 6264 140556 6316
rect 142620 6264 142672 6316
rect 145380 6307 145432 6316
rect 143908 6239 143960 6248
rect 143908 6205 143917 6239
rect 143917 6205 143951 6239
rect 143951 6205 143960 6239
rect 143908 6196 143960 6205
rect 145104 6239 145156 6248
rect 145104 6205 145113 6239
rect 145113 6205 145147 6239
rect 145147 6205 145156 6239
rect 145104 6196 145156 6205
rect 145380 6273 145389 6307
rect 145389 6273 145423 6307
rect 145423 6273 145432 6307
rect 145380 6264 145432 6273
rect 147680 6264 147732 6316
rect 150624 6307 150676 6316
rect 150624 6273 150633 6307
rect 150633 6273 150667 6307
rect 150667 6273 150676 6307
rect 150624 6264 150676 6273
rect 151636 6307 151688 6316
rect 151636 6273 151645 6307
rect 151645 6273 151679 6307
rect 151679 6273 151688 6307
rect 151636 6264 151688 6273
rect 153292 6307 153344 6316
rect 153292 6273 153301 6307
rect 153301 6273 153335 6307
rect 153335 6273 153344 6307
rect 153292 6264 153344 6273
rect 153936 6196 153988 6248
rect 134708 6060 134760 6112
rect 135536 6128 135588 6180
rect 152188 6128 152240 6180
rect 140412 6060 140464 6112
rect 145104 6060 145156 6112
rect 145840 6060 145892 6112
rect 24078 5958 24130 6010
rect 64078 5958 64130 6010
rect 104078 5958 104130 6010
rect 144078 5958 144130 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 6736 5856 6788 5908
rect 8576 5856 8628 5908
rect 10140 5856 10192 5908
rect 10232 5856 10284 5908
rect 13452 5856 13504 5908
rect 21088 5856 21140 5908
rect 27620 5899 27672 5908
rect 4712 5788 4764 5840
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 7472 5652 7524 5704
rect 3608 5584 3660 5636
rect 12256 5788 12308 5840
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 8944 5652 8996 5704
rect 13452 5763 13504 5772
rect 13452 5729 13461 5763
rect 13461 5729 13495 5763
rect 13495 5729 13504 5763
rect 13452 5720 13504 5729
rect 14004 5720 14056 5772
rect 19984 5763 20036 5772
rect 10600 5652 10652 5704
rect 10876 5652 10928 5704
rect 8760 5584 8812 5636
rect 11888 5584 11940 5636
rect 12440 5652 12492 5704
rect 14096 5652 14148 5704
rect 14924 5652 14976 5704
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 21088 5720 21140 5772
rect 12808 5584 12860 5636
rect 16304 5584 16356 5636
rect 19340 5652 19392 5704
rect 20168 5652 20220 5704
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 27620 5865 27629 5899
rect 27629 5865 27663 5899
rect 27663 5865 27672 5899
rect 27620 5856 27672 5865
rect 32404 5899 32456 5908
rect 32404 5865 32413 5899
rect 32413 5865 32447 5899
rect 32447 5865 32456 5899
rect 32404 5856 32456 5865
rect 36084 5899 36136 5908
rect 36084 5865 36093 5899
rect 36093 5865 36127 5899
rect 36127 5865 36136 5899
rect 36084 5856 36136 5865
rect 43996 5899 44048 5908
rect 43996 5865 44005 5899
rect 44005 5865 44039 5899
rect 44039 5865 44048 5899
rect 43996 5856 44048 5865
rect 46112 5856 46164 5908
rect 53748 5856 53800 5908
rect 67088 5856 67140 5908
rect 68100 5856 68152 5908
rect 70676 5856 70728 5908
rect 82544 5856 82596 5908
rect 83372 5856 83424 5908
rect 85212 5899 85264 5908
rect 85212 5865 85221 5899
rect 85221 5865 85255 5899
rect 85255 5865 85264 5899
rect 85212 5856 85264 5865
rect 89720 5856 89772 5908
rect 99472 5856 99524 5908
rect 99656 5856 99708 5908
rect 103888 5856 103940 5908
rect 105084 5899 105136 5908
rect 105084 5865 105093 5899
rect 105093 5865 105127 5899
rect 105127 5865 105136 5899
rect 105084 5856 105136 5865
rect 105360 5856 105412 5908
rect 108948 5856 109000 5908
rect 109132 5856 109184 5908
rect 115020 5856 115072 5908
rect 115112 5856 115164 5908
rect 24584 5788 24636 5840
rect 25044 5763 25096 5772
rect 25044 5729 25053 5763
rect 25053 5729 25087 5763
rect 25087 5729 25096 5763
rect 25044 5720 25096 5729
rect 28632 5763 28684 5772
rect 28632 5729 28641 5763
rect 28641 5729 28675 5763
rect 28675 5729 28684 5763
rect 28632 5720 28684 5729
rect 34336 5788 34388 5840
rect 34612 5788 34664 5840
rect 46756 5788 46808 5840
rect 47124 5788 47176 5840
rect 58992 5788 59044 5840
rect 29736 5763 29788 5772
rect 29736 5729 29745 5763
rect 29745 5729 29779 5763
rect 29779 5729 29788 5763
rect 29736 5720 29788 5729
rect 30564 5720 30616 5772
rect 31944 5720 31996 5772
rect 33600 5720 33652 5772
rect 36728 5720 36780 5772
rect 39120 5763 39172 5772
rect 31760 5652 31812 5704
rect 34888 5652 34940 5704
rect 37740 5695 37792 5704
rect 37740 5661 37749 5695
rect 37749 5661 37783 5695
rect 37783 5661 37792 5695
rect 37740 5652 37792 5661
rect 39120 5729 39129 5763
rect 39129 5729 39163 5763
rect 39163 5729 39172 5763
rect 39120 5720 39172 5729
rect 46572 5763 46624 5772
rect 46572 5729 46581 5763
rect 46581 5729 46615 5763
rect 46615 5729 46624 5763
rect 46572 5720 46624 5729
rect 40132 5695 40184 5704
rect 40132 5661 40141 5695
rect 40141 5661 40175 5695
rect 40175 5661 40184 5695
rect 40132 5652 40184 5661
rect 41972 5695 42024 5704
rect 41972 5661 41981 5695
rect 41981 5661 42015 5695
rect 42015 5661 42024 5695
rect 41972 5652 42024 5661
rect 50528 5763 50580 5772
rect 50528 5729 50537 5763
rect 50537 5729 50571 5763
rect 50571 5729 50580 5763
rect 50528 5720 50580 5729
rect 51632 5763 51684 5772
rect 51632 5729 51641 5763
rect 51641 5729 51675 5763
rect 51675 5729 51684 5763
rect 51632 5720 51684 5729
rect 54576 5763 54628 5772
rect 54576 5729 54585 5763
rect 54585 5729 54619 5763
rect 54619 5729 54628 5763
rect 54576 5720 54628 5729
rect 50160 5652 50212 5704
rect 52920 5695 52972 5704
rect 52920 5661 52929 5695
rect 52929 5661 52963 5695
rect 52963 5661 52972 5695
rect 52920 5652 52972 5661
rect 53840 5652 53892 5704
rect 56324 5720 56376 5772
rect 59268 5763 59320 5772
rect 54760 5652 54812 5704
rect 57704 5695 57756 5704
rect 57704 5661 57713 5695
rect 57713 5661 57747 5695
rect 57747 5661 57756 5695
rect 57704 5652 57756 5661
rect 59268 5729 59277 5763
rect 59277 5729 59311 5763
rect 59311 5729 59320 5763
rect 59268 5720 59320 5729
rect 62028 5720 62080 5772
rect 72884 5788 72936 5840
rect 68836 5763 68888 5772
rect 60372 5695 60424 5704
rect 23296 5584 23348 5636
rect 32864 5584 32916 5636
rect 47216 5584 47268 5636
rect 60372 5661 60381 5695
rect 60381 5661 60415 5695
rect 60415 5661 60424 5695
rect 60372 5652 60424 5661
rect 61844 5695 61896 5704
rect 61844 5661 61853 5695
rect 61853 5661 61887 5695
rect 61887 5661 61896 5695
rect 61844 5652 61896 5661
rect 68836 5729 68845 5763
rect 68845 5729 68879 5763
rect 68879 5729 68888 5763
rect 68836 5720 68888 5729
rect 72608 5763 72660 5772
rect 72608 5729 72617 5763
rect 72617 5729 72651 5763
rect 72651 5729 72660 5763
rect 72608 5720 72660 5729
rect 73160 5720 73212 5772
rect 74448 5720 74500 5772
rect 78128 5720 78180 5772
rect 79140 5763 79192 5772
rect 79140 5729 79149 5763
rect 79149 5729 79183 5763
rect 79183 5729 79192 5763
rect 79140 5720 79192 5729
rect 80980 5720 81032 5772
rect 66444 5695 66496 5704
rect 66444 5661 66453 5695
rect 66453 5661 66487 5695
rect 66487 5661 66496 5695
rect 66444 5652 66496 5661
rect 67456 5695 67508 5704
rect 67456 5661 67465 5695
rect 67465 5661 67499 5695
rect 67499 5661 67508 5695
rect 67456 5652 67508 5661
rect 68744 5695 68796 5704
rect 68744 5661 68753 5695
rect 68753 5661 68787 5695
rect 68787 5661 68796 5695
rect 68744 5652 68796 5661
rect 77576 5695 77628 5704
rect 2780 5516 2832 5568
rect 10232 5516 10284 5568
rect 12716 5516 12768 5568
rect 14556 5516 14608 5568
rect 18880 5516 18932 5568
rect 20260 5516 20312 5568
rect 22836 5516 22888 5568
rect 25228 5516 25280 5568
rect 43260 5516 43312 5568
rect 45652 5516 45704 5568
rect 61200 5584 61252 5636
rect 73712 5584 73764 5636
rect 73804 5584 73856 5636
rect 74724 5584 74776 5636
rect 62856 5559 62908 5568
rect 62856 5525 62865 5559
rect 62865 5525 62899 5559
rect 62899 5525 62908 5559
rect 62856 5516 62908 5525
rect 73160 5516 73212 5568
rect 75460 5559 75512 5568
rect 75460 5525 75469 5559
rect 75469 5525 75503 5559
rect 75503 5525 75512 5559
rect 75460 5516 75512 5525
rect 77576 5661 77585 5695
rect 77585 5661 77619 5695
rect 77619 5661 77628 5695
rect 77576 5652 77628 5661
rect 77668 5652 77720 5704
rect 104164 5788 104216 5840
rect 109592 5788 109644 5840
rect 109868 5788 109920 5840
rect 114468 5788 114520 5840
rect 120632 5856 120684 5908
rect 126612 5856 126664 5908
rect 127072 5856 127124 5908
rect 128268 5856 128320 5908
rect 133512 5856 133564 5908
rect 133604 5856 133656 5908
rect 133788 5856 133840 5908
rect 134064 5856 134116 5908
rect 142160 5899 142212 5908
rect 142160 5865 142169 5899
rect 142169 5865 142203 5899
rect 142203 5865 142212 5899
rect 142160 5856 142212 5865
rect 143264 5899 143316 5908
rect 143264 5865 143273 5899
rect 143273 5865 143307 5899
rect 143307 5865 143316 5899
rect 143264 5856 143316 5865
rect 143908 5856 143960 5908
rect 83372 5763 83424 5772
rect 83372 5729 83381 5763
rect 83381 5729 83415 5763
rect 83415 5729 83424 5763
rect 83372 5720 83424 5729
rect 89628 5763 89680 5772
rect 89628 5729 89637 5763
rect 89637 5729 89671 5763
rect 89671 5729 89680 5763
rect 89628 5720 89680 5729
rect 91192 5720 91244 5772
rect 94688 5720 94740 5772
rect 96804 5720 96856 5772
rect 96988 5720 97040 5772
rect 97724 5720 97776 5772
rect 99104 5720 99156 5772
rect 79048 5627 79100 5636
rect 79048 5593 79057 5627
rect 79057 5593 79091 5627
rect 79091 5593 79100 5627
rect 79048 5584 79100 5593
rect 80428 5584 80480 5636
rect 89720 5627 89772 5636
rect 89720 5593 89729 5627
rect 89729 5593 89763 5627
rect 89763 5593 89772 5627
rect 89720 5584 89772 5593
rect 91376 5559 91428 5568
rect 91376 5525 91385 5559
rect 91385 5525 91419 5559
rect 91419 5525 91428 5559
rect 91376 5516 91428 5525
rect 94780 5652 94832 5704
rect 95700 5695 95752 5704
rect 95700 5661 95709 5695
rect 95709 5661 95743 5695
rect 95743 5661 95752 5695
rect 95700 5652 95752 5661
rect 98184 5652 98236 5704
rect 99288 5652 99340 5704
rect 99472 5695 99524 5704
rect 99472 5661 99481 5695
rect 99481 5661 99515 5695
rect 99515 5661 99524 5695
rect 99472 5652 99524 5661
rect 103888 5720 103940 5772
rect 104072 5763 104124 5772
rect 104072 5729 104081 5763
rect 104081 5729 104115 5763
rect 104115 5729 104124 5763
rect 104072 5720 104124 5729
rect 104348 5720 104400 5772
rect 107476 5720 107528 5772
rect 107936 5720 107988 5772
rect 108764 5763 108816 5772
rect 108764 5729 108773 5763
rect 108773 5729 108807 5763
rect 108807 5729 108816 5763
rect 108764 5720 108816 5729
rect 111616 5720 111668 5772
rect 112260 5763 112312 5772
rect 112260 5729 112269 5763
rect 112269 5729 112303 5763
rect 112303 5729 112312 5763
rect 112260 5720 112312 5729
rect 94504 5584 94556 5636
rect 94872 5584 94924 5636
rect 98644 5516 98696 5568
rect 103060 5516 103112 5568
rect 103152 5516 103204 5568
rect 104256 5584 104308 5636
rect 105636 5584 105688 5636
rect 106372 5652 106424 5704
rect 107660 5695 107712 5704
rect 107660 5661 107669 5695
rect 107669 5661 107703 5695
rect 107703 5661 107712 5695
rect 107660 5652 107712 5661
rect 108948 5652 109000 5704
rect 109868 5652 109920 5704
rect 110696 5695 110748 5704
rect 110696 5661 110705 5695
rect 110705 5661 110739 5695
rect 110739 5661 110748 5695
rect 110696 5652 110748 5661
rect 113088 5695 113140 5704
rect 106740 5584 106792 5636
rect 107936 5584 107988 5636
rect 108396 5516 108448 5568
rect 108488 5516 108540 5568
rect 110236 5584 110288 5636
rect 110880 5584 110932 5636
rect 111432 5584 111484 5636
rect 111616 5584 111668 5636
rect 113088 5661 113097 5695
rect 113097 5661 113131 5695
rect 113131 5661 113140 5695
rect 113088 5652 113140 5661
rect 117044 5720 117096 5772
rect 114744 5652 114796 5704
rect 116124 5652 116176 5704
rect 116308 5695 116360 5704
rect 116308 5661 116317 5695
rect 116317 5661 116351 5695
rect 116351 5661 116360 5695
rect 116308 5652 116360 5661
rect 121828 5788 121880 5840
rect 121368 5720 121420 5772
rect 122656 5720 122708 5772
rect 127440 5788 127492 5840
rect 127532 5788 127584 5840
rect 154396 5788 154448 5840
rect 124772 5720 124824 5772
rect 126336 5720 126388 5772
rect 128176 5720 128228 5772
rect 128820 5763 128872 5772
rect 128820 5729 128829 5763
rect 128829 5729 128863 5763
rect 128863 5729 128872 5763
rect 128820 5720 128872 5729
rect 129280 5720 129332 5772
rect 131764 5763 131816 5772
rect 117688 5584 117740 5636
rect 122012 5652 122064 5704
rect 123024 5652 123076 5704
rect 123484 5652 123536 5704
rect 127532 5652 127584 5704
rect 127624 5695 127676 5704
rect 127624 5661 127633 5695
rect 127633 5661 127667 5695
rect 127667 5661 127676 5695
rect 130660 5695 130712 5704
rect 127624 5652 127676 5661
rect 130660 5661 130669 5695
rect 130669 5661 130703 5695
rect 130703 5661 130712 5695
rect 130660 5652 130712 5661
rect 131764 5729 131773 5763
rect 131773 5729 131807 5763
rect 131807 5729 131816 5763
rect 131764 5720 131816 5729
rect 133144 5763 133196 5772
rect 133144 5729 133153 5763
rect 133153 5729 133187 5763
rect 133187 5729 133196 5763
rect 133144 5720 133196 5729
rect 133604 5720 133656 5772
rect 134616 5720 134668 5772
rect 134892 5720 134944 5772
rect 136640 5720 136692 5772
rect 139860 5720 139912 5772
rect 119620 5516 119672 5568
rect 123944 5584 123996 5636
rect 128912 5627 128964 5636
rect 128544 5516 128596 5568
rect 128912 5593 128921 5627
rect 128921 5593 128955 5627
rect 128955 5593 128964 5627
rect 128912 5584 128964 5593
rect 129372 5584 129424 5636
rect 131580 5584 131632 5636
rect 131948 5627 132000 5636
rect 131948 5593 131957 5627
rect 131957 5593 131991 5627
rect 131991 5593 132000 5627
rect 131948 5584 132000 5593
rect 132224 5652 132276 5704
rect 134156 5584 134208 5636
rect 134616 5627 134668 5636
rect 134616 5593 134625 5627
rect 134625 5593 134659 5627
rect 134659 5593 134668 5627
rect 134616 5584 134668 5593
rect 134800 5652 134852 5704
rect 138756 5695 138808 5704
rect 135536 5584 135588 5636
rect 135904 5584 135956 5636
rect 136180 5516 136232 5568
rect 137652 5584 137704 5636
rect 137560 5516 137612 5568
rect 138756 5661 138765 5695
rect 138765 5661 138799 5695
rect 138799 5661 138808 5695
rect 138756 5652 138808 5661
rect 141148 5720 141200 5772
rect 153660 5720 153712 5772
rect 146116 5652 146168 5704
rect 146392 5652 146444 5704
rect 148784 5652 148836 5704
rect 153292 5652 153344 5704
rect 151360 5584 151412 5636
rect 152924 5584 152976 5636
rect 156512 5516 156564 5568
rect 4078 5414 4130 5466
rect 44078 5414 44130 5466
rect 84078 5414 84130 5466
rect 124078 5414 124130 5466
rect 70492 5312 70544 5364
rect 94504 5312 94556 5364
rect 94688 5312 94740 5364
rect 96068 5312 96120 5364
rect 101220 5312 101272 5364
rect 8024 5244 8076 5296
rect 9312 5244 9364 5296
rect 38476 5244 38528 5296
rect 43720 5244 43772 5296
rect 49608 5244 49660 5296
rect 55956 5244 56008 5296
rect 57980 5287 58032 5296
rect 57980 5253 57989 5287
rect 57989 5253 58023 5287
rect 58023 5253 58032 5287
rect 57980 5244 58032 5253
rect 59176 5244 59228 5296
rect 6920 5176 6972 5228
rect 8484 5176 8536 5228
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 15384 5176 15436 5228
rect 20260 5219 20312 5228
rect 20260 5185 20269 5219
rect 20269 5185 20303 5219
rect 20303 5185 20312 5219
rect 20260 5176 20312 5185
rect 20812 5176 20864 5228
rect 22468 5176 22520 5228
rect 30380 5219 30432 5228
rect 30380 5185 30389 5219
rect 30389 5185 30423 5219
rect 30423 5185 30432 5219
rect 30380 5176 30432 5185
rect 31760 5219 31812 5228
rect 31760 5185 31769 5219
rect 31769 5185 31803 5219
rect 31803 5185 31812 5219
rect 31760 5176 31812 5185
rect 32312 5176 32364 5228
rect 34888 5219 34940 5228
rect 34888 5185 34897 5219
rect 34897 5185 34931 5219
rect 34931 5185 34940 5219
rect 34888 5176 34940 5185
rect 40132 5176 40184 5228
rect 47124 5219 47176 5228
rect 47124 5185 47133 5219
rect 47133 5185 47167 5219
rect 47167 5185 47176 5219
rect 47124 5176 47176 5185
rect 48504 5176 48556 5228
rect 52920 5176 52972 5228
rect 53288 5219 53340 5228
rect 53288 5185 53297 5219
rect 53297 5185 53331 5219
rect 53331 5185 53340 5219
rect 53288 5176 53340 5185
rect 59084 5176 59136 5228
rect 62212 5244 62264 5296
rect 66536 5244 66588 5296
rect 72240 5244 72292 5296
rect 7472 5108 7524 5160
rect 7932 5151 7984 5160
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 13360 5108 13412 5160
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 15292 5108 15344 5160
rect 15936 5151 15988 5160
rect 15936 5117 15945 5151
rect 15945 5117 15979 5151
rect 15979 5117 15988 5151
rect 15936 5108 15988 5117
rect 20444 5108 20496 5160
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 23480 5108 23532 5160
rect 23756 5108 23808 5160
rect 29368 5151 29420 5160
rect 29368 5117 29377 5151
rect 29377 5117 29411 5151
rect 29411 5117 29420 5151
rect 29368 5108 29420 5117
rect 30472 5151 30524 5160
rect 30472 5117 30481 5151
rect 30481 5117 30515 5151
rect 30515 5117 30524 5151
rect 30472 5108 30524 5117
rect 32956 5151 33008 5160
rect 32956 5117 32965 5151
rect 32965 5117 32999 5151
rect 32999 5117 33008 5151
rect 32956 5108 33008 5117
rect 36084 5108 36136 5160
rect 41144 5108 41196 5160
rect 42340 5108 42392 5160
rect 44548 5108 44600 5160
rect 46112 5151 46164 5160
rect 46112 5117 46121 5151
rect 46121 5117 46155 5151
rect 46155 5117 46164 5151
rect 46112 5108 46164 5117
rect 47216 5151 47268 5160
rect 47216 5117 47225 5151
rect 47225 5117 47259 5151
rect 47259 5117 47268 5151
rect 47216 5108 47268 5117
rect 53564 5151 53616 5160
rect 53564 5117 53573 5151
rect 53573 5117 53607 5151
rect 53607 5117 53616 5151
rect 53564 5108 53616 5117
rect 54852 5151 54904 5160
rect 54852 5117 54861 5151
rect 54861 5117 54895 5151
rect 54895 5117 54904 5151
rect 54852 5108 54904 5117
rect 55956 5151 56008 5160
rect 55956 5117 55965 5151
rect 55965 5117 55999 5151
rect 55999 5117 56008 5151
rect 55956 5108 56008 5117
rect 47768 5040 47820 5092
rect 58072 5108 58124 5160
rect 61936 5176 61988 5228
rect 63224 5151 63276 5160
rect 59360 5040 59412 5092
rect 63224 5117 63233 5151
rect 63233 5117 63267 5151
rect 63267 5117 63276 5151
rect 63224 5108 63276 5117
rect 63868 5176 63920 5228
rect 70584 5176 70636 5228
rect 70768 5176 70820 5228
rect 66444 5108 66496 5160
rect 67732 5108 67784 5160
rect 69020 5151 69072 5160
rect 69020 5117 69029 5151
rect 69029 5117 69063 5151
rect 69063 5117 69072 5151
rect 69020 5108 69072 5117
rect 69940 5108 69992 5160
rect 70860 5151 70912 5160
rect 70860 5117 70869 5151
rect 70869 5117 70903 5151
rect 70903 5117 70912 5151
rect 70860 5108 70912 5117
rect 77576 5176 77628 5228
rect 72424 5151 72476 5160
rect 71228 5040 71280 5092
rect 7012 4972 7064 5024
rect 10968 4972 11020 5024
rect 51724 4972 51776 5024
rect 67548 4972 67600 5024
rect 67732 4972 67784 5024
rect 72424 5117 72433 5151
rect 72433 5117 72467 5151
rect 72467 5117 72476 5151
rect 72424 5108 72476 5117
rect 72516 5108 72568 5160
rect 74172 5151 74224 5160
rect 74172 5117 74181 5151
rect 74181 5117 74215 5151
rect 74215 5117 74224 5151
rect 74172 5108 74224 5117
rect 74540 5151 74592 5160
rect 74540 5117 74549 5151
rect 74549 5117 74583 5151
rect 74583 5117 74592 5151
rect 74540 5108 74592 5117
rect 74724 5151 74776 5160
rect 74724 5117 74733 5151
rect 74733 5117 74767 5151
rect 74767 5117 74776 5151
rect 74724 5108 74776 5117
rect 77668 5108 77720 5160
rect 78772 5244 78824 5296
rect 81624 5244 81676 5296
rect 89996 5287 90048 5296
rect 89996 5253 90005 5287
rect 90005 5253 90039 5287
rect 90039 5253 90048 5287
rect 89996 5244 90048 5253
rect 79784 5151 79836 5160
rect 79784 5117 79793 5151
rect 79793 5117 79827 5151
rect 79827 5117 79836 5151
rect 79784 5108 79836 5117
rect 80152 5151 80204 5160
rect 80152 5117 80161 5151
rect 80161 5117 80195 5151
rect 80195 5117 80204 5151
rect 80152 5108 80204 5117
rect 118516 5312 118568 5364
rect 118608 5312 118660 5364
rect 119528 5312 119580 5364
rect 81624 5151 81676 5160
rect 81624 5117 81633 5151
rect 81633 5117 81667 5151
rect 81667 5117 81676 5151
rect 81624 5108 81676 5117
rect 82084 5151 82136 5160
rect 82084 5117 82093 5151
rect 82093 5117 82127 5151
rect 82127 5117 82136 5151
rect 82084 5108 82136 5117
rect 86776 5151 86828 5160
rect 86776 5117 86785 5151
rect 86785 5117 86819 5151
rect 86819 5117 86828 5151
rect 86776 5108 86828 5117
rect 88524 5151 88576 5160
rect 88524 5117 88533 5151
rect 88533 5117 88567 5151
rect 88567 5117 88576 5151
rect 88524 5108 88576 5117
rect 90272 5108 90324 5160
rect 91652 5151 91704 5160
rect 91652 5117 91661 5151
rect 91661 5117 91695 5151
rect 91695 5117 91704 5151
rect 91652 5108 91704 5117
rect 92756 5108 92808 5160
rect 93860 5108 93912 5160
rect 96528 5108 96580 5160
rect 96712 5151 96764 5160
rect 96712 5117 96721 5151
rect 96721 5117 96755 5151
rect 96755 5117 96764 5151
rect 98184 5151 98236 5160
rect 96712 5108 96764 5117
rect 98184 5117 98193 5151
rect 98193 5117 98227 5151
rect 98227 5117 98236 5151
rect 98184 5108 98236 5117
rect 99472 5176 99524 5228
rect 105452 5219 105504 5228
rect 105452 5185 105461 5219
rect 105461 5185 105495 5219
rect 105495 5185 105504 5219
rect 105452 5176 105504 5185
rect 106372 5219 106424 5228
rect 106372 5185 106381 5219
rect 106381 5185 106415 5219
rect 106415 5185 106424 5219
rect 106372 5176 106424 5185
rect 106556 5176 106608 5228
rect 111800 5176 111852 5228
rect 113088 5176 113140 5228
rect 102876 5108 102928 5160
rect 105084 5151 105136 5160
rect 105084 5117 105093 5151
rect 105093 5117 105127 5151
rect 105127 5117 105136 5151
rect 105084 5108 105136 5117
rect 105176 5108 105228 5160
rect 106280 5108 106332 5160
rect 108120 5151 108172 5160
rect 72884 5040 72936 5092
rect 108120 5117 108129 5151
rect 108129 5117 108163 5151
rect 108163 5117 108172 5151
rect 108120 5108 108172 5117
rect 108396 5108 108448 5160
rect 110236 5108 110288 5160
rect 110420 5151 110472 5160
rect 110420 5117 110429 5151
rect 110429 5117 110463 5151
rect 110463 5117 110472 5151
rect 110420 5108 110472 5117
rect 110604 5151 110656 5160
rect 110604 5117 110613 5151
rect 110613 5117 110647 5151
rect 110647 5117 110656 5151
rect 110604 5108 110656 5117
rect 110880 5040 110932 5092
rect 111432 5108 111484 5160
rect 112996 5040 113048 5092
rect 113088 5040 113140 5092
rect 114836 5040 114888 5092
rect 77024 4972 77076 5024
rect 81440 4972 81492 5024
rect 88708 4972 88760 5024
rect 94688 4972 94740 5024
rect 95056 4972 95108 5024
rect 96620 4972 96672 5024
rect 106372 4972 106424 5024
rect 106556 4972 106608 5024
rect 113824 4972 113876 5024
rect 116308 5176 116360 5228
rect 123484 5312 123536 5364
rect 123576 5312 123628 5364
rect 124772 5312 124824 5364
rect 122012 5244 122064 5296
rect 124680 5244 124732 5296
rect 129372 5312 129424 5364
rect 129740 5312 129792 5364
rect 131212 5312 131264 5364
rect 131304 5312 131356 5364
rect 138204 5312 138256 5364
rect 126244 5244 126296 5296
rect 118516 5176 118568 5228
rect 128176 5176 128228 5228
rect 131028 5244 131080 5296
rect 131120 5219 131172 5228
rect 115112 5108 115164 5160
rect 117228 5108 117280 5160
rect 118792 5040 118844 5092
rect 123300 5108 123352 5160
rect 124680 5151 124732 5160
rect 123484 5040 123536 5092
rect 124680 5117 124689 5151
rect 124689 5117 124723 5151
rect 124723 5117 124732 5151
rect 124680 5108 124732 5117
rect 126244 5151 126296 5160
rect 126244 5117 126253 5151
rect 126253 5117 126287 5151
rect 126287 5117 126296 5151
rect 126244 5108 126296 5117
rect 128636 5108 128688 5160
rect 130200 5108 130252 5160
rect 131120 5185 131129 5219
rect 131129 5185 131163 5219
rect 131163 5185 131172 5219
rect 131120 5176 131172 5185
rect 130476 5108 130528 5160
rect 137284 5244 137336 5296
rect 144828 5312 144880 5364
rect 145380 5312 145432 5364
rect 155960 5312 156012 5364
rect 149612 5244 149664 5296
rect 131488 5176 131540 5228
rect 132224 5151 132276 5160
rect 132224 5117 132233 5151
rect 132233 5117 132267 5151
rect 132267 5117 132276 5151
rect 132224 5108 132276 5117
rect 132408 5219 132460 5228
rect 132408 5185 132417 5219
rect 132417 5185 132451 5219
rect 132451 5185 132460 5219
rect 132408 5176 132460 5185
rect 132592 5176 132644 5228
rect 133328 5176 133380 5228
rect 133512 5219 133564 5228
rect 133512 5185 133521 5219
rect 133521 5185 133555 5219
rect 133555 5185 133564 5219
rect 133512 5176 133564 5185
rect 133972 5176 134024 5228
rect 135076 5176 135128 5228
rect 135352 5176 135404 5228
rect 136180 5176 136232 5228
rect 137192 5176 137244 5228
rect 137008 5108 137060 5160
rect 137376 5108 137428 5160
rect 137652 5176 137704 5228
rect 142620 5176 142672 5228
rect 143264 5176 143316 5228
rect 144368 5219 144420 5228
rect 144368 5185 144377 5219
rect 144377 5185 144411 5219
rect 144411 5185 144420 5219
rect 144368 5176 144420 5185
rect 121276 4972 121328 5024
rect 121368 4972 121420 5024
rect 123760 4972 123812 5024
rect 126060 4972 126112 5024
rect 126704 4972 126756 5024
rect 128084 4972 128136 5024
rect 131120 5040 131172 5092
rect 131212 5040 131264 5092
rect 136824 5040 136876 5092
rect 143356 5108 143408 5160
rect 138848 5040 138900 5092
rect 132592 4972 132644 5024
rect 132684 4972 132736 5024
rect 133604 4972 133656 5024
rect 133788 4972 133840 5024
rect 134340 4972 134392 5024
rect 134524 5015 134576 5024
rect 134524 4981 134533 5015
rect 134533 4981 134567 5015
rect 134567 4981 134576 5015
rect 134524 4972 134576 4981
rect 134616 4972 134668 5024
rect 140780 4972 140832 5024
rect 144828 5176 144880 5228
rect 146392 5176 146444 5228
rect 153292 5219 153344 5228
rect 153292 5185 153301 5219
rect 153301 5185 153335 5219
rect 153335 5185 153344 5219
rect 153292 5176 153344 5185
rect 156512 5040 156564 5092
rect 144828 4972 144880 5024
rect 24078 4870 24130 4922
rect 64078 4870 64130 4922
rect 104078 4870 104130 4922
rect 144078 4870 144130 4922
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 15292 4811 15344 4820
rect 15292 4777 15301 4811
rect 15301 4777 15335 4811
rect 15335 4777 15344 4811
rect 15292 4768 15344 4777
rect 18052 4768 18104 4820
rect 19340 4811 19392 4820
rect 19340 4777 19349 4811
rect 19349 4777 19383 4811
rect 19383 4777 19392 4811
rect 19340 4768 19392 4777
rect 20444 4768 20496 4820
rect 21272 4768 21324 4820
rect 36084 4811 36136 4820
rect 36084 4777 36093 4811
rect 36093 4777 36127 4811
rect 36127 4777 36136 4811
rect 36084 4768 36136 4777
rect 37740 4811 37792 4820
rect 37740 4777 37749 4811
rect 37749 4777 37783 4811
rect 37783 4777 37792 4811
rect 37740 4768 37792 4777
rect 43628 4768 43680 4820
rect 46112 4768 46164 4820
rect 54852 4768 54904 4820
rect 61660 4768 61712 4820
rect 63224 4768 63276 4820
rect 67456 4768 67508 4820
rect 71320 4768 71372 4820
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 12532 4675 12584 4684
rect 12532 4641 12541 4675
rect 12541 4641 12575 4675
rect 12575 4641 12584 4675
rect 12532 4632 12584 4641
rect 23572 4632 23624 4684
rect 32312 4632 32364 4684
rect 34980 4632 35032 4684
rect 6276 4564 6328 4616
rect 8576 4564 8628 4616
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 13268 4564 13320 4616
rect 23848 4564 23900 4616
rect 26976 4607 27028 4616
rect 20904 4496 20956 4548
rect 26976 4573 26985 4607
rect 26985 4573 27019 4607
rect 27019 4573 27028 4607
rect 26976 4564 27028 4573
rect 28264 4607 28316 4616
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 30564 4564 30616 4616
rect 30748 4607 30800 4616
rect 30748 4573 30757 4607
rect 30757 4573 30791 4607
rect 30791 4573 30800 4607
rect 30748 4564 30800 4573
rect 33508 4564 33560 4616
rect 33692 4607 33744 4616
rect 33692 4573 33701 4607
rect 33701 4573 33735 4607
rect 33735 4573 33744 4607
rect 33692 4564 33744 4573
rect 33784 4564 33836 4616
rect 40776 4607 40828 4616
rect 40776 4573 40785 4607
rect 40785 4573 40819 4607
rect 40819 4573 40828 4607
rect 40776 4564 40828 4573
rect 42064 4607 42116 4616
rect 42064 4573 42073 4607
rect 42073 4573 42107 4607
rect 42107 4573 42116 4607
rect 42064 4564 42116 4573
rect 42800 4632 42852 4684
rect 47308 4632 47360 4684
rect 52736 4700 52788 4752
rect 51724 4675 51776 4684
rect 51724 4641 51733 4675
rect 51733 4641 51767 4675
rect 51767 4641 51776 4675
rect 51724 4632 51776 4641
rect 54760 4632 54812 4684
rect 56232 4675 56284 4684
rect 56232 4641 56241 4675
rect 56241 4641 56275 4675
rect 56275 4641 56284 4675
rect 56232 4632 56284 4641
rect 59544 4632 59596 4684
rect 70492 4675 70544 4684
rect 70492 4641 70501 4675
rect 70501 4641 70535 4675
rect 70535 4641 70544 4675
rect 70492 4632 70544 4641
rect 77392 4700 77444 4752
rect 73068 4632 73120 4684
rect 82912 4768 82964 4820
rect 88524 4768 88576 4820
rect 88708 4811 88760 4820
rect 88708 4777 88717 4811
rect 88717 4777 88751 4811
rect 88751 4777 88760 4811
rect 88708 4768 88760 4777
rect 88984 4768 89036 4820
rect 102600 4768 102652 4820
rect 79968 4700 80020 4752
rect 81072 4675 81124 4684
rect 81072 4641 81081 4675
rect 81081 4641 81115 4675
rect 81115 4641 81124 4675
rect 81072 4632 81124 4641
rect 83924 4675 83976 4684
rect 83924 4641 83933 4675
rect 83933 4641 83967 4675
rect 83967 4641 83976 4675
rect 83924 4632 83976 4641
rect 84384 4675 84436 4684
rect 84384 4641 84393 4675
rect 84393 4641 84427 4675
rect 84427 4641 84436 4675
rect 84384 4632 84436 4641
rect 85580 4675 85632 4684
rect 85580 4641 85589 4675
rect 85589 4641 85623 4675
rect 85623 4641 85632 4675
rect 85580 4632 85632 4641
rect 86408 4632 86460 4684
rect 89260 4632 89312 4684
rect 44364 4564 44416 4616
rect 45100 4607 45152 4616
rect 45100 4573 45109 4607
rect 45109 4573 45143 4607
rect 45143 4573 45152 4607
rect 45100 4564 45152 4573
rect 48136 4564 48188 4616
rect 48964 4607 49016 4616
rect 48964 4573 48973 4607
rect 48973 4573 49007 4607
rect 49007 4573 49016 4607
rect 48964 4564 49016 4573
rect 52000 4564 52052 4616
rect 54208 4564 54260 4616
rect 58072 4607 58124 4616
rect 52368 4496 52420 4548
rect 58072 4573 58081 4607
rect 58081 4573 58115 4607
rect 58115 4573 58124 4607
rect 58072 4564 58124 4573
rect 61200 4607 61252 4616
rect 61200 4573 61209 4607
rect 61209 4573 61243 4607
rect 61243 4573 61252 4607
rect 61200 4564 61252 4573
rect 70308 4607 70360 4616
rect 70308 4573 70317 4607
rect 70317 4573 70351 4607
rect 70351 4573 70360 4607
rect 70308 4564 70360 4573
rect 71412 4607 71464 4616
rect 71412 4573 71421 4607
rect 71421 4573 71455 4607
rect 71455 4573 71464 4607
rect 71412 4564 71464 4573
rect 72884 4607 72936 4616
rect 72884 4573 72893 4607
rect 72893 4573 72927 4607
rect 72927 4573 72936 4607
rect 72884 4564 72936 4573
rect 74632 4564 74684 4616
rect 79508 4607 79560 4616
rect 79508 4573 79517 4607
rect 79517 4573 79551 4607
rect 79551 4573 79560 4607
rect 79508 4564 79560 4573
rect 88984 4564 89036 4616
rect 74724 4471 74776 4480
rect 74724 4437 74733 4471
rect 74733 4437 74767 4471
rect 74767 4437 74776 4471
rect 74724 4428 74776 4437
rect 85672 4428 85724 4480
rect 92020 4675 92072 4684
rect 92020 4641 92029 4675
rect 92029 4641 92063 4675
rect 92063 4641 92072 4675
rect 92020 4632 92072 4641
rect 92112 4632 92164 4684
rect 90456 4607 90508 4616
rect 90456 4573 90465 4607
rect 90465 4573 90499 4607
rect 90499 4573 90508 4607
rect 90456 4564 90508 4573
rect 91928 4607 91980 4616
rect 91928 4573 91937 4607
rect 91937 4573 91971 4607
rect 91971 4573 91980 4607
rect 91928 4564 91980 4573
rect 93032 4564 93084 4616
rect 96712 4632 96764 4684
rect 95792 4607 95844 4616
rect 91836 4496 91888 4548
rect 95792 4573 95801 4607
rect 95801 4573 95835 4607
rect 95835 4573 95844 4607
rect 95792 4564 95844 4573
rect 99288 4700 99340 4752
rect 103612 4700 103664 4752
rect 102140 4632 102192 4684
rect 106096 4768 106148 4820
rect 106188 4768 106240 4820
rect 111248 4768 111300 4820
rect 111432 4811 111484 4820
rect 111432 4777 111441 4811
rect 111441 4777 111475 4811
rect 111475 4777 111484 4811
rect 111432 4768 111484 4777
rect 102508 4607 102560 4616
rect 102508 4573 102517 4607
rect 102517 4573 102551 4607
rect 102551 4573 102560 4607
rect 102508 4564 102560 4573
rect 106556 4700 106608 4752
rect 108028 4700 108080 4752
rect 118608 4768 118660 4820
rect 118884 4768 118936 4820
rect 124956 4768 125008 4820
rect 126244 4768 126296 4820
rect 130936 4768 130988 4820
rect 104900 4632 104952 4684
rect 105360 4675 105412 4684
rect 105360 4641 105369 4675
rect 105369 4641 105403 4675
rect 105403 4641 105412 4675
rect 105360 4632 105412 4641
rect 105636 4675 105688 4684
rect 105636 4641 105645 4675
rect 105645 4641 105679 4675
rect 105679 4641 105688 4675
rect 105636 4632 105688 4641
rect 104164 4564 104216 4616
rect 106188 4632 106240 4684
rect 113824 4700 113876 4752
rect 113088 4632 113140 4684
rect 107936 4564 107988 4616
rect 108856 4564 108908 4616
rect 112444 4607 112496 4616
rect 112444 4573 112453 4607
rect 112453 4573 112487 4607
rect 112487 4573 112496 4607
rect 112444 4564 112496 4573
rect 113640 4632 113692 4684
rect 118424 4632 118476 4684
rect 119804 4632 119856 4684
rect 120172 4632 120224 4684
rect 120540 4632 120592 4684
rect 123852 4675 123904 4684
rect 114744 4564 114796 4616
rect 114928 4564 114980 4616
rect 117136 4607 117188 4616
rect 117136 4573 117145 4607
rect 117145 4573 117179 4607
rect 117179 4573 117188 4607
rect 117136 4564 117188 4573
rect 119344 4564 119396 4616
rect 123852 4641 123861 4675
rect 123861 4641 123895 4675
rect 123895 4641 123904 4675
rect 123852 4632 123904 4641
rect 125048 4675 125100 4684
rect 124128 4607 124180 4616
rect 94320 4496 94372 4548
rect 96528 4496 96580 4548
rect 106188 4496 106240 4548
rect 102416 4428 102468 4480
rect 102600 4428 102652 4480
rect 104164 4428 104216 4480
rect 104348 4428 104400 4480
rect 106004 4428 106056 4480
rect 106556 4496 106608 4548
rect 108028 4428 108080 4480
rect 109132 4428 109184 4480
rect 109316 4496 109368 4548
rect 112260 4496 112312 4548
rect 113548 4496 113600 4548
rect 113824 4428 113876 4480
rect 113916 4428 113968 4480
rect 119620 4496 119672 4548
rect 114744 4428 114796 4480
rect 116952 4428 117004 4480
rect 118332 4428 118384 4480
rect 121644 4496 121696 4548
rect 124128 4573 124137 4607
rect 124137 4573 124171 4607
rect 124171 4573 124180 4607
rect 124128 4564 124180 4573
rect 125048 4641 125057 4675
rect 125057 4641 125091 4675
rect 125091 4641 125100 4675
rect 125048 4632 125100 4641
rect 126152 4675 126204 4684
rect 126152 4641 126161 4675
rect 126161 4641 126195 4675
rect 126195 4641 126204 4675
rect 126152 4632 126204 4641
rect 126336 4700 126388 4752
rect 137560 4768 137612 4820
rect 137652 4768 137704 4820
rect 138756 4811 138808 4820
rect 127992 4632 128044 4684
rect 129924 4675 129976 4684
rect 129924 4641 129933 4675
rect 129933 4641 129967 4675
rect 129967 4641 129976 4675
rect 129924 4632 129976 4641
rect 131672 4632 131724 4684
rect 133512 4632 133564 4684
rect 138296 4700 138348 4752
rect 138756 4777 138765 4811
rect 138765 4777 138799 4811
rect 138799 4777 138808 4811
rect 138756 4768 138808 4777
rect 139676 4700 139728 4752
rect 134340 4632 134392 4684
rect 136088 4675 136140 4684
rect 136088 4641 136097 4675
rect 136097 4641 136131 4675
rect 136131 4641 136140 4675
rect 136088 4632 136140 4641
rect 126336 4496 126388 4548
rect 126520 4539 126572 4548
rect 126520 4505 126529 4539
rect 126529 4505 126563 4539
rect 126563 4505 126572 4539
rect 126520 4496 126572 4505
rect 126796 4564 126848 4616
rect 131304 4564 131356 4616
rect 137376 4607 137428 4616
rect 123392 4428 123444 4480
rect 125232 4428 125284 4480
rect 126796 4428 126848 4480
rect 127900 4496 127952 4548
rect 137376 4573 137385 4607
rect 137385 4573 137419 4607
rect 137419 4573 137428 4607
rect 137376 4564 137428 4573
rect 137560 4632 137612 4684
rect 141056 4768 141108 4820
rect 148324 4768 148376 4820
rect 155500 4768 155552 4820
rect 141608 4675 141660 4684
rect 141608 4641 141617 4675
rect 141617 4641 141651 4675
rect 141651 4641 141660 4675
rect 141608 4632 141660 4641
rect 140044 4607 140096 4616
rect 140044 4573 140053 4607
rect 140053 4573 140087 4607
rect 140087 4573 140096 4607
rect 140044 4564 140096 4573
rect 142436 4607 142488 4616
rect 142436 4573 142445 4607
rect 142445 4573 142479 4607
rect 142479 4573 142488 4607
rect 142436 4564 142488 4573
rect 148324 4564 148376 4616
rect 133512 4496 133564 4548
rect 136364 4496 136416 4548
rect 128636 4428 128688 4480
rect 132040 4428 132092 4480
rect 134708 4428 134760 4480
rect 136180 4428 136232 4480
rect 136640 4496 136692 4548
rect 140688 4496 140740 4548
rect 141516 4539 141568 4548
rect 141516 4505 141525 4539
rect 141525 4505 141559 4539
rect 141559 4505 141568 4539
rect 141516 4496 141568 4505
rect 137744 4428 137796 4480
rect 137836 4428 137888 4480
rect 145380 4428 145432 4480
rect 4078 4326 4130 4378
rect 44078 4326 44130 4378
rect 84078 4326 84130 4378
rect 124078 4326 124130 4378
rect 56232 4224 56284 4276
rect 75920 4224 75972 4276
rect 88892 4224 88944 4276
rect 92112 4224 92164 4276
rect 94504 4224 94556 4276
rect 100208 4224 100260 4276
rect 30288 4156 30340 4208
rect 34336 4156 34388 4208
rect 45008 4156 45060 4208
rect 4160 4088 4212 4140
rect 3608 4020 3660 4072
rect 5540 4088 5592 4140
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 12440 4131 12492 4140
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 12440 4088 12492 4097
rect 5632 3952 5684 4004
rect 9956 4020 10008 4072
rect 11152 4063 11204 4072
rect 11152 4029 11161 4063
rect 11161 4029 11195 4063
rect 11195 4029 11204 4063
rect 11152 4020 11204 4029
rect 19800 4020 19852 4072
rect 9680 3952 9732 4004
rect 11244 3952 11296 4004
rect 3240 3884 3292 3936
rect 6092 3884 6144 3936
rect 23480 4088 23532 4140
rect 25228 4088 25280 4140
rect 26976 4088 27028 4140
rect 29368 4088 29420 4140
rect 30748 4088 30800 4140
rect 33508 4131 33560 4140
rect 33508 4097 33517 4131
rect 33517 4097 33551 4131
rect 33551 4097 33560 4131
rect 33508 4088 33560 4097
rect 40776 4088 40828 4140
rect 41972 4088 42024 4140
rect 44548 4088 44600 4140
rect 46480 4131 46532 4140
rect 46480 4097 46489 4131
rect 46489 4097 46523 4131
rect 46523 4097 46532 4131
rect 46480 4088 46532 4097
rect 55128 4156 55180 4208
rect 48964 4088 49016 4140
rect 52000 4088 52052 4140
rect 22744 4020 22796 4072
rect 22836 4020 22888 4072
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 30196 4020 30248 4072
rect 33416 4020 33468 4072
rect 43352 4063 43404 4072
rect 43352 4029 43361 4063
rect 43361 4029 43395 4063
rect 43395 4029 43404 4063
rect 43352 4020 43404 4029
rect 44732 4020 44784 4072
rect 52828 4063 52880 4072
rect 52828 4029 52837 4063
rect 52837 4029 52871 4063
rect 52871 4029 52880 4063
rect 52828 4020 52880 4029
rect 48964 3952 49016 4004
rect 55220 4063 55272 4072
rect 55220 4029 55229 4063
rect 55229 4029 55263 4063
rect 55263 4029 55272 4063
rect 58072 4088 58124 4140
rect 60648 4131 60700 4140
rect 55220 4020 55272 4029
rect 58256 4063 58308 4072
rect 58256 4029 58265 4063
rect 58265 4029 58299 4063
rect 58299 4029 58308 4063
rect 58256 4020 58308 4029
rect 60648 4097 60657 4131
rect 60657 4097 60691 4131
rect 60691 4097 60700 4131
rect 60648 4088 60700 4097
rect 68836 4156 68888 4208
rect 107660 4224 107712 4276
rect 109684 4224 109736 4276
rect 118516 4224 118568 4276
rect 118608 4224 118660 4276
rect 118884 4224 118936 4276
rect 102416 4156 102468 4208
rect 108304 4156 108356 4208
rect 109132 4156 109184 4208
rect 119896 4224 119948 4276
rect 119988 4224 120040 4276
rect 122472 4224 122524 4276
rect 123484 4224 123536 4276
rect 63684 4088 63736 4140
rect 67548 4088 67600 4140
rect 60464 4063 60516 4072
rect 26884 3884 26936 3936
rect 44640 3884 44692 3936
rect 49424 3884 49476 3936
rect 60464 4029 60473 4063
rect 60473 4029 60507 4063
rect 60507 4029 60516 4063
rect 60464 4020 60516 4029
rect 63316 4020 63368 4072
rect 67732 4020 67784 4072
rect 67916 4020 67968 4072
rect 70400 4088 70452 4140
rect 71780 4088 71832 4140
rect 73804 4088 73856 4140
rect 79508 4088 79560 4140
rect 80060 4088 80112 4140
rect 81624 4088 81676 4140
rect 82268 4088 82320 4140
rect 84292 4088 84344 4140
rect 85580 4088 85632 4140
rect 86132 4088 86184 4140
rect 58992 3952 59044 4004
rect 59360 3952 59412 4004
rect 65524 3952 65576 4004
rect 70952 4020 71004 4072
rect 72976 4020 73028 4072
rect 72608 3952 72660 4004
rect 72884 3952 72936 4004
rect 59636 3884 59688 3936
rect 61200 3884 61252 3936
rect 71964 3884 72016 3936
rect 78772 4020 78824 4072
rect 80336 4020 80388 4072
rect 80888 4020 80940 4072
rect 83832 4020 83884 4072
rect 86040 4020 86092 4072
rect 86868 4020 86920 4072
rect 75920 3952 75972 4004
rect 87236 3952 87288 4004
rect 77392 3884 77444 3936
rect 83740 3884 83792 3936
rect 83832 3884 83884 3936
rect 84108 3884 84160 3936
rect 87788 4020 87840 4072
rect 90456 4088 90508 4140
rect 92572 4088 92624 4140
rect 91100 4020 91152 4072
rect 93400 4020 93452 4072
rect 94320 4020 94372 4072
rect 94780 4088 94832 4140
rect 95608 4088 95660 4140
rect 99196 4088 99248 4140
rect 100116 4088 100168 4140
rect 102508 4088 102560 4140
rect 105544 4131 105596 4140
rect 105544 4097 105553 4131
rect 105553 4097 105587 4131
rect 105587 4097 105596 4131
rect 105544 4088 105596 4097
rect 105728 4088 105780 4140
rect 110696 4088 110748 4140
rect 112444 4088 112496 4140
rect 98552 4020 98604 4072
rect 100760 4063 100812 4072
rect 100760 4029 100769 4063
rect 100769 4029 100803 4063
rect 100803 4029 100812 4063
rect 100760 4020 100812 4029
rect 106740 4063 106792 4072
rect 90824 3952 90876 4004
rect 93768 3952 93820 4004
rect 94136 3952 94188 4004
rect 98644 3952 98696 4004
rect 106740 4029 106749 4063
rect 106749 4029 106783 4063
rect 106783 4029 106792 4063
rect 106740 4020 106792 4029
rect 107752 4020 107804 4072
rect 110420 4063 110472 4072
rect 110420 4029 110429 4063
rect 110429 4029 110463 4063
rect 110463 4029 110472 4063
rect 110420 4020 110472 4029
rect 115940 4088 115992 4140
rect 114928 4020 114980 4072
rect 92756 3884 92808 3936
rect 94688 3884 94740 3936
rect 98920 3884 98972 3936
rect 101496 3884 101548 3936
rect 102140 3884 102192 3936
rect 113364 3884 113416 3936
rect 113456 3884 113508 3936
rect 115940 3952 115992 4004
rect 117136 4088 117188 4140
rect 118148 4088 118200 4140
rect 123116 4156 123168 4208
rect 123300 4156 123352 4208
rect 126520 4224 126572 4276
rect 126336 4156 126388 4208
rect 126428 4156 126480 4208
rect 126888 4156 126940 4208
rect 128452 4199 128504 4208
rect 128452 4165 128461 4199
rect 128461 4165 128495 4199
rect 128495 4165 128504 4199
rect 128452 4156 128504 4165
rect 128636 4156 128688 4208
rect 130384 4156 130436 4208
rect 131120 4224 131172 4276
rect 133972 4224 134024 4276
rect 136088 4224 136140 4276
rect 136548 4224 136600 4276
rect 137836 4224 137888 4276
rect 131580 4156 131632 4208
rect 137192 4156 137244 4208
rect 137284 4156 137336 4208
rect 145656 4224 145708 4276
rect 138204 4156 138256 4208
rect 139124 4156 139176 4208
rect 121552 4088 121604 4140
rect 122012 4088 122064 4140
rect 116676 4020 116728 4072
rect 119344 4020 119396 4072
rect 123392 4020 123444 4072
rect 125876 4020 125928 4072
rect 127164 4063 127216 4072
rect 125692 3952 125744 4004
rect 127164 4029 127173 4063
rect 127173 4029 127207 4063
rect 127207 4029 127216 4063
rect 127164 4020 127216 4029
rect 131028 4088 131080 4140
rect 128176 4020 128228 4072
rect 132500 4088 132552 4140
rect 133696 4088 133748 4140
rect 134248 4131 134300 4140
rect 134248 4097 134257 4131
rect 134257 4097 134291 4131
rect 134291 4097 134300 4131
rect 134248 4088 134300 4097
rect 132040 4063 132092 4072
rect 132040 4029 132049 4063
rect 132049 4029 132083 4063
rect 132083 4029 132092 4063
rect 132040 4020 132092 4029
rect 132408 4020 132460 4072
rect 135720 4088 135772 4140
rect 134616 4020 134668 4072
rect 134984 4020 135036 4072
rect 136548 4088 136600 4140
rect 136640 4088 136692 4140
rect 140044 4088 140096 4140
rect 140596 4156 140648 4208
rect 143540 4156 143592 4208
rect 140872 4088 140924 4140
rect 141516 4131 141568 4140
rect 141516 4097 141525 4131
rect 141525 4097 141559 4131
rect 141559 4097 141568 4131
rect 141516 4088 141568 4097
rect 136824 4020 136876 4072
rect 138112 4020 138164 4072
rect 115296 3884 115348 3936
rect 119528 3884 119580 3936
rect 125968 3884 126020 3936
rect 133696 3952 133748 4004
rect 134248 3952 134300 4004
rect 135444 3952 135496 4004
rect 136548 3952 136600 4004
rect 131580 3884 131632 3936
rect 131672 3884 131724 3936
rect 134340 3884 134392 3936
rect 134708 3884 134760 3936
rect 137376 3884 137428 3936
rect 137744 3952 137796 4004
rect 138664 3952 138716 4004
rect 139124 4020 139176 4072
rect 139216 4063 139268 4072
rect 139216 4029 139225 4063
rect 139225 4029 139259 4063
rect 139259 4029 139268 4063
rect 139216 4020 139268 4029
rect 139400 4020 139452 4072
rect 152372 4020 152424 4072
rect 138940 3884 138992 3936
rect 140320 3884 140372 3936
rect 151728 3884 151780 3936
rect 24078 3782 24130 3834
rect 64078 3782 64130 3834
rect 104078 3782 104130 3834
rect 144078 3782 144130 3834
rect 8300 3680 8352 3732
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 18972 3680 19024 3732
rect 19800 3723 19852 3732
rect 19800 3689 19809 3723
rect 19809 3689 19843 3723
rect 19843 3689 19852 3723
rect 19800 3680 19852 3689
rect 22836 3723 22888 3732
rect 22836 3689 22845 3723
rect 22845 3689 22879 3723
rect 22879 3689 22888 3723
rect 22836 3680 22888 3689
rect 23848 3723 23900 3732
rect 23848 3689 23857 3723
rect 23857 3689 23891 3723
rect 23891 3689 23900 3723
rect 23848 3680 23900 3689
rect 26056 3680 26108 3732
rect 28264 3680 28316 3732
rect 38292 3680 38344 3732
rect 43444 3723 43496 3732
rect 43444 3689 43453 3723
rect 43453 3689 43487 3723
rect 43487 3689 43496 3723
rect 43444 3680 43496 3689
rect 52368 3680 52420 3732
rect 53104 3680 53156 3732
rect 55588 3723 55640 3732
rect 55588 3689 55597 3723
rect 55597 3689 55631 3723
rect 55631 3689 55640 3723
rect 55588 3680 55640 3689
rect 57704 3680 57756 3732
rect 58808 3680 58860 3732
rect 60372 3680 60424 3732
rect 69020 3680 69072 3732
rect 71412 3680 71464 3732
rect 74172 3680 74224 3732
rect 76656 3680 76708 3732
rect 83280 3680 83332 3732
rect 83740 3680 83792 3732
rect 94504 3680 94556 3732
rect 95792 3680 95844 3732
rect 96160 3680 96212 3732
rect 17040 3612 17092 3664
rect 33048 3612 33100 3664
rect 47400 3612 47452 3664
rect 52092 3612 52144 3664
rect 55220 3612 55272 3664
rect 61292 3612 61344 3664
rect 73344 3612 73396 3664
rect 74724 3612 74776 3664
rect 2320 3544 2372 3596
rect 572 3476 624 3528
rect 2780 3408 2832 3460
rect 8392 3544 8444 3596
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 13912 3544 13964 3596
rect 18052 3544 18104 3596
rect 26332 3544 26384 3596
rect 27160 3587 27212 3596
rect 27160 3553 27169 3587
rect 27169 3553 27203 3587
rect 27203 3553 27212 3587
rect 27160 3544 27212 3553
rect 33784 3544 33836 3596
rect 34520 3544 34572 3596
rect 37648 3544 37700 3596
rect 39856 3544 39908 3596
rect 44640 3587 44692 3596
rect 11612 3476 11664 3528
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 33968 3519 34020 3528
rect 33968 3485 33977 3519
rect 33977 3485 34011 3519
rect 34011 3485 34020 3519
rect 33968 3476 34020 3485
rect 41236 3476 41288 3528
rect 44640 3553 44649 3587
rect 44649 3553 44683 3587
rect 44683 3553 44692 3587
rect 44640 3544 44692 3553
rect 46204 3587 46256 3596
rect 46204 3553 46213 3587
rect 46213 3553 46247 3587
rect 46247 3553 46256 3587
rect 46204 3544 46256 3553
rect 46756 3544 46808 3596
rect 45652 3519 45704 3528
rect 45652 3485 45661 3519
rect 45661 3485 45695 3519
rect 45695 3485 45704 3519
rect 45652 3476 45704 3485
rect 47400 3476 47452 3528
rect 53288 3544 53340 3596
rect 61568 3587 61620 3596
rect 61568 3553 61577 3587
rect 61577 3553 61611 3587
rect 61611 3553 61620 3587
rect 61568 3544 61620 3553
rect 66536 3587 66588 3596
rect 66536 3553 66545 3587
rect 66545 3553 66579 3587
rect 66579 3553 66588 3587
rect 66536 3544 66588 3553
rect 72792 3544 72844 3596
rect 74264 3544 74316 3596
rect 74632 3544 74684 3596
rect 60740 3476 60792 3528
rect 67272 3476 67324 3528
rect 72516 3476 72568 3528
rect 97632 3612 97684 3664
rect 74908 3544 74960 3596
rect 75552 3544 75604 3596
rect 77024 3544 77076 3596
rect 79324 3587 79376 3596
rect 75092 3476 75144 3528
rect 75828 3476 75880 3528
rect 77392 3476 77444 3528
rect 79324 3553 79333 3587
rect 79333 3553 79367 3587
rect 79367 3553 79376 3587
rect 79324 3544 79376 3553
rect 80244 3544 80296 3596
rect 82084 3544 82136 3596
rect 83924 3544 83976 3596
rect 84292 3587 84344 3596
rect 84292 3553 84301 3587
rect 84301 3553 84335 3587
rect 84335 3553 84344 3587
rect 84292 3544 84344 3553
rect 80888 3476 80940 3528
rect 81164 3476 81216 3528
rect 83188 3476 83240 3528
rect 86040 3544 86092 3596
rect 89352 3544 89404 3596
rect 91652 3544 91704 3596
rect 93032 3544 93084 3596
rect 88156 3476 88208 3528
rect 91284 3476 91336 3528
rect 11796 3408 11848 3460
rect 26516 3408 26568 3460
rect 29092 3408 29144 3460
rect 34612 3408 34664 3460
rect 41420 3408 41472 3460
rect 59268 3408 59320 3460
rect 92480 3408 92532 3460
rect 40684 3340 40736 3392
rect 45192 3340 45244 3392
rect 53932 3340 53984 3392
rect 57244 3340 57296 3392
rect 72516 3383 72568 3392
rect 72516 3349 72525 3383
rect 72525 3349 72559 3383
rect 72559 3349 72568 3383
rect 72516 3340 72568 3349
rect 84292 3340 84344 3392
rect 86040 3383 86092 3392
rect 86040 3349 86049 3383
rect 86049 3349 86083 3383
rect 86083 3349 86092 3383
rect 86040 3340 86092 3349
rect 91008 3340 91060 3392
rect 94964 3544 95016 3596
rect 97724 3587 97776 3596
rect 97724 3553 97733 3587
rect 97733 3553 97767 3587
rect 97767 3553 97776 3587
rect 97724 3544 97776 3553
rect 99012 3680 99064 3732
rect 103060 3723 103112 3732
rect 103060 3689 103069 3723
rect 103069 3689 103103 3723
rect 103103 3689 103112 3723
rect 103060 3680 103112 3689
rect 104900 3680 104952 3732
rect 105176 3612 105228 3664
rect 99748 3544 99800 3596
rect 108212 3612 108264 3664
rect 107292 3587 107344 3596
rect 107292 3553 107301 3587
rect 107301 3553 107335 3587
rect 107335 3553 107344 3587
rect 107292 3544 107344 3553
rect 109040 3544 109092 3596
rect 97356 3476 97408 3528
rect 103428 3476 103480 3528
rect 106004 3476 106056 3528
rect 94504 3408 94556 3460
rect 97724 3340 97776 3392
rect 101680 3340 101732 3392
rect 104164 3408 104216 3460
rect 109224 3408 109276 3460
rect 105728 3340 105780 3392
rect 106556 3340 106608 3392
rect 107108 3340 107160 3392
rect 110512 3680 110564 3732
rect 115204 3723 115256 3732
rect 115204 3689 115213 3723
rect 115213 3689 115247 3723
rect 115247 3689 115256 3723
rect 115204 3680 115256 3689
rect 115388 3680 115440 3732
rect 117228 3680 117280 3732
rect 122196 3723 122248 3732
rect 122196 3689 122205 3723
rect 122205 3689 122239 3723
rect 122239 3689 122248 3723
rect 122196 3680 122248 3689
rect 111800 3612 111852 3664
rect 109868 3476 109920 3528
rect 116860 3544 116912 3596
rect 112812 3519 112864 3528
rect 112812 3485 112821 3519
rect 112821 3485 112855 3519
rect 112855 3485 112864 3519
rect 112812 3476 112864 3485
rect 113364 3476 113416 3528
rect 116584 3476 116636 3528
rect 117964 3544 118016 3596
rect 118516 3476 118568 3528
rect 122012 3544 122064 3596
rect 122104 3587 122156 3596
rect 122104 3553 122113 3587
rect 122113 3553 122147 3587
rect 122147 3553 122156 3587
rect 122104 3544 122156 3553
rect 123024 3544 123076 3596
rect 126244 3612 126296 3664
rect 128268 3680 128320 3732
rect 128636 3680 128688 3732
rect 131304 3680 131356 3732
rect 132316 3680 132368 3732
rect 132408 3612 132460 3664
rect 133052 3612 133104 3664
rect 137836 3680 137888 3732
rect 138204 3680 138256 3732
rect 140320 3680 140372 3732
rect 140964 3680 141016 3732
rect 145472 3680 145524 3732
rect 150440 3680 150492 3732
rect 133696 3612 133748 3664
rect 137928 3612 137980 3664
rect 138388 3612 138440 3664
rect 138664 3612 138716 3664
rect 139216 3612 139268 3664
rect 139768 3655 139820 3664
rect 139768 3621 139777 3655
rect 139777 3621 139811 3655
rect 139811 3621 139820 3655
rect 139768 3612 139820 3621
rect 125600 3544 125652 3596
rect 125968 3587 126020 3596
rect 125968 3553 125977 3587
rect 125977 3553 126011 3587
rect 126011 3553 126020 3587
rect 125968 3544 126020 3553
rect 126060 3587 126112 3596
rect 126060 3553 126069 3587
rect 126069 3553 126103 3587
rect 126103 3553 126112 3587
rect 126060 3544 126112 3553
rect 127440 3544 127492 3596
rect 128268 3476 128320 3528
rect 129004 3544 129056 3596
rect 130292 3544 130344 3596
rect 131120 3587 131172 3596
rect 131120 3553 131129 3587
rect 131129 3553 131163 3587
rect 131163 3553 131172 3587
rect 131120 3544 131172 3553
rect 133144 3587 133196 3596
rect 133144 3553 133153 3587
rect 133153 3553 133187 3587
rect 133187 3553 133196 3587
rect 133144 3544 133196 3553
rect 133788 3544 133840 3596
rect 134064 3544 134116 3596
rect 134524 3544 134576 3596
rect 136364 3587 136416 3596
rect 136364 3553 136373 3587
rect 136373 3553 136407 3587
rect 136407 3553 136416 3587
rect 136364 3544 136416 3553
rect 137468 3544 137520 3596
rect 141332 3612 141384 3664
rect 141148 3544 141200 3596
rect 142160 3587 142212 3596
rect 142160 3553 142169 3587
rect 142169 3553 142203 3587
rect 142203 3553 142212 3587
rect 142160 3544 142212 3553
rect 142252 3544 142304 3596
rect 128452 3408 128504 3460
rect 116492 3340 116544 3392
rect 118148 3383 118200 3392
rect 118148 3349 118157 3383
rect 118157 3349 118191 3383
rect 118191 3349 118200 3383
rect 118148 3340 118200 3349
rect 118700 3340 118752 3392
rect 119528 3340 119580 3392
rect 120356 3383 120408 3392
rect 120356 3349 120365 3383
rect 120365 3349 120399 3383
rect 120399 3349 120408 3383
rect 120356 3340 120408 3349
rect 124588 3340 124640 3392
rect 125508 3340 125560 3392
rect 125968 3340 126020 3392
rect 126152 3340 126204 3392
rect 130476 3340 130528 3392
rect 131212 3408 131264 3460
rect 131488 3408 131540 3460
rect 136548 3476 136600 3528
rect 137100 3476 137152 3528
rect 137836 3476 137888 3528
rect 134064 3408 134116 3460
rect 137284 3408 137336 3460
rect 137376 3408 137428 3460
rect 138940 3476 138992 3528
rect 144000 3476 144052 3528
rect 131580 3340 131632 3392
rect 131672 3340 131724 3392
rect 133696 3340 133748 3392
rect 133788 3340 133840 3392
rect 134800 3340 134852 3392
rect 135444 3340 135496 3392
rect 137468 3383 137520 3392
rect 137468 3349 137477 3383
rect 137477 3349 137511 3383
rect 137511 3349 137520 3383
rect 137468 3340 137520 3349
rect 144736 3544 144788 3596
rect 144276 3476 144328 3528
rect 147588 3544 147640 3596
rect 144920 3476 144972 3528
rect 145748 3476 145800 3528
rect 151820 3612 151872 3664
rect 156880 3544 156932 3596
rect 151820 3476 151872 3528
rect 157156 3476 157208 3528
rect 197268 3476 197320 3528
rect 198004 3476 198056 3528
rect 146024 3408 146076 3460
rect 138388 3340 138440 3392
rect 138756 3340 138808 3392
rect 138940 3340 138992 3392
rect 144276 3340 144328 3392
rect 144460 3383 144512 3392
rect 144460 3349 144469 3383
rect 144469 3349 144503 3383
rect 144503 3349 144512 3383
rect 144460 3340 144512 3349
rect 144736 3383 144788 3392
rect 144736 3349 144745 3383
rect 144745 3349 144779 3383
rect 144779 3349 144788 3383
rect 144736 3340 144788 3349
rect 144828 3340 144880 3392
rect 152648 3408 152700 3460
rect 149704 3340 149756 3392
rect 4078 3238 4130 3290
rect 44078 3238 44130 3290
rect 84078 3238 84130 3290
rect 124078 3238 124130 3290
rect 7840 3136 7892 3188
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 11428 3179 11480 3188
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 12532 3179 12584 3188
rect 12532 3145 12541 3179
rect 12541 3145 12575 3179
rect 12575 3145 12584 3179
rect 12532 3136 12584 3145
rect 13452 3136 13504 3188
rect 14924 3179 14976 3188
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 19984 3179 20036 3188
rect 19984 3145 19993 3179
rect 19993 3145 20027 3179
rect 20027 3145 20036 3179
rect 19984 3136 20036 3145
rect 21088 3179 21140 3188
rect 21088 3145 21097 3179
rect 21097 3145 21131 3179
rect 21131 3145 21140 3179
rect 21088 3136 21140 3145
rect 27068 3179 27120 3188
rect 1492 2932 1544 2984
rect 14188 3000 14240 3052
rect 204 2864 256 2916
rect 7104 2932 7156 2984
rect 8852 2975 8904 2984
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 9772 2932 9824 2984
rect 11520 2932 11572 2984
rect 1860 2796 1912 2848
rect 11060 2796 11112 2848
rect 12348 2864 12400 2916
rect 14556 2932 14608 2984
rect 18420 2932 18472 2984
rect 25412 3068 25464 3120
rect 27068 3145 27077 3179
rect 27077 3145 27111 3179
rect 27111 3145 27120 3179
rect 27068 3136 27120 3145
rect 29552 3136 29604 3188
rect 32588 3136 32640 3188
rect 33600 3136 33652 3188
rect 41328 3136 41380 3188
rect 43076 3136 43128 3188
rect 43812 3179 43864 3188
rect 43812 3145 43821 3179
rect 43821 3145 43855 3179
rect 43855 3145 43864 3179
rect 43812 3136 43864 3145
rect 47216 3136 47268 3188
rect 49148 3136 49200 3188
rect 52828 3136 52880 3188
rect 53564 3179 53616 3188
rect 53564 3145 53573 3179
rect 53573 3145 53607 3179
rect 53607 3145 53616 3179
rect 53564 3136 53616 3145
rect 55956 3136 56008 3188
rect 59084 3136 59136 3188
rect 92480 3136 92532 3188
rect 95240 3136 95292 3188
rect 96804 3136 96856 3188
rect 104164 3136 104216 3188
rect 104532 3136 104584 3188
rect 109132 3136 109184 3188
rect 111064 3179 111116 3188
rect 111064 3145 111073 3179
rect 111073 3145 111107 3179
rect 111107 3145 111116 3179
rect 111064 3136 111116 3145
rect 26516 3000 26568 3052
rect 19340 2864 19392 2916
rect 25872 2932 25924 2984
rect 22744 2864 22796 2916
rect 15200 2796 15252 2848
rect 29828 3068 29880 3120
rect 37188 3068 37240 3120
rect 43444 3068 43496 3120
rect 26700 3000 26752 3052
rect 31576 3000 31628 3052
rect 33140 2932 33192 2984
rect 29368 2864 29420 2916
rect 31116 2864 31168 2916
rect 35440 3000 35492 3052
rect 36360 3000 36412 3052
rect 43076 3000 43128 3052
rect 45100 3000 45152 3052
rect 45192 3000 45244 3052
rect 47492 3000 47544 3052
rect 37740 2864 37792 2916
rect 33048 2796 33100 2848
rect 38476 2932 38528 2984
rect 39488 2864 39540 2916
rect 42432 2864 42484 2916
rect 45008 2932 45060 2984
rect 62856 3068 62908 3120
rect 87236 3068 87288 3120
rect 99196 3068 99248 3120
rect 99288 3068 99340 3120
rect 53932 3000 53984 3052
rect 54024 3000 54076 3052
rect 58072 3000 58124 3052
rect 60280 3000 60332 3052
rect 41604 2796 41656 2848
rect 41972 2796 42024 2848
rect 42800 2796 42852 2848
rect 43720 2796 43772 2848
rect 44180 2796 44232 2848
rect 45652 2796 45704 2848
rect 45928 2864 45980 2916
rect 49884 2796 49936 2848
rect 51540 2864 51592 2916
rect 54208 2932 54260 2984
rect 55036 2932 55088 2984
rect 58440 2932 58492 2984
rect 63040 2975 63092 2984
rect 63040 2941 63049 2975
rect 63049 2941 63083 2975
rect 63083 2941 63092 2975
rect 63040 2932 63092 2941
rect 64512 2932 64564 2984
rect 66996 2975 67048 2984
rect 66996 2941 67005 2975
rect 67005 2941 67039 2975
rect 67039 2941 67048 2975
rect 66996 2932 67048 2941
rect 73252 3000 73304 3052
rect 74448 3000 74500 3052
rect 79784 3000 79836 3052
rect 81348 3043 81400 3052
rect 81348 3009 81357 3043
rect 81357 3009 81391 3043
rect 81391 3009 81400 3043
rect 81348 3000 81400 3009
rect 87144 3043 87196 3052
rect 87144 3009 87153 3043
rect 87153 3009 87187 3043
rect 87187 3009 87196 3043
rect 87144 3000 87196 3009
rect 89812 3000 89864 3052
rect 99472 3000 99524 3052
rect 70860 2975 70912 2984
rect 70860 2941 70869 2975
rect 70869 2941 70903 2975
rect 70903 2941 70912 2975
rect 70860 2932 70912 2941
rect 72700 2975 72752 2984
rect 72700 2941 72709 2975
rect 72709 2941 72743 2975
rect 72743 2941 72752 2975
rect 72700 2932 72752 2941
rect 76196 2975 76248 2984
rect 76196 2941 76205 2975
rect 76205 2941 76239 2975
rect 76239 2941 76248 2975
rect 76196 2932 76248 2941
rect 77944 2932 77996 2984
rect 80428 2975 80480 2984
rect 80428 2941 80437 2975
rect 80437 2941 80471 2975
rect 80471 2941 80480 2975
rect 80428 2932 80480 2941
rect 80612 2932 80664 2984
rect 85764 2975 85816 2984
rect 85764 2941 85773 2975
rect 85773 2941 85807 2975
rect 85807 2941 85816 2975
rect 85764 2932 85816 2941
rect 87328 2932 87380 2984
rect 91468 2975 91520 2984
rect 91468 2941 91477 2975
rect 91477 2941 91511 2975
rect 91511 2941 91520 2975
rect 91468 2932 91520 2941
rect 93584 2975 93636 2984
rect 93584 2941 93593 2975
rect 93593 2941 93627 2975
rect 93627 2941 93636 2975
rect 93584 2932 93636 2941
rect 94596 2975 94648 2984
rect 94596 2941 94605 2975
rect 94605 2941 94639 2975
rect 94639 2941 94648 2975
rect 94596 2932 94648 2941
rect 95884 2932 95936 2984
rect 98828 2975 98880 2984
rect 52552 2864 52604 2916
rect 54668 2864 54720 2916
rect 58532 2864 58584 2916
rect 61568 2864 61620 2916
rect 66352 2907 66404 2916
rect 66352 2873 66361 2907
rect 66361 2873 66395 2907
rect 66395 2873 66404 2907
rect 66352 2864 66404 2873
rect 68560 2907 68612 2916
rect 68560 2873 68569 2907
rect 68569 2873 68603 2907
rect 68603 2873 68612 2907
rect 68560 2864 68612 2873
rect 69020 2864 69072 2916
rect 71596 2864 71648 2916
rect 74632 2864 74684 2916
rect 76840 2864 76892 2916
rect 80796 2864 80848 2916
rect 82912 2864 82964 2916
rect 85120 2864 85172 2916
rect 89444 2864 89496 2916
rect 94320 2864 94372 2916
rect 96896 2864 96948 2916
rect 53472 2796 53524 2848
rect 53564 2796 53616 2848
rect 56784 2796 56836 2848
rect 90916 2796 90968 2848
rect 98828 2941 98837 2975
rect 98837 2941 98871 2975
rect 98871 2941 98880 2975
rect 98828 2932 98880 2941
rect 101220 3000 101272 3052
rect 100576 2975 100628 2984
rect 100576 2941 100585 2975
rect 100585 2941 100619 2975
rect 100619 2941 100628 2975
rect 100576 2932 100628 2941
rect 102968 2932 103020 2984
rect 103152 2975 103204 2984
rect 103152 2941 103161 2975
rect 103161 2941 103195 2975
rect 103195 2941 103204 2975
rect 103152 2932 103204 2941
rect 100392 2864 100444 2916
rect 102140 2864 102192 2916
rect 104256 3068 104308 3120
rect 108120 3068 108172 3120
rect 108028 3000 108080 3052
rect 106924 2932 106976 2984
rect 111432 3068 111484 3120
rect 109224 2932 109276 2984
rect 109776 2975 109828 2984
rect 107108 2864 107160 2916
rect 108304 2864 108356 2916
rect 109776 2941 109785 2975
rect 109785 2941 109819 2975
rect 109819 2941 109828 2975
rect 109776 2932 109828 2941
rect 116308 3136 116360 3188
rect 116400 3136 116452 3188
rect 116584 3136 116636 3188
rect 117964 3136 118016 3188
rect 123300 3136 123352 3188
rect 123944 3136 123996 3188
rect 126244 3136 126296 3188
rect 126336 3136 126388 3188
rect 128268 3136 128320 3188
rect 128728 3179 128780 3188
rect 128728 3145 128737 3179
rect 128737 3145 128771 3179
rect 128771 3145 128780 3179
rect 128728 3136 128780 3145
rect 129096 3136 129148 3188
rect 129280 3136 129332 3188
rect 130108 3136 130160 3188
rect 130844 3136 130896 3188
rect 117504 3068 117556 3120
rect 118792 3068 118844 3120
rect 121644 3111 121696 3120
rect 112076 3043 112128 3052
rect 112076 3009 112085 3043
rect 112085 3009 112119 3043
rect 112119 3009 112128 3043
rect 113824 3043 113876 3052
rect 112076 3000 112128 3009
rect 113824 3009 113833 3043
rect 113833 3009 113867 3043
rect 113867 3009 113876 3043
rect 113824 3000 113876 3009
rect 118608 3000 118660 3052
rect 120356 3000 120408 3052
rect 121644 3077 121653 3111
rect 121653 3077 121687 3111
rect 121687 3077 121696 3111
rect 121644 3068 121696 3077
rect 123576 3043 123628 3052
rect 123576 3009 123585 3043
rect 123585 3009 123619 3043
rect 123619 3009 123628 3043
rect 123576 3000 123628 3009
rect 100668 2796 100720 2848
rect 103888 2796 103940 2848
rect 106924 2796 106976 2848
rect 112996 2864 113048 2916
rect 113548 2907 113600 2916
rect 113548 2873 113557 2907
rect 113557 2873 113591 2907
rect 113591 2873 113600 2907
rect 113548 2864 113600 2873
rect 116860 2864 116912 2916
rect 117320 2864 117372 2916
rect 119344 2932 119396 2984
rect 120540 2975 120592 2984
rect 120172 2864 120224 2916
rect 109500 2796 109552 2848
rect 111248 2796 111300 2848
rect 111432 2796 111484 2848
rect 116308 2796 116360 2848
rect 116952 2796 117004 2848
rect 120540 2941 120549 2975
rect 120549 2941 120583 2975
rect 120583 2941 120592 2975
rect 120540 2932 120592 2941
rect 126060 3068 126112 3120
rect 127900 3111 127952 3120
rect 127900 3077 127909 3111
rect 127909 3077 127943 3111
rect 127943 3077 127952 3111
rect 127900 3068 127952 3077
rect 125600 3000 125652 3052
rect 126428 3043 126480 3052
rect 126428 3009 126437 3043
rect 126437 3009 126471 3043
rect 126471 3009 126480 3043
rect 126428 3000 126480 3009
rect 125324 2864 125376 2916
rect 126980 2932 127032 2984
rect 126888 2864 126940 2916
rect 128636 2932 128688 2984
rect 130660 3068 130712 3120
rect 134708 3136 134760 3188
rect 135076 3136 135128 3188
rect 135628 3136 135680 3188
rect 132500 3068 132552 3120
rect 129280 3000 129332 3052
rect 129648 2932 129700 2984
rect 129924 2932 129976 2984
rect 121552 2796 121604 2848
rect 123300 2796 123352 2848
rect 125140 2796 125192 2848
rect 125416 2796 125468 2848
rect 128452 2864 128504 2916
rect 130844 2864 130896 2916
rect 131120 3000 131172 3052
rect 133604 3000 133656 3052
rect 136272 3068 136324 3120
rect 137008 3068 137060 3120
rect 137928 3068 137980 3120
rect 138112 3136 138164 3188
rect 138756 3136 138808 3188
rect 141700 3136 141752 3188
rect 142160 3136 142212 3188
rect 144828 3068 144880 3120
rect 145564 3068 145616 3120
rect 146116 3068 146168 3120
rect 147128 3068 147180 3120
rect 147588 3068 147640 3120
rect 151360 3068 151412 3120
rect 156696 3068 156748 3120
rect 156972 3068 157024 3120
rect 134064 3000 134116 3052
rect 131212 2975 131264 2984
rect 131212 2941 131221 2975
rect 131221 2941 131255 2975
rect 131255 2941 131264 2975
rect 131212 2932 131264 2941
rect 133880 2932 133932 2984
rect 134432 2932 134484 2984
rect 135904 2975 135956 2984
rect 135904 2941 135913 2975
rect 135913 2941 135947 2975
rect 135947 2941 135956 2975
rect 135904 2932 135956 2941
rect 135996 2975 136048 2984
rect 135996 2941 136005 2975
rect 136005 2941 136039 2975
rect 136039 2941 136048 2975
rect 135996 2932 136048 2941
rect 137008 2864 137060 2916
rect 137192 3043 137244 3052
rect 137192 3009 137201 3043
rect 137201 3009 137235 3043
rect 137235 3009 137244 3043
rect 137192 3000 137244 3009
rect 138020 3000 138072 3052
rect 138204 2932 138256 2984
rect 143724 2932 143776 2984
rect 145196 2932 145248 2984
rect 145288 2932 145340 2984
rect 148324 2932 148376 2984
rect 151452 2932 151504 2984
rect 151544 2932 151596 2984
rect 156420 2932 156472 2984
rect 128544 2796 128596 2848
rect 138664 2864 138716 2916
rect 144368 2864 144420 2916
rect 144552 2864 144604 2916
rect 137928 2796 137980 2848
rect 138480 2796 138532 2848
rect 138572 2796 138624 2848
rect 140412 2839 140464 2848
rect 140412 2805 140421 2839
rect 140421 2805 140455 2839
rect 140455 2805 140464 2839
rect 140412 2796 140464 2805
rect 141056 2796 141108 2848
rect 141792 2796 141844 2848
rect 144460 2796 144512 2848
rect 146116 2864 146168 2916
rect 156144 2864 156196 2916
rect 161204 2932 161256 2984
rect 162676 2932 162728 2984
rect 162768 2932 162820 2984
rect 166724 2932 166776 2984
rect 147036 2796 147088 2848
rect 149244 2796 149296 2848
rect 157432 2796 157484 2848
rect 158352 2796 158404 2848
rect 158536 2796 158588 2848
rect 161480 2796 161532 2848
rect 166264 2864 166316 2916
rect 173808 2932 173860 2984
rect 180156 2932 180208 2984
rect 180340 2932 180392 2984
rect 187056 2932 187108 2984
rect 193588 2932 193640 2984
rect 196900 2932 196952 2984
rect 171784 2864 171836 2916
rect 176476 2864 176528 2916
rect 176660 2864 176712 2916
rect 180432 2864 180484 2916
rect 184204 2864 184256 2916
rect 195888 2864 195940 2916
rect 199752 2864 199804 2916
rect 165068 2796 165120 2848
rect 165344 2796 165396 2848
rect 167092 2796 167144 2848
rect 173348 2796 173400 2848
rect 179236 2796 179288 2848
rect 190460 2796 190512 2848
rect 192300 2796 192352 2848
rect 194692 2796 194744 2848
rect 199292 2796 199344 2848
rect 24078 2694 24130 2746
rect 64078 2694 64130 2746
rect 104078 2694 104130 2746
rect 144078 2694 144130 2746
rect 184078 2694 184130 2746
rect 6460 2592 6512 2644
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 8668 2592 8720 2644
rect 11704 2592 11756 2644
rect 13912 2635 13964 2644
rect 13912 2601 13921 2635
rect 13921 2601 13955 2635
rect 13955 2601 13964 2635
rect 13912 2592 13964 2601
rect 15936 2592 15988 2644
rect 17224 2635 17276 2644
rect 17224 2601 17233 2635
rect 17233 2601 17267 2635
rect 17267 2601 17276 2635
rect 17224 2592 17276 2601
rect 20720 2592 20772 2644
rect 22376 2592 22428 2644
rect 24860 2592 24912 2644
rect 25136 2635 25188 2644
rect 25136 2601 25145 2635
rect 25145 2601 25179 2635
rect 25179 2601 25188 2635
rect 25136 2592 25188 2601
rect 27712 2592 27764 2644
rect 33324 2635 33376 2644
rect 33324 2601 33333 2635
rect 33333 2601 33367 2635
rect 33367 2601 33376 2635
rect 33324 2592 33376 2601
rect 36544 2592 36596 2644
rect 43352 2592 43404 2644
rect 44364 2592 44416 2644
rect 45560 2592 45612 2644
rect 46572 2592 46624 2644
rect 47768 2635 47820 2644
rect 47768 2601 47777 2635
rect 47777 2601 47811 2635
rect 47811 2601 47820 2635
rect 47768 2592 47820 2601
rect 51632 2592 51684 2644
rect 51816 2635 51868 2644
rect 51816 2601 51825 2635
rect 51825 2601 51859 2635
rect 51859 2601 51868 2635
rect 51816 2592 51868 2601
rect 52736 2592 52788 2644
rect 54760 2635 54812 2644
rect 54760 2601 54769 2635
rect 54769 2601 54803 2635
rect 54803 2601 54812 2635
rect 54760 2592 54812 2601
rect 55220 2592 55272 2644
rect 55680 2592 55732 2644
rect 59452 2592 59504 2644
rect 75276 2592 75328 2644
rect 83096 2592 83148 2644
rect 88340 2592 88392 2644
rect 92940 2592 92992 2644
rect 34520 2524 34572 2576
rect 47584 2524 47636 2576
rect 62028 2524 62080 2576
rect 69664 2524 69716 2576
rect 85948 2524 86000 2576
rect 1032 2456 1084 2508
rect 5816 2456 5868 2508
rect 6736 2456 6788 2508
rect 8024 2456 8076 2508
rect 10600 2456 10652 2508
rect 12808 2456 12860 2508
rect 13636 2388 13688 2440
rect 12992 2320 13044 2372
rect 15016 2320 15068 2372
rect 17224 2456 17276 2508
rect 20168 2388 20220 2440
rect 23296 2456 23348 2508
rect 24216 2456 24268 2508
rect 25136 2456 25188 2508
rect 28448 2456 28500 2508
rect 33692 2456 33744 2508
rect 34152 2388 34204 2440
rect 43260 2456 43312 2508
rect 45652 2499 45704 2508
rect 38936 2388 38988 2440
rect 40224 2320 40276 2372
rect 45652 2465 45661 2499
rect 45661 2465 45695 2499
rect 45695 2465 45704 2499
rect 45652 2456 45704 2465
rect 45468 2388 45520 2440
rect 48136 2456 48188 2508
rect 48504 2456 48556 2508
rect 54668 2499 54720 2508
rect 49792 2388 49844 2440
rect 50252 2320 50304 2372
rect 54668 2465 54677 2499
rect 54677 2465 54711 2499
rect 54711 2465 54720 2499
rect 54668 2456 54720 2465
rect 55496 2456 55548 2508
rect 57980 2456 58032 2508
rect 60556 2456 60608 2508
rect 63408 2499 63460 2508
rect 63408 2465 63417 2499
rect 63417 2465 63451 2499
rect 63451 2465 63460 2499
rect 63408 2456 63460 2465
rect 67640 2456 67692 2508
rect 68744 2456 68796 2508
rect 71504 2456 71556 2508
rect 73160 2456 73212 2508
rect 74540 2456 74592 2508
rect 77300 2499 77352 2508
rect 77300 2465 77309 2499
rect 77309 2465 77343 2499
rect 77343 2465 77352 2499
rect 77300 2456 77352 2465
rect 78496 2456 78548 2508
rect 80704 2499 80756 2508
rect 80704 2465 80713 2499
rect 80713 2465 80747 2499
rect 80747 2465 80756 2499
rect 80704 2456 80756 2465
rect 81532 2456 81584 2508
rect 85304 2456 85356 2508
rect 89628 2524 89680 2576
rect 90088 2456 90140 2508
rect 95056 2524 95108 2576
rect 95884 2524 95936 2576
rect 96344 2524 96396 2576
rect 99932 2524 99984 2576
rect 110420 2592 110472 2644
rect 110512 2592 110564 2644
rect 114192 2635 114244 2644
rect 104256 2524 104308 2576
rect 105544 2524 105596 2576
rect 109500 2524 109552 2576
rect 94872 2499 94924 2508
rect 56324 2388 56376 2440
rect 57336 2388 57388 2440
rect 62212 2388 62264 2440
rect 64604 2388 64656 2440
rect 66812 2388 66864 2440
rect 68100 2388 68152 2440
rect 71228 2388 71280 2440
rect 72148 2388 72200 2440
rect 76012 2388 76064 2440
rect 78588 2388 78640 2440
rect 79508 2388 79560 2440
rect 82544 2388 82596 2440
rect 88616 2388 88668 2440
rect 89076 2388 89128 2440
rect 89720 2388 89772 2440
rect 94872 2465 94881 2499
rect 94881 2465 94915 2499
rect 94915 2465 94924 2499
rect 94872 2456 94924 2465
rect 97264 2499 97316 2508
rect 97264 2465 97273 2499
rect 97273 2465 97307 2499
rect 97307 2465 97316 2499
rect 97264 2456 97316 2465
rect 98092 2456 98144 2508
rect 92572 2388 92624 2440
rect 92756 2388 92808 2440
rect 60464 2320 60516 2372
rect 94504 2320 94556 2372
rect 95240 2388 95292 2440
rect 97908 2320 97960 2372
rect 54852 2252 54904 2304
rect 56600 2252 56652 2304
rect 59452 2252 59504 2304
rect 63316 2252 63368 2304
rect 81072 2252 81124 2304
rect 98276 2252 98328 2304
rect 99104 2388 99156 2440
rect 102600 2388 102652 2440
rect 103520 2456 103572 2508
rect 104348 2388 104400 2440
rect 106464 2456 106516 2508
rect 111892 2524 111944 2576
rect 114192 2601 114201 2635
rect 114201 2601 114235 2635
rect 114235 2601 114244 2635
rect 114192 2592 114244 2601
rect 118240 2635 118292 2644
rect 118240 2601 118249 2635
rect 118249 2601 118283 2635
rect 118283 2601 118292 2635
rect 118240 2592 118292 2601
rect 118976 2592 119028 2644
rect 123668 2592 123720 2644
rect 115204 2567 115256 2576
rect 115204 2533 115213 2567
rect 115213 2533 115247 2567
rect 115247 2533 115256 2567
rect 115204 2524 115256 2533
rect 110604 2456 110656 2508
rect 108672 2388 108724 2440
rect 108856 2388 108908 2440
rect 109040 2320 109092 2372
rect 109224 2388 109276 2440
rect 110052 2388 110104 2440
rect 112352 2431 112404 2440
rect 112352 2397 112361 2431
rect 112361 2397 112395 2431
rect 112395 2397 112404 2431
rect 112352 2388 112404 2397
rect 113824 2388 113876 2440
rect 116860 2456 116912 2508
rect 117136 2499 117188 2508
rect 117136 2465 117145 2499
rect 117145 2465 117179 2499
rect 117179 2465 117188 2499
rect 117136 2456 117188 2465
rect 117872 2456 117924 2508
rect 118148 2499 118200 2508
rect 118148 2465 118157 2499
rect 118157 2465 118191 2499
rect 118191 2465 118200 2499
rect 118148 2456 118200 2465
rect 120172 2499 120224 2508
rect 120172 2465 120181 2499
rect 120181 2465 120215 2499
rect 120215 2465 120224 2499
rect 120172 2456 120224 2465
rect 124312 2524 124364 2576
rect 125600 2592 125652 2644
rect 125784 2635 125836 2644
rect 125784 2601 125793 2635
rect 125793 2601 125827 2635
rect 125827 2601 125836 2635
rect 125784 2592 125836 2601
rect 126980 2592 127032 2644
rect 129556 2592 129608 2644
rect 129924 2592 129976 2644
rect 131672 2592 131724 2644
rect 132132 2592 132184 2644
rect 132592 2592 132644 2644
rect 133788 2592 133840 2644
rect 124680 2499 124732 2508
rect 124680 2465 124689 2499
rect 124689 2465 124723 2499
rect 124723 2465 124732 2499
rect 124680 2456 124732 2465
rect 125692 2499 125744 2508
rect 125692 2465 125701 2499
rect 125701 2465 125735 2499
rect 125735 2465 125744 2499
rect 125692 2456 125744 2465
rect 128176 2524 128228 2576
rect 132224 2524 132276 2576
rect 132316 2524 132368 2576
rect 134800 2592 134852 2644
rect 138664 2592 138716 2644
rect 138756 2592 138808 2644
rect 139676 2592 139728 2644
rect 139860 2635 139912 2644
rect 139860 2601 139869 2635
rect 139869 2601 139903 2635
rect 139903 2601 139912 2635
rect 139860 2592 139912 2601
rect 139952 2592 140004 2644
rect 144184 2592 144236 2644
rect 144552 2592 144604 2644
rect 147956 2592 148008 2644
rect 128452 2456 128504 2508
rect 129372 2456 129424 2508
rect 129556 2499 129608 2508
rect 129556 2465 129565 2499
rect 129565 2465 129599 2499
rect 129599 2465 129608 2499
rect 129556 2456 129608 2465
rect 130936 2456 130988 2508
rect 131856 2499 131908 2508
rect 131856 2465 131865 2499
rect 131865 2465 131899 2499
rect 131899 2465 131908 2499
rect 131856 2456 131908 2465
rect 133512 2456 133564 2508
rect 134064 2456 134116 2508
rect 135812 2456 135864 2508
rect 100116 2252 100168 2304
rect 107292 2252 107344 2304
rect 107384 2252 107436 2304
rect 109316 2252 109368 2304
rect 110420 2252 110472 2304
rect 111248 2252 111300 2304
rect 111432 2320 111484 2372
rect 116216 2252 116268 2304
rect 116308 2252 116360 2304
rect 118240 2252 118292 2304
rect 118332 2252 118384 2304
rect 120172 2252 120224 2304
rect 125140 2320 125192 2372
rect 127348 2320 127400 2372
rect 127440 2320 127492 2372
rect 128084 2388 128136 2440
rect 130200 2388 130252 2440
rect 133420 2388 133472 2440
rect 134616 2388 134668 2440
rect 135628 2388 135680 2440
rect 129280 2320 129332 2372
rect 130384 2320 130436 2372
rect 135536 2320 135588 2372
rect 135812 2363 135864 2372
rect 135812 2329 135821 2363
rect 135821 2329 135855 2363
rect 135855 2329 135864 2363
rect 135812 2320 135864 2329
rect 136180 2456 136232 2508
rect 137836 2456 137888 2508
rect 138020 2456 138072 2508
rect 138388 2456 138440 2508
rect 136640 2320 136692 2372
rect 137744 2388 137796 2440
rect 140320 2456 140372 2508
rect 144552 2499 144604 2508
rect 144552 2465 144561 2499
rect 144561 2465 144595 2499
rect 144595 2465 144604 2499
rect 144552 2456 144604 2465
rect 145748 2524 145800 2576
rect 150256 2524 150308 2576
rect 157892 2524 157944 2576
rect 157984 2524 158036 2576
rect 162032 2524 162084 2576
rect 162492 2592 162544 2644
rect 164332 2592 164384 2644
rect 165528 2592 165580 2644
rect 171140 2592 171192 2644
rect 171692 2592 171744 2644
rect 163044 2524 163096 2576
rect 129556 2252 129608 2304
rect 129740 2252 129792 2304
rect 129832 2252 129884 2304
rect 130752 2252 130804 2304
rect 131028 2252 131080 2304
rect 137192 2252 137244 2304
rect 138204 2320 138256 2372
rect 146116 2388 146168 2440
rect 146668 2456 146720 2508
rect 155316 2456 155368 2508
rect 155408 2456 155460 2508
rect 156052 2456 156104 2508
rect 157064 2499 157116 2508
rect 157064 2465 157073 2499
rect 157073 2465 157107 2499
rect 157107 2465 157116 2499
rect 157064 2456 157116 2465
rect 157156 2456 157208 2508
rect 157524 2456 157576 2508
rect 147404 2388 147456 2440
rect 149060 2388 149112 2440
rect 158260 2456 158312 2508
rect 161020 2456 161072 2508
rect 137652 2252 137704 2304
rect 139492 2252 139544 2304
rect 144460 2320 144512 2372
rect 144644 2320 144696 2372
rect 145012 2320 145064 2372
rect 153660 2320 153712 2372
rect 157984 2320 158036 2372
rect 158812 2388 158864 2440
rect 159088 2431 159140 2440
rect 159088 2397 159097 2431
rect 159097 2397 159131 2431
rect 159131 2397 159140 2431
rect 159088 2388 159140 2397
rect 161112 2388 161164 2440
rect 161296 2456 161348 2508
rect 162400 2456 162452 2508
rect 162768 2456 162820 2508
rect 163228 2456 163280 2508
rect 167460 2524 167512 2576
rect 163688 2456 163740 2508
rect 161480 2388 161532 2440
rect 161572 2388 161624 2440
rect 164424 2388 164476 2440
rect 167276 2456 167328 2508
rect 169760 2524 169812 2576
rect 175740 2592 175792 2644
rect 175924 2635 175976 2644
rect 175924 2601 175933 2635
rect 175933 2601 175967 2635
rect 175967 2601 175976 2635
rect 175924 2592 175976 2601
rect 165436 2388 165488 2440
rect 167736 2456 167788 2508
rect 169116 2456 169168 2508
rect 169300 2456 169352 2508
rect 173348 2456 173400 2508
rect 173992 2499 174044 2508
rect 173992 2465 174001 2499
rect 174001 2465 174035 2499
rect 174035 2465 174044 2499
rect 173992 2456 174044 2465
rect 167552 2388 167604 2440
rect 176752 2524 176804 2576
rect 174912 2499 174964 2508
rect 174912 2465 174921 2499
rect 174921 2465 174955 2499
rect 174955 2465 174964 2499
rect 175832 2499 175884 2508
rect 174912 2456 174964 2465
rect 175832 2465 175841 2499
rect 175841 2465 175875 2499
rect 175875 2465 175884 2499
rect 175832 2456 175884 2465
rect 178132 2592 178184 2644
rect 184388 2592 184440 2644
rect 185124 2592 185176 2644
rect 176292 2388 176344 2440
rect 177028 2456 177080 2508
rect 181076 2456 181128 2508
rect 184572 2456 184624 2508
rect 184480 2388 184532 2440
rect 185676 2524 185728 2576
rect 186872 2524 186924 2576
rect 189356 2567 189408 2576
rect 185952 2456 186004 2508
rect 186044 2431 186096 2440
rect 146392 2252 146444 2304
rect 153016 2252 153068 2304
rect 160928 2252 160980 2304
rect 163136 2252 163188 2304
rect 163320 2252 163372 2304
rect 164884 2252 164936 2304
rect 167092 2252 167144 2304
rect 167184 2252 167236 2304
rect 177764 2252 177816 2304
rect 179604 2252 179656 2304
rect 181260 2320 181312 2372
rect 182548 2320 182600 2372
rect 184940 2320 184992 2372
rect 185124 2363 185176 2372
rect 185124 2329 185133 2363
rect 185133 2329 185167 2363
rect 185167 2329 185176 2363
rect 185124 2320 185176 2329
rect 186044 2397 186053 2431
rect 186053 2397 186087 2431
rect 186087 2397 186096 2431
rect 186044 2388 186096 2397
rect 187424 2431 187476 2440
rect 187424 2397 187433 2431
rect 187433 2397 187467 2431
rect 187467 2397 187476 2431
rect 187424 2388 187476 2397
rect 189356 2533 189365 2567
rect 189365 2533 189399 2567
rect 189399 2533 189408 2567
rect 189356 2524 189408 2533
rect 190184 2524 190236 2576
rect 192760 2592 192812 2644
rect 193864 2635 193916 2644
rect 193864 2601 193873 2635
rect 193873 2601 193907 2635
rect 193907 2601 193916 2635
rect 193864 2592 193916 2601
rect 194048 2592 194100 2644
rect 194968 2635 195020 2644
rect 194968 2601 194977 2635
rect 194977 2601 195011 2635
rect 195011 2601 195020 2635
rect 194968 2592 195020 2601
rect 195060 2592 195112 2644
rect 196440 2592 196492 2644
rect 189724 2456 189776 2508
rect 190552 2499 190604 2508
rect 190552 2465 190561 2499
rect 190561 2465 190595 2499
rect 190595 2465 190604 2499
rect 190552 2456 190604 2465
rect 190736 2456 190788 2508
rect 186596 2320 186648 2372
rect 191012 2320 191064 2372
rect 193220 2456 193272 2508
rect 194048 2456 194100 2508
rect 196900 2499 196952 2508
rect 192760 2388 192812 2440
rect 196900 2465 196909 2499
rect 196909 2465 196943 2499
rect 196943 2465 196952 2499
rect 196900 2456 196952 2465
rect 192668 2320 192720 2372
rect 193496 2320 193548 2372
rect 187332 2252 187384 2304
rect 187516 2252 187568 2304
rect 193312 2252 193364 2304
rect 4078 2150 4130 2202
rect 44078 2150 44130 2202
rect 84078 2150 84130 2202
rect 124078 2150 124130 2202
rect 164078 2150 164130 2202
rect 5724 2048 5776 2100
rect 6368 2048 6420 2100
rect 7472 2048 7524 2100
rect 8944 2091 8996 2100
rect 8944 2057 8953 2091
rect 8953 2057 8987 2091
rect 8987 2057 8996 2091
rect 8944 2048 8996 2057
rect 9956 2091 10008 2100
rect 9956 2057 9965 2091
rect 9965 2057 9999 2091
rect 9999 2057 10008 2091
rect 9956 2048 10008 2057
rect 11152 2048 11204 2100
rect 13544 2048 13596 2100
rect 13820 2091 13872 2100
rect 13820 2057 13829 2091
rect 13829 2057 13863 2091
rect 13863 2057 13872 2091
rect 13820 2048 13872 2057
rect 16672 2048 16724 2100
rect 19432 2048 19484 2100
rect 20536 2091 20588 2100
rect 20536 2057 20545 2091
rect 20545 2057 20579 2091
rect 20579 2057 20588 2091
rect 20536 2048 20588 2057
rect 23572 2048 23624 2100
rect 25044 2048 25096 2100
rect 27896 2048 27948 2100
rect 30472 2048 30524 2100
rect 32312 2091 32364 2100
rect 32312 2057 32321 2091
rect 32321 2057 32355 2091
rect 32355 2057 32364 2091
rect 32312 2048 32364 2057
rect 32772 2048 32824 2100
rect 34980 2091 35032 2100
rect 34980 2057 34989 2091
rect 34989 2057 35023 2091
rect 35023 2057 35032 2091
rect 34980 2048 35032 2057
rect 37924 2048 37976 2100
rect 39396 2091 39448 2100
rect 39396 2057 39405 2091
rect 39405 2057 39439 2091
rect 39439 2057 39448 2091
rect 39396 2048 39448 2057
rect 41144 2091 41196 2100
rect 41144 2057 41153 2091
rect 41153 2057 41187 2091
rect 41187 2057 41196 2091
rect 41144 2048 41196 2057
rect 42340 2091 42392 2100
rect 42340 2057 42349 2091
rect 42349 2057 42383 2091
rect 42383 2057 42392 2091
rect 42340 2048 42392 2057
rect 44272 2048 44324 2100
rect 44456 2091 44508 2100
rect 44456 2057 44465 2091
rect 44465 2057 44499 2091
rect 44499 2057 44508 2091
rect 44456 2048 44508 2057
rect 46204 2048 46256 2100
rect 47308 2091 47360 2100
rect 47308 2057 47317 2091
rect 47317 2057 47351 2091
rect 47351 2057 47360 2091
rect 47308 2048 47360 2057
rect 49700 2048 49752 2100
rect 54852 2048 54904 2100
rect 24768 1980 24820 2032
rect 30196 1980 30248 2032
rect 33416 1980 33468 2032
rect 57336 2048 57388 2100
rect 59544 2048 59596 2100
rect 67732 2048 67784 2100
rect 69664 2048 69716 2100
rect 93216 2048 93268 2100
rect 94504 2048 94556 2100
rect 100208 2091 100260 2100
rect 15844 1912 15896 1964
rect 4528 1844 4580 1896
rect 5356 1844 5408 1896
rect 6276 1776 6328 1828
rect 9312 1844 9364 1896
rect 10140 1844 10192 1896
rect 11060 1844 11112 1896
rect 13268 1844 13320 1896
rect 11888 1776 11940 1828
rect 15384 1844 15436 1896
rect 16672 1844 16724 1896
rect 21640 1912 21692 1964
rect 24584 1912 24636 1964
rect 17592 1776 17644 1828
rect 21088 1776 21140 1828
rect 22836 1776 22888 1828
rect 29736 1912 29788 1964
rect 30288 1912 30340 1964
rect 28080 1844 28132 1896
rect 28908 1776 28960 1828
rect 31944 1912 31996 1964
rect 41420 1912 41472 1964
rect 21456 1708 21508 1760
rect 23756 1708 23808 1760
rect 27620 1708 27672 1760
rect 32864 1776 32916 1828
rect 37740 1887 37792 1896
rect 37740 1853 37749 1887
rect 37749 1853 37783 1887
rect 37783 1853 37792 1887
rect 37740 1844 37792 1853
rect 35900 1776 35952 1828
rect 36728 1708 36780 1760
rect 42892 1844 42944 1896
rect 43444 1844 43496 1896
rect 41512 1776 41564 1828
rect 46388 1844 46440 1896
rect 47676 1844 47728 1896
rect 50712 1844 50764 1896
rect 53564 1844 53616 1896
rect 58900 1980 58952 2032
rect 57704 1912 57756 1964
rect 54024 1887 54076 1896
rect 54024 1853 54033 1887
rect 54033 1853 54067 1887
rect 54067 1853 54076 1887
rect 54024 1844 54076 1853
rect 55128 1887 55180 1896
rect 55128 1853 55137 1887
rect 55137 1853 55171 1887
rect 55171 1853 55180 1887
rect 55128 1844 55180 1853
rect 62304 1980 62356 2032
rect 62028 1912 62080 1964
rect 65984 1980 66036 2032
rect 54668 1776 54720 1828
rect 62120 1844 62172 1896
rect 71872 1980 71924 2032
rect 81440 1980 81492 2032
rect 81992 1980 82044 2032
rect 83004 1980 83056 2032
rect 83280 1980 83332 2032
rect 89720 1980 89772 2032
rect 100208 2057 100217 2091
rect 100217 2057 100251 2091
rect 100251 2057 100260 2091
rect 100208 2048 100260 2057
rect 105268 2048 105320 2100
rect 108396 2048 108448 2100
rect 108764 2048 108816 2100
rect 108948 2048 109000 2100
rect 109316 2048 109368 2100
rect 109408 2048 109460 2100
rect 113916 2048 113968 2100
rect 114008 2048 114060 2100
rect 116216 2091 116268 2100
rect 116216 2057 116225 2091
rect 116225 2057 116259 2091
rect 116259 2057 116268 2091
rect 116216 2048 116268 2057
rect 117596 2048 117648 2100
rect 118608 2048 118660 2100
rect 69848 1912 69900 1964
rect 66260 1887 66312 1896
rect 62948 1776 63000 1828
rect 43536 1708 43588 1760
rect 47032 1708 47084 1760
rect 66260 1853 66269 1887
rect 66269 1853 66303 1887
rect 66303 1853 66312 1887
rect 66260 1844 66312 1853
rect 68928 1887 68980 1896
rect 68928 1853 68937 1887
rect 68937 1853 68971 1887
rect 68971 1853 68980 1887
rect 68928 1844 68980 1853
rect 70584 1887 70636 1896
rect 70584 1853 70593 1887
rect 70593 1853 70627 1887
rect 70627 1853 70636 1887
rect 70584 1844 70636 1853
rect 72424 1887 72476 1896
rect 72424 1853 72433 1887
rect 72433 1853 72467 1887
rect 72467 1853 72476 1887
rect 72424 1844 72476 1853
rect 73528 1844 73580 1896
rect 81716 1912 81768 1964
rect 78220 1887 78272 1896
rect 78220 1853 78229 1887
rect 78229 1853 78263 1887
rect 78263 1853 78272 1887
rect 78220 1844 78272 1853
rect 80152 1887 80204 1896
rect 80152 1853 80161 1887
rect 80161 1853 80195 1887
rect 80195 1853 80204 1887
rect 80152 1844 80204 1853
rect 82176 1844 82228 1896
rect 93032 1912 93084 1964
rect 84660 1844 84712 1896
rect 85856 1887 85908 1896
rect 85856 1853 85865 1887
rect 85865 1853 85899 1887
rect 85899 1853 85908 1887
rect 85856 1844 85908 1853
rect 88432 1844 88484 1896
rect 88800 1887 88852 1896
rect 88800 1853 88809 1887
rect 88809 1853 88843 1887
rect 88843 1853 88852 1887
rect 88800 1844 88852 1853
rect 91376 1887 91428 1896
rect 91376 1853 91385 1887
rect 91385 1853 91419 1887
rect 91419 1853 91428 1887
rect 91376 1844 91428 1853
rect 92848 1887 92900 1896
rect 92848 1853 92857 1887
rect 92857 1853 92891 1887
rect 92891 1853 92900 1887
rect 92848 1844 92900 1853
rect 96252 1912 96304 1964
rect 105452 1980 105504 2032
rect 108120 1980 108172 2032
rect 110880 1980 110932 2032
rect 110972 1980 111024 2032
rect 113364 1980 113416 2032
rect 95976 1844 96028 1896
rect 97080 1844 97132 1896
rect 63776 1776 63828 1828
rect 66168 1776 66220 1828
rect 69572 1776 69624 1828
rect 70768 1776 70820 1828
rect 77760 1776 77812 1828
rect 89904 1776 89956 1828
rect 92940 1776 92992 1828
rect 96436 1776 96488 1828
rect 98184 1776 98236 1828
rect 98276 1776 98328 1828
rect 100852 1912 100904 1964
rect 106648 1912 106700 1964
rect 107752 1912 107804 1964
rect 66904 1708 66956 1760
rect 78128 1708 78180 1760
rect 79876 1708 79928 1760
rect 81624 1751 81676 1760
rect 81624 1717 81633 1751
rect 81633 1717 81667 1751
rect 81667 1717 81676 1751
rect 81624 1708 81676 1717
rect 83372 1751 83424 1760
rect 83372 1717 83381 1751
rect 83381 1717 83415 1751
rect 83415 1717 83424 1751
rect 83372 1708 83424 1717
rect 85580 1708 85632 1760
rect 87328 1708 87380 1760
rect 93216 1708 93268 1760
rect 96988 1708 97040 1760
rect 100668 1776 100720 1828
rect 101128 1887 101180 1896
rect 101128 1853 101137 1887
rect 101137 1853 101171 1887
rect 101171 1853 101180 1887
rect 102784 1887 102836 1896
rect 101128 1844 101180 1853
rect 102784 1853 102793 1887
rect 102793 1853 102827 1887
rect 102827 1853 102836 1887
rect 102784 1844 102836 1853
rect 104256 1776 104308 1828
rect 105268 1887 105320 1896
rect 105268 1853 105277 1887
rect 105277 1853 105311 1887
rect 105311 1853 105320 1887
rect 105268 1844 105320 1853
rect 107844 1844 107896 1896
rect 106740 1776 106792 1828
rect 108212 1776 108264 1828
rect 108488 1887 108540 1896
rect 108488 1853 108497 1887
rect 108497 1853 108531 1887
rect 108531 1853 108540 1887
rect 108488 1844 108540 1853
rect 109960 1844 110012 1896
rect 110788 1844 110840 1896
rect 110420 1776 110472 1828
rect 111708 1776 111760 1828
rect 112076 1887 112128 1896
rect 112076 1853 112085 1887
rect 112085 1853 112119 1887
rect 112119 1853 112128 1887
rect 119988 1980 120040 2032
rect 120264 2091 120316 2100
rect 120264 2057 120273 2091
rect 120273 2057 120307 2091
rect 120307 2057 120316 2091
rect 120264 2048 120316 2057
rect 124496 2048 124548 2100
rect 124864 2048 124916 2100
rect 125324 2048 125376 2100
rect 126520 2048 126572 2100
rect 126796 2048 126848 2100
rect 127808 2048 127860 2100
rect 132868 2091 132920 2100
rect 122840 1980 122892 2032
rect 113548 1955 113600 1964
rect 113548 1921 113557 1955
rect 113557 1921 113591 1955
rect 113591 1921 113600 1955
rect 113548 1912 113600 1921
rect 113824 1912 113876 1964
rect 117136 1912 117188 1964
rect 112076 1844 112128 1853
rect 113640 1844 113692 1896
rect 114468 1844 114520 1896
rect 115112 1887 115164 1896
rect 115112 1853 115121 1887
rect 115121 1853 115155 1887
rect 115155 1853 115164 1887
rect 115112 1844 115164 1853
rect 115204 1844 115256 1896
rect 118332 1912 118384 1964
rect 118056 1844 118108 1896
rect 128176 1912 128228 1964
rect 118608 1844 118660 1896
rect 119896 1844 119948 1896
rect 119160 1819 119212 1828
rect 119160 1785 119169 1819
rect 119169 1785 119203 1819
rect 119203 1785 119212 1819
rect 119160 1776 119212 1785
rect 120080 1819 120132 1828
rect 120080 1785 120089 1819
rect 120089 1785 120123 1819
rect 120123 1785 120132 1819
rect 120080 1776 120132 1785
rect 123024 1776 123076 1828
rect 123944 1844 123996 1896
rect 124956 1776 125008 1828
rect 125784 1887 125836 1896
rect 125784 1853 125793 1887
rect 125793 1853 125827 1887
rect 125827 1853 125836 1887
rect 125784 1844 125836 1853
rect 126796 1887 126848 1896
rect 126796 1853 126805 1887
rect 126805 1853 126839 1887
rect 126839 1853 126848 1887
rect 126796 1844 126848 1853
rect 126888 1887 126940 1896
rect 126888 1853 126897 1887
rect 126897 1853 126931 1887
rect 126931 1853 126940 1887
rect 126888 1844 126940 1853
rect 131028 1980 131080 2032
rect 131304 1980 131356 2032
rect 131764 1980 131816 2032
rect 132868 2057 132877 2091
rect 132877 2057 132911 2091
rect 132911 2057 132920 2091
rect 132868 2048 132920 2057
rect 133972 2048 134024 2100
rect 134064 2048 134116 2100
rect 136732 2048 136784 2100
rect 137560 2048 137612 2100
rect 137652 2048 137704 2100
rect 138572 2048 138624 2100
rect 139584 2048 139636 2100
rect 143356 2048 143408 2100
rect 137744 1980 137796 2032
rect 137836 1980 137888 2032
rect 144184 1980 144236 2032
rect 130292 1887 130344 1896
rect 130292 1853 130301 1887
rect 130301 1853 130335 1887
rect 130335 1853 130344 1887
rect 130292 1844 130344 1853
rect 125324 1776 125376 1828
rect 104532 1708 104584 1760
rect 104624 1708 104676 1760
rect 108764 1708 108816 1760
rect 110604 1708 110656 1760
rect 114284 1708 114336 1760
rect 114376 1708 114428 1760
rect 116032 1708 116084 1760
rect 116124 1708 116176 1760
rect 121920 1708 121972 1760
rect 124680 1708 124732 1760
rect 125048 1751 125100 1760
rect 125048 1717 125057 1751
rect 125057 1717 125091 1751
rect 125091 1717 125100 1751
rect 125048 1708 125100 1717
rect 129188 1776 129240 1828
rect 131212 1844 131264 1896
rect 138204 1912 138256 1964
rect 133696 1844 133748 1896
rect 133880 1844 133932 1896
rect 130752 1776 130804 1828
rect 131672 1776 131724 1828
rect 134616 1844 134668 1896
rect 134800 1887 134852 1896
rect 134800 1853 134809 1887
rect 134809 1853 134843 1887
rect 134843 1853 134852 1887
rect 134800 1844 134852 1853
rect 135352 1844 135404 1896
rect 135812 1844 135864 1896
rect 134248 1776 134300 1828
rect 135996 1844 136048 1896
rect 137284 1844 137336 1896
rect 140044 1912 140096 1964
rect 140136 1912 140188 1964
rect 144276 1912 144328 1964
rect 144460 1980 144512 2032
rect 147128 2048 147180 2100
rect 147312 2048 147364 2100
rect 148876 2048 148928 2100
rect 146944 1980 146996 2032
rect 147404 1980 147456 2032
rect 150072 1980 150124 2032
rect 153476 2048 153528 2100
rect 159364 2048 159416 2100
rect 159456 2048 159508 2100
rect 160836 2091 160888 2100
rect 153844 1980 153896 2032
rect 155684 1980 155736 2032
rect 128176 1708 128228 1760
rect 129556 1708 129608 1760
rect 134156 1708 134208 1760
rect 134616 1708 134668 1760
rect 138020 1776 138072 1828
rect 139216 1844 139268 1896
rect 138848 1776 138900 1828
rect 139676 1776 139728 1828
rect 140872 1776 140924 1828
rect 144736 1844 144788 1896
rect 145472 1844 145524 1896
rect 145564 1844 145616 1896
rect 145288 1776 145340 1828
rect 150900 1912 150952 1964
rect 155224 1912 155276 1964
rect 159548 1980 159600 2032
rect 160836 2057 160845 2091
rect 160845 2057 160879 2091
rect 160879 2057 160888 2091
rect 160836 2048 160888 2057
rect 160928 2048 160980 2100
rect 162400 2048 162452 2100
rect 163228 1980 163280 2032
rect 164332 1980 164384 2032
rect 164516 2048 164568 2100
rect 155960 1912 156012 1964
rect 158720 1955 158772 1964
rect 158720 1921 158729 1955
rect 158729 1921 158763 1955
rect 158763 1921 158772 1955
rect 158720 1912 158772 1921
rect 159732 1955 159784 1964
rect 159732 1921 159741 1955
rect 159741 1921 159775 1955
rect 159775 1921 159784 1955
rect 159732 1912 159784 1921
rect 159824 1912 159876 1964
rect 162216 1912 162268 1964
rect 146852 1776 146904 1828
rect 160560 1844 160612 1896
rect 160744 1887 160796 1896
rect 160744 1853 160753 1887
rect 160753 1853 160787 1887
rect 160787 1853 160796 1887
rect 160744 1844 160796 1853
rect 161112 1844 161164 1896
rect 161572 1844 161624 1896
rect 161756 1887 161808 1896
rect 161756 1853 161765 1887
rect 161765 1853 161799 1887
rect 161799 1853 161808 1887
rect 161756 1844 161808 1853
rect 149612 1776 149664 1828
rect 136180 1708 136232 1760
rect 136640 1708 136692 1760
rect 137100 1708 137152 1760
rect 138112 1708 138164 1760
rect 138296 1708 138348 1760
rect 140136 1708 140188 1760
rect 140228 1708 140280 1760
rect 145104 1708 145156 1760
rect 145196 1708 145248 1760
rect 155960 1708 156012 1760
rect 156052 1708 156104 1760
rect 159364 1776 159416 1828
rect 161480 1776 161532 1828
rect 163044 1844 163096 1896
rect 164240 1844 164292 1896
rect 163596 1776 163648 1828
rect 163688 1776 163740 1828
rect 164700 1955 164752 1964
rect 164700 1921 164709 1955
rect 164709 1921 164743 1955
rect 164743 1921 164752 1955
rect 165252 1980 165304 2032
rect 165620 1980 165672 2032
rect 165712 2023 165764 2032
rect 165712 1989 165721 2023
rect 165721 1989 165755 2023
rect 165755 1989 165764 2023
rect 167092 2048 167144 2100
rect 168564 2091 168616 2100
rect 165712 1980 165764 1989
rect 167184 1980 167236 2032
rect 164700 1912 164752 1921
rect 167000 1912 167052 1964
rect 167552 1980 167604 2032
rect 168564 2057 168573 2091
rect 168573 2057 168607 2091
rect 168607 2057 168616 2091
rect 168564 2048 168616 2057
rect 168656 2048 168708 2100
rect 173992 2048 174044 2100
rect 175740 2048 175792 2100
rect 177764 2048 177816 2100
rect 177856 2048 177908 2100
rect 179604 2048 179656 2100
rect 181996 2091 182048 2100
rect 171232 1980 171284 2032
rect 176476 1980 176528 2032
rect 178224 1980 178276 2032
rect 180340 1980 180392 2032
rect 181996 2057 182005 2091
rect 182005 2057 182039 2091
rect 182039 2057 182048 2091
rect 181996 2048 182048 2057
rect 184848 2048 184900 2100
rect 185400 2091 185452 2100
rect 185400 2057 185409 2091
rect 185409 2057 185443 2091
rect 185443 2057 185452 2091
rect 185400 2048 185452 2057
rect 186320 2048 186372 2100
rect 186412 2048 186464 2100
rect 189264 2048 189316 2100
rect 192944 2091 192996 2100
rect 192944 2057 192953 2091
rect 192953 2057 192987 2091
rect 192987 2057 192996 2091
rect 192944 2048 192996 2057
rect 195060 2048 195112 2100
rect 195888 2048 195940 2100
rect 186228 1980 186280 2032
rect 186596 1980 186648 2032
rect 189448 1980 189500 2032
rect 176844 1912 176896 1964
rect 165436 1844 165488 1896
rect 168380 1844 168432 1896
rect 169484 1844 169536 1896
rect 169668 1844 169720 1896
rect 169944 1844 169996 1896
rect 171876 1844 171928 1896
rect 172980 1887 173032 1896
rect 172980 1853 172989 1887
rect 172989 1853 173023 1887
rect 173023 1853 173032 1887
rect 172980 1844 173032 1853
rect 173072 1844 173124 1896
rect 173624 1844 173676 1896
rect 173808 1887 173860 1896
rect 173808 1853 173817 1887
rect 173817 1853 173851 1887
rect 173851 1853 173860 1887
rect 173808 1844 173860 1853
rect 176200 1844 176252 1896
rect 176292 1844 176344 1896
rect 178224 1844 178276 1896
rect 181076 1912 181128 1964
rect 186044 1912 186096 1964
rect 179328 1844 179380 1896
rect 161940 1708 161992 1760
rect 162032 1708 162084 1760
rect 169760 1708 169812 1760
rect 172428 1708 172480 1760
rect 172980 1708 173032 1760
rect 176016 1708 176068 1760
rect 176108 1708 176160 1760
rect 179512 1844 179564 1896
rect 180708 1844 180760 1896
rect 181628 1776 181680 1828
rect 183468 1708 183520 1760
rect 183744 1844 183796 1896
rect 184940 1844 184992 1896
rect 187700 1912 187752 1964
rect 191472 1912 191524 1964
rect 191932 1912 191984 1964
rect 194692 1955 194744 1964
rect 190460 1844 190512 1896
rect 185768 1776 185820 1828
rect 186320 1776 186372 1828
rect 189264 1776 189316 1828
rect 190644 1887 190696 1896
rect 190644 1853 190653 1887
rect 190653 1853 190687 1887
rect 190687 1853 190696 1887
rect 190644 1844 190696 1853
rect 193312 1844 193364 1896
rect 194692 1921 194701 1955
rect 194701 1921 194735 1955
rect 194735 1921 194744 1955
rect 194692 1912 194744 1921
rect 197268 1776 197320 1828
rect 185308 1708 185360 1760
rect 185952 1708 186004 1760
rect 189816 1708 189868 1760
rect 195152 1708 195204 1760
rect 24078 1606 24130 1658
rect 64078 1606 64130 1658
rect 104078 1606 104130 1658
rect 144078 1606 144130 1658
rect 184078 1606 184130 1658
rect 5908 1504 5960 1556
rect 7196 1504 7248 1556
rect 7932 1504 7984 1556
rect 16580 1504 16632 1556
rect 16856 1547 16908 1556
rect 16856 1513 16865 1547
rect 16865 1513 16899 1547
rect 16899 1513 16908 1547
rect 16856 1504 16908 1513
rect 21916 1504 21968 1556
rect 22008 1504 22060 1556
rect 24952 1504 25004 1556
rect 25320 1504 25372 1556
rect 28540 1547 28592 1556
rect 28540 1513 28549 1547
rect 28549 1513 28583 1547
rect 28583 1513 28592 1547
rect 28540 1504 28592 1513
rect 32956 1547 33008 1556
rect 32956 1513 32965 1547
rect 32965 1513 32999 1547
rect 32999 1513 33008 1547
rect 32956 1504 33008 1513
rect 33876 1504 33928 1556
rect 35992 1504 36044 1556
rect 39120 1547 39172 1556
rect 39120 1513 39129 1547
rect 39129 1513 39163 1547
rect 39163 1513 39172 1547
rect 39120 1504 39172 1513
rect 43536 1504 43588 1556
rect 43628 1504 43680 1556
rect 45376 1504 45428 1556
rect 50344 1504 50396 1556
rect 52552 1504 52604 1556
rect 53840 1504 53892 1556
rect 54116 1547 54168 1556
rect 54116 1513 54125 1547
rect 54125 1513 54159 1547
rect 54159 1513 54168 1547
rect 54116 1504 54168 1513
rect 62488 1504 62540 1556
rect 75368 1504 75420 1556
rect 79968 1547 80020 1556
rect 79968 1513 79977 1547
rect 79977 1513 80011 1547
rect 80011 1513 80020 1547
rect 79968 1504 80020 1513
rect 14096 1436 14148 1488
rect 3976 1368 4028 1420
rect 4988 1300 5040 1352
rect 7564 1368 7616 1420
rect 16304 1368 16356 1420
rect 20628 1436 20680 1488
rect 18880 1368 18932 1420
rect 19800 1300 19852 1352
rect 21456 1411 21508 1420
rect 21456 1377 21465 1411
rect 21465 1377 21499 1411
rect 21499 1377 21508 1411
rect 32404 1436 32456 1488
rect 21456 1368 21508 1377
rect 21916 1300 21968 1352
rect 22560 1300 22612 1352
rect 23664 1232 23716 1284
rect 30656 1368 30708 1420
rect 33048 1368 33100 1420
rect 38108 1436 38160 1488
rect 34980 1300 35032 1352
rect 41604 1368 41656 1420
rect 43076 1436 43128 1488
rect 51172 1436 51224 1488
rect 47492 1368 47544 1420
rect 49884 1368 49936 1420
rect 52920 1368 52972 1420
rect 58624 1368 58676 1420
rect 63500 1436 63552 1488
rect 65064 1436 65116 1488
rect 79048 1436 79100 1488
rect 59820 1368 59872 1420
rect 61476 1411 61528 1420
rect 61476 1377 61485 1411
rect 61485 1377 61519 1411
rect 61519 1377 61528 1411
rect 61476 1368 61528 1377
rect 64236 1368 64288 1420
rect 66168 1368 66220 1420
rect 69480 1368 69532 1420
rect 70308 1368 70360 1420
rect 72608 1411 72660 1420
rect 55956 1300 56008 1352
rect 72608 1377 72617 1411
rect 72617 1377 72651 1411
rect 72651 1377 72660 1411
rect 72608 1368 72660 1377
rect 75460 1411 75512 1420
rect 75460 1377 75469 1411
rect 75469 1377 75503 1411
rect 75503 1377 75512 1411
rect 75460 1368 75512 1377
rect 76380 1368 76432 1420
rect 81440 1504 81492 1556
rect 82176 1504 82228 1556
rect 83280 1504 83332 1556
rect 86316 1504 86368 1556
rect 91192 1547 91244 1556
rect 84660 1411 84712 1420
rect 84660 1377 84669 1411
rect 84669 1377 84703 1411
rect 84703 1377 84712 1411
rect 84660 1368 84712 1377
rect 85672 1368 85724 1420
rect 91192 1513 91201 1547
rect 91201 1513 91235 1547
rect 91235 1513 91244 1547
rect 91192 1504 91244 1513
rect 95516 1504 95568 1556
rect 96988 1547 97040 1556
rect 96988 1513 96997 1547
rect 96997 1513 97031 1547
rect 97031 1513 97040 1547
rect 96988 1504 97040 1513
rect 92756 1436 92808 1488
rect 93032 1436 93084 1488
rect 87420 1411 87472 1420
rect 87420 1377 87429 1411
rect 87429 1377 87463 1411
rect 87463 1377 87472 1411
rect 87420 1368 87472 1377
rect 89628 1368 89680 1420
rect 90180 1411 90232 1420
rect 90180 1377 90189 1411
rect 90189 1377 90223 1411
rect 90223 1377 90232 1411
rect 90180 1368 90232 1377
rect 90364 1411 90416 1420
rect 90364 1377 90373 1411
rect 90373 1377 90407 1411
rect 90407 1377 90416 1411
rect 90364 1368 90416 1377
rect 92112 1368 92164 1420
rect 93124 1411 93176 1420
rect 93124 1377 93133 1411
rect 93133 1377 93167 1411
rect 93167 1377 93176 1411
rect 93124 1368 93176 1377
rect 86408 1300 86460 1352
rect 95240 1436 95292 1488
rect 95148 1368 95200 1420
rect 98920 1436 98972 1488
rect 104624 1504 104676 1556
rect 105728 1547 105780 1556
rect 105728 1513 105737 1547
rect 105737 1513 105771 1547
rect 105771 1513 105780 1547
rect 105728 1504 105780 1513
rect 99288 1436 99340 1488
rect 104716 1436 104768 1488
rect 109040 1504 109092 1556
rect 102232 1368 102284 1420
rect 99288 1232 99340 1284
rect 105544 1368 105596 1420
rect 109500 1504 109552 1556
rect 109684 1547 109736 1556
rect 109684 1513 109693 1547
rect 109693 1513 109727 1547
rect 109727 1513 109736 1547
rect 109684 1504 109736 1513
rect 109776 1504 109828 1556
rect 114376 1504 114428 1556
rect 115756 1504 115808 1556
rect 117688 1504 117740 1556
rect 119160 1504 119212 1556
rect 120448 1504 120500 1556
rect 121092 1504 121144 1556
rect 121828 1504 121880 1556
rect 123760 1504 123812 1556
rect 127900 1504 127952 1556
rect 128084 1504 128136 1556
rect 140320 1504 140372 1556
rect 141240 1547 141292 1556
rect 141240 1513 141249 1547
rect 141249 1513 141283 1547
rect 141283 1513 141292 1547
rect 141240 1504 141292 1513
rect 141700 1504 141752 1556
rect 143080 1504 143132 1556
rect 146208 1504 146260 1556
rect 146852 1504 146904 1556
rect 147404 1504 147456 1556
rect 150348 1547 150400 1556
rect 150348 1513 150357 1547
rect 150357 1513 150391 1547
rect 150391 1513 150400 1547
rect 150348 1504 150400 1513
rect 152464 1547 152516 1556
rect 152464 1513 152473 1547
rect 152473 1513 152507 1547
rect 152507 1513 152516 1547
rect 152464 1504 152516 1513
rect 154028 1504 154080 1556
rect 105820 1368 105872 1420
rect 106832 1411 106884 1420
rect 104532 1300 104584 1352
rect 106832 1377 106841 1411
rect 106841 1377 106875 1411
rect 106875 1377 106884 1411
rect 106832 1368 106884 1377
rect 109408 1368 109460 1420
rect 108304 1232 108356 1284
rect 99196 1207 99248 1216
rect 99196 1173 99205 1207
rect 99205 1173 99239 1207
rect 99239 1173 99248 1207
rect 99196 1164 99248 1173
rect 108580 1164 108632 1216
rect 110604 1411 110656 1420
rect 110604 1377 110613 1411
rect 110613 1377 110647 1411
rect 110647 1377 110656 1411
rect 110604 1368 110656 1377
rect 110696 1411 110748 1420
rect 110696 1377 110705 1411
rect 110705 1377 110739 1411
rect 110739 1377 110748 1411
rect 110696 1368 110748 1377
rect 112352 1368 112404 1420
rect 112536 1343 112588 1352
rect 112536 1309 112545 1343
rect 112545 1309 112579 1343
rect 112579 1309 112588 1343
rect 112536 1300 112588 1309
rect 118884 1436 118936 1488
rect 115296 1411 115348 1420
rect 115296 1377 115305 1411
rect 115305 1377 115339 1411
rect 115339 1377 115348 1411
rect 115296 1368 115348 1377
rect 118056 1368 118108 1420
rect 118792 1368 118844 1420
rect 122196 1436 122248 1488
rect 122288 1436 122340 1488
rect 124680 1436 124732 1488
rect 125232 1436 125284 1488
rect 129188 1436 129240 1488
rect 129464 1436 129516 1488
rect 121368 1411 121420 1420
rect 121368 1377 121377 1411
rect 121377 1377 121411 1411
rect 121411 1377 121420 1411
rect 121368 1368 121420 1377
rect 123760 1368 123812 1420
rect 124864 1411 124916 1420
rect 116492 1300 116544 1352
rect 119344 1300 119396 1352
rect 123392 1300 123444 1352
rect 124864 1377 124873 1411
rect 124873 1377 124907 1411
rect 124907 1377 124916 1411
rect 124864 1368 124916 1377
rect 125048 1368 125100 1420
rect 125140 1300 125192 1352
rect 128084 1368 128136 1420
rect 128452 1411 128504 1420
rect 128452 1377 128461 1411
rect 128461 1377 128495 1411
rect 128495 1377 128504 1411
rect 128452 1368 128504 1377
rect 129648 1368 129700 1420
rect 127808 1300 127860 1352
rect 132408 1411 132460 1420
rect 132408 1377 132417 1411
rect 132417 1377 132451 1411
rect 132451 1377 132460 1411
rect 132408 1368 132460 1377
rect 133236 1368 133288 1420
rect 133420 1411 133472 1420
rect 133420 1377 133429 1411
rect 133429 1377 133463 1411
rect 133463 1377 133472 1411
rect 133420 1368 133472 1377
rect 134064 1368 134116 1420
rect 112168 1232 112220 1284
rect 118148 1232 118200 1284
rect 127532 1232 127584 1284
rect 127900 1232 127952 1284
rect 129096 1232 129148 1284
rect 129280 1232 129332 1284
rect 117044 1164 117096 1216
rect 120540 1164 120592 1216
rect 125232 1164 125284 1216
rect 125968 1164 126020 1216
rect 127440 1164 127492 1216
rect 127624 1164 127676 1216
rect 134984 1300 135036 1352
rect 135444 1436 135496 1488
rect 135628 1436 135680 1488
rect 136180 1436 136232 1488
rect 136364 1479 136416 1488
rect 136364 1445 136373 1479
rect 136373 1445 136407 1479
rect 136407 1445 136416 1479
rect 136364 1436 136416 1445
rect 136824 1436 136876 1488
rect 137836 1436 137888 1488
rect 137928 1436 137980 1488
rect 138848 1436 138900 1488
rect 135260 1411 135312 1420
rect 135260 1377 135269 1411
rect 135269 1377 135303 1411
rect 135303 1377 135312 1411
rect 135260 1368 135312 1377
rect 137008 1368 137060 1420
rect 137192 1368 137244 1420
rect 138572 1368 138624 1420
rect 138940 1411 138992 1420
rect 138940 1377 138949 1411
rect 138949 1377 138983 1411
rect 138983 1377 138992 1411
rect 138940 1368 138992 1377
rect 139032 1411 139084 1420
rect 139032 1377 139041 1411
rect 139041 1377 139075 1411
rect 139075 1377 139084 1411
rect 139032 1368 139084 1377
rect 139676 1368 139728 1420
rect 142988 1436 143040 1488
rect 141148 1411 141200 1420
rect 141148 1377 141157 1411
rect 141157 1377 141191 1411
rect 141191 1377 141200 1411
rect 141148 1368 141200 1377
rect 141516 1368 141568 1420
rect 143816 1368 143868 1420
rect 144920 1436 144972 1488
rect 145104 1479 145156 1488
rect 145104 1445 145113 1479
rect 145113 1445 145147 1479
rect 145147 1445 145156 1479
rect 145104 1436 145156 1445
rect 144644 1368 144696 1420
rect 137100 1300 137152 1352
rect 137284 1300 137336 1352
rect 145472 1368 145524 1420
rect 146668 1411 146720 1420
rect 133420 1232 133472 1284
rect 141516 1232 141568 1284
rect 133696 1164 133748 1216
rect 138848 1164 138900 1216
rect 139124 1164 139176 1216
rect 140688 1164 140740 1216
rect 144644 1232 144696 1284
rect 142896 1164 142948 1216
rect 145012 1164 145064 1216
rect 146668 1377 146677 1411
rect 146677 1377 146711 1411
rect 146711 1377 146720 1411
rect 146668 1368 146720 1377
rect 146944 1436 146996 1488
rect 148784 1436 148836 1488
rect 155684 1504 155736 1556
rect 161020 1547 161072 1556
rect 159824 1479 159876 1488
rect 149060 1368 149112 1420
rect 150256 1411 150308 1420
rect 150256 1377 150265 1411
rect 150265 1377 150299 1411
rect 150299 1377 150308 1411
rect 150256 1368 150308 1377
rect 153844 1368 153896 1420
rect 155040 1300 155092 1352
rect 156328 1368 156380 1420
rect 157248 1368 157300 1420
rect 159824 1445 159833 1479
rect 159833 1445 159867 1479
rect 159867 1445 159876 1479
rect 159824 1436 159876 1445
rect 161020 1513 161029 1547
rect 161029 1513 161063 1547
rect 161063 1513 161072 1547
rect 161020 1504 161072 1513
rect 161204 1504 161256 1556
rect 162492 1504 162544 1556
rect 162124 1436 162176 1488
rect 160652 1368 160704 1420
rect 163688 1504 163740 1556
rect 164516 1479 164568 1488
rect 164516 1445 164525 1479
rect 164525 1445 164559 1479
rect 164559 1445 164568 1479
rect 164516 1436 164568 1445
rect 164976 1504 165028 1556
rect 165252 1436 165304 1488
rect 165528 1479 165580 1488
rect 165528 1445 165537 1479
rect 165537 1445 165571 1479
rect 165571 1445 165580 1479
rect 165528 1436 165580 1445
rect 162768 1411 162820 1420
rect 162768 1377 162777 1411
rect 162777 1377 162811 1411
rect 162811 1377 162820 1411
rect 162768 1368 162820 1377
rect 163596 1368 163648 1420
rect 164976 1368 165028 1420
rect 165068 1368 165120 1420
rect 167920 1368 167972 1420
rect 169300 1504 169352 1556
rect 170036 1504 170088 1556
rect 168104 1436 168156 1488
rect 169944 1436 169996 1488
rect 169392 1368 169444 1420
rect 174912 1504 174964 1556
rect 171324 1479 171376 1488
rect 171324 1445 171333 1479
rect 171333 1445 171367 1479
rect 171367 1445 171376 1479
rect 171324 1436 171376 1445
rect 171232 1411 171284 1420
rect 171232 1377 171241 1411
rect 171241 1377 171275 1411
rect 171275 1377 171284 1411
rect 171232 1368 171284 1377
rect 173072 1436 173124 1488
rect 173624 1436 173676 1488
rect 174452 1436 174504 1488
rect 172428 1411 172480 1420
rect 172428 1377 172437 1411
rect 172437 1377 172471 1411
rect 172471 1377 172480 1411
rect 172428 1368 172480 1377
rect 173256 1368 173308 1420
rect 173348 1411 173400 1420
rect 173348 1377 173357 1411
rect 173357 1377 173391 1411
rect 173391 1377 173400 1411
rect 173348 1368 173400 1377
rect 173532 1368 173584 1420
rect 175740 1504 175792 1556
rect 176568 1504 176620 1556
rect 178316 1504 178368 1556
rect 179328 1504 179380 1556
rect 182272 1504 182324 1556
rect 183560 1504 183612 1556
rect 184756 1504 184808 1556
rect 185492 1504 185544 1556
rect 187884 1504 187936 1556
rect 188988 1504 189040 1556
rect 155500 1300 155552 1352
rect 156052 1300 156104 1352
rect 159088 1300 159140 1352
rect 162032 1300 162084 1352
rect 162400 1300 162452 1352
rect 164332 1300 164384 1352
rect 164884 1300 164936 1352
rect 166908 1300 166960 1352
rect 167368 1343 167420 1352
rect 167368 1309 167377 1343
rect 167377 1309 167411 1343
rect 167411 1309 167420 1343
rect 167368 1300 167420 1309
rect 167460 1300 167512 1352
rect 176108 1368 176160 1420
rect 176844 1436 176896 1488
rect 186136 1436 186188 1488
rect 186320 1436 186372 1488
rect 188804 1436 188856 1488
rect 188896 1436 188948 1488
rect 191380 1504 191432 1556
rect 194968 1504 195020 1556
rect 175372 1300 175424 1352
rect 177488 1368 177540 1420
rect 178132 1411 178184 1420
rect 178132 1377 178141 1411
rect 178141 1377 178175 1411
rect 178175 1377 178184 1411
rect 178132 1368 178184 1377
rect 181260 1411 181312 1420
rect 180524 1300 180576 1352
rect 181260 1377 181269 1411
rect 181269 1377 181303 1411
rect 181303 1377 181312 1411
rect 181260 1368 181312 1377
rect 183192 1300 183244 1352
rect 186688 1368 186740 1420
rect 186872 1368 186924 1420
rect 187148 1368 187200 1420
rect 186228 1300 186280 1352
rect 145748 1232 145800 1284
rect 175188 1232 175240 1284
rect 175464 1232 175516 1284
rect 147864 1164 147916 1216
rect 148232 1164 148284 1216
rect 160100 1164 160152 1216
rect 162308 1164 162360 1216
rect 162768 1164 162820 1216
rect 162860 1164 162912 1216
rect 186596 1232 186648 1284
rect 188436 1368 188488 1420
rect 193312 1411 193364 1420
rect 193312 1377 193321 1411
rect 193321 1377 193355 1411
rect 193355 1377 193364 1411
rect 193312 1368 193364 1377
rect 195060 1368 195112 1420
rect 195152 1411 195204 1420
rect 195152 1377 195161 1411
rect 195161 1377 195195 1411
rect 195195 1377 195204 1411
rect 195152 1368 195204 1377
rect 198464 1368 198516 1420
rect 191380 1300 191432 1352
rect 196716 1300 196768 1352
rect 195796 1232 195848 1284
rect 176476 1164 176528 1216
rect 178776 1164 178828 1216
rect 181352 1207 181404 1216
rect 181352 1173 181361 1207
rect 181361 1173 181395 1207
rect 181395 1173 181404 1207
rect 181352 1164 181404 1173
rect 181628 1164 181680 1216
rect 182272 1164 182324 1216
rect 4078 1062 4130 1114
rect 44078 1062 44130 1114
rect 84078 1062 84130 1114
rect 124078 1062 124130 1114
rect 164078 1062 164130 1114
rect 108120 960 108172 1012
rect 112168 960 112220 1012
rect 117780 960 117832 1012
rect 108028 892 108080 944
rect 113456 892 113508 944
rect 106740 824 106792 876
rect 115664 892 115716 944
rect 118884 892 118936 944
rect 123944 892 123996 944
rect 126244 892 126296 944
rect 130016 892 130068 944
rect 130108 892 130160 944
rect 133052 892 133104 944
rect 115112 824 115164 876
rect 127624 824 127676 876
rect 127992 824 128044 876
rect 132500 824 132552 876
rect 133788 960 133840 1012
rect 134800 960 134852 1012
rect 134892 960 134944 1012
rect 137284 960 137336 1012
rect 149704 960 149756 1012
rect 152924 960 152976 1012
rect 162860 960 162912 1012
rect 162952 960 163004 1012
rect 166080 960 166132 1012
rect 140504 892 140556 944
rect 140688 892 140740 944
rect 144552 892 144604 944
rect 156880 892 156932 944
rect 160468 892 160520 944
rect 160560 892 160612 944
rect 162032 892 162084 944
rect 168288 892 168340 944
rect 169116 960 169168 1012
rect 172704 892 172756 944
rect 181444 892 181496 944
rect 181536 892 181588 944
rect 143816 824 143868 876
rect 148232 824 148284 876
rect 119712 756 119764 808
rect 132408 756 132460 808
rect 121368 688 121420 740
rect 115296 552 115348 604
rect 137100 756 137152 808
rect 142896 756 142948 808
rect 142988 756 143040 808
rect 152740 824 152792 876
rect 155960 824 156012 876
rect 167000 824 167052 876
rect 169024 824 169076 876
rect 175280 824 175332 876
rect 175832 824 175884 876
rect 181812 824 181864 876
rect 142528 688 142580 740
rect 143724 688 143776 740
rect 144644 688 144696 740
rect 144920 688 144972 740
rect 163412 756 163464 808
rect 163780 756 163832 808
rect 171140 756 171192 808
rect 188068 756 188120 808
rect 164792 688 164844 740
rect 169576 688 169628 740
rect 155592 620 155644 672
rect 156052 620 156104 672
rect 165620 620 165672 672
rect 166264 620 166316 672
rect 173900 620 173952 672
rect 140596 552 140648 604
rect 143632 552 143684 604
rect 149244 552 149296 604
rect 151452 552 151504 604
rect 171324 552 171376 604
rect 130936 484 130988 536
rect 156972 484 157024 536
rect 160652 484 160704 536
rect 166540 484 166592 536
rect 167368 484 167420 536
rect 128452 416 128504 468
rect 155408 416 155460 468
rect 156236 416 156288 468
rect 161756 416 161808 468
rect 173532 416 173584 468
rect 119896 348 119948 400
rect 150808 348 150860 400
rect 155040 348 155092 400
rect 177856 348 177908 400
rect 129372 280 129424 332
rect 137652 280 137704 332
rect 156512 280 156564 332
rect 157524 280 157576 332
rect 129648 212 129700 264
rect 157800 212 157852 264
rect 130292 144 130344 196
rect 159088 144 159140 196
rect 159272 280 159324 332
rect 178316 280 178368 332
rect 159548 212 159600 264
rect 166908 212 166960 264
rect 170036 212 170088 264
rect 160652 144 160704 196
rect 160744 144 160796 196
rect 179604 144 179656 196
rect 129004 76 129056 128
rect 132868 76 132920 128
rect 133144 76 133196 128
rect 163044 76 163096 128
rect 163228 76 163280 128
rect 168472 76 168524 128
rect 131120 8 131172 60
rect 162584 8 162636 60
rect 162768 8 162820 60
rect 172152 8 172204 60
<< metal2 >>
rect 202 10200 258 11400
rect 570 10200 626 11400
rect 1030 10200 1086 11400
rect 1490 10200 1546 11400
rect 1858 10200 1914 11400
rect 2318 10200 2374 11400
rect 2778 10200 2834 11400
rect 3238 10200 3294 11400
rect 3606 10200 3662 11400
rect 4066 10200 4122 11400
rect 4526 10200 4582 11400
rect 4986 10200 5042 11400
rect 5354 10200 5410 11400
rect 5814 10200 5870 11400
rect 6274 10200 6330 11400
rect 6734 10200 6790 11400
rect 7102 10200 7158 11400
rect 7562 10200 7618 11400
rect 8022 10200 8078 11400
rect 8390 10200 8446 11400
rect 8850 10200 8906 11400
rect 9310 10200 9366 11400
rect 9770 10200 9826 11400
rect 10138 10200 10194 11400
rect 10598 10200 10654 11400
rect 11058 10200 11114 11400
rect 11518 10200 11574 11400
rect 11886 10200 11942 11400
rect 12346 10200 12402 11400
rect 12806 10200 12862 11400
rect 13266 10200 13322 11400
rect 13634 10200 13690 11400
rect 14094 10200 14150 11400
rect 14554 10200 14610 11400
rect 15014 10200 15070 11400
rect 15382 10200 15438 11400
rect 15842 10200 15898 11400
rect 16302 10200 16358 11400
rect 16670 10200 16726 11400
rect 17130 10200 17186 11400
rect 17590 10200 17646 11400
rect 18050 10200 18106 11400
rect 18418 10200 18474 11400
rect 18878 10200 18934 11400
rect 19338 10200 19394 11400
rect 19798 10200 19854 11400
rect 20166 10200 20222 11400
rect 20626 10200 20682 11400
rect 21086 10200 21142 11400
rect 21546 10200 21602 11400
rect 21914 10200 21970 11400
rect 22374 10200 22430 11400
rect 22834 10200 22890 11400
rect 23294 10200 23350 11400
rect 23662 10200 23718 11400
rect 24122 10200 24178 11400
rect 24582 10200 24638 11400
rect 24950 10200 25006 11400
rect 25410 10200 25466 11400
rect 25870 10200 25926 11400
rect 26330 10200 26386 11400
rect 26698 10200 26754 11400
rect 27158 10200 27214 11400
rect 27618 10200 27674 11400
rect 28078 10200 28134 11400
rect 28446 10200 28502 11400
rect 28906 10200 28962 11400
rect 29366 10200 29422 11400
rect 29826 10200 29882 11400
rect 30194 10200 30250 11400
rect 30654 10200 30710 11400
rect 31114 10200 31170 11400
rect 31574 10200 31630 11400
rect 31942 10200 31998 11400
rect 32402 10200 32458 11400
rect 32862 10200 32918 11400
rect 33230 10200 33286 11400
rect 33690 10200 33746 11400
rect 34150 10200 34206 11400
rect 34610 10200 34666 11400
rect 34978 10200 35034 11400
rect 35438 10200 35494 11400
rect 35898 10200 35954 11400
rect 36358 10200 36414 11400
rect 36726 10200 36782 11400
rect 37186 10200 37242 11400
rect 37646 10200 37702 11400
rect 38106 10200 38162 11400
rect 38474 10200 38530 11400
rect 38934 10200 38990 11400
rect 39394 10200 39450 11400
rect 39854 10200 39910 11400
rect 40222 10200 40278 11400
rect 40682 10200 40738 11400
rect 41142 10200 41198 11400
rect 41510 10200 41566 11400
rect 41970 10200 42026 11400
rect 42430 10200 42486 11400
rect 42890 10200 42946 11400
rect 43258 10200 43314 11400
rect 43718 10200 43774 11400
rect 44178 10200 44234 11400
rect 44638 10200 44694 11400
rect 45006 10200 45062 11400
rect 45466 10200 45522 11400
rect 45926 10200 45982 11400
rect 46386 10200 46442 11400
rect 46754 10200 46810 11400
rect 47214 10200 47270 11400
rect 47674 10200 47730 11400
rect 48134 10200 48190 11400
rect 48502 10200 48558 11400
rect 48962 10200 49018 11400
rect 49422 10200 49478 11400
rect 49790 10200 49846 11400
rect 50250 10200 50306 11400
rect 50710 10200 50766 11400
rect 51170 10200 51226 11400
rect 51538 10200 51594 11400
rect 51998 10200 52054 11400
rect 52458 10200 52514 11400
rect 52918 10200 52974 11400
rect 53286 10200 53342 11400
rect 53746 10200 53802 11400
rect 54206 10200 54262 11400
rect 54666 10200 54722 11400
rect 55034 10200 55090 11400
rect 55494 10200 55550 11400
rect 55954 10200 56010 11400
rect 56322 10200 56378 11400
rect 56782 10200 56838 11400
rect 57242 10200 57298 11400
rect 57702 10200 57758 11400
rect 58070 10200 58126 11400
rect 58530 10200 58586 11400
rect 58990 10200 59046 11400
rect 59450 10200 59506 11400
rect 59818 10200 59874 11400
rect 60278 10200 60334 11400
rect 60738 10200 60794 11400
rect 61198 10200 61254 11400
rect 61566 10200 61622 11400
rect 62026 10200 62082 11400
rect 62486 10200 62542 11400
rect 62946 10200 63002 11400
rect 63314 10200 63370 11400
rect 63774 10200 63830 11400
rect 64234 10200 64290 11400
rect 64602 10200 64658 11400
rect 65062 10200 65118 11400
rect 65522 10200 65578 11400
rect 65982 10200 66038 11400
rect 66350 10200 66406 11400
rect 66810 10200 66866 11400
rect 67270 10200 67326 11400
rect 67730 10200 67786 11400
rect 68098 10200 68154 11400
rect 68558 10200 68614 11400
rect 69018 10200 69074 11400
rect 69478 10200 69534 11400
rect 69846 10200 69902 11400
rect 70306 10200 70362 11400
rect 70766 10200 70822 11400
rect 71226 10200 71282 11400
rect 71594 10200 71650 11400
rect 72054 10200 72110 11400
rect 72514 10200 72570 11400
rect 72882 10200 72938 11400
rect 73342 10200 73398 11400
rect 73802 10200 73858 11400
rect 74262 10200 74318 11400
rect 74630 10200 74686 11400
rect 75090 10200 75146 11400
rect 75550 10200 75606 11400
rect 76010 10200 76066 11400
rect 76378 10200 76434 11400
rect 76838 10200 76894 11400
rect 77298 10200 77354 11400
rect 77758 10200 77814 11400
rect 78126 10200 78182 11400
rect 78586 10200 78642 11400
rect 79046 10200 79102 11400
rect 79506 10200 79562 11400
rect 79874 10200 79930 11400
rect 80334 10200 80390 11400
rect 80794 10200 80850 11400
rect 81162 10200 81218 11400
rect 81622 10200 81678 11400
rect 82082 10200 82138 11400
rect 82176 10464 82228 10470
rect 82176 10406 82228 10412
rect 216 9586 244 10200
rect 204 9580 256 9586
rect 204 9522 256 9528
rect 584 6730 612 10200
rect 1044 9722 1072 10200
rect 1032 9716 1084 9722
rect 1032 9658 1084 9664
rect 1504 9518 1532 10200
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 572 6724 624 6730
rect 572 6666 624 6672
rect 1872 6390 1900 10200
rect 2332 6662 2360 10200
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 1860 6384 1912 6390
rect 1860 6326 1912 6332
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1964 5914 1992 6190
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2792 5574 2820 10200
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2780 5568 2832 5574
rect 2976 5545 3004 6802
rect 3252 6118 3280 10200
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 8498 3372 9454
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3344 7410 3372 7754
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3620 5642 3648 10200
rect 4080 10010 4108 10200
rect 3988 9982 4108 10010
rect 3988 6730 4016 9982
rect 4076 9820 4132 9840
rect 4076 9744 4132 9764
rect 4066 9208 4122 9217
rect 4066 9143 4122 9152
rect 4080 9110 4108 9143
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 4540 8906 4568 10200
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4076 8732 4132 8752
rect 4076 8656 4132 8676
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4076 7644 4132 7664
rect 4076 7568 4132 7588
rect 4356 7410 4384 7822
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6458 3832 6598
rect 4076 6556 4132 6576
rect 4076 6480 4132 6500
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 4632 6322 4660 8910
rect 5000 8498 5028 10200
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5368 7886 5396 10200
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4724 5846 4752 6734
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 2780 5510 2832 5516
rect 2962 5536 3018 5545
rect 2962 5471 3018 5480
rect 4076 5468 4132 5488
rect 4076 5392 4132 5412
rect 4076 4380 4132 4400
rect 4076 4304 4132 4324
rect 5552 4146 5580 9454
rect 5828 8974 5856 10200
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 204 2916 256 2922
rect 204 2858 256 2864
rect 216 800 244 2858
rect 584 800 612 3470
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1032 2508 1084 2514
rect 1032 2450 1084 2456
rect 1044 800 1072 2450
rect 1504 800 1532 2926
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 800 1900 2790
rect 2332 800 2360 3538
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2792 800 2820 3402
rect 3252 800 3280 3878
rect 3620 800 3648 4014
rect 4076 3292 4132 3312
rect 4076 3216 4132 3236
rect 4076 2204 4132 2224
rect 4076 2128 4132 2148
rect 4066 1864 4122 1873
rect 4172 1850 4200 4082
rect 5644 4010 5672 8366
rect 5736 6866 5764 8366
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5736 2106 5764 4626
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5724 2100 5776 2106
rect 5724 2042 5776 2048
rect 4122 1822 4200 1850
rect 4528 1896 4580 1902
rect 4528 1838 4580 1844
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 4066 1799 4122 1808
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 3988 898 4016 1362
rect 4076 1116 4132 1136
rect 4076 1040 4132 1060
rect 3988 870 4108 898
rect 4080 800 4108 870
rect 4540 800 4568 1838
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5000 800 5028 1294
rect 5368 800 5396 1838
rect 5828 800 5856 2450
rect 5920 1562 5948 8978
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6104 3942 6132 7890
rect 6288 4622 6316 10200
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6380 2106 6408 7278
rect 6748 6798 6776 10200
rect 7116 9602 7144 10200
rect 7024 9574 7144 9602
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6932 9178 6960 9454
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 8498 6868 8910
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7024 7478 7052 9574
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7116 9178 7144 9454
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7392 8090 7420 8298
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6932 6390 6960 7210
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6736 6248 6788 6254
rect 6920 6248 6972 6254
rect 6736 6190 6788 6196
rect 6840 6196 6920 6202
rect 6840 6190 6972 6196
rect 6748 5914 6776 6190
rect 6840 6174 6960 6190
rect 6840 6118 6868 6174
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6472 2650 6500 5714
rect 6932 5234 6960 6054
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7024 4690 7052 4966
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6276 1828 6328 1834
rect 6276 1770 6328 1776
rect 5908 1556 5960 1562
rect 5908 1498 5960 1504
rect 6288 800 6316 1770
rect 6748 800 6776 2450
rect 7116 800 7144 2926
rect 7208 1562 7236 6802
rect 7300 6458 7328 7754
rect 7484 7410 7512 7822
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7576 6338 7604 10200
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7852 6662 7880 8434
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7484 6310 7604 6338
rect 7484 5710 7512 6310
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 2106 7512 5102
rect 7576 2650 7604 6190
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7852 3194 7880 6122
rect 8036 5302 8064 10200
rect 8404 6322 8432 10200
rect 8864 7868 8892 10200
rect 8772 7840 8892 7868
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 8496 5234 8524 6734
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 7944 1562 7972 5102
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 3738 8340 4626
rect 8588 4622 8616 5850
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 7196 1556 7248 1562
rect 7196 1498 7248 1504
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 7576 800 7604 1362
rect 8036 800 8064 2450
rect 8404 800 8432 3538
rect 8680 2650 8708 6802
rect 8772 6390 8800 7840
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8772 4146 8800 5578
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8864 3074 8892 7278
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8956 3194 8984 5646
rect 9324 5302 9352 10200
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9692 6866 9720 7822
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9784 6798 9812 10200
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5778 9720 6054
rect 10152 5914 10180 10200
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 10244 5574 10272 5850
rect 10612 5710 10640 10200
rect 11072 7478 11100 10200
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 9042 11284 9318
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11164 7410 11192 8230
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9692 4146 9720 4558
rect 10888 4146 10916 5646
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10980 4690 11008 4966
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9692 3738 9720 3946
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8864 3046 8984 3074
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8864 800 8892 2926
rect 8956 2106 8984 3046
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 9312 1896 9364 1902
rect 9312 1838 9364 1844
rect 9324 800 9352 1838
rect 9784 800 9812 2926
rect 9968 2106 9996 4014
rect 11072 2854 11100 7278
rect 11348 6730 11376 9522
rect 11532 8566 11560 10200
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 10140 1896 10192 1902
rect 10140 1838 10192 1844
rect 10152 800 10180 1838
rect 10612 800 10640 2450
rect 11164 2106 11192 4014
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11256 3602 11284 3946
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11440 3194 11468 8366
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11532 7954 11560 8298
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11624 3534 11652 8978
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11060 1896 11112 1902
rect 11060 1838 11112 1844
rect 11072 800 11100 1838
rect 11532 800 11560 2926
rect 11716 2650 11744 6802
rect 11808 3466 11836 7890
rect 11900 5642 11928 10200
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12268 5846 12296 8774
rect 12360 6798 12388 10200
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12452 7410 12480 7822
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 12452 4146 12480 5646
rect 12820 5642 12848 10200
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 12544 3194 12572 4626
rect 12728 3534 12756 5510
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11888 1828 11940 1834
rect 11888 1770 11940 1776
rect 11900 800 11928 1770
rect 12360 800 12388 2858
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12820 800 12848 2450
rect 13004 2378 13032 7278
rect 13280 4622 13308 10200
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13464 5914 13492 7346
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13372 4826 13400 5102
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13464 3194 13492 5714
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 12992 2372 13044 2378
rect 12992 2314 13044 2320
rect 13556 2106 13584 6190
rect 13648 5234 13676 10200
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13740 6186 13768 7278
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 14016 5778 14044 6734
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14108 5710 14136 10200
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14384 8498 14412 8910
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13268 1896 13320 1902
rect 13268 1838 13320 1844
rect 13280 800 13308 1838
rect 13648 800 13676 2382
rect 13832 2106 13860 5102
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 2650 13952 3538
rect 14200 3058 14228 7210
rect 14568 5574 14596 10200
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14844 7410 14872 7822
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 15028 6390 15056 10200
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 9178 15332 9454
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14936 3194 14964 5646
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 13820 2100 13872 2106
rect 13820 2042 13872 2048
rect 14096 1488 14148 1494
rect 14096 1430 14148 1436
rect 14108 800 14136 1430
rect 14568 800 14596 2926
rect 15212 2854 15240 8978
rect 15396 5234 15424 10200
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15580 6322 15608 7822
rect 15856 7818 15884 10200
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 16316 5642 16344 10200
rect 16684 7410 16712 10200
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16776 8498 16804 8910
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15304 4826 15332 5102
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15948 2650 15976 5102
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 15028 800 15056 2314
rect 15844 1964 15896 1970
rect 15844 1906 15896 1912
rect 15384 1896 15436 1902
rect 15384 1838 15436 1844
rect 15396 800 15424 1838
rect 15856 800 15884 1906
rect 16592 1562 16620 6802
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16684 2106 16712 6190
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 16672 1896 16724 1902
rect 16672 1838 16724 1844
rect 16580 1556 16632 1562
rect 16580 1498 16632 1504
rect 16304 1420 16356 1426
rect 16304 1362 16356 1368
rect 16316 800 16344 1362
rect 16684 800 16712 1838
rect 16868 1562 16896 7890
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16960 7002 16988 7822
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 17052 3670 17080 9454
rect 17144 6390 17172 10200
rect 17604 7546 17632 10200
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 18064 7460 18092 10200
rect 17972 7432 18092 7460
rect 17224 7268 17276 7274
rect 17224 7210 17276 7216
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 17236 2650 17264 7210
rect 17972 6798 18000 7432
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 7002 18092 7278
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18432 6322 18460 10200
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 18064 4826 18092 6190
rect 18892 5574 18920 10200
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18984 3738 19012 8366
rect 19352 6390 19380 10200
rect 19812 8566 19840 10200
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 4826 19380 5646
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 16856 1556 16908 1562
rect 16856 1498 16908 1504
rect 17236 1306 17264 2450
rect 17592 1828 17644 1834
rect 17592 1770 17644 1776
rect 17144 1278 17264 1306
rect 17144 800 17172 1278
rect 17604 800 17632 1770
rect 18064 800 18092 3538
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18432 800 18460 2926
rect 19340 2916 19392 2922
rect 19340 2858 19392 2864
rect 18880 1420 18932 1426
rect 18880 1362 18932 1368
rect 18892 800 18920 1362
rect 19352 800 19380 2858
rect 19444 2106 19472 6190
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19812 3738 19840 4014
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19996 3194 20024 5714
rect 20180 5710 20208 10200
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20456 8498 20484 8910
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20456 7410 20484 7822
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 5234 20300 5510
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20456 4826 20484 5102
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 19812 800 19840 1294
rect 20180 800 20208 2382
rect 20548 2106 20576 7210
rect 20640 6322 20668 10200
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20824 5234 20852 6190
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20732 2650 20760 5102
rect 20916 4554 20944 6326
rect 21100 5914 21128 10200
rect 21560 6118 21588 10200
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21744 6866 21772 7822
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21928 6798 21956 10200
rect 22388 7478 22416 10200
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21916 6180 21968 6186
rect 21916 6122 21968 6128
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 21100 3194 21128 5714
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21284 4826 21312 5646
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20536 2100 20588 2106
rect 20536 2042 20588 2048
rect 21640 1964 21692 1970
rect 21640 1906 21692 1912
rect 21088 1828 21140 1834
rect 21088 1770 21140 1776
rect 20628 1488 20680 1494
rect 20628 1430 20680 1436
rect 20640 800 20668 1430
rect 21100 800 21128 1770
rect 21456 1760 21508 1766
rect 21456 1702 21508 1708
rect 21468 1426 21496 1702
rect 21456 1420 21508 1426
rect 21456 1362 21508 1368
rect 21652 1034 21680 1906
rect 21928 1562 21956 6122
rect 22020 1562 22048 7278
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22388 2650 22416 6802
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22480 5234 22508 6054
rect 22848 5574 22876 10200
rect 23308 5642 23336 10200
rect 23676 8650 23704 10200
rect 24136 9466 24164 10200
rect 24136 9438 24256 9466
rect 24076 9276 24132 9296
rect 24076 9200 24132 9220
rect 23676 8622 23796 8650
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23584 6866 23612 7822
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23676 6322 23704 7142
rect 23768 6798 23796 8622
rect 24076 8188 24132 8208
rect 24076 8112 24132 8132
rect 24228 7274 24256 9438
rect 24216 7268 24268 7274
rect 24216 7210 24268 7216
rect 24076 7100 24132 7120
rect 24076 7024 24132 7044
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 24076 6012 24132 6032
rect 24076 5936 24132 5956
rect 24596 5846 24624 10200
rect 24964 8650 24992 10200
rect 24964 8622 25084 8650
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24964 8090 24992 8366
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24872 7410 24900 7822
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 23296 5636 23348 5642
rect 23296 5578 23348 5584
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 23492 4146 23520 5102
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 22744 4072 22796 4078
rect 22744 4014 22796 4020
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22756 2922 22784 4014
rect 22848 3738 22876 4014
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 23296 2508 23348 2514
rect 23296 2450 23348 2456
rect 22836 1828 22888 1834
rect 22836 1770 22888 1776
rect 21916 1556 21968 1562
rect 21916 1498 21968 1504
rect 22008 1556 22060 1562
rect 22008 1498 22060 1504
rect 21916 1352 21968 1358
rect 21916 1294 21968 1300
rect 22560 1352 22612 1358
rect 22560 1294 22612 1300
rect 21560 1006 21680 1034
rect 21560 800 21588 1006
rect 21928 800 21956 1294
rect 22572 898 22600 1294
rect 22388 870 22600 898
rect 22388 800 22416 870
rect 22848 800 22876 1770
rect 23308 800 23336 2450
rect 23584 2106 23612 4626
rect 23572 2100 23624 2106
rect 23572 2042 23624 2048
rect 23768 1766 23796 5102
rect 24076 4924 24132 4944
rect 24076 4848 24132 4868
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23860 3738 23888 4558
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24076 3836 24132 3856
rect 24076 3760 24132 3780
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 24076 2748 24132 2768
rect 24076 2672 24132 2692
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 23756 1760 23808 1766
rect 23756 1702 23808 1708
rect 24076 1660 24132 1680
rect 24076 1584 24132 1604
rect 24228 1306 24256 2450
rect 24780 2038 24808 4014
rect 24872 2650 24900 6190
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 24768 2032 24820 2038
rect 24768 1974 24820 1980
rect 24584 1964 24636 1970
rect 24584 1906 24636 1912
rect 23664 1284 23716 1290
rect 23664 1226 23716 1232
rect 24136 1278 24256 1306
rect 23676 800 23704 1226
rect 24136 800 24164 1278
rect 24596 800 24624 1906
rect 24964 1562 24992 6802
rect 25056 6322 25084 8622
rect 25136 7812 25188 7818
rect 25136 7754 25188 7760
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25044 5772 25096 5778
rect 25044 5714 25096 5720
rect 25056 2106 25084 5714
rect 25148 2650 25176 7754
rect 25424 7478 25452 10200
rect 25884 7886 25912 10200
rect 26056 8424 26108 8430
rect 26056 8366 26108 8372
rect 25872 7880 25924 7886
rect 25872 7822 25924 7828
rect 25412 7472 25464 7478
rect 25412 7414 25464 7420
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 25240 4146 25268 5510
rect 25228 4140 25280 4146
rect 25228 4082 25280 4088
rect 25136 2644 25188 2650
rect 25136 2586 25188 2592
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25044 2100 25096 2106
rect 25044 2042 25096 2048
rect 24952 1556 25004 1562
rect 24952 1498 25004 1504
rect 25148 1306 25176 2450
rect 25332 1562 25360 6938
rect 26068 3738 26096 8366
rect 26344 6322 26372 10200
rect 26712 6798 26740 10200
rect 27068 9104 27120 9110
rect 27068 9046 27120 9052
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26884 6384 26936 6390
rect 26884 6326 26936 6332
rect 26332 6316 26384 6322
rect 26332 6258 26384 6264
rect 26896 3942 26924 6326
rect 26976 4616 27028 4622
rect 26976 4558 27028 4564
rect 26988 4146 27016 4558
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 26332 3596 26384 3602
rect 26332 3538 26384 3544
rect 25412 3120 25464 3126
rect 25412 3062 25464 3068
rect 25320 1556 25372 1562
rect 25320 1498 25372 1504
rect 24964 1278 25176 1306
rect 24964 800 24992 1278
rect 25424 800 25452 3062
rect 25872 2984 25924 2990
rect 25872 2926 25924 2932
rect 25884 800 25912 2926
rect 26344 800 26372 3538
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 26528 3058 26556 3402
rect 27080 3194 27108 9046
rect 27172 6458 27200 10200
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 27356 7954 27384 8230
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 27264 6866 27292 7142
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 27632 6390 27660 10200
rect 27896 9376 27948 9382
rect 27896 9318 27948 9324
rect 27908 9042 27936 9318
rect 27896 9036 27948 9042
rect 27896 8978 27948 8984
rect 28092 8566 28120 10200
rect 28080 8560 28132 8566
rect 28080 8502 28132 8508
rect 28460 6866 28488 10200
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 28448 6860 28500 6866
rect 28448 6802 28500 6808
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27632 5914 27660 6190
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 27160 3596 27212 3602
rect 27160 3538 27212 3544
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 26712 800 26740 2994
rect 27172 800 27200 3538
rect 27724 2650 27752 6802
rect 27896 6248 27948 6254
rect 27896 6190 27948 6196
rect 27712 2644 27764 2650
rect 27712 2586 27764 2592
rect 27908 2106 27936 6190
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28276 3738 28304 4558
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 27896 2100 27948 2106
rect 27896 2042 27948 2048
rect 28080 1896 28132 1902
rect 28080 1838 28132 1844
rect 27620 1760 27672 1766
rect 27620 1702 27672 1708
rect 27632 800 27660 1702
rect 28092 800 28120 1838
rect 28460 800 28488 2450
rect 28552 1562 28580 7142
rect 28632 6792 28684 6798
rect 28632 6734 28684 6740
rect 28644 5778 28672 6734
rect 28920 6662 28948 10200
rect 29276 8968 29328 8974
rect 29276 8910 29328 8916
rect 29288 8498 29316 8910
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29092 8424 29144 8430
rect 29092 8366 29144 8372
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 28632 5772 28684 5778
rect 28632 5714 28684 5720
rect 29104 3466 29132 8366
rect 29380 6390 29408 10200
rect 29552 8016 29604 8022
rect 29552 7958 29604 7964
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29472 7410 29500 7822
rect 29460 7404 29512 7410
rect 29460 7346 29512 7352
rect 29368 6384 29420 6390
rect 29368 6326 29420 6332
rect 29368 5160 29420 5166
rect 29368 5102 29420 5108
rect 29380 4146 29408 5102
rect 29368 4140 29420 4146
rect 29368 4082 29420 4088
rect 29092 3460 29144 3466
rect 29092 3402 29144 3408
rect 29564 3194 29592 7958
rect 29644 6792 29696 6798
rect 29644 6734 29696 6740
rect 29656 6322 29684 6734
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 29840 6118 29868 10200
rect 30208 6730 30236 10200
rect 30288 7812 30340 7818
rect 30288 7754 30340 7760
rect 30300 6866 30328 7754
rect 30564 7336 30616 7342
rect 30564 7278 30616 7284
rect 30576 7002 30604 7278
rect 30564 6996 30616 7002
rect 30564 6938 30616 6944
rect 30288 6860 30340 6866
rect 30288 6802 30340 6808
rect 30196 6724 30248 6730
rect 30196 6666 30248 6672
rect 30668 6202 30696 10200
rect 31128 8974 31156 10200
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31588 8566 31616 10200
rect 31576 8560 31628 8566
rect 31576 8502 31628 8508
rect 31852 7880 31904 7886
rect 31852 7822 31904 7828
rect 31864 7410 31892 7822
rect 31852 7404 31904 7410
rect 31852 7346 31904 7352
rect 30300 6174 30696 6202
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 29736 5772 29788 5778
rect 29736 5714 29788 5720
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29368 2916 29420 2922
rect 29368 2858 29420 2864
rect 28908 1828 28960 1834
rect 28908 1770 28960 1776
rect 28540 1556 28592 1562
rect 28540 1498 28592 1504
rect 28920 800 28948 1770
rect 29380 800 29408 2858
rect 29748 1970 29776 5714
rect 30300 4214 30328 6174
rect 30380 6112 30432 6118
rect 30380 6054 30432 6060
rect 30392 5234 30420 6054
rect 31956 5778 31984 10200
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 32220 8968 32272 8974
rect 32220 8910 32272 8916
rect 32140 7954 32168 8910
rect 32232 8498 32260 8910
rect 32220 8492 32272 8498
rect 32220 8434 32272 8440
rect 32128 7948 32180 7954
rect 32128 7890 32180 7896
rect 32416 6882 32444 10200
rect 32588 8016 32640 8022
rect 32588 7958 32640 7964
rect 32324 6854 32444 6882
rect 30564 5772 30616 5778
rect 30564 5714 30616 5720
rect 31944 5772 31996 5778
rect 31944 5714 31996 5720
rect 30380 5228 30432 5234
rect 30380 5170 30432 5176
rect 30472 5160 30524 5166
rect 30472 5102 30524 5108
rect 30288 4208 30340 4214
rect 30288 4150 30340 4156
rect 30196 4072 30248 4078
rect 30196 4014 30248 4020
rect 29828 3120 29880 3126
rect 29828 3062 29880 3068
rect 29736 1964 29788 1970
rect 29736 1906 29788 1912
rect 29840 800 29868 3062
rect 30208 2038 30236 4014
rect 30484 2106 30512 5102
rect 30576 4622 30604 5714
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 31772 5234 31800 5646
rect 32324 5234 32352 6854
rect 32404 6248 32456 6254
rect 32404 6190 32456 6196
rect 32416 5914 32444 6190
rect 32404 5908 32456 5914
rect 32404 5850 32456 5856
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 32312 5228 32364 5234
rect 32312 5170 32364 5176
rect 32312 4684 32364 4690
rect 32312 4626 32364 4632
rect 30564 4616 30616 4622
rect 30564 4558 30616 4564
rect 30748 4616 30800 4622
rect 30748 4558 30800 4564
rect 30760 4146 30788 4558
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 31116 2916 31168 2922
rect 31116 2858 31168 2864
rect 30472 2100 30524 2106
rect 30472 2042 30524 2048
rect 30196 2032 30248 2038
rect 30196 1974 30248 1980
rect 30288 1964 30340 1970
rect 30288 1906 30340 1912
rect 30300 1034 30328 1906
rect 30656 1420 30708 1426
rect 30656 1362 30708 1368
rect 30208 1006 30328 1034
rect 30208 800 30236 1006
rect 30668 800 30696 1362
rect 31128 800 31156 2858
rect 31588 800 31616 2994
rect 32324 2106 32352 4626
rect 32600 3194 32628 7958
rect 32772 6180 32824 6186
rect 32772 6122 32824 6128
rect 32588 3188 32640 3194
rect 32588 3130 32640 3136
rect 32784 2106 32812 6122
rect 32876 5642 32904 10200
rect 33244 8786 33272 10200
rect 33244 8758 33364 8786
rect 33232 8492 33284 8498
rect 33232 8434 33284 8440
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 32864 5636 32916 5642
rect 32864 5578 32916 5584
rect 32956 5160 33008 5166
rect 32956 5102 33008 5108
rect 32312 2100 32364 2106
rect 32312 2042 32364 2048
rect 32772 2100 32824 2106
rect 32772 2042 32824 2048
rect 31944 1964 31996 1970
rect 31944 1906 31996 1912
rect 31956 800 31984 1906
rect 32864 1828 32916 1834
rect 32864 1770 32916 1776
rect 32404 1488 32456 1494
rect 32404 1430 32456 1436
rect 32416 800 32444 1430
rect 32876 800 32904 1770
rect 32968 1562 32996 5102
rect 33060 3670 33088 8366
rect 33244 6662 33272 8434
rect 33336 7410 33364 8758
rect 33324 7404 33376 7410
rect 33324 7346 33376 7352
rect 33324 6860 33376 6866
rect 33324 6802 33376 6808
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 33048 3664 33100 3670
rect 33048 3606 33100 3612
rect 33140 2984 33192 2990
rect 33192 2944 33272 2972
rect 33140 2926 33192 2932
rect 33048 2848 33100 2854
rect 33048 2790 33100 2796
rect 32956 1556 33008 1562
rect 32956 1498 33008 1504
rect 33060 1426 33088 2790
rect 33048 1420 33100 1426
rect 33048 1362 33100 1368
rect 33244 800 33272 2944
rect 33336 2650 33364 6802
rect 33600 5772 33652 5778
rect 33600 5714 33652 5720
rect 33508 4616 33560 4622
rect 33508 4558 33560 4564
rect 33520 4146 33548 4558
rect 33508 4140 33560 4146
rect 33508 4082 33560 4088
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 33324 2644 33376 2650
rect 33324 2586 33376 2592
rect 33428 2038 33456 4014
rect 33612 3194 33640 5714
rect 33704 4622 33732 10200
rect 34164 8498 34192 10200
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 33968 6860 34020 6866
rect 33968 6802 34020 6808
rect 33876 6248 33928 6254
rect 33876 6190 33928 6196
rect 33692 4616 33744 4622
rect 33692 4558 33744 4564
rect 33784 4616 33836 4622
rect 33784 4558 33836 4564
rect 33796 3602 33824 4558
rect 33784 3596 33836 3602
rect 33784 3538 33836 3544
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 33692 2508 33744 2514
rect 33692 2450 33744 2456
rect 33416 2032 33468 2038
rect 33416 1974 33468 1980
rect 33704 800 33732 2450
rect 33888 1562 33916 6190
rect 33980 3534 34008 6802
rect 34624 5846 34652 10200
rect 34888 8288 34940 8294
rect 34888 8230 34940 8236
rect 34900 7954 34928 8230
rect 34888 7948 34940 7954
rect 34888 7890 34940 7896
rect 34992 7886 35020 10200
rect 34980 7880 35032 7886
rect 34980 7822 35032 7828
rect 35452 6390 35480 10200
rect 35912 6866 35940 10200
rect 35992 8356 36044 8362
rect 35992 8298 36044 8304
rect 35900 6860 35952 6866
rect 35900 6802 35952 6808
rect 35440 6384 35492 6390
rect 35440 6326 35492 6332
rect 34336 5840 34388 5846
rect 34336 5782 34388 5788
rect 34612 5840 34664 5846
rect 34612 5782 34664 5788
rect 34348 4214 34376 5782
rect 34888 5704 34940 5710
rect 34888 5646 34940 5652
rect 34900 5234 34928 5646
rect 34888 5228 34940 5234
rect 34888 5170 34940 5176
rect 34980 4684 35032 4690
rect 34980 4626 35032 4632
rect 34336 4208 34388 4214
rect 34336 4150 34388 4156
rect 34520 3596 34572 3602
rect 34520 3538 34572 3544
rect 33968 3528 34020 3534
rect 33968 3470 34020 3476
rect 34532 2582 34560 3538
rect 34612 3460 34664 3466
rect 34612 3402 34664 3408
rect 34520 2576 34572 2582
rect 34520 2518 34572 2524
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 33876 1556 33928 1562
rect 33876 1498 33928 1504
rect 34164 800 34192 2382
rect 34624 800 34652 3402
rect 34992 2106 35020 4626
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 34980 2100 35032 2106
rect 34980 2042 35032 2048
rect 34980 1352 35032 1358
rect 34980 1294 35032 1300
rect 34992 800 35020 1294
rect 35452 800 35480 2994
rect 35900 1828 35952 1834
rect 35900 1770 35952 1776
rect 35912 800 35940 1770
rect 36004 1562 36032 8298
rect 36372 6458 36400 10200
rect 36360 6452 36412 6458
rect 36360 6394 36412 6400
rect 36084 6248 36136 6254
rect 36084 6190 36136 6196
rect 36544 6248 36596 6254
rect 36544 6190 36596 6196
rect 36096 5914 36124 6190
rect 36084 5908 36136 5914
rect 36084 5850 36136 5856
rect 36084 5160 36136 5166
rect 36084 5102 36136 5108
rect 36096 4826 36124 5102
rect 36084 4820 36136 4826
rect 36084 4762 36136 4768
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 35992 1556 36044 1562
rect 35992 1498 36044 1504
rect 36372 800 36400 2994
rect 36556 2650 36584 6190
rect 36740 5778 36768 10200
rect 37200 6730 37228 10200
rect 37556 8424 37608 8430
rect 37556 8366 37608 8372
rect 37568 8090 37596 8366
rect 37556 8084 37608 8090
rect 37556 8026 37608 8032
rect 37188 6724 37240 6730
rect 37188 6666 37240 6672
rect 37660 6390 37688 10200
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 37924 7336 37976 7342
rect 37924 7278 37976 7284
rect 37752 6866 37780 7278
rect 37740 6860 37792 6866
rect 37740 6802 37792 6808
rect 37832 6792 37884 6798
rect 37832 6734 37884 6740
rect 37648 6384 37700 6390
rect 37648 6326 37700 6332
rect 37844 6322 37872 6734
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 36728 5772 36780 5778
rect 36728 5714 36780 5720
rect 37740 5704 37792 5710
rect 37740 5646 37792 5652
rect 37752 4826 37780 5646
rect 37740 4820 37792 4826
rect 37740 4762 37792 4768
rect 37648 3596 37700 3602
rect 37648 3538 37700 3544
rect 37188 3120 37240 3126
rect 37188 3062 37240 3068
rect 36544 2644 36596 2650
rect 36544 2586 36596 2592
rect 36728 1760 36780 1766
rect 36728 1702 36780 1708
rect 36740 800 36768 1702
rect 37200 800 37228 3062
rect 37660 800 37688 3538
rect 37740 2916 37792 2922
rect 37740 2858 37792 2864
rect 37752 1902 37780 2858
rect 37936 2106 37964 7278
rect 38120 6848 38148 10200
rect 38292 9036 38344 9042
rect 38292 8978 38344 8984
rect 38200 6860 38252 6866
rect 38120 6820 38200 6848
rect 38200 6802 38252 6808
rect 38304 3738 38332 8978
rect 38488 5302 38516 10200
rect 38948 7818 38976 10200
rect 39408 8974 39436 10200
rect 39120 8968 39172 8974
rect 39120 8910 39172 8916
rect 39396 8968 39448 8974
rect 39396 8910 39448 8916
rect 39132 8498 39160 8910
rect 39120 8492 39172 8498
rect 39120 8434 39172 8440
rect 38936 7812 38988 7818
rect 38936 7754 38988 7760
rect 39396 6248 39448 6254
rect 39396 6190 39448 6196
rect 39120 5772 39172 5778
rect 39120 5714 39172 5720
rect 38476 5296 38528 5302
rect 38476 5238 38528 5244
rect 38292 3732 38344 3738
rect 38292 3674 38344 3680
rect 38476 2984 38528 2990
rect 38476 2926 38528 2932
rect 37924 2100 37976 2106
rect 37924 2042 37976 2048
rect 37740 1896 37792 1902
rect 37740 1838 37792 1844
rect 38108 1488 38160 1494
rect 38108 1430 38160 1436
rect 38120 800 38148 1430
rect 38488 800 38516 2926
rect 38936 2440 38988 2446
rect 38936 2382 38988 2388
rect 38948 800 38976 2382
rect 39132 1562 39160 5714
rect 39408 2106 39436 6190
rect 39868 6186 39896 10200
rect 40236 8906 40264 10200
rect 40224 8900 40276 8906
rect 40224 8842 40276 8848
rect 39948 7336 40000 7342
rect 39948 7278 40000 7284
rect 39960 6866 39988 7278
rect 39948 6860 40000 6866
rect 39948 6802 40000 6808
rect 40696 6798 40724 10200
rect 40960 9512 41012 9518
rect 40960 9454 41012 9460
rect 40868 9376 40920 9382
rect 40868 9318 40920 9324
rect 40880 9042 40908 9318
rect 40868 9036 40920 9042
rect 40868 8978 40920 8984
rect 40972 8498 41000 9454
rect 40960 8492 41012 8498
rect 40960 8434 41012 8440
rect 41156 7478 41184 10200
rect 41328 9104 41380 9110
rect 41328 9046 41380 9052
rect 41144 7472 41196 7478
rect 41144 7414 41196 7420
rect 40684 6792 40736 6798
rect 40684 6734 40736 6740
rect 39856 6180 39908 6186
rect 39856 6122 39908 6128
rect 40132 5704 40184 5710
rect 40132 5646 40184 5652
rect 40144 5234 40172 5646
rect 40132 5228 40184 5234
rect 40132 5170 40184 5176
rect 41144 5160 41196 5166
rect 41144 5102 41196 5108
rect 40776 4616 40828 4622
rect 40776 4558 40828 4564
rect 40788 4146 40816 4558
rect 40776 4140 40828 4146
rect 40776 4082 40828 4088
rect 39856 3596 39908 3602
rect 39856 3538 39908 3544
rect 39488 2916 39540 2922
rect 39488 2858 39540 2864
rect 39396 2100 39448 2106
rect 39396 2042 39448 2048
rect 39120 1556 39172 1562
rect 39120 1498 39172 1504
rect 39500 1442 39528 2858
rect 39408 1414 39528 1442
rect 39408 800 39436 1414
rect 39868 800 39896 3538
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 40224 2372 40276 2378
rect 40224 2314 40276 2320
rect 40236 800 40264 2314
rect 40696 800 40724 3334
rect 41156 2106 41184 5102
rect 41236 3528 41288 3534
rect 41236 3470 41288 3476
rect 41144 2100 41196 2106
rect 41144 2042 41196 2048
rect 41248 1442 41276 3470
rect 41340 3194 41368 9046
rect 41420 8492 41472 8498
rect 41420 8434 41472 8440
rect 41432 6730 41460 8434
rect 41524 7750 41552 10200
rect 41984 8650 42012 10200
rect 41984 8622 42104 8650
rect 41972 8424 42024 8430
rect 41972 8366 42024 8372
rect 41984 8090 42012 8366
rect 41972 8084 42024 8090
rect 41972 8026 42024 8032
rect 41880 7880 41932 7886
rect 41880 7822 41932 7828
rect 41512 7744 41564 7750
rect 41512 7686 41564 7692
rect 41892 7410 41920 7822
rect 41880 7404 41932 7410
rect 41880 7346 41932 7352
rect 41420 6724 41472 6730
rect 41420 6666 41472 6672
rect 41972 5704 42024 5710
rect 41972 5646 42024 5652
rect 41984 4146 42012 5646
rect 42076 4622 42104 8622
rect 42444 6934 42472 10200
rect 42904 9330 42932 10200
rect 42720 9302 42932 9330
rect 42720 8974 42748 9302
rect 42708 8968 42760 8974
rect 42708 8910 42760 8916
rect 42892 7336 42944 7342
rect 42892 7278 42944 7284
rect 42432 6928 42484 6934
rect 42432 6870 42484 6876
rect 42904 6866 42932 7278
rect 43076 7268 43128 7274
rect 43076 7210 43128 7216
rect 42892 6860 42944 6866
rect 42892 6802 42944 6808
rect 42616 6792 42668 6798
rect 42616 6734 42668 6740
rect 42628 6322 42656 6734
rect 42616 6316 42668 6322
rect 42616 6258 42668 6264
rect 42340 5160 42392 5166
rect 42340 5102 42392 5108
rect 42064 4616 42116 4622
rect 42064 4558 42116 4564
rect 41972 4140 42024 4146
rect 41972 4082 42024 4088
rect 41420 3460 41472 3466
rect 41420 3402 41472 3408
rect 41328 3188 41380 3194
rect 41328 3130 41380 3136
rect 41432 1970 41460 3402
rect 41604 2848 41656 2854
rect 41604 2790 41656 2796
rect 41972 2848 42024 2854
rect 41972 2790 42024 2796
rect 41420 1964 41472 1970
rect 41420 1906 41472 1912
rect 41512 1828 41564 1834
rect 41512 1770 41564 1776
rect 41156 1414 41276 1442
rect 41156 800 41184 1414
rect 41524 800 41552 1770
rect 41616 1426 41644 2790
rect 41604 1420 41656 1426
rect 41604 1362 41656 1368
rect 41984 800 42012 2790
rect 42352 2106 42380 5102
rect 42800 4684 42852 4690
rect 42800 4626 42852 4632
rect 42432 2916 42484 2922
rect 42432 2858 42484 2864
rect 42340 2100 42392 2106
rect 42340 2042 42392 2048
rect 42444 800 42472 2858
rect 42812 2854 42840 4626
rect 43088 3194 43116 7210
rect 43272 5574 43300 10200
rect 43732 9586 43760 10200
rect 44076 9820 44132 9840
rect 44076 9744 44132 9764
rect 43720 9580 43772 9586
rect 43720 9522 43772 9528
rect 43628 9444 43680 9450
rect 43628 9386 43680 9392
rect 43444 9036 43496 9042
rect 43444 8978 43496 8984
rect 43260 5568 43312 5574
rect 43260 5510 43312 5516
rect 43352 4072 43404 4078
rect 43352 4014 43404 4020
rect 43076 3188 43128 3194
rect 43076 3130 43128 3136
rect 43076 3052 43128 3058
rect 43076 2994 43128 3000
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42892 1896 42944 1902
rect 42892 1838 42944 1844
rect 42904 800 42932 1838
rect 43088 1494 43116 2994
rect 43364 2650 43392 4014
rect 43456 3738 43484 8978
rect 43536 8424 43588 8430
rect 43536 8366 43588 8372
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 43444 3120 43496 3126
rect 43444 3062 43496 3068
rect 43352 2644 43404 2650
rect 43352 2586 43404 2592
rect 43260 2508 43312 2514
rect 43260 2450 43312 2456
rect 43076 1488 43128 1494
rect 43076 1430 43128 1436
rect 43272 800 43300 2450
rect 43456 1902 43484 3062
rect 43548 1986 43576 8366
rect 43640 4826 43668 9386
rect 43812 9104 43864 9110
rect 43812 9046 43864 9052
rect 43720 8968 43772 8974
rect 43720 8910 43772 8916
rect 43732 8498 43760 8910
rect 43720 8492 43772 8498
rect 43720 8434 43772 8440
rect 43720 6384 43772 6390
rect 43720 6326 43772 6332
rect 43732 5302 43760 6326
rect 43720 5296 43772 5302
rect 43720 5238 43772 5244
rect 43628 4820 43680 4826
rect 43628 4762 43680 4768
rect 43824 3194 43852 9046
rect 44192 8974 44220 10200
rect 44180 8968 44232 8974
rect 44180 8910 44232 8916
rect 44076 8732 44132 8752
rect 44076 8656 44132 8676
rect 44364 8288 44416 8294
rect 44364 8230 44416 8236
rect 44376 7954 44404 8230
rect 44364 7948 44416 7954
rect 44364 7890 44416 7896
rect 44456 7948 44508 7954
rect 44456 7890 44508 7896
rect 44076 7644 44132 7664
rect 44076 7568 44132 7588
rect 44076 6556 44132 6576
rect 44076 6480 44132 6500
rect 43996 6248 44048 6254
rect 43996 6190 44048 6196
rect 44272 6248 44324 6254
rect 44272 6190 44324 6196
rect 44008 5914 44036 6190
rect 43996 5908 44048 5914
rect 43996 5850 44048 5856
rect 44076 5468 44132 5488
rect 44076 5392 44132 5412
rect 44076 4380 44132 4400
rect 44076 4304 44132 4324
rect 44076 3292 44132 3312
rect 44076 3216 44132 3236
rect 43812 3188 43864 3194
rect 43812 3130 43864 3136
rect 43720 2848 43772 2854
rect 43720 2790 43772 2796
rect 44180 2848 44232 2854
rect 44180 2790 44232 2796
rect 43548 1958 43668 1986
rect 43444 1896 43496 1902
rect 43444 1838 43496 1844
rect 43536 1760 43588 1766
rect 43536 1702 43588 1708
rect 43548 1562 43576 1702
rect 43640 1562 43668 1958
rect 43536 1556 43588 1562
rect 43536 1498 43588 1504
rect 43628 1556 43680 1562
rect 43628 1498 43680 1504
rect 43732 800 43760 2790
rect 44076 2204 44132 2224
rect 44076 2128 44132 2148
rect 44076 1116 44132 1136
rect 44076 1040 44132 1060
rect 44192 800 44220 2790
rect 44284 2106 44312 6190
rect 44364 4616 44416 4622
rect 44364 4558 44416 4564
rect 44376 2650 44404 4558
rect 44364 2644 44416 2650
rect 44364 2586 44416 2592
rect 44468 2106 44496 7890
rect 44652 6390 44680 10200
rect 44640 6384 44692 6390
rect 44640 6326 44692 6332
rect 44548 5160 44600 5166
rect 44548 5102 44600 5108
rect 44560 4146 44588 5102
rect 45020 4214 45048 10200
rect 45376 7336 45428 7342
rect 45376 7278 45428 7284
rect 45100 4616 45152 4622
rect 45100 4558 45152 4564
rect 45008 4208 45060 4214
rect 45008 4150 45060 4156
rect 44548 4140 44600 4146
rect 44548 4082 44600 4088
rect 44732 4072 44784 4078
rect 44732 4014 44784 4020
rect 44640 3936 44692 3942
rect 44640 3878 44692 3884
rect 44652 3602 44680 3878
rect 44640 3596 44692 3602
rect 44640 3538 44692 3544
rect 44744 2122 44772 4014
rect 45112 3058 45140 4558
rect 45192 3392 45244 3398
rect 45192 3334 45244 3340
rect 45204 3058 45232 3334
rect 45100 3052 45152 3058
rect 45100 2994 45152 3000
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45008 2984 45060 2990
rect 45008 2926 45060 2932
rect 44272 2100 44324 2106
rect 44272 2042 44324 2048
rect 44456 2100 44508 2106
rect 44456 2042 44508 2048
rect 44652 2094 44772 2122
rect 44652 800 44680 2094
rect 45020 800 45048 2926
rect 45388 1562 45416 7278
rect 45480 6118 45508 10200
rect 45560 6860 45612 6866
rect 45560 6802 45612 6808
rect 45468 6112 45520 6118
rect 45468 6054 45520 6060
rect 45572 2650 45600 6802
rect 45940 6798 45968 10200
rect 46112 9376 46164 9382
rect 46112 9318 46164 9324
rect 46124 7342 46152 9318
rect 46400 8566 46428 10200
rect 46388 8560 46440 8566
rect 46388 8502 46440 8508
rect 46480 8424 46532 8430
rect 46480 8366 46532 8372
rect 46112 7336 46164 7342
rect 46112 7278 46164 7284
rect 45928 6792 45980 6798
rect 45928 6734 45980 6740
rect 46112 6248 46164 6254
rect 46112 6190 46164 6196
rect 46124 5914 46152 6190
rect 46112 5908 46164 5914
rect 46112 5850 46164 5856
rect 45652 5568 45704 5574
rect 45652 5510 45704 5516
rect 45664 3534 45692 5510
rect 46112 5160 46164 5166
rect 46112 5102 46164 5108
rect 46124 4826 46152 5102
rect 46112 4820 46164 4826
rect 46112 4762 46164 4768
rect 46492 4146 46520 8366
rect 46768 5846 46796 10200
rect 46940 9376 46992 9382
rect 46940 9318 46992 9324
rect 46952 8974 46980 9318
rect 46940 8968 46992 8974
rect 46940 8910 46992 8916
rect 47032 6248 47084 6254
rect 47032 6190 47084 6196
rect 46756 5840 46808 5846
rect 46756 5782 46808 5788
rect 46572 5772 46624 5778
rect 46572 5714 46624 5720
rect 46480 4140 46532 4146
rect 46480 4082 46532 4088
rect 46204 3596 46256 3602
rect 46204 3538 46256 3544
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 45928 2916 45980 2922
rect 45928 2858 45980 2864
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 45560 2644 45612 2650
rect 45560 2586 45612 2592
rect 45664 2514 45692 2790
rect 45652 2508 45704 2514
rect 45652 2450 45704 2456
rect 45468 2440 45520 2446
rect 45468 2382 45520 2388
rect 45376 1556 45428 1562
rect 45376 1498 45428 1504
rect 45480 800 45508 2382
rect 45940 800 45968 2858
rect 46216 2106 46244 3538
rect 46584 2650 46612 5714
rect 46756 3596 46808 3602
rect 46756 3538 46808 3544
rect 46572 2644 46624 2650
rect 46572 2586 46624 2592
rect 46204 2100 46256 2106
rect 46204 2042 46256 2048
rect 46388 1896 46440 1902
rect 46388 1838 46440 1844
rect 46400 800 46428 1838
rect 46768 800 46796 3538
rect 47044 1766 47072 6190
rect 47124 5840 47176 5846
rect 47124 5782 47176 5788
rect 47136 5234 47164 5782
rect 47228 5642 47256 10200
rect 47584 8968 47636 8974
rect 47584 8910 47636 8916
rect 47596 8498 47624 8910
rect 47584 8492 47636 8498
rect 47584 8434 47636 8440
rect 47308 8016 47360 8022
rect 47308 7958 47360 7964
rect 47320 6866 47348 7958
rect 47400 7948 47452 7954
rect 47400 7890 47452 7896
rect 47308 6860 47360 6866
rect 47308 6802 47360 6808
rect 47216 5636 47268 5642
rect 47216 5578 47268 5584
rect 47124 5228 47176 5234
rect 47124 5170 47176 5176
rect 47216 5160 47268 5166
rect 47216 5102 47268 5108
rect 47228 3194 47256 5102
rect 47308 4684 47360 4690
rect 47308 4626 47360 4632
rect 47216 3188 47268 3194
rect 47216 3130 47268 3136
rect 47320 2106 47348 4626
rect 47412 3670 47440 7890
rect 47584 6860 47636 6866
rect 47584 6802 47636 6808
rect 47400 3664 47452 3670
rect 47400 3606 47452 3612
rect 47400 3528 47452 3534
rect 47400 3470 47452 3476
rect 47308 2100 47360 2106
rect 47308 2042 47360 2048
rect 47412 1850 47440 3470
rect 47492 3052 47544 3058
rect 47492 2994 47544 3000
rect 47228 1822 47440 1850
rect 47032 1760 47084 1766
rect 47032 1702 47084 1708
rect 47228 800 47256 1822
rect 47504 1426 47532 2994
rect 47596 2582 47624 6802
rect 47688 6798 47716 10200
rect 47676 6792 47728 6798
rect 47676 6734 47728 6740
rect 47768 5092 47820 5098
rect 47768 5034 47820 5040
rect 47780 2650 47808 5034
rect 48148 4622 48176 10200
rect 48516 8634 48544 10200
rect 48976 9058 49004 10200
rect 48976 9042 49096 9058
rect 48976 9036 49108 9042
rect 48976 9030 49056 9036
rect 49056 8978 49108 8984
rect 48504 8628 48556 8634
rect 48504 8570 48556 8576
rect 48964 8356 49016 8362
rect 48964 8298 49016 8304
rect 48976 6866 49004 8298
rect 49240 7880 49292 7886
rect 49240 7822 49292 7828
rect 49252 7410 49280 7822
rect 49240 7404 49292 7410
rect 49240 7346 49292 7352
rect 49332 7404 49384 7410
rect 49332 7346 49384 7352
rect 49344 6934 49372 7346
rect 49332 6928 49384 6934
rect 49332 6870 49384 6876
rect 48964 6860 49016 6866
rect 48964 6802 49016 6808
rect 49148 6860 49200 6866
rect 49148 6802 49200 6808
rect 48504 6248 48556 6254
rect 48504 6190 48556 6196
rect 48516 5234 48544 6190
rect 48504 5228 48556 5234
rect 48504 5170 48556 5176
rect 48136 4616 48188 4622
rect 48136 4558 48188 4564
rect 48964 4616 49016 4622
rect 48964 4558 49016 4564
rect 48976 4146 49004 4558
rect 48964 4140 49016 4146
rect 48964 4082 49016 4088
rect 48964 4004 49016 4010
rect 48964 3946 49016 3952
rect 47768 2644 47820 2650
rect 47768 2586 47820 2592
rect 47584 2576 47636 2582
rect 47584 2518 47636 2524
rect 48136 2508 48188 2514
rect 48136 2450 48188 2456
rect 48504 2508 48556 2514
rect 48504 2450 48556 2456
rect 47676 1896 47728 1902
rect 47676 1838 47728 1844
rect 47492 1420 47544 1426
rect 47492 1362 47544 1368
rect 47688 800 47716 1838
rect 48148 800 48176 2450
rect 48516 800 48544 2450
rect 48976 800 49004 3946
rect 49160 3194 49188 6802
rect 49436 6322 49464 10200
rect 49804 6338 49832 10200
rect 50264 10146 50292 10200
rect 49424 6316 49476 6322
rect 49424 6258 49476 6264
rect 49620 6310 49832 6338
rect 50172 10118 50292 10146
rect 49620 5302 49648 6310
rect 49700 6248 49752 6254
rect 49700 6190 49752 6196
rect 49608 5296 49660 5302
rect 49608 5238 49660 5244
rect 49424 3936 49476 3942
rect 49424 3878 49476 3884
rect 49148 3188 49200 3194
rect 49148 3130 49200 3136
rect 49436 800 49464 3878
rect 49712 2106 49740 6190
rect 50172 5710 50200 10118
rect 50344 7336 50396 7342
rect 50344 7278 50396 7284
rect 50160 5704 50212 5710
rect 50160 5646 50212 5652
rect 49884 2848 49936 2854
rect 49884 2790 49936 2796
rect 49792 2440 49844 2446
rect 49792 2382 49844 2388
rect 49700 2100 49752 2106
rect 49700 2042 49752 2048
rect 49804 800 49832 2382
rect 49896 1426 49924 2790
rect 50252 2372 50304 2378
rect 50252 2314 50304 2320
rect 49884 1420 49936 1426
rect 49884 1362 49936 1368
rect 50264 800 50292 2314
rect 50356 1562 50384 7278
rect 50436 6656 50488 6662
rect 50436 6598 50488 6604
rect 50448 6118 50476 6598
rect 50724 6458 50752 10200
rect 51184 7818 51212 10200
rect 51172 7812 51224 7818
rect 51172 7754 51224 7760
rect 51552 7478 51580 10200
rect 51724 7880 51776 7886
rect 51724 7822 51776 7828
rect 51540 7472 51592 7478
rect 51540 7414 51592 7420
rect 51736 7410 51764 7822
rect 51724 7404 51776 7410
rect 51724 7346 51776 7352
rect 51816 7336 51868 7342
rect 51816 7278 51868 7284
rect 50712 6452 50764 6458
rect 50712 6394 50764 6400
rect 50436 6112 50488 6118
rect 50436 6054 50488 6060
rect 50528 6112 50580 6118
rect 50528 6054 50580 6060
rect 50540 5778 50568 6054
rect 50528 5772 50580 5778
rect 50528 5714 50580 5720
rect 51632 5772 51684 5778
rect 51632 5714 51684 5720
rect 51540 2916 51592 2922
rect 51540 2858 51592 2864
rect 50712 1896 50764 1902
rect 50712 1838 50764 1844
rect 50344 1556 50396 1562
rect 50344 1498 50396 1504
rect 50724 800 50752 1838
rect 51172 1488 51224 1494
rect 51172 1430 51224 1436
rect 51184 800 51212 1430
rect 51552 800 51580 2858
rect 51644 2650 51672 5714
rect 51724 5024 51776 5030
rect 51724 4966 51776 4972
rect 51736 4690 51764 4966
rect 51724 4684 51776 4690
rect 51724 4626 51776 4632
rect 51828 2650 51856 7278
rect 52012 4622 52040 10200
rect 52092 8424 52144 8430
rect 52092 8366 52144 8372
rect 52000 4616 52052 4622
rect 52000 4558 52052 4564
rect 52000 4140 52052 4146
rect 52000 4082 52052 4088
rect 51632 2644 51684 2650
rect 51632 2586 51684 2592
rect 51816 2644 51868 2650
rect 51816 2586 51868 2592
rect 52012 800 52040 4082
rect 52104 3670 52132 8366
rect 52472 6934 52500 10200
rect 52552 7880 52604 7886
rect 52552 7822 52604 7828
rect 52460 6928 52512 6934
rect 52460 6870 52512 6876
rect 52564 6866 52592 7822
rect 52552 6860 52604 6866
rect 52552 6802 52604 6808
rect 52644 6860 52696 6866
rect 52644 6802 52696 6808
rect 52368 4548 52420 4554
rect 52368 4490 52420 4496
rect 52380 3738 52408 4490
rect 52368 3732 52420 3738
rect 52368 3674 52420 3680
rect 52092 3664 52144 3670
rect 52092 3606 52144 3612
rect 52472 2922 52592 2938
rect 52472 2916 52604 2922
rect 52472 2910 52552 2916
rect 52472 800 52500 2910
rect 52552 2858 52604 2864
rect 52552 1556 52604 1562
rect 52656 1544 52684 6802
rect 52932 6390 52960 10200
rect 53104 8900 53156 8906
rect 53104 8842 53156 8848
rect 53012 6792 53064 6798
rect 53012 6734 53064 6740
rect 52920 6384 52972 6390
rect 52920 6326 52972 6332
rect 53024 6322 53052 6734
rect 53012 6316 53064 6322
rect 53012 6258 53064 6264
rect 52920 5704 52972 5710
rect 52920 5646 52972 5652
rect 52932 5234 52960 5646
rect 52920 5228 52972 5234
rect 52920 5170 52972 5176
rect 52736 4752 52788 4758
rect 52736 4694 52788 4700
rect 52748 2650 52776 4694
rect 52828 4072 52880 4078
rect 52828 4014 52880 4020
rect 52840 3194 52868 4014
rect 53116 3738 53144 8842
rect 53300 5234 53328 10200
rect 53760 5914 53788 10200
rect 54116 8356 54168 8362
rect 54116 8298 54168 8304
rect 54128 7410 54156 8298
rect 54116 7404 54168 7410
rect 54116 7346 54168 7352
rect 54116 6248 54168 6254
rect 54116 6190 54168 6196
rect 53748 5908 53800 5914
rect 53748 5850 53800 5856
rect 53840 5704 53892 5710
rect 53840 5646 53892 5652
rect 53288 5228 53340 5234
rect 53288 5170 53340 5176
rect 53564 5160 53616 5166
rect 53564 5102 53616 5108
rect 53104 3732 53156 3738
rect 53104 3674 53156 3680
rect 53288 3596 53340 3602
rect 53288 3538 53340 3544
rect 52828 3188 52880 3194
rect 52828 3130 52880 3136
rect 52736 2644 52788 2650
rect 52736 2586 52788 2592
rect 52604 1516 52684 1544
rect 52552 1498 52604 1504
rect 52920 1420 52972 1426
rect 52920 1362 52972 1368
rect 52932 800 52960 1362
rect 53300 800 53328 3538
rect 53576 3194 53604 5102
rect 53564 3188 53616 3194
rect 53564 3130 53616 3136
rect 53484 3046 53788 3074
rect 53484 2854 53512 3046
rect 53472 2848 53524 2854
rect 53472 2790 53524 2796
rect 53564 2848 53616 2854
rect 53564 2790 53616 2796
rect 53576 1902 53604 2790
rect 53564 1896 53616 1902
rect 53564 1838 53616 1844
rect 53760 800 53788 3046
rect 53852 1562 53880 5646
rect 53932 3392 53984 3398
rect 53932 3334 53984 3340
rect 53944 3058 53972 3334
rect 53932 3052 53984 3058
rect 53932 2994 53984 3000
rect 54024 3052 54076 3058
rect 54024 2994 54076 3000
rect 54036 1902 54064 2994
rect 54024 1896 54076 1902
rect 54024 1838 54076 1844
rect 54128 1562 54156 6190
rect 54220 4622 54248 10200
rect 54680 8514 54708 10200
rect 55048 8786 55076 10200
rect 55048 8758 55168 8786
rect 54680 8486 54800 8514
rect 54668 8424 54720 8430
rect 54668 8366 54720 8372
rect 54680 8090 54708 8366
rect 54668 8084 54720 8090
rect 54668 8026 54720 8032
rect 54576 6112 54628 6118
rect 54576 6054 54628 6060
rect 54588 5778 54616 6054
rect 54576 5772 54628 5778
rect 54576 5714 54628 5720
rect 54772 5710 54800 8486
rect 55140 7936 55168 8758
rect 55140 7908 55260 7936
rect 55232 7478 55260 7908
rect 55220 7472 55272 7478
rect 55220 7414 55272 7420
rect 55508 6100 55536 10200
rect 55864 8968 55916 8974
rect 55864 8910 55916 8916
rect 55876 8090 55904 8910
rect 55864 8084 55916 8090
rect 55864 8026 55916 8032
rect 55680 7472 55732 7478
rect 55680 7414 55732 7420
rect 55588 7336 55640 7342
rect 55588 7278 55640 7284
rect 55140 6072 55536 6100
rect 54760 5704 54812 5710
rect 54760 5646 54812 5652
rect 54852 5160 54904 5166
rect 54852 5102 54904 5108
rect 54864 4826 54892 5102
rect 54852 4820 54904 4826
rect 54852 4762 54904 4768
rect 54760 4684 54812 4690
rect 54760 4626 54812 4632
rect 54208 4616 54260 4622
rect 54208 4558 54260 4564
rect 54208 2984 54260 2990
rect 54208 2926 54260 2932
rect 53840 1556 53892 1562
rect 53840 1498 53892 1504
rect 54116 1556 54168 1562
rect 54116 1498 54168 1504
rect 54220 800 54248 2926
rect 54668 2916 54720 2922
rect 54668 2858 54720 2864
rect 54680 2514 54708 2858
rect 54772 2650 54800 4626
rect 55140 4214 55168 6072
rect 55128 4208 55180 4214
rect 55128 4150 55180 4156
rect 55220 4072 55272 4078
rect 55220 4014 55272 4020
rect 55232 3670 55260 4014
rect 55600 3738 55628 7278
rect 55588 3732 55640 3738
rect 55588 3674 55640 3680
rect 55220 3664 55272 3670
rect 55220 3606 55272 3612
rect 55036 2984 55088 2990
rect 55036 2926 55088 2932
rect 54760 2644 54812 2650
rect 54760 2586 54812 2592
rect 54668 2508 54720 2514
rect 54668 2450 54720 2456
rect 54852 2304 54904 2310
rect 54852 2246 54904 2252
rect 54864 2106 54892 2246
rect 54852 2100 54904 2106
rect 54852 2042 54904 2048
rect 54668 1828 54720 1834
rect 54668 1770 54720 1776
rect 54680 800 54708 1770
rect 55048 800 55076 2926
rect 55692 2650 55720 7414
rect 55968 5302 55996 10200
rect 56336 5778 56364 10200
rect 56600 6860 56652 6866
rect 56600 6802 56652 6808
rect 56324 5772 56376 5778
rect 56324 5714 56376 5720
rect 55956 5296 56008 5302
rect 55956 5238 56008 5244
rect 55956 5160 56008 5166
rect 55956 5102 56008 5108
rect 55968 3194 55996 5102
rect 56232 4684 56284 4690
rect 56232 4626 56284 4632
rect 56244 4282 56272 4626
rect 56232 4276 56284 4282
rect 56232 4218 56284 4224
rect 55956 3188 56008 3194
rect 55956 3130 56008 3136
rect 55220 2644 55272 2650
rect 55220 2586 55272 2592
rect 55680 2644 55732 2650
rect 55680 2586 55732 2592
rect 55128 1896 55180 1902
rect 55232 1850 55260 2586
rect 55496 2508 55548 2514
rect 55496 2450 55548 2456
rect 55180 1844 55260 1850
rect 55128 1838 55260 1844
rect 55140 1822 55260 1838
rect 55508 800 55536 2450
rect 56324 2440 56376 2446
rect 56324 2382 56376 2388
rect 55956 1352 56008 1358
rect 55956 1294 56008 1300
rect 55968 800 55996 1294
rect 56336 800 56364 2382
rect 56612 2310 56640 6802
rect 56796 6118 56824 10200
rect 57256 6390 57284 10200
rect 57716 6798 57744 10200
rect 57336 6792 57388 6798
rect 57336 6734 57388 6740
rect 57704 6792 57756 6798
rect 57704 6734 57756 6740
rect 57244 6384 57296 6390
rect 57244 6326 57296 6332
rect 57348 6322 57376 6734
rect 57336 6316 57388 6322
rect 57336 6258 57388 6264
rect 56784 6112 56836 6118
rect 56784 6054 56836 6060
rect 57704 5704 57756 5710
rect 57704 5646 57756 5652
rect 57716 3738 57744 5646
rect 57980 5296 58032 5302
rect 57980 5238 58032 5244
rect 57704 3732 57756 3738
rect 57704 3674 57756 3680
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 56784 2848 56836 2854
rect 56784 2790 56836 2796
rect 56600 2304 56652 2310
rect 56600 2246 56652 2252
rect 56796 800 56824 2790
rect 57256 800 57284 3334
rect 57992 2514 58020 5238
rect 58084 5166 58112 10200
rect 58544 8378 58572 10200
rect 58544 8350 58664 8378
rect 58532 8288 58584 8294
rect 58532 8230 58584 8236
rect 58544 7954 58572 8230
rect 58532 7948 58584 7954
rect 58532 7890 58584 7896
rect 58256 7744 58308 7750
rect 58256 7686 58308 7692
rect 58072 5160 58124 5166
rect 58072 5102 58124 5108
rect 58072 4616 58124 4622
rect 58072 4558 58124 4564
rect 58084 4146 58112 4558
rect 58072 4140 58124 4146
rect 58072 4082 58124 4088
rect 58268 4078 58296 7686
rect 58440 7336 58492 7342
rect 58440 7278 58492 7284
rect 58256 4072 58308 4078
rect 58256 4014 58308 4020
rect 58072 3052 58124 3058
rect 58072 2994 58124 3000
rect 57980 2508 58032 2514
rect 57980 2450 58032 2456
rect 57336 2440 57388 2446
rect 57336 2382 57388 2388
rect 57348 2106 57376 2382
rect 57336 2100 57388 2106
rect 57336 2042 57388 2048
rect 57704 1964 57756 1970
rect 57704 1906 57756 1912
rect 57716 800 57744 1906
rect 58084 800 58112 2994
rect 58452 2990 58480 7278
rect 58636 6866 58664 8350
rect 58624 6860 58676 6866
rect 58624 6802 58676 6808
rect 58808 6860 58860 6866
rect 58808 6802 58860 6808
rect 58624 6656 58676 6662
rect 58624 6598 58676 6604
rect 58440 2984 58492 2990
rect 58440 2926 58492 2932
rect 58532 2916 58584 2922
rect 58532 2858 58584 2864
rect 58544 800 58572 2858
rect 58636 1426 58664 6598
rect 58820 3738 58848 6802
rect 58900 6656 58952 6662
rect 58900 6598 58952 6604
rect 58808 3732 58860 3738
rect 58808 3674 58860 3680
rect 58912 2038 58940 6598
rect 59004 5846 59032 10200
rect 59360 9376 59412 9382
rect 59360 9318 59412 9324
rect 59372 7410 59400 9318
rect 59464 7410 59492 10200
rect 59544 8968 59596 8974
rect 59544 8910 59596 8916
rect 59556 8498 59584 8910
rect 59544 8492 59596 8498
rect 59544 8434 59596 8440
rect 59636 8424 59688 8430
rect 59636 8366 59688 8372
rect 59360 7404 59412 7410
rect 59360 7346 59412 7352
rect 59452 7404 59504 7410
rect 59452 7346 59504 7352
rect 59452 6248 59504 6254
rect 59452 6190 59504 6196
rect 59176 6112 59228 6118
rect 59176 6054 59228 6060
rect 58992 5840 59044 5846
rect 58992 5782 59044 5788
rect 59188 5302 59216 6054
rect 59268 5772 59320 5778
rect 59268 5714 59320 5720
rect 59176 5296 59228 5302
rect 59176 5238 59228 5244
rect 59084 5228 59136 5234
rect 59084 5170 59136 5176
rect 58992 4004 59044 4010
rect 58992 3946 59044 3952
rect 58900 2032 58952 2038
rect 58900 1974 58952 1980
rect 58624 1420 58676 1426
rect 58624 1362 58676 1368
rect 59004 800 59032 3946
rect 59096 3194 59124 5170
rect 59280 3466 59308 5714
rect 59360 5092 59412 5098
rect 59360 5034 59412 5040
rect 59372 4010 59400 5034
rect 59360 4004 59412 4010
rect 59360 3946 59412 3952
rect 59268 3460 59320 3466
rect 59268 3402 59320 3408
rect 59084 3188 59136 3194
rect 59084 3130 59136 3136
rect 59464 2650 59492 6190
rect 59544 4684 59596 4690
rect 59544 4626 59596 4632
rect 59452 2644 59504 2650
rect 59452 2586 59504 2592
rect 59452 2304 59504 2310
rect 59452 2246 59504 2252
rect 59464 800 59492 2246
rect 59556 2106 59584 4626
rect 59648 3942 59676 8366
rect 59832 6118 59860 10200
rect 60292 7206 60320 10200
rect 60464 9036 60516 9042
rect 60464 8978 60516 8984
rect 60476 8566 60504 8978
rect 60556 8968 60608 8974
rect 60556 8910 60608 8916
rect 60464 8560 60516 8566
rect 60464 8502 60516 8508
rect 60280 7200 60332 7206
rect 60280 7142 60332 7148
rect 59820 6112 59872 6118
rect 59820 6054 59872 6060
rect 60372 5704 60424 5710
rect 60372 5646 60424 5652
rect 59636 3936 59688 3942
rect 59636 3878 59688 3884
rect 60384 3738 60412 5646
rect 60464 4072 60516 4078
rect 60464 4014 60516 4020
rect 60372 3732 60424 3738
rect 60372 3674 60424 3680
rect 60280 3052 60332 3058
rect 60280 2994 60332 3000
rect 59544 2100 59596 2106
rect 59544 2042 59596 2048
rect 59820 1420 59872 1426
rect 59820 1362 59872 1368
rect 59832 800 59860 1362
rect 60292 800 60320 2994
rect 60476 2378 60504 4014
rect 60568 2514 60596 8910
rect 60752 8022 60780 10200
rect 61212 9042 61240 10200
rect 61580 9518 61608 10200
rect 61292 9512 61344 9518
rect 61292 9454 61344 9460
rect 61476 9512 61528 9518
rect 61476 9454 61528 9460
rect 61568 9512 61620 9518
rect 61568 9454 61620 9460
rect 61304 9178 61332 9454
rect 61292 9172 61344 9178
rect 61292 9114 61344 9120
rect 61200 9036 61252 9042
rect 61200 8978 61252 8984
rect 61108 8968 61160 8974
rect 61108 8910 61160 8916
rect 60832 8492 60884 8498
rect 60832 8434 60884 8440
rect 60740 8016 60792 8022
rect 60740 7958 60792 7964
rect 60844 6458 60872 8434
rect 61120 7954 61148 8910
rect 61108 7948 61160 7954
rect 61108 7890 61160 7896
rect 61292 7948 61344 7954
rect 61292 7890 61344 7896
rect 60832 6452 60884 6458
rect 60832 6394 60884 6400
rect 61200 5636 61252 5642
rect 61200 5578 61252 5584
rect 61212 4622 61240 5578
rect 61200 4616 61252 4622
rect 61200 4558 61252 4564
rect 60648 4140 60700 4146
rect 60648 4082 60700 4088
rect 60660 4049 60688 4082
rect 60646 4040 60702 4049
rect 60646 3975 60702 3984
rect 61200 3936 61252 3942
rect 61200 3878 61252 3884
rect 60740 3528 60792 3534
rect 60740 3470 60792 3476
rect 60556 2508 60608 2514
rect 60556 2450 60608 2456
rect 60464 2372 60516 2378
rect 60464 2314 60516 2320
rect 60752 800 60780 3470
rect 61212 800 61240 3878
rect 61304 3670 61332 7890
rect 61292 3664 61344 3670
rect 61292 3606 61344 3612
rect 61488 1426 61516 9454
rect 62040 7834 62068 10200
rect 62040 7818 62160 7834
rect 62040 7812 62172 7818
rect 62040 7806 62120 7812
rect 62120 7754 62172 7760
rect 62500 7342 62528 10200
rect 62672 9376 62724 9382
rect 62672 9318 62724 9324
rect 62580 8968 62632 8974
rect 62580 8910 62632 8916
rect 61568 7336 61620 7342
rect 61568 7278 61620 7284
rect 62488 7336 62540 7342
rect 62488 7278 62540 7284
rect 61580 3602 61608 7278
rect 62592 6866 62620 8910
rect 62684 7410 62712 9318
rect 62960 7410 62988 10200
rect 63328 7970 63356 10200
rect 63684 8424 63736 8430
rect 63684 8366 63736 8372
rect 63328 7942 63540 7970
rect 63040 7880 63092 7886
rect 63040 7822 63092 7828
rect 62672 7404 62724 7410
rect 62672 7346 62724 7352
rect 62948 7404 63000 7410
rect 62948 7346 63000 7352
rect 62580 6860 62632 6866
rect 62580 6802 62632 6808
rect 61660 6792 61712 6798
rect 61660 6734 61712 6740
rect 61672 4826 61700 6734
rect 62304 6656 62356 6662
rect 62304 6598 62356 6604
rect 62120 6384 62172 6390
rect 62120 6326 62172 6332
rect 61844 6180 61896 6186
rect 61844 6122 61896 6128
rect 61856 5710 61884 6122
rect 61936 6112 61988 6118
rect 61936 6054 61988 6060
rect 61844 5704 61896 5710
rect 61844 5646 61896 5652
rect 61948 5234 61976 6054
rect 62028 5772 62080 5778
rect 62028 5714 62080 5720
rect 61936 5228 61988 5234
rect 61936 5170 61988 5176
rect 61660 4820 61712 4826
rect 61660 4762 61712 4768
rect 61568 3596 61620 3602
rect 61568 3538 61620 3544
rect 61568 2916 61620 2922
rect 61568 2858 61620 2864
rect 61476 1420 61528 1426
rect 61476 1362 61528 1368
rect 61580 800 61608 2858
rect 62040 2582 62068 5714
rect 62028 2576 62080 2582
rect 62028 2518 62080 2524
rect 62028 1964 62080 1970
rect 62028 1906 62080 1912
rect 62040 800 62068 1906
rect 62132 1902 62160 6326
rect 62212 5296 62264 5302
rect 62212 5238 62264 5244
rect 62224 2446 62252 5238
rect 62212 2440 62264 2446
rect 62212 2382 62264 2388
rect 62316 2038 62344 6598
rect 62856 5568 62908 5574
rect 62856 5510 62908 5516
rect 62868 3126 62896 5510
rect 62856 3120 62908 3126
rect 62856 3062 62908 3068
rect 63052 2990 63080 7822
rect 63512 7818 63540 7942
rect 63500 7812 63552 7818
rect 63500 7754 63552 7760
rect 63408 7472 63460 7478
rect 63408 7414 63460 7420
rect 63316 7336 63368 7342
rect 63316 7278 63368 7284
rect 63224 5160 63276 5166
rect 63224 5102 63276 5108
rect 63236 4826 63264 5102
rect 63224 4820 63276 4826
rect 63224 4762 63276 4768
rect 63328 4078 63356 7278
rect 63316 4072 63368 4078
rect 63316 4014 63368 4020
rect 63040 2984 63092 2990
rect 63040 2926 63092 2932
rect 63420 2514 63448 7414
rect 63500 6656 63552 6662
rect 63500 6598 63552 6604
rect 63408 2508 63460 2514
rect 63408 2450 63460 2456
rect 63316 2304 63368 2310
rect 63316 2246 63368 2252
rect 62304 2032 62356 2038
rect 62304 1974 62356 1980
rect 62120 1896 62172 1902
rect 62120 1838 62172 1844
rect 62948 1828 63000 1834
rect 62948 1770 63000 1776
rect 62488 1556 62540 1562
rect 62488 1498 62540 1504
rect 62500 800 62528 1498
rect 62960 800 62988 1770
rect 63328 800 63356 2246
rect 63512 1494 63540 6598
rect 63696 4146 63724 8366
rect 63788 6866 63816 10200
rect 64076 9276 64132 9296
rect 64076 9200 64132 9220
rect 63960 8288 64012 8294
rect 63960 8230 64012 8236
rect 63972 8022 64000 8230
rect 64076 8188 64132 8208
rect 64076 8112 64132 8132
rect 63960 8016 64012 8022
rect 63960 7958 64012 7964
rect 64076 7100 64132 7120
rect 64076 7024 64132 7044
rect 64248 6866 64276 10200
rect 64512 7880 64564 7886
rect 64512 7822 64564 7828
rect 63776 6860 63828 6866
rect 63776 6802 63828 6808
rect 64052 6860 64104 6866
rect 64052 6802 64104 6808
rect 64236 6860 64288 6866
rect 64236 6802 64288 6808
rect 64064 6322 64092 6802
rect 64052 6316 64104 6322
rect 64052 6258 64104 6264
rect 63868 6248 63920 6254
rect 63868 6190 63920 6196
rect 63880 5234 63908 6190
rect 64076 6012 64132 6032
rect 64076 5936 64132 5956
rect 63868 5228 63920 5234
rect 63868 5170 63920 5176
rect 64076 4924 64132 4944
rect 64076 4848 64132 4868
rect 63684 4140 63736 4146
rect 63684 4082 63736 4088
rect 64076 3836 64132 3856
rect 64076 3760 64132 3780
rect 64524 2990 64552 7822
rect 64616 6254 64644 10200
rect 64696 9376 64748 9382
rect 64696 9318 64748 9324
rect 64708 9178 64736 9318
rect 64696 9172 64748 9178
rect 64696 9114 64748 9120
rect 64972 8288 65024 8294
rect 64972 8230 65024 8236
rect 64984 8022 65012 8230
rect 64972 8016 65024 8022
rect 64972 7958 65024 7964
rect 64788 7880 64840 7886
rect 64788 7822 64840 7828
rect 64800 7342 64828 7822
rect 65076 7342 65104 10200
rect 64788 7336 64840 7342
rect 64788 7278 64840 7284
rect 65064 7336 65116 7342
rect 65064 7278 65116 7284
rect 64696 7200 64748 7206
rect 64696 7142 64748 7148
rect 64708 6254 64736 7142
rect 65536 6798 65564 10200
rect 65708 9376 65760 9382
rect 65708 9318 65760 9324
rect 65720 9042 65748 9318
rect 65708 9036 65760 9042
rect 65708 8978 65760 8984
rect 65996 7290 66024 10200
rect 66076 8968 66128 8974
rect 66076 8910 66128 8916
rect 66088 8498 66116 8910
rect 66076 8492 66128 8498
rect 66076 8434 66128 8440
rect 66364 7290 66392 10200
rect 65996 7274 66300 7290
rect 65996 7268 66312 7274
rect 65996 7262 66260 7268
rect 66364 7262 66484 7290
rect 66260 7210 66312 7216
rect 66352 7200 66404 7206
rect 66352 7142 66404 7148
rect 66364 6866 66392 7142
rect 66352 6860 66404 6866
rect 66352 6802 66404 6808
rect 65524 6792 65576 6798
rect 65524 6734 65576 6740
rect 66456 6730 66484 7262
rect 66824 6798 66852 10200
rect 67088 8492 67140 8498
rect 67088 8434 67140 8440
rect 66812 6792 66864 6798
rect 66812 6734 66864 6740
rect 66444 6724 66496 6730
rect 66444 6666 66496 6672
rect 66260 6656 66312 6662
rect 66260 6598 66312 6604
rect 64604 6248 64656 6254
rect 64604 6190 64656 6196
rect 64696 6248 64748 6254
rect 64696 6190 64748 6196
rect 65524 4004 65576 4010
rect 65524 3946 65576 3952
rect 64512 2984 64564 2990
rect 64512 2926 64564 2932
rect 64076 2748 64132 2768
rect 64076 2672 64132 2692
rect 64604 2440 64656 2446
rect 64604 2382 64656 2388
rect 63776 1828 63828 1834
rect 63776 1770 63828 1776
rect 63500 1488 63552 1494
rect 63500 1430 63552 1436
rect 63788 800 63816 1770
rect 64076 1660 64132 1680
rect 64076 1584 64132 1604
rect 64236 1420 64288 1426
rect 64236 1362 64288 1368
rect 64248 800 64276 1362
rect 64616 800 64644 2382
rect 65064 1488 65116 1494
rect 65064 1430 65116 1436
rect 65076 800 65104 1430
rect 65536 800 65564 3946
rect 65984 2032 66036 2038
rect 65984 1974 66036 1980
rect 65996 800 66024 1974
rect 66272 1902 66300 6598
rect 66996 6384 67048 6390
rect 66996 6326 67048 6332
rect 66904 6248 66956 6254
rect 66904 6190 66956 6196
rect 66444 5704 66496 5710
rect 66444 5646 66496 5652
rect 66456 5166 66484 5646
rect 66536 5296 66588 5302
rect 66536 5238 66588 5244
rect 66444 5160 66496 5166
rect 66444 5102 66496 5108
rect 66548 3602 66576 5238
rect 66536 3596 66588 3602
rect 66536 3538 66588 3544
rect 66352 2916 66404 2922
rect 66352 2858 66404 2864
rect 66260 1896 66312 1902
rect 66260 1838 66312 1844
rect 66168 1828 66220 1834
rect 66168 1770 66220 1776
rect 66180 1426 66208 1770
rect 66168 1420 66220 1426
rect 66168 1362 66220 1368
rect 66364 800 66392 2858
rect 66812 2440 66864 2446
rect 66812 2382 66864 2388
rect 66824 800 66852 2382
rect 66916 1766 66944 6190
rect 67008 2990 67036 6326
rect 67100 5914 67128 8434
rect 67284 8022 67312 10200
rect 67272 8016 67324 8022
rect 67272 7958 67324 7964
rect 67180 6860 67232 6866
rect 67180 6802 67232 6808
rect 67192 6322 67220 6802
rect 67744 6662 67772 10200
rect 67824 8968 67876 8974
rect 67824 8910 67876 8916
rect 67836 7954 67864 8910
rect 67824 7948 67876 7954
rect 67824 7890 67876 7896
rect 67916 7880 67968 7886
rect 67916 7822 67968 7828
rect 67640 6656 67692 6662
rect 67640 6598 67692 6604
rect 67732 6656 67784 6662
rect 67732 6598 67784 6604
rect 67180 6316 67232 6322
rect 67180 6258 67232 6264
rect 67088 5908 67140 5914
rect 67088 5850 67140 5856
rect 67456 5704 67508 5710
rect 67456 5646 67508 5652
rect 67468 4826 67496 5646
rect 67548 5024 67600 5030
rect 67548 4966 67600 4972
rect 67456 4820 67508 4826
rect 67456 4762 67508 4768
rect 67560 4146 67588 4966
rect 67548 4140 67600 4146
rect 67548 4082 67600 4088
rect 67272 3528 67324 3534
rect 67272 3470 67324 3476
rect 66996 2984 67048 2990
rect 66996 2926 67048 2932
rect 66904 1760 66956 1766
rect 66904 1702 66956 1708
rect 67284 800 67312 3470
rect 67652 2514 67680 6598
rect 67732 6112 67784 6118
rect 67732 6054 67784 6060
rect 67744 5166 67772 6054
rect 67732 5160 67784 5166
rect 67732 5102 67784 5108
rect 67732 5024 67784 5030
rect 67732 4966 67784 4972
rect 67744 4078 67772 4966
rect 67928 4078 67956 7822
rect 68112 5914 68140 10200
rect 68468 7472 68520 7478
rect 68468 7414 68520 7420
rect 68100 5908 68152 5914
rect 68100 5850 68152 5856
rect 68480 5114 68508 7414
rect 68572 7410 68600 10200
rect 69032 8514 69060 10200
rect 69032 8486 69152 8514
rect 69020 8356 69072 8362
rect 69020 8298 69072 8304
rect 68836 7880 68888 7886
rect 68836 7822 68888 7828
rect 68560 7404 68612 7410
rect 68560 7346 68612 7352
rect 68848 7342 68876 7822
rect 68836 7336 68888 7342
rect 68742 7304 68798 7313
rect 68836 7278 68888 7284
rect 68928 7336 68980 7342
rect 68928 7278 68980 7284
rect 68742 7239 68798 7248
rect 68756 5710 68784 7239
rect 68836 6656 68888 6662
rect 68836 6598 68888 6604
rect 68848 6390 68876 6598
rect 68836 6384 68888 6390
rect 68836 6326 68888 6332
rect 68836 5772 68888 5778
rect 68836 5714 68888 5720
rect 68744 5704 68796 5710
rect 68744 5646 68796 5652
rect 68480 5086 68784 5114
rect 67732 4072 67784 4078
rect 67732 4014 67784 4020
rect 67916 4072 67968 4078
rect 67916 4014 67968 4020
rect 68560 2916 68612 2922
rect 68560 2858 68612 2864
rect 67640 2508 67692 2514
rect 67640 2450 67692 2456
rect 68100 2440 68152 2446
rect 68100 2382 68152 2388
rect 67732 2100 67784 2106
rect 67732 2042 67784 2048
rect 67744 800 67772 2042
rect 68112 800 68140 2382
rect 68572 800 68600 2858
rect 68756 2514 68784 5086
rect 68848 4214 68876 5714
rect 68836 4208 68888 4214
rect 68836 4150 68888 4156
rect 68744 2508 68796 2514
rect 68744 2450 68796 2456
rect 68940 1902 68968 7278
rect 69032 6866 69060 8298
rect 69020 6860 69072 6866
rect 69020 6802 69072 6808
rect 69020 6656 69072 6662
rect 69020 6598 69072 6604
rect 69032 6254 69060 6598
rect 69020 6248 69072 6254
rect 69020 6190 69072 6196
rect 69124 6118 69152 8486
rect 69492 6882 69520 10200
rect 69492 6854 69612 6882
rect 69480 6792 69532 6798
rect 69480 6734 69532 6740
rect 69112 6112 69164 6118
rect 69112 6054 69164 6060
rect 69020 5160 69072 5166
rect 69020 5102 69072 5108
rect 69032 3738 69060 5102
rect 69020 3732 69072 3738
rect 69020 3674 69072 3680
rect 69020 2916 69072 2922
rect 69020 2858 69072 2864
rect 68928 1896 68980 1902
rect 68928 1838 68980 1844
rect 69032 800 69060 2858
rect 69492 1426 69520 6734
rect 69584 6322 69612 6854
rect 69860 6798 69888 10200
rect 70320 9058 70348 10200
rect 70492 9376 70544 9382
rect 70492 9318 70544 9324
rect 70228 9030 70348 9058
rect 69940 8968 69992 8974
rect 69940 8910 69992 8916
rect 69848 6792 69900 6798
rect 69848 6734 69900 6740
rect 69572 6316 69624 6322
rect 69572 6258 69624 6264
rect 69952 5166 69980 8910
rect 70124 7880 70176 7886
rect 70124 7822 70176 7828
rect 70136 6662 70164 7822
rect 70228 6730 70256 9030
rect 70308 8968 70360 8974
rect 70308 8910 70360 8916
rect 70320 6866 70348 8910
rect 70504 7342 70532 9318
rect 70492 7336 70544 7342
rect 70492 7278 70544 7284
rect 70308 6860 70360 6866
rect 70308 6802 70360 6808
rect 70216 6724 70268 6730
rect 70216 6666 70268 6672
rect 70124 6656 70176 6662
rect 70124 6598 70176 6604
rect 70400 6248 70452 6254
rect 70400 6190 70452 6196
rect 70676 6248 70728 6254
rect 70676 6190 70728 6196
rect 69940 5160 69992 5166
rect 69940 5102 69992 5108
rect 70308 4616 70360 4622
rect 70306 4584 70308 4593
rect 70360 4584 70362 4593
rect 70306 4519 70362 4528
rect 70412 4146 70440 6190
rect 70688 5914 70716 6190
rect 70676 5908 70728 5914
rect 70676 5850 70728 5856
rect 70492 5364 70544 5370
rect 70492 5306 70544 5312
rect 70504 4690 70532 5306
rect 70780 5234 70808 10200
rect 70952 8900 71004 8906
rect 70952 8842 71004 8848
rect 70964 8430 70992 8842
rect 70952 8424 71004 8430
rect 70952 8366 71004 8372
rect 70952 6384 71004 6390
rect 70952 6326 71004 6332
rect 70584 5228 70636 5234
rect 70584 5170 70636 5176
rect 70768 5228 70820 5234
rect 70768 5170 70820 5176
rect 70492 4684 70544 4690
rect 70492 4626 70544 4632
rect 70400 4140 70452 4146
rect 70400 4082 70452 4088
rect 69664 2576 69716 2582
rect 69664 2518 69716 2524
rect 69676 2106 69704 2518
rect 69664 2100 69716 2106
rect 69664 2042 69716 2048
rect 69848 1964 69900 1970
rect 69848 1906 69900 1912
rect 69572 1828 69624 1834
rect 69572 1770 69624 1776
rect 69480 1420 69532 1426
rect 69480 1362 69532 1368
rect 69584 898 69612 1770
rect 69492 870 69612 898
rect 69492 800 69520 870
rect 69860 800 69888 1906
rect 70596 1902 70624 5170
rect 70860 5160 70912 5166
rect 70860 5102 70912 5108
rect 70872 2990 70900 5102
rect 70964 4078 70992 6326
rect 71240 5098 71268 10200
rect 71608 9602 71636 10200
rect 71608 9574 71728 9602
rect 71412 9512 71464 9518
rect 71412 9454 71464 9460
rect 71320 8424 71372 8430
rect 71320 8366 71372 8372
rect 71228 5092 71280 5098
rect 71228 5034 71280 5040
rect 71332 4826 71360 8366
rect 71424 7954 71452 9454
rect 71596 9444 71648 9450
rect 71596 9386 71648 9392
rect 71608 8430 71636 9386
rect 71596 8424 71648 8430
rect 71596 8366 71648 8372
rect 71700 8004 71728 9574
rect 71780 8016 71832 8022
rect 71700 7976 71780 8004
rect 71780 7958 71832 7964
rect 71412 7948 71464 7954
rect 71412 7890 71464 7896
rect 71964 7880 72016 7886
rect 71964 7822 72016 7828
rect 71504 6656 71556 6662
rect 71504 6598 71556 6604
rect 71320 4820 71372 4826
rect 71320 4762 71372 4768
rect 71412 4616 71464 4622
rect 71412 4558 71464 4564
rect 70952 4072 71004 4078
rect 70952 4014 71004 4020
rect 71424 3738 71452 4558
rect 71412 3732 71464 3738
rect 71412 3674 71464 3680
rect 70860 2984 70912 2990
rect 70860 2926 70912 2932
rect 71516 2514 71544 6598
rect 71780 6248 71832 6254
rect 71780 6190 71832 6196
rect 71872 6248 71924 6254
rect 71872 6190 71924 6196
rect 71792 4146 71820 6190
rect 71780 4140 71832 4146
rect 71780 4082 71832 4088
rect 71596 2916 71648 2922
rect 71596 2858 71648 2864
rect 71504 2508 71556 2514
rect 71504 2450 71556 2456
rect 71228 2440 71280 2446
rect 71228 2382 71280 2388
rect 70584 1896 70636 1902
rect 70584 1838 70636 1844
rect 70768 1828 70820 1834
rect 70768 1770 70820 1776
rect 70308 1420 70360 1426
rect 70308 1362 70360 1368
rect 70320 800 70348 1362
rect 70780 800 70808 1770
rect 71240 800 71268 2382
rect 71608 800 71636 2858
rect 71884 2038 71912 6190
rect 71976 3942 72004 7822
rect 72068 6390 72096 10200
rect 72240 8968 72292 8974
rect 72240 8910 72292 8916
rect 72056 6384 72108 6390
rect 72056 6326 72108 6332
rect 72252 5302 72280 8910
rect 72240 5296 72292 5302
rect 72240 5238 72292 5244
rect 72528 5166 72556 10200
rect 72792 6656 72844 6662
rect 72792 6598 72844 6604
rect 72700 6384 72752 6390
rect 72700 6326 72752 6332
rect 72608 5772 72660 5778
rect 72608 5714 72660 5720
rect 72424 5160 72476 5166
rect 72424 5102 72476 5108
rect 72516 5160 72568 5166
rect 72516 5102 72568 5108
rect 71964 3936 72016 3942
rect 71964 3878 72016 3884
rect 72148 2440 72200 2446
rect 72148 2382 72200 2388
rect 71872 2032 71924 2038
rect 71872 1974 71924 1980
rect 72160 1170 72188 2382
rect 72436 1902 72464 5102
rect 72620 4706 72648 5714
rect 72528 4678 72648 4706
rect 72528 3534 72556 4678
rect 72608 4004 72660 4010
rect 72608 3946 72660 3952
rect 72516 3528 72568 3534
rect 72516 3470 72568 3476
rect 72516 3392 72568 3398
rect 72516 3334 72568 3340
rect 72424 1896 72476 1902
rect 72424 1838 72476 1844
rect 72068 1142 72188 1170
rect 72068 800 72096 1142
rect 72528 800 72556 3334
rect 72620 1426 72648 3946
rect 72712 2990 72740 6326
rect 72804 3602 72832 6598
rect 72896 5846 72924 10200
rect 73160 9648 73212 9654
rect 73160 9590 73212 9596
rect 73068 8424 73120 8430
rect 73068 8366 73120 8372
rect 72976 7336 73028 7342
rect 72976 7278 73028 7284
rect 72884 5840 72936 5846
rect 72884 5782 72936 5788
rect 72884 5092 72936 5098
rect 72884 5034 72936 5040
rect 72896 4622 72924 5034
rect 72884 4616 72936 4622
rect 72884 4558 72936 4564
rect 72988 4078 73016 7278
rect 73080 4690 73108 8366
rect 73172 5778 73200 9590
rect 73252 6724 73304 6730
rect 73252 6666 73304 6672
rect 73160 5772 73212 5778
rect 73160 5714 73212 5720
rect 73160 5568 73212 5574
rect 73160 5510 73212 5516
rect 73068 4684 73120 4690
rect 73068 4626 73120 4632
rect 72976 4072 73028 4078
rect 72976 4014 73028 4020
rect 72884 4004 72936 4010
rect 72884 3946 72936 3952
rect 72792 3596 72844 3602
rect 72792 3538 72844 3544
rect 72700 2984 72752 2990
rect 72700 2926 72752 2932
rect 72608 1420 72660 1426
rect 72608 1362 72660 1368
rect 72896 800 72924 3946
rect 73172 2514 73200 5510
rect 73264 3058 73292 6666
rect 73356 6322 73384 10200
rect 73436 9444 73488 9450
rect 73436 9386 73488 9392
rect 73448 7954 73476 9386
rect 73712 9376 73764 9382
rect 73712 9318 73764 9324
rect 73724 9042 73752 9318
rect 73712 9036 73764 9042
rect 73712 8978 73764 8984
rect 73436 7948 73488 7954
rect 73436 7890 73488 7896
rect 73528 7880 73580 7886
rect 73528 7822 73580 7828
rect 73344 6316 73396 6322
rect 73344 6258 73396 6264
rect 73344 3664 73396 3670
rect 73344 3606 73396 3612
rect 73252 3052 73304 3058
rect 73252 2994 73304 3000
rect 73160 2508 73212 2514
rect 73160 2450 73212 2456
rect 73356 800 73384 3606
rect 73540 1902 73568 7822
rect 73712 6452 73764 6458
rect 73712 6394 73764 6400
rect 73724 5642 73752 6394
rect 73816 5642 73844 10200
rect 73988 9376 74040 9382
rect 73988 9318 74040 9324
rect 74000 7410 74028 9318
rect 73988 7404 74040 7410
rect 73988 7346 74040 7352
rect 74276 6866 74304 10200
rect 74448 9172 74500 9178
rect 74448 9114 74500 9120
rect 74460 8430 74488 9114
rect 74448 8424 74500 8430
rect 74448 8366 74500 8372
rect 74644 7342 74672 10200
rect 75104 8498 75132 10200
rect 75184 10192 75236 10198
rect 75184 10134 75236 10140
rect 75196 8974 75224 10134
rect 75368 9648 75420 9654
rect 75368 9590 75420 9596
rect 75276 9036 75328 9042
rect 75276 8978 75328 8984
rect 75184 8968 75236 8974
rect 75184 8910 75236 8916
rect 75092 8492 75144 8498
rect 75092 8434 75144 8440
rect 75288 8090 75316 8978
rect 75380 8430 75408 9590
rect 75460 9036 75512 9042
rect 75460 8978 75512 8984
rect 75368 8424 75420 8430
rect 75368 8366 75420 8372
rect 75276 8084 75328 8090
rect 75276 8026 75328 8032
rect 75276 7948 75328 7954
rect 75276 7890 75328 7896
rect 74632 7336 74684 7342
rect 74632 7278 74684 7284
rect 74908 7336 74960 7342
rect 74908 7278 74960 7284
rect 74540 7200 74592 7206
rect 74540 7142 74592 7148
rect 74264 6860 74316 6866
rect 74264 6802 74316 6808
rect 74552 6798 74580 7142
rect 74540 6792 74592 6798
rect 74540 6734 74592 6740
rect 74448 5772 74500 5778
rect 74448 5714 74500 5720
rect 73712 5636 73764 5642
rect 73712 5578 73764 5584
rect 73804 5636 73856 5642
rect 73804 5578 73856 5584
rect 74172 5160 74224 5166
rect 74172 5102 74224 5108
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 73528 1896 73580 1902
rect 73528 1838 73580 1844
rect 73816 800 73844 4082
rect 74184 3738 74212 5102
rect 74172 3732 74224 3738
rect 74172 3674 74224 3680
rect 74264 3596 74316 3602
rect 74264 3538 74316 3544
rect 74276 800 74304 3538
rect 74460 3058 74488 5714
rect 74724 5636 74776 5642
rect 74724 5578 74776 5584
rect 74736 5166 74764 5578
rect 74540 5160 74592 5166
rect 74540 5102 74592 5108
rect 74724 5160 74776 5166
rect 74724 5102 74776 5108
rect 74448 3052 74500 3058
rect 74448 2994 74500 3000
rect 74552 2514 74580 5102
rect 74632 4616 74684 4622
rect 74632 4558 74684 4564
rect 74644 3602 74672 4558
rect 74724 4480 74776 4486
rect 74724 4422 74776 4428
rect 74736 3670 74764 4422
rect 74724 3664 74776 3670
rect 74724 3606 74776 3612
rect 74920 3602 74948 7278
rect 74632 3596 74684 3602
rect 74632 3538 74684 3544
rect 74908 3596 74960 3602
rect 74908 3538 74960 3544
rect 75092 3528 75144 3534
rect 75092 3470 75144 3476
rect 74632 2916 74684 2922
rect 74632 2858 74684 2864
rect 74540 2508 74592 2514
rect 74540 2450 74592 2456
rect 74644 800 74672 2858
rect 75104 800 75132 3470
rect 75288 2650 75316 7890
rect 75472 5930 75500 8978
rect 75564 7818 75592 10200
rect 75828 8560 75880 8566
rect 76024 8548 76052 10200
rect 76392 9466 76420 10200
rect 76392 9438 76512 9466
rect 76380 9376 76432 9382
rect 76380 9318 76432 9324
rect 75880 8520 76052 8548
rect 75828 8502 75880 8508
rect 75828 7880 75880 7886
rect 75828 7822 75880 7828
rect 75552 7812 75604 7818
rect 75552 7754 75604 7760
rect 75380 5902 75500 5930
rect 75276 2644 75328 2650
rect 75276 2586 75328 2592
rect 75380 1562 75408 5902
rect 75460 5568 75512 5574
rect 75460 5510 75512 5516
rect 75368 1556 75420 1562
rect 75368 1498 75420 1504
rect 75472 1426 75500 5510
rect 75552 3596 75604 3602
rect 75552 3538 75604 3544
rect 75460 1420 75512 1426
rect 75460 1362 75512 1368
rect 75564 800 75592 3538
rect 75840 3534 75868 7822
rect 76392 7410 76420 9318
rect 76380 7404 76432 7410
rect 76380 7346 76432 7352
rect 76484 6866 76512 9438
rect 76852 9058 76880 10200
rect 77312 9602 77340 10200
rect 77220 9574 77340 9602
rect 77220 9110 77248 9574
rect 76760 9030 76880 9058
rect 77208 9104 77260 9110
rect 77208 9046 77260 9052
rect 76760 7342 76788 9030
rect 77392 8968 77444 8974
rect 77392 8910 77444 8916
rect 76840 8900 76892 8906
rect 76840 8842 76892 8848
rect 76852 8430 76880 8842
rect 77404 8634 77432 8910
rect 77392 8628 77444 8634
rect 77392 8570 77444 8576
rect 76840 8424 76892 8430
rect 76840 8366 76892 8372
rect 77024 7880 77076 7886
rect 77024 7822 77076 7828
rect 76748 7336 76800 7342
rect 76748 7278 76800 7284
rect 76472 6860 76524 6866
rect 76472 6802 76524 6808
rect 76196 6656 76248 6662
rect 76196 6598 76248 6604
rect 75920 4276 75972 4282
rect 75920 4218 75972 4224
rect 75932 4010 75960 4218
rect 75920 4004 75972 4010
rect 75920 3946 75972 3952
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76208 2990 76236 6598
rect 76656 6248 76708 6254
rect 76656 6190 76708 6196
rect 76668 3738 76696 6190
rect 77036 6118 77064 7822
rect 77300 6316 77352 6322
rect 77300 6258 77352 6264
rect 77024 6112 77076 6118
rect 77024 6054 77076 6060
rect 77024 5024 77076 5030
rect 77024 4966 77076 4972
rect 76656 3732 76708 3738
rect 76656 3674 76708 3680
rect 77036 3602 77064 4966
rect 77024 3596 77076 3602
rect 77024 3538 77076 3544
rect 76196 2984 76248 2990
rect 76196 2926 76248 2932
rect 76840 2916 76892 2922
rect 76840 2858 76892 2864
rect 76012 2440 76064 2446
rect 76012 2382 76064 2388
rect 76024 800 76052 2382
rect 76380 1420 76432 1426
rect 76380 1362 76432 1368
rect 76392 800 76420 1362
rect 76852 800 76880 2858
rect 77312 2514 77340 6258
rect 77772 6254 77800 10200
rect 77852 9920 77904 9926
rect 77852 9862 77904 9868
rect 77864 9042 77892 9862
rect 77852 9036 77904 9042
rect 77852 8978 77904 8984
rect 77944 7336 77996 7342
rect 77944 7278 77996 7284
rect 77760 6248 77812 6254
rect 77760 6190 77812 6196
rect 77576 5704 77628 5710
rect 77576 5646 77628 5652
rect 77668 5704 77720 5710
rect 77668 5646 77720 5652
rect 77588 5234 77616 5646
rect 77576 5228 77628 5234
rect 77576 5170 77628 5176
rect 77680 5166 77708 5646
rect 77668 5160 77720 5166
rect 77668 5102 77720 5108
rect 77392 4752 77444 4758
rect 77392 4694 77444 4700
rect 77404 3942 77432 4694
rect 77392 3936 77444 3942
rect 77392 3878 77444 3884
rect 77392 3528 77444 3534
rect 77392 3470 77444 3476
rect 77300 2508 77352 2514
rect 77300 2450 77352 2456
rect 77404 1034 77432 3470
rect 77956 2990 77984 7278
rect 78140 5778 78168 10200
rect 78220 9376 78272 9382
rect 78220 9318 78272 9324
rect 78232 7954 78260 9318
rect 78404 8356 78456 8362
rect 78404 8298 78456 8304
rect 78220 7948 78272 7954
rect 78220 7890 78272 7896
rect 78220 6384 78272 6390
rect 78220 6326 78272 6332
rect 78128 5772 78180 5778
rect 78128 5714 78180 5720
rect 77944 2984 77996 2990
rect 77944 2926 77996 2932
rect 78232 1902 78260 6326
rect 78416 6254 78444 8298
rect 78496 7880 78548 7886
rect 78496 7822 78548 7828
rect 78404 6248 78456 6254
rect 78404 6190 78456 6196
rect 78508 2514 78536 7822
rect 78600 7342 78628 10200
rect 78588 7336 78640 7342
rect 78588 7278 78640 7284
rect 79060 6322 79088 10200
rect 79520 7818 79548 10200
rect 79508 7812 79560 7818
rect 79508 7754 79560 7760
rect 79324 6384 79376 6390
rect 79324 6326 79376 6332
rect 79048 6316 79100 6322
rect 79048 6258 79100 6264
rect 79140 5772 79192 5778
rect 79140 5714 79192 5720
rect 79048 5636 79100 5642
rect 79048 5578 79100 5584
rect 78772 5296 78824 5302
rect 78772 5238 78824 5244
rect 78784 4078 78812 5238
rect 78772 4072 78824 4078
rect 78772 4014 78824 4020
rect 79060 3641 79088 5578
rect 79046 3632 79102 3641
rect 79046 3567 79102 3576
rect 78496 2508 78548 2514
rect 78496 2450 78548 2456
rect 78588 2440 78640 2446
rect 79152 2417 79180 5714
rect 79336 3602 79364 6326
rect 79888 6254 79916 10200
rect 80244 8560 80296 8566
rect 80244 8502 80296 8508
rect 79876 6248 79928 6254
rect 79876 6190 79928 6196
rect 80060 6248 80112 6254
rect 80060 6190 80112 6196
rect 79784 5160 79836 5166
rect 79784 5102 79836 5108
rect 79508 4616 79560 4622
rect 79508 4558 79560 4564
rect 79520 4146 79548 4558
rect 79508 4140 79560 4146
rect 79508 4082 79560 4088
rect 79324 3596 79376 3602
rect 79324 3538 79376 3544
rect 79796 3058 79824 5102
rect 79968 4752 80020 4758
rect 79968 4694 80020 4700
rect 79784 3052 79836 3058
rect 79784 2994 79836 3000
rect 79508 2440 79560 2446
rect 78588 2382 78640 2388
rect 79138 2408 79194 2417
rect 78220 1896 78272 1902
rect 78220 1838 78272 1844
rect 77760 1828 77812 1834
rect 77760 1770 77812 1776
rect 77312 1006 77432 1034
rect 77312 800 77340 1006
rect 77772 800 77800 1770
rect 78128 1760 78180 1766
rect 78128 1702 78180 1708
rect 78140 800 78168 1702
rect 78600 800 78628 2382
rect 79508 2382 79560 2388
rect 79138 2343 79194 2352
rect 79048 1488 79100 1494
rect 79048 1430 79100 1436
rect 79060 800 79088 1430
rect 79520 800 79548 2382
rect 79876 1760 79928 1766
rect 79876 1702 79928 1708
rect 79888 800 79916 1702
rect 79980 1562 80008 4694
rect 80072 4146 80100 6190
rect 80152 5160 80204 5166
rect 80152 5102 80204 5108
rect 80060 4140 80112 4146
rect 80060 4082 80112 4088
rect 80164 1902 80192 5102
rect 80256 3602 80284 8502
rect 80348 8022 80376 10200
rect 80704 9376 80756 9382
rect 80704 9318 80756 9324
rect 80716 8498 80744 9318
rect 80704 8492 80756 8498
rect 80704 8434 80756 8440
rect 80336 8016 80388 8022
rect 80336 7958 80388 7964
rect 80612 7880 80664 7886
rect 80612 7822 80664 7828
rect 80428 5636 80480 5642
rect 80428 5578 80480 5584
rect 80336 4072 80388 4078
rect 80336 4014 80388 4020
rect 80244 3596 80296 3602
rect 80244 3538 80296 3544
rect 80152 1896 80204 1902
rect 80152 1838 80204 1844
rect 79968 1556 80020 1562
rect 79968 1498 80020 1504
rect 80348 800 80376 4014
rect 80440 2990 80468 5578
rect 80624 2990 80652 7822
rect 80704 7472 80756 7478
rect 80704 7414 80756 7420
rect 80428 2984 80480 2990
rect 80428 2926 80480 2932
rect 80612 2984 80664 2990
rect 80612 2926 80664 2932
rect 80716 2514 80744 7414
rect 80808 6662 80836 10200
rect 80980 8288 81032 8294
rect 80980 8230 81032 8236
rect 80992 7954 81020 8230
rect 80980 7948 81032 7954
rect 80980 7890 81032 7896
rect 81176 7410 81204 10200
rect 81532 8968 81584 8974
rect 81532 8910 81584 8916
rect 81256 8084 81308 8090
rect 81256 8026 81308 8032
rect 81164 7404 81216 7410
rect 81164 7346 81216 7352
rect 80796 6656 80848 6662
rect 80796 6598 80848 6604
rect 80980 5772 81032 5778
rect 80980 5714 81032 5720
rect 80888 4072 80940 4078
rect 80888 4014 80940 4020
rect 80900 3534 80928 4014
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 80796 2916 80848 2922
rect 80796 2858 80848 2864
rect 80704 2508 80756 2514
rect 80704 2450 80756 2456
rect 80808 800 80836 2858
rect 80992 1465 81020 5714
rect 81072 4684 81124 4690
rect 81072 4626 81124 4632
rect 81084 2310 81112 4626
rect 81164 3528 81216 3534
rect 81164 3470 81216 3476
rect 81072 2304 81124 2310
rect 81072 2246 81124 2252
rect 80978 1456 81034 1465
rect 80978 1391 81034 1400
rect 81176 800 81204 3470
rect 81268 2961 81296 8026
rect 81544 7342 81572 8910
rect 81532 7336 81584 7342
rect 81532 7278 81584 7284
rect 81348 7268 81400 7274
rect 81348 7210 81400 7216
rect 81360 3058 81388 7210
rect 81532 6792 81584 6798
rect 81532 6734 81584 6740
rect 81440 6248 81492 6254
rect 81440 6190 81492 6196
rect 81452 5030 81480 6190
rect 81440 5024 81492 5030
rect 81440 4966 81492 4972
rect 81348 3052 81400 3058
rect 81348 2994 81400 3000
rect 81254 2952 81310 2961
rect 81254 2887 81310 2896
rect 81544 2514 81572 6734
rect 81636 5302 81664 10200
rect 81900 7812 81952 7818
rect 81900 7754 81952 7760
rect 81912 6254 81940 7754
rect 81992 6384 82044 6390
rect 81992 6326 82044 6332
rect 81716 6248 81768 6254
rect 81900 6248 81952 6254
rect 81716 6190 81768 6196
rect 81806 6216 81862 6225
rect 81624 5296 81676 5302
rect 81624 5238 81676 5244
rect 81624 5160 81676 5166
rect 81624 5102 81676 5108
rect 81636 4146 81664 5102
rect 81624 4140 81676 4146
rect 81624 4082 81676 4088
rect 81532 2508 81584 2514
rect 81532 2450 81584 2456
rect 81440 2032 81492 2038
rect 81440 1974 81492 1980
rect 81452 1562 81480 1974
rect 81728 1970 81756 6190
rect 81900 6190 81952 6196
rect 81806 6151 81808 6160
rect 81860 6151 81862 6160
rect 81808 6122 81860 6128
rect 82004 2038 82032 6326
rect 82096 5166 82124 10200
rect 82188 8566 82216 10406
rect 82542 10200 82598 11400
rect 82910 10200 82966 11400
rect 83370 10200 83426 11400
rect 83830 10200 83886 11400
rect 84290 10200 84346 11400
rect 84658 10200 84714 11400
rect 85118 10200 85174 11400
rect 85578 10200 85634 11400
rect 86038 10200 86094 11400
rect 86406 10200 86462 11400
rect 86866 10200 86922 11400
rect 87326 10200 87382 11400
rect 87786 10200 87842 11400
rect 88154 10200 88210 11400
rect 88614 10200 88670 11400
rect 89074 10200 89130 11400
rect 89442 10200 89498 11400
rect 89902 10200 89958 11400
rect 90362 10200 90418 11400
rect 90822 10200 90878 11400
rect 91190 10200 91246 11400
rect 91650 10200 91706 11400
rect 92110 10200 92166 11400
rect 92570 10200 92626 11400
rect 92938 10200 92994 11400
rect 93398 10200 93454 11400
rect 93858 10200 93914 11400
rect 94318 10200 94374 11400
rect 94686 10200 94742 11400
rect 95146 10200 95202 11400
rect 95606 10200 95662 11400
rect 96066 10200 96122 11400
rect 96434 10200 96490 11400
rect 96894 10200 96950 11400
rect 97354 10200 97410 11400
rect 97722 10200 97778 11400
rect 97816 10328 97868 10334
rect 97816 10270 97868 10276
rect 82268 8628 82320 8634
rect 82268 8570 82320 8576
rect 82176 8560 82228 8566
rect 82176 8502 82228 8508
rect 82174 6216 82230 6225
rect 82174 6151 82176 6160
rect 82228 6151 82230 6160
rect 82176 6122 82228 6128
rect 82084 5160 82136 5166
rect 82084 5102 82136 5108
rect 82280 4146 82308 8570
rect 82556 5914 82584 10200
rect 82636 9376 82688 9382
rect 82636 9318 82688 9324
rect 82728 9376 82780 9382
rect 82728 9318 82780 9324
rect 82648 6866 82676 9318
rect 82740 8022 82768 9318
rect 82820 8832 82872 8838
rect 82820 8774 82872 8780
rect 82832 8634 82860 8774
rect 82820 8628 82872 8634
rect 82820 8570 82872 8576
rect 82924 8498 82952 10200
rect 82912 8492 82964 8498
rect 82912 8434 82964 8440
rect 83096 8084 83148 8090
rect 83096 8026 83148 8032
rect 82728 8016 82780 8022
rect 82728 7958 82780 7964
rect 83004 7948 83056 7954
rect 83004 7890 83056 7896
rect 83016 7546 83044 7890
rect 83004 7540 83056 7546
rect 83004 7482 83056 7488
rect 82636 6860 82688 6866
rect 82636 6802 82688 6808
rect 83004 6792 83056 6798
rect 83004 6734 83056 6740
rect 82912 6248 82964 6254
rect 82912 6190 82964 6196
rect 82544 5908 82596 5914
rect 82544 5850 82596 5856
rect 82924 4826 82952 6190
rect 82912 4820 82964 4826
rect 82912 4762 82964 4768
rect 82268 4140 82320 4146
rect 82268 4082 82320 4088
rect 82084 3596 82136 3602
rect 82084 3538 82136 3544
rect 81992 2032 82044 2038
rect 81992 1974 82044 1980
rect 81716 1964 81768 1970
rect 81716 1906 81768 1912
rect 81624 1760 81676 1766
rect 81624 1702 81676 1708
rect 81440 1556 81492 1562
rect 81440 1498 81492 1504
rect 81636 800 81664 1702
rect 82096 800 82124 3538
rect 82912 2916 82964 2922
rect 82912 2858 82964 2864
rect 82544 2440 82596 2446
rect 82544 2382 82596 2388
rect 82176 1896 82228 1902
rect 82176 1838 82228 1844
rect 82188 1562 82216 1838
rect 82176 1556 82228 1562
rect 82176 1498 82228 1504
rect 82556 800 82584 2382
rect 82924 800 82952 2858
rect 83016 2038 83044 6734
rect 83108 2650 83136 8026
rect 83280 7948 83332 7954
rect 83280 7890 83332 7896
rect 83188 7336 83240 7342
rect 83188 7278 83240 7284
rect 83200 3534 83228 7278
rect 83292 3738 83320 7890
rect 83384 6866 83412 10200
rect 83844 9654 83872 10200
rect 84076 9820 84132 9840
rect 84076 9744 84132 9764
rect 83832 9648 83884 9654
rect 83832 9590 83884 9596
rect 83556 8968 83608 8974
rect 83556 8910 83608 8916
rect 83568 8498 83596 8910
rect 84076 8732 84132 8752
rect 84076 8656 84132 8676
rect 83924 8628 83976 8634
rect 83924 8570 83976 8576
rect 83556 8492 83608 8498
rect 83556 8434 83608 8440
rect 83832 7540 83884 7546
rect 83832 7482 83884 7488
rect 83372 6860 83424 6866
rect 83372 6802 83424 6808
rect 83464 6656 83516 6662
rect 83464 6598 83516 6604
rect 83476 6254 83504 6598
rect 83464 6248 83516 6254
rect 83464 6190 83516 6196
rect 83372 5908 83424 5914
rect 83372 5850 83424 5856
rect 83384 5778 83412 5850
rect 83372 5772 83424 5778
rect 83372 5714 83424 5720
rect 83844 4078 83872 7482
rect 83936 5284 83964 8570
rect 84076 7644 84132 7664
rect 84076 7568 84132 7588
rect 84304 6798 84332 10200
rect 84384 8356 84436 8362
rect 84384 8298 84436 8304
rect 84292 6792 84344 6798
rect 84292 6734 84344 6740
rect 84076 6556 84132 6576
rect 84076 6480 84132 6500
rect 84076 5468 84132 5488
rect 84076 5392 84132 5412
rect 83936 5256 84056 5284
rect 83924 4684 83976 4690
rect 83924 4626 83976 4632
rect 83832 4072 83884 4078
rect 83832 4014 83884 4020
rect 83740 3936 83792 3942
rect 83740 3878 83792 3884
rect 83832 3936 83884 3942
rect 83832 3878 83884 3884
rect 83752 3738 83780 3878
rect 83280 3732 83332 3738
rect 83280 3674 83332 3680
rect 83740 3732 83792 3738
rect 83740 3674 83792 3680
rect 83188 3528 83240 3534
rect 83188 3470 83240 3476
rect 83096 2644 83148 2650
rect 83096 2586 83148 2592
rect 83004 2032 83056 2038
rect 83004 1974 83056 1980
rect 83280 2032 83332 2038
rect 83280 1974 83332 1980
rect 83292 1562 83320 1974
rect 83372 1760 83424 1766
rect 83372 1702 83424 1708
rect 83280 1556 83332 1562
rect 83280 1498 83332 1504
rect 83384 800 83412 1702
rect 83844 800 83872 3878
rect 83936 3602 83964 4626
rect 84028 4570 84056 5256
rect 84396 4690 84424 8298
rect 84672 8294 84700 10200
rect 84660 8288 84712 8294
rect 84660 8230 84712 8236
rect 85132 6866 85160 10200
rect 85592 9602 85620 10200
rect 86052 9926 86080 10200
rect 86040 9920 86092 9926
rect 86040 9862 86092 9868
rect 85856 9716 85908 9722
rect 85856 9658 85908 9664
rect 85592 9574 85804 9602
rect 85580 9376 85632 9382
rect 85580 9318 85632 9324
rect 85672 9376 85724 9382
rect 85672 9318 85724 9324
rect 85488 9104 85540 9110
rect 85488 9046 85540 9052
rect 85500 8022 85528 9046
rect 85488 8016 85540 8022
rect 85488 7958 85540 7964
rect 85304 7880 85356 7886
rect 85304 7822 85356 7828
rect 85120 6860 85172 6866
rect 85120 6802 85172 6808
rect 84660 6656 84712 6662
rect 84660 6598 84712 6604
rect 84384 4684 84436 4690
rect 84384 4626 84436 4632
rect 84028 4542 84240 4570
rect 84076 4380 84132 4400
rect 84076 4304 84132 4324
rect 84212 4162 84240 4542
rect 84120 4134 84240 4162
rect 84292 4140 84344 4146
rect 84120 3942 84148 4134
rect 84292 4082 84344 4088
rect 84108 3936 84160 3942
rect 84108 3878 84160 3884
rect 84304 3602 84332 4082
rect 83924 3596 83976 3602
rect 83924 3538 83976 3544
rect 84292 3596 84344 3602
rect 84292 3538 84344 3544
rect 84292 3392 84344 3398
rect 84292 3334 84344 3340
rect 84076 3292 84132 3312
rect 84076 3216 84132 3236
rect 84076 2204 84132 2224
rect 84076 2128 84132 2148
rect 84076 1116 84132 1136
rect 84076 1040 84132 1060
rect 84304 800 84332 3334
rect 84672 1902 84700 6598
rect 85212 6248 85264 6254
rect 85212 6190 85264 6196
rect 85224 5914 85252 6190
rect 85212 5908 85264 5914
rect 85212 5850 85264 5856
rect 85120 2916 85172 2922
rect 85120 2858 85172 2864
rect 84660 1896 84712 1902
rect 84660 1838 84712 1844
rect 84660 1420 84712 1426
rect 84660 1362 84712 1368
rect 84672 800 84700 1362
rect 85132 800 85160 2858
rect 85316 2514 85344 7822
rect 85592 7342 85620 9318
rect 85684 8430 85712 9318
rect 85672 8424 85724 8430
rect 85672 8366 85724 8372
rect 85672 8288 85724 8294
rect 85672 8230 85724 8236
rect 85684 7954 85712 8230
rect 85672 7948 85724 7954
rect 85672 7890 85724 7896
rect 85776 7750 85804 9574
rect 85868 8974 85896 9658
rect 85948 9648 86000 9654
rect 85948 9590 86000 9596
rect 85960 9042 85988 9590
rect 86132 9580 86184 9586
rect 86132 9522 86184 9528
rect 85948 9036 86000 9042
rect 85948 8978 86000 8984
rect 85856 8968 85908 8974
rect 85856 8910 85908 8916
rect 85948 8424 86000 8430
rect 85948 8366 86000 8372
rect 85764 7744 85816 7750
rect 85764 7686 85816 7692
rect 85580 7336 85632 7342
rect 85580 7278 85632 7284
rect 85856 7336 85908 7342
rect 85856 7278 85908 7284
rect 85764 6248 85816 6254
rect 85764 6190 85816 6196
rect 85580 4684 85632 4690
rect 85580 4626 85632 4632
rect 85592 4146 85620 4626
rect 85672 4480 85724 4486
rect 85672 4422 85724 4428
rect 85580 4140 85632 4146
rect 85580 4082 85632 4088
rect 85304 2508 85356 2514
rect 85304 2450 85356 2456
rect 85580 1760 85632 1766
rect 85580 1702 85632 1708
rect 85592 800 85620 1702
rect 85684 1426 85712 4422
rect 85776 2990 85804 6190
rect 85764 2984 85816 2990
rect 85764 2926 85816 2932
rect 85868 1902 85896 7278
rect 85960 2582 85988 8366
rect 86144 4146 86172 9522
rect 86316 7880 86368 7886
rect 86316 7822 86368 7828
rect 86132 4140 86184 4146
rect 86132 4082 86184 4088
rect 86040 4072 86092 4078
rect 86040 4014 86092 4020
rect 86052 3602 86080 4014
rect 86040 3596 86092 3602
rect 86040 3538 86092 3544
rect 86040 3392 86092 3398
rect 86040 3334 86092 3340
rect 85948 2576 86000 2582
rect 85948 2518 86000 2524
rect 85856 1896 85908 1902
rect 85856 1838 85908 1844
rect 85672 1420 85724 1426
rect 85672 1362 85724 1368
rect 86052 800 86080 3334
rect 86328 1562 86356 7822
rect 86420 4690 86448 10200
rect 86880 6254 86908 10200
rect 87236 9444 87288 9450
rect 87236 9386 87288 9392
rect 86960 9172 87012 9178
rect 86960 9114 87012 9120
rect 86972 8498 87000 9114
rect 86960 8492 87012 8498
rect 86960 8434 87012 8440
rect 87248 8430 87276 9386
rect 87236 8424 87288 8430
rect 87236 8366 87288 8372
rect 86960 7812 87012 7818
rect 86960 7754 87012 7760
rect 86972 6934 87000 7754
rect 87340 7478 87368 10200
rect 87800 7546 87828 10200
rect 87788 7540 87840 7546
rect 87788 7482 87840 7488
rect 87328 7472 87380 7478
rect 87328 7414 87380 7420
rect 87328 7336 87380 7342
rect 87328 7278 87380 7284
rect 86960 6928 87012 6934
rect 86960 6870 87012 6876
rect 86868 6248 86920 6254
rect 86868 6190 86920 6196
rect 87144 6248 87196 6254
rect 87144 6190 87196 6196
rect 86776 5160 86828 5166
rect 86776 5102 86828 5108
rect 86408 4684 86460 4690
rect 86408 4626 86460 4632
rect 86788 1873 86816 5102
rect 86868 4072 86920 4078
rect 86868 4014 86920 4020
rect 86774 1864 86830 1873
rect 86774 1799 86830 1808
rect 86316 1556 86368 1562
rect 86316 1498 86368 1504
rect 86408 1352 86460 1358
rect 86408 1294 86460 1300
rect 86420 800 86448 1294
rect 86880 800 86908 4014
rect 87156 3058 87184 6190
rect 87236 4004 87288 4010
rect 87236 3946 87288 3952
rect 87248 3126 87276 3946
rect 87236 3120 87288 3126
rect 87236 3062 87288 3068
rect 87144 3052 87196 3058
rect 87144 2994 87196 3000
rect 87340 2990 87368 7278
rect 88168 6254 88196 10200
rect 88628 8838 88656 10200
rect 88616 8832 88668 8838
rect 88616 8774 88668 8780
rect 88340 8424 88392 8430
rect 88340 8366 88392 8372
rect 88892 8424 88944 8430
rect 88892 8366 88944 8372
rect 87420 6248 87472 6254
rect 87420 6190 87472 6196
rect 88156 6248 88208 6254
rect 88156 6190 88208 6196
rect 87328 2984 87380 2990
rect 87328 2926 87380 2932
rect 87328 1760 87380 1766
rect 87328 1702 87380 1708
rect 87340 800 87368 1702
rect 87432 1426 87460 6190
rect 87788 4072 87840 4078
rect 87788 4014 87840 4020
rect 87420 1420 87472 1426
rect 87420 1362 87472 1368
rect 87800 800 87828 4014
rect 88156 3528 88208 3534
rect 88156 3470 88208 3476
rect 88168 800 88196 3470
rect 88352 2650 88380 8366
rect 88800 7812 88852 7818
rect 88800 7754 88852 7760
rect 88432 6384 88484 6390
rect 88432 6326 88484 6332
rect 88340 2644 88392 2650
rect 88340 2586 88392 2592
rect 88444 1902 88472 6326
rect 88524 5160 88576 5166
rect 88524 5102 88576 5108
rect 88536 4826 88564 5102
rect 88708 5024 88760 5030
rect 88708 4966 88760 4972
rect 88720 4826 88748 4966
rect 88524 4820 88576 4826
rect 88524 4762 88576 4768
rect 88708 4820 88760 4826
rect 88708 4762 88760 4768
rect 88616 2440 88668 2446
rect 88616 2382 88668 2388
rect 88432 1896 88484 1902
rect 88432 1838 88484 1844
rect 88628 800 88656 2382
rect 88812 1902 88840 7754
rect 88904 4282 88932 8366
rect 89088 6236 89116 10200
rect 89456 9518 89484 10200
rect 89444 9512 89496 9518
rect 89444 9454 89496 9460
rect 89260 8968 89312 8974
rect 89260 8910 89312 8916
rect 89272 7410 89300 8910
rect 89352 7880 89404 7886
rect 89352 7822 89404 7828
rect 89260 7404 89312 7410
rect 89260 7346 89312 7352
rect 89260 6384 89312 6390
rect 89260 6326 89312 6332
rect 89168 6248 89220 6254
rect 89088 6208 89168 6236
rect 89168 6190 89220 6196
rect 88984 4820 89036 4826
rect 88984 4762 89036 4768
rect 88996 4622 89024 4762
rect 89272 4690 89300 6326
rect 89260 4684 89312 4690
rect 89260 4626 89312 4632
rect 88984 4616 89036 4622
rect 88984 4558 89036 4564
rect 88892 4276 88944 4282
rect 88892 4218 88944 4224
rect 89364 3602 89392 7822
rect 89916 6866 89944 10200
rect 90376 9058 90404 10200
rect 90284 9030 90404 9058
rect 90284 8294 90312 9030
rect 90364 8968 90416 8974
rect 90364 8910 90416 8916
rect 90272 8288 90324 8294
rect 90272 8230 90324 8236
rect 90088 7404 90140 7410
rect 90088 7346 90140 7352
rect 89904 6860 89956 6866
rect 89904 6802 89956 6808
rect 89812 6316 89864 6322
rect 89812 6258 89864 6264
rect 89720 5908 89772 5914
rect 89720 5850 89772 5856
rect 89628 5772 89680 5778
rect 89628 5714 89680 5720
rect 89352 3596 89404 3602
rect 89352 3538 89404 3544
rect 89640 3369 89668 5714
rect 89732 5642 89760 5850
rect 89720 5636 89772 5642
rect 89720 5578 89772 5584
rect 89626 3360 89682 3369
rect 89626 3295 89682 3304
rect 89824 3058 89852 6258
rect 89996 5296 90048 5302
rect 89994 5264 89996 5273
rect 90048 5264 90050 5273
rect 89994 5199 90050 5208
rect 89812 3052 89864 3058
rect 89812 2994 89864 3000
rect 89444 2916 89496 2922
rect 89444 2858 89496 2864
rect 89076 2440 89128 2446
rect 89076 2382 89128 2388
rect 88800 1896 88852 1902
rect 88800 1838 88852 1844
rect 89088 800 89116 2382
rect 89456 800 89484 2858
rect 89628 2576 89680 2582
rect 89628 2518 89680 2524
rect 89640 1426 89668 2518
rect 90100 2514 90128 7346
rect 90376 6866 90404 8910
rect 90836 8362 90864 10200
rect 91100 8628 91152 8634
rect 91100 8570 91152 8576
rect 90824 8356 90876 8362
rect 90824 8298 90876 8304
rect 90916 7948 90968 7954
rect 90916 7890 90968 7896
rect 90364 6860 90416 6866
rect 90364 6802 90416 6808
rect 90180 6656 90232 6662
rect 90180 6598 90232 6604
rect 90088 2508 90140 2514
rect 90088 2450 90140 2456
rect 89720 2440 89772 2446
rect 89720 2382 89772 2388
rect 89732 2038 89760 2382
rect 89720 2032 89772 2038
rect 89720 1974 89772 1980
rect 89904 1828 89956 1834
rect 89904 1770 89956 1776
rect 89628 1420 89680 1426
rect 89628 1362 89680 1368
rect 89916 800 89944 1770
rect 90192 1426 90220 6598
rect 90272 5160 90324 5166
rect 90272 5102 90324 5108
rect 90284 2553 90312 5102
rect 90456 4616 90508 4622
rect 90456 4558 90508 4564
rect 90468 4146 90496 4558
rect 90456 4140 90508 4146
rect 90456 4082 90508 4088
rect 90824 4004 90876 4010
rect 90824 3946 90876 3952
rect 90270 2544 90326 2553
rect 90270 2479 90326 2488
rect 90180 1420 90232 1426
rect 90180 1362 90232 1368
rect 90364 1420 90416 1426
rect 90364 1362 90416 1368
rect 90376 800 90404 1362
rect 90836 800 90864 3946
rect 90928 2854 90956 7890
rect 91008 7880 91060 7886
rect 91008 7822 91060 7828
rect 91020 3398 91048 7822
rect 91112 4078 91140 8570
rect 91204 7274 91232 10200
rect 91376 8288 91428 8294
rect 91376 8230 91428 8236
rect 91388 7954 91416 8230
rect 91664 8090 91692 10200
rect 91836 8968 91888 8974
rect 91836 8910 91888 8916
rect 91652 8084 91704 8090
rect 91652 8026 91704 8032
rect 91376 7948 91428 7954
rect 91376 7890 91428 7896
rect 91468 7336 91520 7342
rect 91468 7278 91520 7284
rect 91744 7336 91796 7342
rect 91744 7278 91796 7284
rect 91192 7268 91244 7274
rect 91192 7210 91244 7216
rect 91192 5772 91244 5778
rect 91192 5714 91244 5720
rect 91100 4072 91152 4078
rect 91100 4014 91152 4020
rect 91008 3392 91060 3398
rect 91008 3334 91060 3340
rect 90916 2848 90968 2854
rect 90916 2790 90968 2796
rect 91204 1562 91232 5714
rect 91376 5568 91428 5574
rect 91376 5510 91428 5516
rect 91284 3528 91336 3534
rect 91284 3470 91336 3476
rect 91192 1556 91244 1562
rect 91192 1498 91244 1504
rect 91296 1442 91324 3470
rect 91388 1902 91416 5510
rect 91480 2990 91508 7278
rect 91756 7002 91784 7278
rect 91744 6996 91796 7002
rect 91744 6938 91796 6944
rect 91652 6656 91704 6662
rect 91652 6598 91704 6604
rect 91560 6248 91612 6254
rect 91560 6190 91612 6196
rect 91572 6118 91600 6190
rect 91560 6112 91612 6118
rect 91560 6054 91612 6060
rect 91664 5166 91692 6598
rect 91744 6384 91796 6390
rect 91744 6326 91796 6332
rect 91756 6186 91784 6326
rect 91744 6180 91796 6186
rect 91744 6122 91796 6128
rect 91652 5160 91704 5166
rect 91652 5102 91704 5108
rect 91848 4554 91876 8910
rect 92124 6866 92152 10200
rect 92584 8786 92612 10200
rect 92400 8758 92612 8786
rect 92400 8566 92428 8758
rect 92388 8560 92440 8566
rect 92388 8502 92440 8508
rect 92572 7880 92624 7886
rect 92952 7834 92980 10200
rect 93412 8498 93440 10200
rect 93400 8492 93452 8498
rect 93400 8434 93452 8440
rect 93676 8492 93728 8498
rect 93676 8434 93728 8440
rect 92572 7822 92624 7828
rect 92112 6860 92164 6866
rect 92112 6802 92164 6808
rect 91926 5536 91982 5545
rect 91926 5471 91982 5480
rect 91940 4622 91968 5471
rect 92020 4684 92072 4690
rect 92020 4626 92072 4632
rect 92112 4684 92164 4690
rect 92112 4626 92164 4632
rect 91928 4616 91980 4622
rect 91928 4558 91980 4564
rect 91836 4548 91888 4554
rect 91836 4490 91888 4496
rect 91652 3596 91704 3602
rect 91652 3538 91704 3544
rect 91468 2984 91520 2990
rect 91468 2926 91520 2932
rect 91376 1896 91428 1902
rect 91376 1838 91428 1844
rect 91204 1414 91324 1442
rect 91204 800 91232 1414
rect 91664 800 91692 3538
rect 92032 2009 92060 4626
rect 92124 4282 92152 4626
rect 92112 4276 92164 4282
rect 92112 4218 92164 4224
rect 92584 4146 92612 7822
rect 92860 7818 92980 7834
rect 92848 7812 92980 7818
rect 92900 7806 92980 7812
rect 92848 7754 92900 7760
rect 93306 7440 93362 7449
rect 93306 7375 93362 7384
rect 93320 7342 93348 7375
rect 92848 7336 92900 7342
rect 92848 7278 92900 7284
rect 93308 7336 93360 7342
rect 93308 7278 93360 7284
rect 92756 5160 92808 5166
rect 92756 5102 92808 5108
rect 92572 4140 92624 4146
rect 92572 4082 92624 4088
rect 92768 3942 92796 5102
rect 92756 3936 92808 3942
rect 92756 3878 92808 3884
rect 92480 3460 92532 3466
rect 92480 3402 92532 3408
rect 92492 3194 92520 3402
rect 92480 3188 92532 3194
rect 92480 3130 92532 3136
rect 92572 2440 92624 2446
rect 92572 2382 92624 2388
rect 92756 2440 92808 2446
rect 92756 2382 92808 2388
rect 92018 2000 92074 2009
rect 92018 1935 92074 1944
rect 92112 1420 92164 1426
rect 92112 1362 92164 1368
rect 92124 800 92152 1362
rect 92584 800 92612 2382
rect 92768 1494 92796 2382
rect 92860 1902 92888 7278
rect 93584 6656 93636 6662
rect 93584 6598 93636 6604
rect 92940 6248 92992 6254
rect 92940 6190 92992 6196
rect 93124 6248 93176 6254
rect 93124 6190 93176 6196
rect 92952 2650 92980 6190
rect 93032 4616 93084 4622
rect 93032 4558 93084 4564
rect 93044 3602 93072 4558
rect 93032 3596 93084 3602
rect 93032 3538 93084 3544
rect 92940 2644 92992 2650
rect 92940 2586 92992 2592
rect 93032 1964 93084 1970
rect 93032 1906 93084 1912
rect 92848 1896 92900 1902
rect 92848 1838 92900 1844
rect 92940 1828 92992 1834
rect 92940 1770 92992 1776
rect 92756 1488 92808 1494
rect 92756 1430 92808 1436
rect 92952 800 92980 1770
rect 93044 1494 93072 1906
rect 93032 1488 93084 1494
rect 93032 1430 93084 1436
rect 93136 1426 93164 6190
rect 93400 4072 93452 4078
rect 93400 4014 93452 4020
rect 93216 2100 93268 2106
rect 93216 2042 93268 2048
rect 93228 1766 93256 2042
rect 93216 1760 93268 1766
rect 93216 1702 93268 1708
rect 93124 1420 93176 1426
rect 93124 1362 93176 1368
rect 93412 800 93440 4014
rect 93596 2990 93624 6598
rect 93584 2984 93636 2990
rect 93584 2926 93636 2932
rect 93688 1329 93716 8434
rect 93768 8424 93820 8430
rect 93768 8366 93820 8372
rect 93780 7585 93808 8366
rect 93766 7576 93822 7585
rect 93766 7511 93822 7520
rect 93872 6254 93900 10200
rect 94332 10010 94360 10200
rect 94240 9982 94360 10010
rect 94240 7410 94268 9982
rect 94320 9920 94372 9926
rect 94320 9862 94372 9868
rect 94332 9586 94360 9862
rect 94320 9580 94372 9586
rect 94320 9522 94372 9528
rect 94596 8084 94648 8090
rect 94596 8026 94648 8032
rect 94608 7954 94636 8026
rect 94596 7948 94648 7954
rect 94596 7890 94648 7896
rect 94596 7744 94648 7750
rect 94596 7686 94648 7692
rect 94504 7472 94556 7478
rect 94504 7414 94556 7420
rect 94228 7404 94280 7410
rect 94228 7346 94280 7352
rect 93860 6248 93912 6254
rect 93860 6190 93912 6196
rect 94516 5642 94544 7414
rect 94504 5636 94556 5642
rect 94504 5578 94556 5584
rect 94504 5364 94556 5370
rect 94504 5306 94556 5312
rect 93860 5160 93912 5166
rect 93860 5102 93912 5108
rect 93872 4128 93900 5102
rect 94320 4548 94372 4554
rect 94320 4490 94372 4496
rect 93780 4100 93900 4128
rect 93780 4010 93808 4100
rect 94332 4078 94360 4490
rect 94516 4282 94544 5306
rect 94504 4276 94556 4282
rect 94504 4218 94556 4224
rect 94320 4072 94372 4078
rect 93872 4010 94176 4026
rect 94320 4014 94372 4020
rect 93768 4004 93820 4010
rect 93768 3946 93820 3952
rect 93872 4004 94188 4010
rect 93872 3998 94136 4004
rect 93674 1320 93730 1329
rect 93674 1255 93730 1264
rect 93872 800 93900 3998
rect 94136 3946 94188 3952
rect 94504 3732 94556 3738
rect 94504 3674 94556 3680
rect 94516 3466 94544 3674
rect 94504 3460 94556 3466
rect 94504 3402 94556 3408
rect 94608 2990 94636 7686
rect 94700 5778 94728 10200
rect 95160 9042 95188 10200
rect 95424 9512 95476 9518
rect 95424 9454 95476 9460
rect 95148 9036 95200 9042
rect 95148 8978 95200 8984
rect 95436 8974 95464 9454
rect 95424 8968 95476 8974
rect 95424 8910 95476 8916
rect 95516 7948 95568 7954
rect 95516 7890 95568 7896
rect 95148 6860 95200 6866
rect 95148 6802 95200 6808
rect 95160 6390 95188 6802
rect 95148 6384 95200 6390
rect 95148 6326 95200 6332
rect 94964 6248 95016 6254
rect 94964 6190 95016 6196
rect 95148 6248 95200 6254
rect 95148 6190 95200 6196
rect 94688 5772 94740 5778
rect 94688 5714 94740 5720
rect 94780 5704 94832 5710
rect 94780 5646 94832 5652
rect 94688 5364 94740 5370
rect 94688 5306 94740 5312
rect 94700 5030 94728 5306
rect 94688 5024 94740 5030
rect 94688 4966 94740 4972
rect 94792 4146 94820 5646
rect 94872 5636 94924 5642
rect 94872 5578 94924 5584
rect 94780 4140 94832 4146
rect 94780 4082 94832 4088
rect 94688 3936 94740 3942
rect 94688 3878 94740 3884
rect 94596 2984 94648 2990
rect 94596 2926 94648 2932
rect 94320 2916 94372 2922
rect 94320 2858 94372 2864
rect 94332 800 94360 2858
rect 94504 2372 94556 2378
rect 94504 2314 94556 2320
rect 94516 2106 94544 2314
rect 94504 2100 94556 2106
rect 94504 2042 94556 2048
rect 94700 800 94728 3878
rect 94884 2514 94912 5578
rect 94976 3602 95004 6190
rect 95056 5024 95108 5030
rect 95056 4966 95108 4972
rect 94964 3596 95016 3602
rect 94964 3538 95016 3544
rect 95068 2582 95096 4966
rect 95056 2576 95108 2582
rect 95056 2518 95108 2524
rect 94872 2508 94924 2514
rect 94872 2450 94924 2456
rect 95160 1426 95188 6190
rect 95240 3188 95292 3194
rect 95240 3130 95292 3136
rect 95252 2446 95280 3130
rect 95240 2440 95292 2446
rect 95240 2382 95292 2388
rect 95528 1562 95556 7890
rect 95620 7818 95648 10200
rect 95700 10124 95752 10130
rect 95700 10066 95752 10072
rect 95608 7812 95660 7818
rect 95608 7754 95660 7760
rect 95712 5710 95740 10066
rect 96080 10010 96108 10200
rect 95896 9982 96108 10010
rect 95792 7812 95844 7818
rect 95792 7754 95844 7760
rect 95804 7342 95832 7754
rect 95792 7336 95844 7342
rect 95792 7278 95844 7284
rect 95896 7002 95924 9982
rect 96068 9920 96120 9926
rect 96068 9862 96120 9868
rect 96080 9518 96108 9862
rect 96068 9512 96120 9518
rect 96068 9454 96120 9460
rect 95976 9444 96028 9450
rect 95976 9386 96028 9392
rect 95884 6996 95936 7002
rect 95884 6938 95936 6944
rect 95700 5704 95752 5710
rect 95700 5646 95752 5652
rect 95792 4616 95844 4622
rect 95792 4558 95844 4564
rect 95608 4140 95660 4146
rect 95608 4082 95660 4088
rect 95516 1556 95568 1562
rect 95516 1498 95568 1504
rect 95240 1488 95292 1494
rect 95240 1430 95292 1436
rect 95148 1420 95200 1426
rect 95148 1362 95200 1368
rect 95252 1306 95280 1430
rect 95160 1278 95280 1306
rect 95160 800 95188 1278
rect 95620 800 95648 4082
rect 95804 3738 95832 4558
rect 95792 3732 95844 3738
rect 95792 3674 95844 3680
rect 95884 2984 95936 2990
rect 95884 2926 95936 2932
rect 95896 2582 95924 2926
rect 95884 2576 95936 2582
rect 95884 2518 95936 2524
rect 95988 1902 96016 9386
rect 96068 7948 96120 7954
rect 96068 7890 96120 7896
rect 96080 5522 96108 7890
rect 96158 7440 96214 7449
rect 96158 7375 96214 7384
rect 96172 7342 96200 7375
rect 96160 7336 96212 7342
rect 96160 7278 96212 7284
rect 96448 6882 96476 10200
rect 96908 9466 96936 10200
rect 96816 9438 96936 9466
rect 96712 8628 96764 8634
rect 96712 8570 96764 8576
rect 96620 8424 96672 8430
rect 96620 8366 96672 8372
rect 96528 6996 96580 7002
rect 96528 6938 96580 6944
rect 96356 6866 96476 6882
rect 96344 6860 96476 6866
rect 96396 6854 96476 6860
rect 96344 6802 96396 6808
rect 96252 6792 96304 6798
rect 96252 6734 96304 6740
rect 96080 5494 96200 5522
rect 96068 5364 96120 5370
rect 96068 5306 96120 5312
rect 95976 1896 96028 1902
rect 95976 1838 96028 1844
rect 96080 800 96108 5306
rect 96172 3738 96200 5494
rect 96160 3732 96212 3738
rect 96160 3674 96212 3680
rect 96264 1970 96292 6734
rect 96540 5250 96568 6938
rect 96356 5222 96568 5250
rect 96356 2582 96384 5222
rect 96528 5160 96580 5166
rect 96528 5102 96580 5108
rect 96540 4554 96568 5102
rect 96632 5030 96660 8366
rect 96724 6866 96752 8570
rect 96712 6860 96764 6866
rect 96712 6802 96764 6808
rect 96816 6254 96844 9438
rect 96896 9376 96948 9382
rect 96896 9318 96948 9324
rect 96988 9376 97040 9382
rect 96988 9318 97040 9324
rect 96908 7410 96936 9318
rect 97000 7954 97028 9318
rect 97080 9036 97132 9042
rect 97080 8978 97132 8984
rect 97092 8945 97120 8978
rect 97078 8936 97134 8945
rect 97078 8871 97134 8880
rect 97368 8514 97396 10200
rect 97540 10056 97592 10062
rect 97540 9998 97592 10004
rect 97448 8832 97500 8838
rect 97448 8774 97500 8780
rect 97276 8498 97396 8514
rect 97264 8492 97396 8498
rect 97316 8486 97396 8492
rect 97264 8434 97316 8440
rect 97080 8424 97132 8430
rect 97080 8366 97132 8372
rect 96988 7948 97040 7954
rect 96988 7890 97040 7896
rect 96896 7404 96948 7410
rect 96896 7346 96948 7352
rect 96804 6248 96856 6254
rect 96804 6190 96856 6196
rect 96896 6180 96948 6186
rect 96896 6122 96948 6128
rect 96908 6089 96936 6122
rect 96988 6112 97040 6118
rect 96894 6080 96950 6089
rect 96988 6054 97040 6060
rect 96894 6015 96950 6024
rect 97000 5778 97028 6054
rect 96804 5772 96856 5778
rect 96804 5714 96856 5720
rect 96988 5772 97040 5778
rect 96988 5714 97040 5720
rect 96712 5160 96764 5166
rect 96712 5102 96764 5108
rect 96620 5024 96672 5030
rect 96620 4966 96672 4972
rect 96724 4690 96752 5102
rect 96712 4684 96764 4690
rect 96712 4626 96764 4632
rect 96528 4548 96580 4554
rect 96528 4490 96580 4496
rect 96816 3194 96844 5714
rect 96804 3188 96856 3194
rect 96804 3130 96856 3136
rect 96896 2916 96948 2922
rect 96896 2858 96948 2864
rect 96344 2576 96396 2582
rect 96344 2518 96396 2524
rect 96252 1964 96304 1970
rect 96252 1906 96304 1912
rect 96436 1828 96488 1834
rect 96436 1770 96488 1776
rect 96448 800 96476 1770
rect 96908 800 96936 2858
rect 97092 1902 97120 8366
rect 97460 6866 97488 8774
rect 97552 8430 97580 9998
rect 97540 8424 97592 8430
rect 97540 8366 97592 8372
rect 97448 6860 97500 6866
rect 97448 6802 97500 6808
rect 97632 6656 97684 6662
rect 97632 6598 97684 6604
rect 97644 6361 97672 6598
rect 97630 6352 97686 6361
rect 97540 6316 97592 6322
rect 97630 6287 97686 6296
rect 97540 6258 97592 6264
rect 97356 6248 97408 6254
rect 97552 6225 97580 6258
rect 97356 6190 97408 6196
rect 97538 6216 97594 6225
rect 97368 4570 97396 6190
rect 97538 6151 97594 6160
rect 97736 5778 97764 10200
rect 97828 8974 97856 10270
rect 98182 10200 98238 11400
rect 98642 10200 98698 11400
rect 99102 10200 99158 11400
rect 99470 10200 99526 11400
rect 99930 10200 99986 11400
rect 100390 10200 100446 11400
rect 100850 10200 100906 11400
rect 101218 10200 101274 11400
rect 101678 10200 101734 11400
rect 102138 10200 102194 11400
rect 102598 10200 102654 11400
rect 102966 10200 103022 11400
rect 103426 10200 103482 11400
rect 103886 10200 103942 11400
rect 104254 10200 104310 11400
rect 104714 10200 104770 11400
rect 105174 10200 105230 11400
rect 105634 10200 105690 11400
rect 106002 10200 106058 11400
rect 106462 10200 106518 11400
rect 106922 10200 106978 11400
rect 107382 10200 107438 11400
rect 107750 10200 107806 11400
rect 108210 10200 108266 11400
rect 108670 10200 108726 11400
rect 109130 10200 109186 11400
rect 109498 10200 109554 11400
rect 109958 10200 110014 11400
rect 110418 10200 110474 11400
rect 110878 10200 110934 11400
rect 111246 10200 111302 11400
rect 111706 10200 111762 11400
rect 112166 10200 112222 11400
rect 112534 10200 112590 11400
rect 112994 10200 113050 11400
rect 113454 10200 113510 11400
rect 113914 10200 113970 11400
rect 114282 10200 114338 11400
rect 114742 10200 114798 11400
rect 115202 10200 115258 11400
rect 115662 10200 115718 11400
rect 116030 10200 116086 11400
rect 116490 10200 116546 11400
rect 116950 10200 117006 11400
rect 117410 10200 117466 11400
rect 117778 10200 117834 11400
rect 118238 10200 118294 11400
rect 118698 10200 118754 11400
rect 119158 10200 119214 11400
rect 119526 10200 119582 11400
rect 119804 10396 119856 10402
rect 119804 10338 119856 10344
rect 119712 10260 119764 10266
rect 119712 10202 119764 10208
rect 98000 9512 98052 9518
rect 98000 9454 98052 9460
rect 97908 9444 97960 9450
rect 97908 9386 97960 9392
rect 97920 9042 97948 9386
rect 97908 9036 97960 9042
rect 97908 8978 97960 8984
rect 97816 8968 97868 8974
rect 97816 8910 97868 8916
rect 98012 8514 98040 9454
rect 98092 8968 98144 8974
rect 98092 8910 98144 8916
rect 97920 8486 98040 8514
rect 97920 8090 97948 8486
rect 98000 8356 98052 8362
rect 98000 8298 98052 8304
rect 98012 8090 98040 8298
rect 97908 8084 97960 8090
rect 97908 8026 97960 8032
rect 98000 8084 98052 8090
rect 98000 8026 98052 8032
rect 97908 6928 97960 6934
rect 97908 6870 97960 6876
rect 97816 6656 97868 6662
rect 97816 6598 97868 6604
rect 97724 5772 97776 5778
rect 97724 5714 97776 5720
rect 97276 4542 97396 4570
rect 97276 2514 97304 4542
rect 97632 3664 97684 3670
rect 97632 3606 97684 3612
rect 97356 3528 97408 3534
rect 97644 3505 97672 3606
rect 97724 3596 97776 3602
rect 97828 3584 97856 6598
rect 97776 3556 97856 3584
rect 97724 3538 97776 3544
rect 97356 3470 97408 3476
rect 97630 3496 97686 3505
rect 97264 2508 97316 2514
rect 97264 2450 97316 2456
rect 97080 1896 97132 1902
rect 97080 1838 97132 1844
rect 96988 1760 97040 1766
rect 96988 1702 97040 1708
rect 97000 1562 97028 1702
rect 96988 1556 97040 1562
rect 96988 1498 97040 1504
rect 97368 800 97396 3470
rect 97630 3431 97686 3440
rect 97724 3392 97776 3398
rect 97724 3334 97776 3340
rect 97736 800 97764 3334
rect 97920 2378 97948 6870
rect 98000 6724 98052 6730
rect 98000 6666 98052 6672
rect 98012 6254 98040 6666
rect 98000 6248 98052 6254
rect 98000 6190 98052 6196
rect 98104 2514 98132 8910
rect 98196 7342 98224 10200
rect 98656 9518 98684 10200
rect 98644 9512 98696 9518
rect 98644 9454 98696 9460
rect 99116 9058 99144 10200
rect 99380 9512 99432 9518
rect 99380 9454 99432 9460
rect 99196 9376 99248 9382
rect 99196 9318 99248 9324
rect 99208 9110 99236 9318
rect 99288 9172 99340 9178
rect 99288 9114 99340 9120
rect 98472 9030 99144 9058
rect 99196 9104 99248 9110
rect 99196 9046 99248 9052
rect 98472 7954 98500 9030
rect 99104 8968 99156 8974
rect 99104 8910 99156 8916
rect 98552 8560 98604 8566
rect 98552 8502 98604 8508
rect 98460 7948 98512 7954
rect 98460 7890 98512 7896
rect 98368 7880 98420 7886
rect 98368 7822 98420 7828
rect 98276 7472 98328 7478
rect 98276 7414 98328 7420
rect 98184 7336 98236 7342
rect 98184 7278 98236 7284
rect 98288 6769 98316 7414
rect 98274 6760 98330 6769
rect 98274 6695 98330 6704
rect 98184 5704 98236 5710
rect 98184 5646 98236 5652
rect 98196 5166 98224 5646
rect 98184 5160 98236 5166
rect 98184 5102 98236 5108
rect 98092 2508 98144 2514
rect 98092 2450 98144 2456
rect 97908 2372 97960 2378
rect 97908 2314 97960 2320
rect 98276 2304 98328 2310
rect 98276 2246 98328 2252
rect 98288 1834 98316 2246
rect 98184 1828 98236 1834
rect 98184 1770 98236 1776
rect 98276 1828 98328 1834
rect 98276 1770 98328 1776
rect 98196 800 98224 1770
rect 202 -400 258 800
rect 570 -400 626 800
rect 1030 -400 1086 800
rect 1490 -400 1546 800
rect 1858 -400 1914 800
rect 2318 -400 2374 800
rect 2778 -400 2834 800
rect 3238 -400 3294 800
rect 3606 -400 3662 800
rect 4066 -400 4122 800
rect 4526 -400 4582 800
rect 4986 -400 5042 800
rect 5354 -400 5410 800
rect 5814 -400 5870 800
rect 6274 -400 6330 800
rect 6734 -400 6790 800
rect 7102 -400 7158 800
rect 7562 -400 7618 800
rect 8022 -400 8078 800
rect 8390 -400 8446 800
rect 8850 -400 8906 800
rect 9310 -400 9366 800
rect 9770 -400 9826 800
rect 10138 -400 10194 800
rect 10598 -400 10654 800
rect 11058 -400 11114 800
rect 11518 -400 11574 800
rect 11886 -400 11942 800
rect 12346 -400 12402 800
rect 12806 -400 12862 800
rect 13266 -400 13322 800
rect 13634 -400 13690 800
rect 14094 -400 14150 800
rect 14554 -400 14610 800
rect 15014 -400 15070 800
rect 15382 -400 15438 800
rect 15842 -400 15898 800
rect 16302 -400 16358 800
rect 16670 -400 16726 800
rect 17130 -400 17186 800
rect 17590 -400 17646 800
rect 18050 -400 18106 800
rect 18418 -400 18474 800
rect 18878 -400 18934 800
rect 19338 -400 19394 800
rect 19798 -400 19854 800
rect 20166 -400 20222 800
rect 20626 -400 20682 800
rect 21086 -400 21142 800
rect 21546 -400 21602 800
rect 21914 -400 21970 800
rect 22374 -400 22430 800
rect 22834 -400 22890 800
rect 23294 -400 23350 800
rect 23662 -400 23718 800
rect 24122 -400 24178 800
rect 24582 -400 24638 800
rect 24950 -400 25006 800
rect 25410 -400 25466 800
rect 25870 -400 25926 800
rect 26330 -400 26386 800
rect 26698 -400 26754 800
rect 27158 -400 27214 800
rect 27618 -400 27674 800
rect 28078 -400 28134 800
rect 28446 -400 28502 800
rect 28906 -400 28962 800
rect 29366 -400 29422 800
rect 29826 -400 29882 800
rect 30194 -400 30250 800
rect 30654 -400 30710 800
rect 31114 -400 31170 800
rect 31574 -400 31630 800
rect 31942 -400 31998 800
rect 32402 -400 32458 800
rect 32862 -400 32918 800
rect 33230 -400 33286 800
rect 33690 -400 33746 800
rect 34150 -400 34206 800
rect 34610 -400 34666 800
rect 34978 -400 35034 800
rect 35438 -400 35494 800
rect 35898 -400 35954 800
rect 36358 -400 36414 800
rect 36726 -400 36782 800
rect 37186 -400 37242 800
rect 37646 -400 37702 800
rect 38106 -400 38162 800
rect 38474 -400 38530 800
rect 38934 -400 38990 800
rect 39394 -400 39450 800
rect 39854 -400 39910 800
rect 40222 -400 40278 800
rect 40682 -400 40738 800
rect 41142 -400 41198 800
rect 41510 -400 41566 800
rect 41970 -400 42026 800
rect 42430 -400 42486 800
rect 42890 -400 42946 800
rect 43258 -400 43314 800
rect 43718 -400 43774 800
rect 44178 -400 44234 800
rect 44638 -400 44694 800
rect 45006 -400 45062 800
rect 45466 -400 45522 800
rect 45926 -400 45982 800
rect 46386 -400 46442 800
rect 46754 -400 46810 800
rect 47214 -400 47270 800
rect 47674 -400 47730 800
rect 48134 -400 48190 800
rect 48502 -400 48558 800
rect 48962 -400 49018 800
rect 49422 -400 49478 800
rect 49790 -400 49846 800
rect 50250 -400 50306 800
rect 50710 -400 50766 800
rect 51170 -400 51226 800
rect 51538 -400 51594 800
rect 51998 -400 52054 800
rect 52458 -400 52514 800
rect 52918 -400 52974 800
rect 53286 -400 53342 800
rect 53746 -400 53802 800
rect 54206 -400 54262 800
rect 54666 -400 54722 800
rect 55034 -400 55090 800
rect 55494 -400 55550 800
rect 55954 -400 56010 800
rect 56322 -400 56378 800
rect 56782 -400 56838 800
rect 57242 -400 57298 800
rect 57702 -400 57758 800
rect 58070 -400 58126 800
rect 58530 -400 58586 800
rect 58990 -400 59046 800
rect 59450 -400 59506 800
rect 59818 -400 59874 800
rect 60278 -400 60334 800
rect 60738 -400 60794 800
rect 61198 -400 61254 800
rect 61566 -400 61622 800
rect 62026 -400 62082 800
rect 62486 -400 62542 800
rect 62946 -400 63002 800
rect 63314 -400 63370 800
rect 63774 -400 63830 800
rect 64234 -400 64290 800
rect 64602 -400 64658 800
rect 65062 -400 65118 800
rect 65522 -400 65578 800
rect 65982 -400 66038 800
rect 66350 -400 66406 800
rect 66810 -400 66866 800
rect 67270 -400 67326 800
rect 67730 -400 67786 800
rect 68098 -400 68154 800
rect 68558 -400 68614 800
rect 69018 -400 69074 800
rect 69478 -400 69534 800
rect 69846 -400 69902 800
rect 70306 -400 70362 800
rect 70766 -400 70822 800
rect 71226 -400 71282 800
rect 71594 -400 71650 800
rect 72054 -400 72110 800
rect 72514 -400 72570 800
rect 72882 -400 72938 800
rect 73342 -400 73398 800
rect 73802 -400 73858 800
rect 74262 -400 74318 800
rect 74630 -400 74686 800
rect 75090 -400 75146 800
rect 75550 -400 75606 800
rect 76010 -400 76066 800
rect 76378 -400 76434 800
rect 76838 -400 76894 800
rect 77298 -400 77354 800
rect 77758 -400 77814 800
rect 78126 -400 78182 800
rect 78586 -400 78642 800
rect 79046 -400 79102 800
rect 79506 -400 79562 800
rect 79874 -400 79930 800
rect 80334 -400 80390 800
rect 80794 -400 80850 800
rect 81162 -400 81218 800
rect 81622 -400 81678 800
rect 82082 -400 82138 800
rect 82542 -400 82598 800
rect 82910 -400 82966 800
rect 83370 -400 83426 800
rect 83830 -400 83886 800
rect 84290 -400 84346 800
rect 84658 -400 84714 800
rect 85118 -400 85174 800
rect 85578 -400 85634 800
rect 86038 -400 86094 800
rect 86406 -400 86462 800
rect 86866 -400 86922 800
rect 87326 -400 87382 800
rect 87786 -400 87842 800
rect 88154 -400 88210 800
rect 88614 -400 88670 800
rect 89074 -400 89130 800
rect 89442 -400 89498 800
rect 89902 -400 89958 800
rect 90362 -400 90418 800
rect 90822 -400 90878 800
rect 91190 -400 91246 800
rect 91650 -400 91706 800
rect 92110 -400 92166 800
rect 92570 -400 92626 800
rect 92938 -400 92994 800
rect 93398 -400 93454 800
rect 93858 -400 93914 800
rect 94318 -400 94374 800
rect 94686 -400 94742 800
rect 95146 -400 95202 800
rect 95606 -400 95662 800
rect 96066 -400 96122 800
rect 96434 -400 96490 800
rect 96894 -400 96950 800
rect 97354 -400 97410 800
rect 97722 -400 97778 800
rect 98182 -400 98238 800
rect 98380 241 98408 7822
rect 98460 7472 98512 7478
rect 98458 7440 98460 7449
rect 98512 7440 98514 7449
rect 98458 7375 98514 7384
rect 98564 4078 98592 8502
rect 99116 8430 99144 8910
rect 99104 8424 99156 8430
rect 99104 8366 99156 8372
rect 99300 8294 99328 9114
rect 99288 8288 99340 8294
rect 99288 8230 99340 8236
rect 98828 7948 98880 7954
rect 98828 7890 98880 7896
rect 98840 7834 98868 7890
rect 98656 7818 98868 7834
rect 98644 7812 98868 7818
rect 98696 7806 98868 7812
rect 98644 7754 98696 7760
rect 99392 7732 99420 9454
rect 99484 8362 99512 10200
rect 99944 9926 99972 10200
rect 99932 9920 99984 9926
rect 99932 9862 99984 9868
rect 99564 9376 99616 9382
rect 99564 9318 99616 9324
rect 99576 8634 99604 9318
rect 99932 8968 99984 8974
rect 99932 8910 99984 8916
rect 99564 8628 99616 8634
rect 99564 8570 99616 8576
rect 99472 8356 99524 8362
rect 99472 8298 99524 8304
rect 99944 8022 99972 8910
rect 99932 8016 99984 8022
rect 99932 7958 99984 7964
rect 99472 7880 99524 7886
rect 99472 7822 99524 7828
rect 99564 7880 99616 7886
rect 99564 7822 99616 7828
rect 99300 7704 99420 7732
rect 99194 6896 99250 6905
rect 99194 6831 99250 6840
rect 99208 6662 99236 6831
rect 99300 6798 99328 7704
rect 99484 7546 99512 7822
rect 99472 7540 99524 7546
rect 99472 7482 99524 7488
rect 99380 7336 99432 7342
rect 99380 7278 99432 7284
rect 99392 7002 99420 7278
rect 99472 7200 99524 7206
rect 99472 7142 99524 7148
rect 99484 7002 99512 7142
rect 99380 6996 99432 7002
rect 99380 6938 99432 6944
rect 99472 6996 99524 7002
rect 99472 6938 99524 6944
rect 99576 6866 99604 7822
rect 99656 7404 99708 7410
rect 99656 7346 99708 7352
rect 99564 6860 99616 6866
rect 99564 6802 99616 6808
rect 99288 6792 99340 6798
rect 99288 6734 99340 6740
rect 99196 6656 99248 6662
rect 99196 6598 99248 6604
rect 99288 6384 99340 6390
rect 99286 6352 99288 6361
rect 99340 6352 99342 6361
rect 99286 6287 99342 6296
rect 98644 6248 98696 6254
rect 98644 6190 98696 6196
rect 98828 6248 98880 6254
rect 99472 6248 99524 6254
rect 98828 6190 98880 6196
rect 99286 6216 99342 6225
rect 98656 5574 98684 6190
rect 98644 5568 98696 5574
rect 98644 5510 98696 5516
rect 98552 4072 98604 4078
rect 98552 4014 98604 4020
rect 98644 4004 98696 4010
rect 98644 3946 98696 3952
rect 98656 800 98684 3946
rect 98840 2990 98868 6190
rect 99286 6151 99342 6160
rect 99470 6216 99472 6225
rect 99524 6216 99526 6225
rect 99470 6151 99526 6160
rect 99300 6118 99328 6151
rect 99012 6112 99064 6118
rect 99012 6054 99064 6060
rect 99288 6112 99340 6118
rect 99288 6054 99340 6060
rect 98920 3936 98972 3942
rect 98920 3878 98972 3884
rect 98828 2984 98880 2990
rect 98828 2926 98880 2932
rect 98932 1494 98960 3878
rect 99024 3738 99052 6054
rect 99470 5944 99526 5953
rect 99668 5914 99696 7346
rect 100404 7342 100432 10200
rect 100864 9042 100892 10200
rect 100852 9036 100904 9042
rect 100852 8978 100904 8984
rect 100944 7744 100996 7750
rect 100944 7686 100996 7692
rect 100956 7410 100984 7686
rect 100760 7404 100812 7410
rect 100760 7346 100812 7352
rect 100944 7404 100996 7410
rect 100944 7346 100996 7352
rect 100392 7336 100444 7342
rect 100392 7278 100444 7284
rect 99746 6896 99802 6905
rect 99746 6831 99748 6840
rect 99800 6831 99802 6840
rect 99748 6802 99800 6808
rect 99746 6760 99802 6769
rect 99746 6695 99802 6704
rect 99470 5879 99472 5888
rect 99524 5879 99526 5888
rect 99656 5908 99708 5914
rect 99472 5850 99524 5856
rect 99656 5850 99708 5856
rect 99286 5808 99342 5817
rect 99104 5772 99156 5778
rect 99286 5743 99342 5752
rect 99104 5714 99156 5720
rect 99116 4128 99144 5714
rect 99300 5710 99328 5743
rect 99288 5704 99340 5710
rect 99288 5646 99340 5652
rect 99472 5704 99524 5710
rect 99472 5646 99524 5652
rect 99484 5234 99512 5646
rect 99472 5228 99524 5234
rect 99472 5170 99524 5176
rect 99288 4752 99340 4758
rect 99288 4694 99340 4700
rect 99196 4140 99248 4146
rect 99116 4100 99196 4128
rect 99196 4082 99248 4088
rect 99012 3732 99064 3738
rect 99012 3674 99064 3680
rect 99300 3126 99328 4694
rect 99760 3602 99788 6695
rect 100116 6384 100168 6390
rect 100116 6326 100168 6332
rect 99932 6316 99984 6322
rect 99984 6276 100064 6304
rect 99932 6258 99984 6264
rect 100036 6118 100064 6276
rect 100024 6112 100076 6118
rect 100128 6089 100156 6326
rect 100576 6316 100628 6322
rect 100576 6258 100628 6264
rect 100024 6054 100076 6060
rect 100114 6080 100170 6089
rect 100114 6015 100170 6024
rect 100208 4276 100260 4282
rect 100208 4218 100260 4224
rect 100116 4140 100168 4146
rect 100116 4082 100168 4088
rect 99748 3596 99800 3602
rect 99748 3538 99800 3544
rect 99196 3120 99248 3126
rect 99196 3062 99248 3068
rect 99288 3120 99340 3126
rect 99288 3062 99340 3068
rect 99104 2440 99156 2446
rect 99104 2382 99156 2388
rect 98920 1488 98972 1494
rect 98920 1430 98972 1436
rect 99116 800 99144 2382
rect 99208 1222 99236 3062
rect 99472 3052 99524 3058
rect 99472 2994 99524 3000
rect 99288 1488 99340 1494
rect 99288 1430 99340 1436
rect 99300 1290 99328 1430
rect 99288 1284 99340 1290
rect 99288 1226 99340 1232
rect 99196 1216 99248 1222
rect 99196 1158 99248 1164
rect 99484 800 99512 2994
rect 99932 2576 99984 2582
rect 99932 2518 99984 2524
rect 99944 800 99972 2518
rect 100128 2310 100156 4082
rect 100116 2304 100168 2310
rect 100116 2246 100168 2252
rect 100220 2106 100248 4218
rect 100588 2990 100616 6258
rect 100772 4078 100800 7346
rect 101232 6118 101260 10200
rect 101496 7336 101548 7342
rect 101496 7278 101548 7284
rect 101220 6112 101272 6118
rect 101220 6054 101272 6060
rect 101218 5400 101274 5409
rect 101218 5335 101220 5344
rect 101272 5335 101274 5344
rect 101220 5306 101272 5312
rect 100760 4072 100812 4078
rect 100760 4014 100812 4020
rect 101508 3942 101536 7278
rect 101692 6730 101720 10200
rect 102048 8968 102100 8974
rect 102048 8910 102100 8916
rect 102060 8498 102088 8910
rect 102048 8492 102100 8498
rect 102048 8434 102100 8440
rect 102152 7954 102180 10200
rect 102612 8838 102640 10200
rect 102600 8832 102652 8838
rect 102600 8774 102652 8780
rect 102232 8288 102284 8294
rect 102232 8230 102284 8236
rect 102244 7954 102272 8230
rect 102140 7948 102192 7954
rect 102140 7890 102192 7896
rect 102232 7948 102284 7954
rect 102232 7890 102284 7896
rect 102784 7472 102836 7478
rect 102784 7414 102836 7420
rect 102232 7200 102284 7206
rect 102232 7142 102284 7148
rect 101680 6724 101732 6730
rect 101680 6666 101732 6672
rect 102140 4684 102192 4690
rect 102140 4626 102192 4632
rect 102152 3942 102180 4626
rect 101496 3936 101548 3942
rect 101496 3878 101548 3884
rect 102140 3936 102192 3942
rect 102140 3878 102192 3884
rect 101680 3392 101732 3398
rect 101680 3334 101732 3340
rect 101220 3052 101272 3058
rect 101220 2994 101272 3000
rect 100576 2984 100628 2990
rect 100576 2926 100628 2932
rect 100392 2916 100444 2922
rect 100392 2858 100444 2864
rect 100208 2100 100260 2106
rect 100208 2042 100260 2048
rect 100404 800 100432 2858
rect 100668 2848 100720 2854
rect 100668 2790 100720 2796
rect 100680 1834 100708 2790
rect 101126 2136 101182 2145
rect 101126 2071 101182 2080
rect 100852 1964 100904 1970
rect 100852 1906 100904 1912
rect 100668 1828 100720 1834
rect 100668 1770 100720 1776
rect 100864 800 100892 1906
rect 101140 1902 101168 2071
rect 101128 1896 101180 1902
rect 101128 1838 101180 1844
rect 101232 800 101260 2994
rect 101692 800 101720 3334
rect 102140 2916 102192 2922
rect 102140 2858 102192 2864
rect 102152 800 102180 2858
rect 102244 1426 102272 7142
rect 102692 6724 102744 6730
rect 102692 6666 102744 6672
rect 102704 5953 102732 6666
rect 102690 5944 102746 5953
rect 102690 5879 102746 5888
rect 102600 4820 102652 4826
rect 102600 4762 102652 4768
rect 102508 4616 102560 4622
rect 102508 4558 102560 4564
rect 102416 4480 102468 4486
rect 102416 4422 102468 4428
rect 102428 4214 102456 4422
rect 102416 4208 102468 4214
rect 102416 4150 102468 4156
rect 102520 4146 102548 4558
rect 102612 4486 102640 4762
rect 102600 4480 102652 4486
rect 102600 4422 102652 4428
rect 102508 4140 102560 4146
rect 102508 4082 102560 4088
rect 102600 2440 102652 2446
rect 102600 2382 102652 2388
rect 102232 1420 102284 1426
rect 102232 1362 102284 1368
rect 102612 800 102640 2382
rect 102796 1902 102824 7414
rect 102980 6225 103008 10200
rect 103060 8968 103112 8974
rect 103060 8910 103112 8916
rect 103072 6866 103100 8910
rect 103440 7886 103468 10200
rect 103520 8628 103572 8634
rect 103520 8570 103572 8576
rect 103428 7880 103480 7886
rect 103428 7822 103480 7828
rect 103060 6860 103112 6866
rect 103060 6802 103112 6808
rect 102966 6216 103022 6225
rect 102966 6151 103022 6160
rect 103060 5568 103112 5574
rect 103060 5510 103112 5516
rect 103152 5568 103204 5574
rect 103152 5510 103204 5516
rect 102876 5160 102928 5166
rect 102876 5102 102928 5108
rect 102888 4729 102916 5102
rect 102874 4720 102930 4729
rect 102874 4655 102930 4664
rect 103072 3738 103100 5510
rect 103060 3732 103112 3738
rect 103060 3674 103112 3680
rect 103164 2990 103192 5510
rect 103428 3528 103480 3534
rect 103428 3470 103480 3476
rect 102968 2984 103020 2990
rect 102968 2926 103020 2932
rect 103152 2984 103204 2990
rect 103152 2926 103204 2932
rect 102784 1896 102836 1902
rect 102784 1838 102836 1844
rect 102980 800 103008 2926
rect 103440 800 103468 3470
rect 103532 2514 103560 8570
rect 103900 8004 103928 10200
rect 104076 9276 104132 9296
rect 104076 9200 104132 9220
rect 104076 8188 104132 8208
rect 104076 8112 104132 8132
rect 103900 7976 104020 8004
rect 103886 7848 103942 7857
rect 103886 7783 103888 7792
rect 103940 7783 103942 7792
rect 103888 7754 103940 7760
rect 103612 7336 103664 7342
rect 103612 7278 103664 7284
rect 103624 4758 103652 7278
rect 103888 6248 103940 6254
rect 103888 6190 103940 6196
rect 103900 5914 103928 6190
rect 103888 5908 103940 5914
rect 103888 5850 103940 5856
rect 103888 5772 103940 5778
rect 103992 5760 104020 7976
rect 104072 7948 104124 7954
rect 104072 7890 104124 7896
rect 104084 7410 104112 7890
rect 104072 7404 104124 7410
rect 104072 7346 104124 7352
rect 104076 7100 104132 7120
rect 104076 7024 104132 7044
rect 104076 6012 104132 6032
rect 104076 5936 104132 5956
rect 104164 5840 104216 5846
rect 104164 5782 104216 5788
rect 104072 5772 104124 5778
rect 103992 5732 104072 5760
rect 103888 5714 103940 5720
rect 104072 5714 104124 5720
rect 103900 5658 103928 5714
rect 104176 5658 104204 5782
rect 103900 5630 104204 5658
rect 104268 5642 104296 10200
rect 104440 9988 104492 9994
rect 104440 9930 104492 9936
rect 104452 6798 104480 9930
rect 104622 8936 104678 8945
rect 104622 8871 104678 8880
rect 104532 8424 104584 8430
rect 104532 8366 104584 8372
rect 104440 6792 104492 6798
rect 104440 6734 104492 6740
rect 104346 5808 104402 5817
rect 104346 5743 104348 5752
rect 104400 5743 104402 5752
rect 104348 5714 104400 5720
rect 104256 5636 104308 5642
rect 104256 5578 104308 5584
rect 104076 4924 104132 4944
rect 104076 4848 104132 4868
rect 103612 4752 103664 4758
rect 103612 4694 103664 4700
rect 104164 4616 104216 4622
rect 104164 4558 104216 4564
rect 104176 4486 104204 4558
rect 104164 4480 104216 4486
rect 104164 4422 104216 4428
rect 104348 4480 104400 4486
rect 104348 4422 104400 4428
rect 104076 3836 104132 3856
rect 104076 3760 104132 3780
rect 104164 3460 104216 3466
rect 104164 3402 104216 3408
rect 104176 3194 104204 3402
rect 104164 3188 104216 3194
rect 104164 3130 104216 3136
rect 104256 3120 104308 3126
rect 104256 3062 104308 3068
rect 103888 2848 103940 2854
rect 103888 2790 103940 2796
rect 103520 2508 103572 2514
rect 103520 2450 103572 2456
rect 103900 800 103928 2790
rect 104076 2748 104132 2768
rect 104076 2672 104132 2692
rect 104268 2582 104296 3062
rect 104256 2576 104308 2582
rect 104256 2518 104308 2524
rect 104360 2446 104388 4422
rect 104544 3194 104572 8366
rect 104532 3188 104584 3194
rect 104532 3130 104584 3136
rect 104636 2689 104664 8871
rect 104728 6322 104756 10200
rect 104808 7744 104860 7750
rect 104808 7686 104860 7692
rect 104820 7206 104848 7686
rect 104808 7200 104860 7206
rect 104808 7142 104860 7148
rect 105084 6792 105136 6798
rect 105084 6734 105136 6740
rect 104716 6316 104768 6322
rect 104716 6258 104768 6264
rect 105096 5914 105124 6734
rect 105188 6338 105216 10200
rect 105648 10062 105676 10200
rect 105636 10056 105688 10062
rect 105636 9998 105688 10004
rect 105636 9444 105688 9450
rect 105636 9386 105688 9392
rect 105648 9178 105676 9386
rect 105636 9172 105688 9178
rect 105636 9114 105688 9120
rect 105728 9172 105780 9178
rect 105728 9114 105780 9120
rect 105268 8560 105320 8566
rect 105268 8502 105320 8508
rect 105280 8129 105308 8502
rect 105740 8430 105768 9114
rect 105728 8424 105780 8430
rect 105728 8366 105780 8372
rect 105266 8120 105322 8129
rect 105266 8055 105322 8064
rect 105360 7948 105412 7954
rect 105360 7890 105412 7896
rect 105372 7721 105400 7890
rect 105358 7712 105414 7721
rect 105358 7647 105414 7656
rect 106016 7478 106044 10200
rect 106096 10056 106148 10062
rect 106096 9998 106148 10004
rect 106108 8430 106136 9998
rect 106096 8424 106148 8430
rect 106096 8366 106148 8372
rect 106280 7812 106332 7818
rect 106280 7754 106332 7760
rect 106004 7472 106056 7478
rect 106004 7414 106056 7420
rect 105912 7336 105964 7342
rect 105912 7278 105964 7284
rect 105636 6996 105688 7002
rect 105636 6938 105688 6944
rect 105188 6310 105584 6338
rect 105556 6254 105584 6310
rect 105360 6248 105412 6254
rect 105360 6190 105412 6196
rect 105544 6248 105596 6254
rect 105544 6190 105596 6196
rect 105372 5914 105400 6190
rect 105648 6100 105676 6938
rect 105924 6934 105952 7278
rect 105912 6928 105964 6934
rect 106292 6882 106320 7754
rect 106372 7336 106424 7342
rect 106372 7278 106424 7284
rect 105912 6870 105964 6876
rect 106108 6854 106320 6882
rect 106108 6730 106136 6854
rect 106280 6792 106332 6798
rect 106280 6734 106332 6740
rect 106096 6724 106148 6730
rect 106096 6666 106148 6672
rect 106292 6322 106320 6734
rect 106280 6316 106332 6322
rect 106280 6258 106332 6264
rect 105556 6072 105676 6100
rect 105084 5908 105136 5914
rect 105084 5850 105136 5856
rect 105360 5908 105412 5914
rect 105360 5850 105412 5856
rect 105174 5400 105230 5409
rect 105174 5335 105230 5344
rect 105188 5166 105216 5335
rect 105452 5228 105504 5234
rect 105452 5170 105504 5176
rect 105084 5160 105136 5166
rect 105082 5128 105084 5137
rect 105176 5160 105228 5166
rect 105136 5128 105138 5137
rect 105176 5102 105228 5108
rect 105082 5063 105138 5072
rect 104900 4684 104952 4690
rect 104900 4626 104952 4632
rect 105360 4684 105412 4690
rect 105360 4626 105412 4632
rect 104912 3738 104940 4626
rect 105372 4321 105400 4626
rect 105358 4312 105414 4321
rect 105358 4247 105414 4256
rect 105464 4185 105492 5170
rect 105450 4176 105506 4185
rect 105556 4146 105584 6072
rect 106384 5794 106412 7278
rect 106476 7274 106504 10200
rect 106936 9110 106964 10200
rect 106924 9104 106976 9110
rect 106924 9046 106976 9052
rect 107292 8832 107344 8838
rect 107292 8774 107344 8780
rect 106740 7880 106792 7886
rect 106740 7822 106792 7828
rect 106464 7268 106516 7274
rect 106464 7210 106516 7216
rect 106556 6928 106608 6934
rect 106556 6870 106608 6876
rect 106568 6390 106596 6870
rect 106648 6724 106700 6730
rect 106648 6666 106700 6672
rect 106556 6384 106608 6390
rect 106556 6326 106608 6332
rect 106660 6118 106688 6666
rect 106556 6112 106608 6118
rect 106556 6054 106608 6060
rect 106648 6112 106700 6118
rect 106648 6054 106700 6060
rect 106384 5766 106504 5794
rect 106372 5704 106424 5710
rect 106372 5646 106424 5652
rect 105636 5636 105688 5642
rect 105636 5578 105688 5584
rect 105648 4690 105676 5578
rect 106384 5234 106412 5646
rect 106372 5228 106424 5234
rect 106372 5170 106424 5176
rect 106280 5160 106332 5166
rect 106280 5102 106332 5108
rect 106292 4865 106320 5102
rect 106372 5024 106424 5030
rect 106370 4992 106372 5001
rect 106424 4992 106426 5001
rect 106370 4927 106426 4936
rect 106278 4856 106334 4865
rect 106108 4826 106228 4842
rect 106096 4820 106240 4826
rect 106148 4814 106188 4820
rect 106096 4762 106148 4768
rect 106278 4791 106334 4800
rect 106188 4762 106240 4768
rect 105636 4684 105688 4690
rect 105636 4626 105688 4632
rect 106188 4684 106240 4690
rect 106188 4626 106240 4632
rect 106200 4554 106228 4626
rect 106188 4548 106240 4554
rect 106188 4490 106240 4496
rect 106004 4480 106056 4486
rect 105924 4440 106004 4468
rect 105924 4321 105952 4440
rect 106004 4422 106056 4428
rect 105910 4312 105966 4321
rect 105910 4247 105966 4256
rect 105450 4111 105506 4120
rect 105544 4140 105596 4146
rect 105728 4140 105780 4146
rect 105544 4082 105596 4088
rect 105648 4100 105728 4128
rect 104900 3732 104952 3738
rect 104900 3674 104952 3680
rect 105176 3664 105228 3670
rect 105176 3606 105228 3612
rect 104622 2680 104678 2689
rect 104622 2615 104678 2624
rect 104348 2440 104400 2446
rect 104348 2382 104400 2388
rect 104256 1828 104308 1834
rect 104256 1770 104308 1776
rect 104076 1660 104132 1680
rect 104076 1584 104132 1604
rect 104268 800 104296 1770
rect 104532 1760 104584 1766
rect 104532 1702 104584 1708
rect 104624 1760 104676 1766
rect 104624 1702 104676 1708
rect 104544 1358 104572 1702
rect 104636 1562 104664 1702
rect 104624 1556 104676 1562
rect 104624 1498 104676 1504
rect 104716 1488 104768 1494
rect 104716 1430 104768 1436
rect 104532 1352 104584 1358
rect 104532 1294 104584 1300
rect 104728 800 104756 1430
rect 105188 800 105216 3606
rect 105544 2576 105596 2582
rect 105544 2518 105596 2524
rect 105450 2136 105506 2145
rect 105268 2100 105320 2106
rect 105450 2071 105506 2080
rect 105268 2042 105320 2048
rect 105280 1902 105308 2042
rect 105464 2038 105492 2071
rect 105452 2032 105504 2038
rect 105452 1974 105504 1980
rect 105268 1896 105320 1902
rect 105268 1838 105320 1844
rect 105556 1426 105584 2518
rect 105544 1420 105596 1426
rect 105544 1362 105596 1368
rect 105648 800 105676 4100
rect 105728 4082 105780 4088
rect 106004 3528 106056 3534
rect 105818 3496 105874 3505
rect 106004 3470 106056 3476
rect 105818 3431 105874 3440
rect 105728 3392 105780 3398
rect 105728 3334 105780 3340
rect 105740 1562 105768 3334
rect 105728 1556 105780 1562
rect 105728 1498 105780 1504
rect 105832 1426 105860 3431
rect 105820 1420 105872 1426
rect 105820 1362 105872 1368
rect 106016 800 106044 3470
rect 106476 2514 106504 5766
rect 106568 5234 106596 6054
rect 106752 5760 106780 7822
rect 106832 6724 106884 6730
rect 106832 6666 106884 6672
rect 106844 6458 106872 6666
rect 106832 6452 106884 6458
rect 106832 6394 106884 6400
rect 106752 5732 106872 5760
rect 106740 5636 106792 5642
rect 106740 5578 106792 5584
rect 106646 5400 106702 5409
rect 106646 5335 106702 5344
rect 106556 5228 106608 5234
rect 106556 5170 106608 5176
rect 106556 5024 106608 5030
rect 106660 5001 106688 5335
rect 106556 4966 106608 4972
rect 106646 4992 106702 5001
rect 106568 4758 106596 4966
rect 106646 4927 106702 4936
rect 106646 4856 106702 4865
rect 106646 4791 106702 4800
rect 106556 4752 106608 4758
rect 106556 4694 106608 4700
rect 106556 4548 106608 4554
rect 106556 4490 106608 4496
rect 106568 4457 106596 4490
rect 106554 4448 106610 4457
rect 106554 4383 106610 4392
rect 106660 3505 106688 4791
rect 106752 4078 106780 5578
rect 106740 4072 106792 4078
rect 106740 4014 106792 4020
rect 106646 3496 106702 3505
rect 106646 3431 106702 3440
rect 106556 3392 106608 3398
rect 106556 3334 106608 3340
rect 106464 2508 106516 2514
rect 106464 2450 106516 2456
rect 106568 1442 106596 3334
rect 106646 2272 106702 2281
rect 106646 2207 106702 2216
rect 106660 1970 106688 2207
rect 106648 1964 106700 1970
rect 106648 1906 106700 1912
rect 106740 1828 106792 1834
rect 106740 1770 106792 1776
rect 106476 1414 106596 1442
rect 106476 800 106504 1414
rect 106752 882 106780 1770
rect 106844 1426 106872 5732
rect 107014 5128 107070 5137
rect 107014 5063 107070 5072
rect 106922 4992 106978 5001
rect 106922 4927 106978 4936
rect 106936 2990 106964 4927
rect 106924 2984 106976 2990
rect 106924 2926 106976 2932
rect 106924 2848 106976 2854
rect 107028 2825 107056 5063
rect 107304 3602 107332 8774
rect 107396 8106 107424 10200
rect 107396 8078 107700 8106
rect 107566 7984 107622 7993
rect 107672 7954 107700 8078
rect 107764 8022 107792 10200
rect 107936 9920 107988 9926
rect 107936 9862 107988 9868
rect 107948 9042 107976 9862
rect 108224 9586 108252 10200
rect 108212 9580 108264 9586
rect 108212 9522 108264 9528
rect 107936 9036 107988 9042
rect 107936 8978 107988 8984
rect 108302 8392 108358 8401
rect 108302 8327 108358 8336
rect 107752 8016 107804 8022
rect 107752 7958 107804 7964
rect 107566 7919 107568 7928
rect 107620 7919 107622 7928
rect 107660 7948 107712 7954
rect 107568 7890 107620 7896
rect 107660 7890 107712 7896
rect 107752 7880 107804 7886
rect 107752 7822 107804 7828
rect 107474 7168 107530 7177
rect 107474 7103 107530 7112
rect 107488 5778 107516 7103
rect 107568 6112 107620 6118
rect 107568 6054 107620 6060
rect 107660 6112 107712 6118
rect 107660 6054 107712 6060
rect 107476 5772 107528 5778
rect 107476 5714 107528 5720
rect 107580 4865 107608 6054
rect 107672 5710 107700 6054
rect 107660 5704 107712 5710
rect 107660 5646 107712 5652
rect 107566 4856 107622 4865
rect 107566 4791 107622 4800
rect 107660 4276 107712 4282
rect 107660 4218 107712 4224
rect 107672 3913 107700 4218
rect 107764 4078 107792 7822
rect 107844 7472 107896 7478
rect 107844 7414 107896 7420
rect 108028 7472 108080 7478
rect 108028 7414 108080 7420
rect 107752 4072 107804 4078
rect 107752 4014 107804 4020
rect 107658 3904 107714 3913
rect 107658 3839 107714 3848
rect 107292 3596 107344 3602
rect 107292 3538 107344 3544
rect 107108 3392 107160 3398
rect 107108 3334 107160 3340
rect 107120 2922 107148 3334
rect 107108 2916 107160 2922
rect 107108 2858 107160 2864
rect 106924 2790 106976 2796
rect 107014 2816 107070 2825
rect 106832 1420 106884 1426
rect 106832 1362 106884 1368
rect 106740 876 106792 882
rect 106740 818 106792 824
rect 106936 800 106964 2790
rect 107014 2751 107070 2760
rect 107292 2304 107344 2310
rect 107292 2246 107344 2252
rect 107384 2304 107436 2310
rect 107384 2246 107436 2252
rect 107304 1737 107332 2246
rect 107290 1728 107346 1737
rect 107290 1663 107346 1672
rect 107396 800 107424 2246
rect 107752 1964 107804 1970
rect 107752 1906 107804 1912
rect 107764 800 107792 1906
rect 107856 1902 107884 7414
rect 108040 7002 108068 7414
rect 108120 7336 108172 7342
rect 108120 7278 108172 7284
rect 108028 6996 108080 7002
rect 108028 6938 108080 6944
rect 108132 6905 108160 7278
rect 108118 6896 108174 6905
rect 108118 6831 108174 6840
rect 108028 6248 108080 6254
rect 108028 6190 108080 6196
rect 108212 6248 108264 6254
rect 108212 6190 108264 6196
rect 107936 5772 107988 5778
rect 107936 5714 107988 5720
rect 107948 5642 107976 5714
rect 107936 5636 107988 5642
rect 107936 5578 107988 5584
rect 108040 4842 108068 6190
rect 108120 5160 108172 5166
rect 108118 5128 108120 5137
rect 108172 5128 108174 5137
rect 108118 5063 108174 5072
rect 108040 4814 108160 4842
rect 108028 4752 108080 4758
rect 107934 4720 107990 4729
rect 108028 4694 108080 4700
rect 107934 4655 107990 4664
rect 107948 4622 107976 4655
rect 107936 4616 107988 4622
rect 107936 4558 107988 4564
rect 108040 4486 108068 4694
rect 108028 4480 108080 4486
rect 108028 4422 108080 4428
rect 108132 3126 108160 4814
rect 108224 3670 108252 6190
rect 108316 4214 108344 8327
rect 108396 6452 108448 6458
rect 108396 6394 108448 6400
rect 108408 6254 108436 6394
rect 108684 6390 108712 10200
rect 108856 8628 108908 8634
rect 108856 8570 108908 8576
rect 108764 8492 108816 8498
rect 108764 8434 108816 8440
rect 108776 6497 108804 8434
rect 108868 6798 108896 8570
rect 109144 8566 109172 10200
rect 109224 8968 109276 8974
rect 109224 8910 109276 8916
rect 109132 8560 109184 8566
rect 109132 8502 109184 8508
rect 109236 8498 109264 8910
rect 109224 8492 109276 8498
rect 109224 8434 109276 8440
rect 109224 7948 109276 7954
rect 109224 7890 109276 7896
rect 109040 7744 109092 7750
rect 109040 7686 109092 7692
rect 108856 6792 108908 6798
rect 108856 6734 108908 6740
rect 108762 6488 108818 6497
rect 108762 6423 108818 6432
rect 108580 6384 108632 6390
rect 108580 6326 108632 6332
rect 108672 6384 108724 6390
rect 108672 6326 108724 6332
rect 108396 6248 108448 6254
rect 108396 6190 108448 6196
rect 108394 5672 108450 5681
rect 108394 5607 108450 5616
rect 108408 5574 108436 5607
rect 108396 5568 108448 5574
rect 108396 5510 108448 5516
rect 108488 5568 108540 5574
rect 108488 5510 108540 5516
rect 108396 5160 108448 5166
rect 108396 5102 108448 5108
rect 108408 5001 108436 5102
rect 108394 4992 108450 5001
rect 108394 4927 108450 4936
rect 108304 4208 108356 4214
rect 108304 4150 108356 4156
rect 108212 3664 108264 3670
rect 108212 3606 108264 3612
rect 108120 3120 108172 3126
rect 108120 3062 108172 3068
rect 108028 3052 108080 3058
rect 108028 2994 108080 3000
rect 107844 1896 107896 1902
rect 107844 1838 107896 1844
rect 108040 950 108068 2994
rect 108304 2916 108356 2922
rect 108304 2858 108356 2864
rect 108120 2032 108172 2038
rect 108120 1974 108172 1980
rect 108132 1018 108160 1974
rect 108212 1828 108264 1834
rect 108212 1770 108264 1776
rect 108120 1012 108172 1018
rect 108120 954 108172 960
rect 108028 944 108080 950
rect 108028 886 108080 892
rect 108224 800 108252 1770
rect 108316 1290 108344 2858
rect 108394 2136 108450 2145
rect 108394 2071 108396 2080
rect 108448 2071 108450 2080
rect 108396 2042 108448 2048
rect 108500 1902 108528 5510
rect 108488 1896 108540 1902
rect 108488 1838 108540 1844
rect 108304 1284 108356 1290
rect 108304 1226 108356 1232
rect 108592 1222 108620 6326
rect 108948 5908 109000 5914
rect 108948 5850 109000 5856
rect 108762 5808 108818 5817
rect 108762 5743 108764 5752
rect 108816 5743 108818 5752
rect 108764 5714 108816 5720
rect 108960 5710 108988 5850
rect 108948 5704 109000 5710
rect 108948 5646 109000 5652
rect 108856 4616 108908 4622
rect 108856 4558 108908 4564
rect 108868 2446 108896 4558
rect 109052 3602 109080 7686
rect 109130 6488 109186 6497
rect 109130 6423 109186 6432
rect 109144 5914 109172 6423
rect 109236 5953 109264 7890
rect 109408 7404 109460 7410
rect 109408 7346 109460 7352
rect 109420 7206 109448 7346
rect 109316 7200 109368 7206
rect 109316 7142 109368 7148
rect 109408 7200 109460 7206
rect 109408 7142 109460 7148
rect 109222 5944 109278 5953
rect 109132 5908 109184 5914
rect 109222 5879 109278 5888
rect 109132 5850 109184 5856
rect 109328 4554 109356 7142
rect 109512 6798 109540 10200
rect 109972 8650 110000 10200
rect 110328 9648 110380 9654
rect 110328 9590 110380 9596
rect 109880 8622 110000 8650
rect 109684 8356 109736 8362
rect 109684 8298 109736 8304
rect 109696 7410 109724 8298
rect 109684 7404 109736 7410
rect 109684 7346 109736 7352
rect 109880 7342 109908 8622
rect 109960 8492 110012 8498
rect 109960 8434 110012 8440
rect 109868 7336 109920 7342
rect 109868 7278 109920 7284
rect 109590 7032 109646 7041
rect 109590 6967 109646 6976
rect 109500 6792 109552 6798
rect 109500 6734 109552 6740
rect 109604 6254 109632 6967
rect 109868 6316 109920 6322
rect 109868 6258 109920 6264
rect 109592 6248 109644 6254
rect 109592 6190 109644 6196
rect 109776 6248 109828 6254
rect 109776 6190 109828 6196
rect 109590 6080 109646 6089
rect 109590 6015 109646 6024
rect 109604 5846 109632 6015
rect 109592 5840 109644 5846
rect 109592 5782 109644 5788
rect 109316 4548 109368 4554
rect 109316 4490 109368 4496
rect 109132 4480 109184 4486
rect 109132 4422 109184 4428
rect 109144 4214 109172 4422
rect 109684 4276 109736 4282
rect 109684 4218 109736 4224
rect 109132 4208 109184 4214
rect 109696 4185 109724 4218
rect 109132 4150 109184 4156
rect 109682 4176 109738 4185
rect 109682 4111 109738 4120
rect 109590 4040 109646 4049
rect 109590 3975 109646 3984
rect 109604 3777 109632 3975
rect 109590 3768 109646 3777
rect 109590 3703 109646 3712
rect 109040 3596 109092 3602
rect 109040 3538 109092 3544
rect 109224 3460 109276 3466
rect 109224 3402 109276 3408
rect 109236 3233 109264 3402
rect 109222 3224 109278 3233
rect 109132 3188 109184 3194
rect 109222 3159 109278 3168
rect 109132 3130 109184 3136
rect 108672 2440 108724 2446
rect 108672 2382 108724 2388
rect 108856 2440 108908 2446
rect 108856 2382 108908 2388
rect 108580 1216 108632 1222
rect 108580 1158 108632 1164
rect 108684 800 108712 2382
rect 109040 2372 109092 2378
rect 109040 2314 109092 2320
rect 109052 2281 109080 2314
rect 108762 2272 108818 2281
rect 108762 2207 108818 2216
rect 109038 2272 109094 2281
rect 109038 2207 109094 2216
rect 108776 2106 108804 2207
rect 108764 2100 108816 2106
rect 108948 2100 109000 2106
rect 108764 2042 108816 2048
rect 108868 2060 108948 2088
rect 108868 1850 108896 2060
rect 108948 2042 109000 2048
rect 108776 1822 108896 1850
rect 108776 1766 108804 1822
rect 108764 1760 108816 1766
rect 108764 1702 108816 1708
rect 109038 1592 109094 1601
rect 109038 1527 109040 1536
rect 109092 1527 109094 1536
rect 109040 1498 109092 1504
rect 109144 800 109172 3130
rect 109788 2990 109816 6190
rect 109880 5846 109908 6258
rect 109868 5840 109920 5846
rect 109868 5782 109920 5788
rect 109868 5704 109920 5710
rect 109868 5646 109920 5652
rect 109880 3534 109908 5646
rect 109868 3528 109920 3534
rect 109868 3470 109920 3476
rect 109224 2984 109276 2990
rect 109776 2984 109828 2990
rect 109276 2932 109540 2938
rect 109224 2926 109540 2932
rect 109776 2926 109828 2932
rect 109236 2910 109540 2926
rect 109512 2854 109540 2910
rect 109500 2848 109552 2854
rect 109500 2790 109552 2796
rect 109500 2576 109552 2582
rect 109500 2518 109552 2524
rect 109224 2440 109276 2446
rect 109224 2382 109276 2388
rect 109236 2145 109264 2382
rect 109316 2304 109368 2310
rect 109316 2246 109368 2252
rect 109222 2136 109278 2145
rect 109328 2106 109356 2246
rect 109512 2145 109540 2518
rect 109498 2136 109554 2145
rect 109222 2071 109278 2080
rect 109316 2100 109368 2106
rect 109316 2042 109368 2048
rect 109408 2100 109460 2106
rect 109498 2071 109554 2080
rect 109408 2042 109460 2048
rect 109420 1426 109448 2042
rect 109972 1986 110000 8434
rect 110144 8424 110196 8430
rect 110144 8366 110196 8372
rect 110052 6384 110104 6390
rect 110052 6326 110104 6332
rect 110064 2446 110092 6326
rect 110052 2440 110104 2446
rect 110052 2382 110104 2388
rect 109972 1958 110092 1986
rect 109960 1896 110012 1902
rect 109960 1838 110012 1844
rect 109682 1728 109738 1737
rect 109682 1663 109738 1672
rect 109696 1562 109724 1663
rect 109774 1592 109830 1601
rect 109500 1556 109552 1562
rect 109500 1498 109552 1504
rect 109684 1556 109736 1562
rect 109774 1527 109776 1536
rect 109684 1498 109736 1504
rect 109828 1527 109830 1536
rect 109776 1498 109828 1504
rect 109408 1420 109460 1426
rect 109408 1362 109460 1368
rect 109512 800 109540 1498
rect 109972 800 110000 1838
rect 98366 232 98422 241
rect 98366 167 98422 176
rect 98642 -400 98698 800
rect 99102 -400 99158 800
rect 99470 -400 99526 800
rect 99930 -400 99986 800
rect 100390 -400 100446 800
rect 100850 -400 100906 800
rect 101218 -400 101274 800
rect 101678 -400 101734 800
rect 102138 -400 102194 800
rect 102598 -400 102654 800
rect 102966 -400 103022 800
rect 103426 -400 103482 800
rect 103886 -400 103942 800
rect 104254 -400 104310 800
rect 104714 -400 104770 800
rect 105174 -400 105230 800
rect 105634 -400 105690 800
rect 106002 -400 106058 800
rect 106462 -400 106518 800
rect 106922 -400 106978 800
rect 107382 -400 107438 800
rect 107750 -400 107806 800
rect 108210 -400 108266 800
rect 108670 -400 108726 800
rect 109130 -400 109186 800
rect 109498 -400 109554 800
rect 109958 -400 110014 800
rect 110064 785 110092 1958
rect 110156 1601 110184 8366
rect 110236 5636 110288 5642
rect 110236 5578 110288 5584
rect 110248 5166 110276 5578
rect 110236 5160 110288 5166
rect 110236 5102 110288 5108
rect 110340 4049 110368 9590
rect 110432 9466 110460 10200
rect 110432 9438 110552 9466
rect 110420 9376 110472 9382
rect 110420 9318 110472 9324
rect 110432 7954 110460 9318
rect 110420 7948 110472 7954
rect 110420 7890 110472 7896
rect 110524 7274 110552 9438
rect 110788 9172 110840 9178
rect 110788 9114 110840 9120
rect 110800 7750 110828 9114
rect 110788 7744 110840 7750
rect 110788 7686 110840 7692
rect 110512 7268 110564 7274
rect 110512 7210 110564 7216
rect 110604 6656 110656 6662
rect 110604 6598 110656 6604
rect 110788 6656 110840 6662
rect 110788 6598 110840 6604
rect 110616 6458 110644 6598
rect 110604 6452 110656 6458
rect 110604 6394 110656 6400
rect 110696 5704 110748 5710
rect 110696 5646 110748 5652
rect 110420 5160 110472 5166
rect 110420 5102 110472 5108
rect 110604 5160 110656 5166
rect 110604 5102 110656 5108
rect 110432 5001 110460 5102
rect 110418 4992 110474 5001
rect 110418 4927 110474 4936
rect 110510 4856 110566 4865
rect 110510 4791 110566 4800
rect 110418 4448 110474 4457
rect 110418 4383 110474 4392
rect 110432 4078 110460 4383
rect 110420 4072 110472 4078
rect 110326 4040 110382 4049
rect 110420 4014 110472 4020
rect 110326 3975 110382 3984
rect 110524 3738 110552 4791
rect 110512 3732 110564 3738
rect 110512 3674 110564 3680
rect 110510 2816 110566 2825
rect 110510 2751 110566 2760
rect 110524 2650 110552 2751
rect 110420 2644 110472 2650
rect 110420 2586 110472 2592
rect 110512 2644 110564 2650
rect 110512 2586 110564 2592
rect 110432 2530 110460 2586
rect 110432 2502 110552 2530
rect 110616 2514 110644 5102
rect 110708 4146 110736 5646
rect 110696 4140 110748 4146
rect 110696 4082 110748 4088
rect 110420 2304 110472 2310
rect 110420 2246 110472 2252
rect 110432 1834 110460 2246
rect 110420 1828 110472 1834
rect 110420 1770 110472 1776
rect 110524 1714 110552 2502
rect 110604 2508 110656 2514
rect 110604 2450 110656 2456
rect 110800 1902 110828 6598
rect 110892 5642 110920 10200
rect 111260 9738 111288 10200
rect 111720 9738 111748 10200
rect 110984 9710 111288 9738
rect 111628 9710 111748 9738
rect 110984 8090 111012 9710
rect 111248 9580 111300 9586
rect 111248 9522 111300 9528
rect 111260 9042 111288 9522
rect 111524 9512 111576 9518
rect 111524 9454 111576 9460
rect 111248 9036 111300 9042
rect 111248 8978 111300 8984
rect 111156 8832 111208 8838
rect 111156 8774 111208 8780
rect 110972 8084 111024 8090
rect 110972 8026 111024 8032
rect 111064 8084 111116 8090
rect 111064 8026 111116 8032
rect 111076 7478 111104 8026
rect 111064 7472 111116 7478
rect 111064 7414 111116 7420
rect 111064 6860 111116 6866
rect 111064 6802 111116 6808
rect 110880 5636 110932 5642
rect 110880 5578 110932 5584
rect 110880 5092 110932 5098
rect 110880 5034 110932 5040
rect 110892 4865 110920 5034
rect 110878 4856 110934 4865
rect 110878 4791 110934 4800
rect 111076 4185 111104 6802
rect 111062 4176 111118 4185
rect 111062 4111 111118 4120
rect 111062 3904 111118 3913
rect 111062 3839 111118 3848
rect 111076 3194 111104 3839
rect 111064 3188 111116 3194
rect 111064 3130 111116 3136
rect 111168 2938 111196 8774
rect 111340 7200 111392 7206
rect 111340 7142 111392 7148
rect 111248 6384 111300 6390
rect 111248 6326 111300 6332
rect 111260 6089 111288 6326
rect 111246 6080 111302 6089
rect 111246 6015 111302 6024
rect 111248 4820 111300 4826
rect 111248 4762 111300 4768
rect 111260 4457 111288 4762
rect 111246 4448 111302 4457
rect 111246 4383 111302 4392
rect 111168 2910 111288 2938
rect 111260 2854 111288 2910
rect 111248 2848 111300 2854
rect 111248 2790 111300 2796
rect 111352 2530 111380 7142
rect 111432 6248 111484 6254
rect 111432 6190 111484 6196
rect 111444 5642 111472 6190
rect 111432 5636 111484 5642
rect 111432 5578 111484 5584
rect 111432 5160 111484 5166
rect 111432 5102 111484 5108
rect 111444 4826 111472 5102
rect 111432 4820 111484 4826
rect 111432 4762 111484 4768
rect 111432 3120 111484 3126
rect 111432 3062 111484 3068
rect 111444 2854 111472 3062
rect 111432 2848 111484 2854
rect 111432 2790 111484 2796
rect 111352 2502 111472 2530
rect 111444 2378 111472 2502
rect 111432 2372 111484 2378
rect 111432 2314 111484 2320
rect 111248 2304 111300 2310
rect 110970 2272 111026 2281
rect 111248 2246 111300 2252
rect 110970 2207 111026 2216
rect 110984 2038 111012 2207
rect 110880 2032 110932 2038
rect 110880 1974 110932 1980
rect 110972 2032 111024 2038
rect 110972 1974 111024 1980
rect 110788 1896 110840 1902
rect 110788 1838 110840 1844
rect 110432 1686 110552 1714
rect 110604 1760 110656 1766
rect 110604 1702 110656 1708
rect 110142 1592 110198 1601
rect 110142 1527 110198 1536
rect 110432 800 110460 1686
rect 110616 1426 110644 1702
rect 110694 1456 110750 1465
rect 110604 1420 110656 1426
rect 110694 1391 110696 1400
rect 110604 1362 110656 1368
rect 110748 1391 110750 1400
rect 110696 1362 110748 1368
rect 110892 800 110920 1974
rect 111260 800 111288 2246
rect 111536 2145 111564 9454
rect 111628 5778 111656 9710
rect 111708 9648 111760 9654
rect 111708 9590 111760 9596
rect 111720 8430 111748 9590
rect 111708 8424 111760 8430
rect 111708 8366 111760 8372
rect 111892 8424 111944 8430
rect 111892 8366 111944 8372
rect 111708 7336 111760 7342
rect 111708 7278 111760 7284
rect 111616 5772 111668 5778
rect 111616 5714 111668 5720
rect 111616 5636 111668 5642
rect 111616 5578 111668 5584
rect 111628 4729 111656 5578
rect 111614 4720 111670 4729
rect 111614 4655 111670 4664
rect 111720 3913 111748 7278
rect 111800 5228 111852 5234
rect 111800 5170 111852 5176
rect 111706 3904 111762 3913
rect 111706 3839 111762 3848
rect 111812 3670 111840 5170
rect 111800 3664 111852 3670
rect 111800 3606 111852 3612
rect 111904 2582 111932 8366
rect 112180 8362 112208 10200
rect 112168 8356 112220 8362
rect 112168 8298 112220 8304
rect 112076 7880 112128 7886
rect 112076 7822 112128 7828
rect 111984 7744 112036 7750
rect 111984 7686 112036 7692
rect 111892 2576 111944 2582
rect 111892 2518 111944 2524
rect 111522 2136 111578 2145
rect 111522 2071 111578 2080
rect 111708 1828 111760 1834
rect 111708 1770 111760 1776
rect 111720 800 111748 1770
rect 111996 1465 112024 7686
rect 112088 7410 112116 7822
rect 112168 7540 112220 7546
rect 112168 7482 112220 7488
rect 112076 7404 112128 7410
rect 112076 7346 112128 7352
rect 112074 3224 112130 3233
rect 112074 3159 112130 3168
rect 112088 3058 112116 3159
rect 112076 3052 112128 3058
rect 112076 2994 112128 3000
rect 112076 1896 112128 1902
rect 112074 1864 112076 1873
rect 112128 1864 112130 1873
rect 112074 1799 112130 1808
rect 111982 1456 112038 1465
rect 111982 1391 112038 1400
rect 112180 1290 112208 7482
rect 112260 6656 112312 6662
rect 112260 6598 112312 6604
rect 112272 5778 112300 6598
rect 112548 6254 112576 10200
rect 112812 8288 112864 8294
rect 112812 8230 112864 8236
rect 112536 6248 112588 6254
rect 112536 6190 112588 6196
rect 112260 5772 112312 5778
rect 112260 5714 112312 5720
rect 112444 4616 112496 4622
rect 112444 4558 112496 4564
rect 112260 4548 112312 4554
rect 112260 4490 112312 4496
rect 112272 1873 112300 4490
rect 112456 4146 112484 4558
rect 112444 4140 112496 4146
rect 112444 4082 112496 4088
rect 112824 3534 112852 8230
rect 113008 5098 113036 10200
rect 113468 8401 113496 10200
rect 113928 9738 113956 10200
rect 113744 9710 113956 9738
rect 113454 8392 113510 8401
rect 113454 8327 113510 8336
rect 113456 8288 113508 8294
rect 113456 8230 113508 8236
rect 113468 7410 113496 8230
rect 113456 7404 113508 7410
rect 113456 7346 113508 7352
rect 113548 6112 113600 6118
rect 113548 6054 113600 6060
rect 113088 5704 113140 5710
rect 113088 5646 113140 5652
rect 113100 5234 113128 5646
rect 113088 5228 113140 5234
rect 113088 5170 113140 5176
rect 112996 5092 113048 5098
rect 112996 5034 113048 5040
rect 113088 5092 113140 5098
rect 113088 5034 113140 5040
rect 113100 4690 113128 5034
rect 113088 4684 113140 4690
rect 113088 4626 113140 4632
rect 113560 4554 113588 6054
rect 113640 4684 113692 4690
rect 113640 4626 113692 4632
rect 113548 4548 113600 4554
rect 113548 4490 113600 4496
rect 113652 4457 113680 4626
rect 113638 4448 113694 4457
rect 113638 4383 113694 4392
rect 113454 4040 113510 4049
rect 113454 3975 113510 3984
rect 113468 3942 113496 3975
rect 113364 3936 113416 3942
rect 113364 3878 113416 3884
rect 113456 3936 113508 3942
rect 113456 3878 113508 3884
rect 113376 3534 113404 3878
rect 113744 3777 113772 9710
rect 113916 9580 113968 9586
rect 113916 9522 113968 9528
rect 113928 7410 113956 9522
rect 114192 7812 114244 7818
rect 114192 7754 114244 7760
rect 114006 7576 114062 7585
rect 114006 7511 114062 7520
rect 113916 7404 113968 7410
rect 113916 7346 113968 7352
rect 113824 5024 113876 5030
rect 113824 4966 113876 4972
rect 113836 4758 113864 4966
rect 113824 4752 113876 4758
rect 113824 4694 113876 4700
rect 113824 4480 113876 4486
rect 113916 4480 113968 4486
rect 113876 4440 113916 4468
rect 113824 4422 113876 4428
rect 113916 4422 113968 4428
rect 113730 3768 113786 3777
rect 113730 3703 113786 3712
rect 112812 3528 112864 3534
rect 112812 3470 112864 3476
rect 113364 3528 113416 3534
rect 113364 3470 113416 3476
rect 112442 3360 112498 3369
rect 112442 3295 112498 3304
rect 112352 2440 112404 2446
rect 112350 2408 112352 2417
rect 112404 2408 112406 2417
rect 112350 2343 112406 2352
rect 112258 1864 112314 1873
rect 112258 1799 112314 1808
rect 112456 1442 112484 3295
rect 113822 3088 113878 3097
rect 113822 3023 113824 3032
rect 113876 3023 113878 3032
rect 113824 2994 113876 3000
rect 113546 2952 113602 2961
rect 112996 2916 113048 2922
rect 113546 2887 113548 2896
rect 112996 2858 113048 2864
rect 113600 2887 113602 2896
rect 113548 2858 113600 2864
rect 112352 1420 112404 1426
rect 112456 1414 112576 1442
rect 112352 1362 112404 1368
rect 112168 1284 112220 1290
rect 112168 1226 112220 1232
rect 112168 1012 112220 1018
rect 112168 954 112220 960
rect 112180 800 112208 954
rect 112364 898 112392 1362
rect 112548 1358 112576 1414
rect 112536 1352 112588 1358
rect 112536 1294 112588 1300
rect 112364 870 112576 898
rect 112548 800 112576 870
rect 113008 800 113036 2858
rect 113824 2440 113876 2446
rect 113824 2382 113876 2388
rect 113364 2032 113416 2038
rect 113364 1974 113416 1980
rect 113546 2000 113602 2009
rect 113376 1850 113404 1974
rect 113836 1970 113864 2382
rect 114020 2106 114048 7511
rect 114204 6338 114232 7754
rect 114296 7177 114324 10200
rect 114652 9376 114704 9382
rect 114652 9318 114704 9324
rect 114664 8498 114692 9318
rect 114652 8492 114704 8498
rect 114652 8434 114704 8440
rect 114466 8120 114522 8129
rect 114466 8055 114522 8064
rect 114376 7404 114428 7410
rect 114376 7346 114428 7352
rect 114282 7168 114338 7177
rect 114282 7103 114338 7112
rect 114388 6474 114416 7346
rect 114480 6798 114508 8055
rect 114468 6792 114520 6798
rect 114756 6780 114784 10200
rect 115216 9602 115244 10200
rect 115032 9574 115244 9602
rect 114468 6734 114520 6740
rect 114572 6752 114784 6780
rect 114836 6792 114888 6798
rect 114466 6488 114522 6497
rect 114388 6446 114466 6474
rect 114466 6423 114522 6432
rect 114466 6352 114522 6361
rect 114204 6310 114466 6338
rect 114466 6287 114522 6296
rect 114572 5930 114600 6752
rect 114836 6734 114888 6740
rect 114848 6225 114876 6734
rect 114834 6216 114890 6225
rect 114834 6151 114890 6160
rect 114480 5902 114600 5930
rect 115032 5914 115060 9574
rect 115204 9512 115256 9518
rect 115204 9454 115256 9460
rect 115112 6860 115164 6866
rect 115112 6802 115164 6808
rect 115124 5914 115152 6802
rect 115020 5908 115072 5914
rect 114480 5846 114508 5902
rect 115020 5850 115072 5856
rect 115112 5908 115164 5914
rect 115112 5850 115164 5856
rect 114468 5840 114520 5846
rect 114468 5782 114520 5788
rect 114744 5704 114796 5710
rect 114742 5672 114744 5681
rect 114796 5672 114798 5681
rect 114742 5607 114798 5616
rect 115112 5160 115164 5166
rect 114940 5120 115112 5148
rect 114940 5114 114968 5120
rect 114848 5098 114968 5114
rect 115112 5102 115164 5108
rect 114836 5092 114968 5098
rect 114888 5086 114968 5092
rect 114836 5034 114888 5040
rect 114744 4616 114796 4622
rect 114744 4558 114796 4564
rect 114928 4616 114980 4622
rect 114928 4558 114980 4564
rect 114756 4486 114784 4558
rect 114744 4480 114796 4486
rect 114744 4422 114796 4428
rect 114940 4078 114968 4558
rect 114928 4072 114980 4078
rect 114928 4014 114980 4020
rect 115216 3738 115244 9454
rect 115296 7336 115348 7342
rect 115296 7278 115348 7284
rect 115308 3942 115336 7278
rect 115676 6866 115704 10200
rect 115848 7948 115900 7954
rect 115848 7890 115900 7896
rect 115664 6860 115716 6866
rect 115664 6802 115716 6808
rect 115756 6724 115808 6730
rect 115756 6666 115808 6672
rect 115296 3936 115348 3942
rect 115296 3878 115348 3884
rect 115386 3904 115442 3913
rect 115386 3839 115442 3848
rect 115400 3738 115428 3839
rect 115204 3732 115256 3738
rect 115204 3674 115256 3680
rect 115388 3732 115440 3738
rect 115388 3674 115440 3680
rect 114190 3496 114246 3505
rect 114190 3431 114246 3440
rect 114204 2650 114232 3431
rect 114192 2644 114244 2650
rect 114192 2586 114244 2592
rect 115204 2576 115256 2582
rect 115202 2544 115204 2553
rect 115256 2544 115258 2553
rect 115202 2479 115258 2488
rect 113916 2100 113968 2106
rect 113916 2042 113968 2048
rect 114008 2100 114060 2106
rect 114008 2042 114060 2048
rect 113546 1935 113548 1944
rect 113600 1935 113602 1944
rect 113824 1964 113876 1970
rect 113548 1906 113600 1912
rect 113824 1906 113876 1912
rect 113640 1896 113692 1902
rect 113376 1844 113640 1850
rect 113376 1838 113692 1844
rect 113376 1822 113680 1838
rect 113456 944 113508 950
rect 113456 886 113508 892
rect 113468 800 113496 886
rect 113928 800 113956 2042
rect 114468 1896 114520 1902
rect 115112 1896 115164 1902
rect 114520 1856 114784 1884
rect 114468 1838 114520 1844
rect 114284 1760 114336 1766
rect 114284 1702 114336 1708
rect 114376 1760 114428 1766
rect 114376 1702 114428 1708
rect 114296 800 114324 1702
rect 114388 1562 114416 1702
rect 114376 1556 114428 1562
rect 114376 1498 114428 1504
rect 114756 800 114784 1856
rect 115112 1838 115164 1844
rect 115204 1896 115256 1902
rect 115204 1838 115256 1844
rect 115124 882 115152 1838
rect 115112 876 115164 882
rect 115112 818 115164 824
rect 115216 800 115244 1838
rect 115768 1562 115796 6666
rect 115860 3233 115888 7890
rect 116044 6390 116072 10200
rect 116308 7880 116360 7886
rect 116308 7822 116360 7828
rect 116320 6866 116348 7822
rect 116308 6860 116360 6866
rect 116308 6802 116360 6808
rect 116032 6384 116084 6390
rect 116504 6372 116532 10200
rect 116584 9376 116636 9382
rect 116584 9318 116636 9324
rect 116596 7410 116624 9318
rect 116584 7404 116636 7410
rect 116584 7346 116636 7352
rect 116032 6326 116084 6332
rect 116136 6344 116532 6372
rect 116136 5710 116164 6344
rect 116400 6248 116452 6254
rect 116400 6190 116452 6196
rect 116124 5704 116176 5710
rect 116124 5646 116176 5652
rect 116308 5704 116360 5710
rect 116308 5646 116360 5652
rect 116320 5234 116348 5646
rect 116308 5228 116360 5234
rect 116308 5170 116360 5176
rect 115940 4140 115992 4146
rect 115992 4100 116164 4128
rect 115940 4082 115992 4088
rect 115940 4004 115992 4010
rect 115940 3946 115992 3952
rect 115952 3505 115980 3946
rect 115938 3496 115994 3505
rect 115938 3431 115994 3440
rect 115846 3224 115902 3233
rect 115846 3159 115902 3168
rect 116136 1766 116164 4100
rect 116412 3194 116440 6190
rect 116964 5409 116992 10200
rect 117228 8900 117280 8906
rect 117228 8842 117280 8848
rect 117240 8242 117268 8842
rect 117240 8214 117360 8242
rect 117044 5772 117096 5778
rect 117044 5714 117096 5720
rect 116950 5400 117006 5409
rect 116950 5335 117006 5344
rect 116952 4480 117004 4486
rect 116950 4448 116952 4457
rect 117004 4448 117006 4457
rect 116950 4383 117006 4392
rect 116676 4072 116728 4078
rect 116676 4014 116728 4020
rect 116584 3528 116636 3534
rect 116584 3470 116636 3476
rect 116492 3392 116544 3398
rect 116490 3360 116492 3369
rect 116544 3360 116546 3369
rect 116490 3295 116546 3304
rect 116596 3194 116624 3470
rect 116308 3188 116360 3194
rect 116308 3130 116360 3136
rect 116400 3188 116452 3194
rect 116400 3130 116452 3136
rect 116584 3188 116636 3194
rect 116584 3130 116636 3136
rect 116320 2854 116348 3130
rect 116688 2961 116716 4014
rect 116858 3904 116914 3913
rect 116858 3839 116914 3848
rect 116872 3602 116900 3839
rect 116860 3596 116912 3602
rect 116860 3538 116912 3544
rect 116674 2952 116730 2961
rect 116674 2887 116730 2896
rect 116860 2916 116912 2922
rect 116860 2858 116912 2864
rect 116308 2848 116360 2854
rect 116872 2825 116900 2858
rect 116952 2848 117004 2854
rect 116308 2790 116360 2796
rect 116858 2816 116914 2825
rect 116952 2790 117004 2796
rect 116858 2751 116914 2760
rect 116860 2508 116912 2514
rect 116860 2450 116912 2456
rect 116216 2304 116268 2310
rect 116308 2304 116360 2310
rect 116216 2246 116268 2252
rect 116306 2272 116308 2281
rect 116360 2272 116362 2281
rect 116228 2106 116256 2246
rect 116306 2207 116362 2216
rect 116216 2100 116268 2106
rect 116216 2042 116268 2048
rect 116032 1760 116084 1766
rect 116032 1702 116084 1708
rect 116124 1760 116176 1766
rect 116124 1702 116176 1708
rect 115756 1556 115808 1562
rect 115756 1498 115808 1504
rect 115296 1420 115348 1426
rect 115296 1362 115348 1368
rect 110050 776 110106 785
rect 110050 711 110106 720
rect 110418 -400 110474 800
rect 110878 -400 110934 800
rect 111246 -400 111302 800
rect 111706 -400 111762 800
rect 112166 -400 112222 800
rect 112534 -400 112590 800
rect 112994 -400 113050 800
rect 113454 -400 113510 800
rect 113914 -400 113970 800
rect 114282 -400 114338 800
rect 114742 -400 114798 800
rect 115202 -400 115258 800
rect 115308 610 115336 1362
rect 115664 944 115716 950
rect 115664 886 115716 892
rect 115676 800 115704 886
rect 116044 800 116072 1702
rect 116492 1352 116544 1358
rect 116492 1294 116544 1300
rect 116504 800 116532 1294
rect 116872 1193 116900 2450
rect 116858 1184 116914 1193
rect 116858 1119 116914 1128
rect 116964 800 116992 2790
rect 117056 1222 117084 5714
rect 117228 5160 117280 5166
rect 117228 5102 117280 5108
rect 117136 4616 117188 4622
rect 117136 4558 117188 4564
rect 117148 4146 117176 4558
rect 117136 4140 117188 4146
rect 117136 4082 117188 4088
rect 117240 3738 117268 5102
rect 117332 4434 117360 8214
rect 117424 4593 117452 10200
rect 117502 9208 117558 9217
rect 117502 9143 117558 9152
rect 117516 6186 117544 9143
rect 117792 6882 117820 10200
rect 118252 7750 118280 10200
rect 118424 8832 118476 8838
rect 118424 8774 118476 8780
rect 118240 7744 118292 7750
rect 118240 7686 118292 7692
rect 118056 7404 118108 7410
rect 118056 7346 118108 7352
rect 117608 6854 117820 6882
rect 117504 6180 117556 6186
rect 117504 6122 117556 6128
rect 117608 4865 117636 6854
rect 118068 6089 118096 7346
rect 118148 6792 118200 6798
rect 118148 6734 118200 6740
rect 118054 6080 118110 6089
rect 118054 6015 118110 6024
rect 117688 5636 117740 5642
rect 117688 5578 117740 5584
rect 117594 4856 117650 4865
rect 117594 4791 117650 4800
rect 117410 4584 117466 4593
rect 117410 4519 117466 4528
rect 117332 4406 117636 4434
rect 117228 3732 117280 3738
rect 117228 3674 117280 3680
rect 117318 3360 117374 3369
rect 117318 3295 117374 3304
rect 117502 3360 117558 3369
rect 117502 3295 117558 3304
rect 117332 2922 117360 3295
rect 117516 3126 117544 3295
rect 117504 3120 117556 3126
rect 117504 3062 117556 3068
rect 117320 2916 117372 2922
rect 117320 2858 117372 2864
rect 117136 2508 117188 2514
rect 117136 2450 117188 2456
rect 117148 2281 117176 2450
rect 117134 2272 117190 2281
rect 117134 2207 117190 2216
rect 117608 2106 117636 4406
rect 117596 2100 117648 2106
rect 117596 2042 117648 2048
rect 117136 1964 117188 1970
rect 117136 1906 117188 1912
rect 117148 1850 117176 1906
rect 117148 1822 117452 1850
rect 117044 1216 117096 1222
rect 117044 1158 117096 1164
rect 117424 800 117452 1822
rect 117700 1562 117728 5578
rect 118160 4842 118188 6734
rect 118332 6656 118384 6662
rect 118332 6598 118384 6604
rect 117792 4814 118188 4842
rect 117688 1556 117740 1562
rect 117688 1498 117740 1504
rect 117792 1018 117820 4814
rect 118344 4486 118372 6598
rect 118436 4690 118464 8774
rect 118712 8514 118740 10200
rect 118712 8486 118832 8514
rect 118700 8356 118752 8362
rect 118700 8298 118752 8304
rect 118712 7954 118740 8298
rect 118700 7948 118752 7954
rect 118700 7890 118752 7896
rect 118804 7313 118832 8486
rect 119068 7880 119120 7886
rect 119068 7822 119120 7828
rect 118790 7304 118846 7313
rect 118790 7239 118846 7248
rect 118606 7168 118662 7177
rect 118606 7103 118662 7112
rect 118620 6118 118648 7103
rect 118700 6792 118752 6798
rect 118700 6734 118752 6740
rect 118884 6792 118936 6798
rect 118884 6734 118936 6740
rect 118712 6322 118740 6734
rect 118700 6316 118752 6322
rect 118700 6258 118752 6264
rect 118896 6225 118924 6734
rect 119080 6322 119108 7822
rect 119068 6316 119120 6322
rect 119068 6258 119120 6264
rect 118882 6216 118938 6225
rect 118882 6151 118938 6160
rect 118608 6112 118660 6118
rect 118608 6054 118660 6060
rect 118514 5400 118570 5409
rect 118514 5335 118516 5344
rect 118568 5335 118570 5344
rect 118608 5364 118660 5370
rect 118516 5306 118568 5312
rect 118608 5306 118660 5312
rect 118620 5250 118648 5306
rect 118528 5234 118648 5250
rect 118516 5228 118648 5234
rect 118568 5222 118648 5228
rect 118516 5170 118568 5176
rect 118792 5092 118844 5098
rect 118792 5034 118844 5040
rect 118608 4820 118660 4826
rect 118608 4762 118660 4768
rect 118424 4684 118476 4690
rect 118424 4626 118476 4632
rect 118332 4480 118384 4486
rect 118332 4422 118384 4428
rect 118620 4282 118648 4762
rect 118516 4276 118568 4282
rect 118516 4218 118568 4224
rect 118608 4276 118660 4282
rect 118608 4218 118660 4224
rect 118148 4140 118200 4146
rect 118148 4082 118200 4088
rect 117964 3596 118016 3602
rect 117964 3538 118016 3544
rect 117976 3194 118004 3538
rect 118160 3398 118188 4082
rect 118528 4049 118556 4218
rect 118514 4040 118570 4049
rect 118514 3975 118570 3984
rect 118514 3768 118570 3777
rect 118514 3703 118570 3712
rect 118528 3534 118556 3703
rect 118516 3528 118568 3534
rect 118516 3470 118568 3476
rect 118148 3392 118200 3398
rect 118700 3392 118752 3398
rect 118148 3334 118200 3340
rect 118698 3360 118700 3369
rect 118752 3360 118754 3369
rect 118698 3295 118754 3304
rect 118330 3224 118386 3233
rect 117964 3188 118016 3194
rect 118330 3159 118386 3168
rect 117964 3130 118016 3136
rect 118344 3074 118372 3159
rect 118804 3126 118832 5034
rect 118884 4820 118936 4826
rect 118884 4762 118936 4768
rect 118896 4282 118924 4762
rect 118974 4448 119030 4457
rect 118974 4383 119030 4392
rect 118884 4276 118936 4282
rect 118884 4218 118936 4224
rect 118792 3120 118844 3126
rect 118344 3058 118648 3074
rect 118792 3062 118844 3068
rect 118344 3052 118660 3058
rect 118344 3046 118608 3052
rect 118608 2994 118660 3000
rect 118606 2952 118662 2961
rect 118606 2887 118662 2896
rect 118238 2680 118294 2689
rect 118238 2615 118240 2624
rect 118292 2615 118294 2624
rect 118240 2586 118292 2592
rect 117872 2508 117924 2514
rect 117872 2450 117924 2456
rect 118148 2508 118200 2514
rect 118148 2450 118200 2456
rect 117780 1012 117832 1018
rect 117780 954 117832 960
rect 117884 898 117912 2450
rect 118056 1896 118108 1902
rect 118056 1838 118108 1844
rect 118068 1426 118096 1838
rect 118056 1420 118108 1426
rect 118056 1362 118108 1368
rect 118160 1290 118188 2450
rect 118240 2304 118292 2310
rect 118240 2246 118292 2252
rect 118332 2304 118384 2310
rect 118332 2246 118384 2252
rect 118148 1284 118200 1290
rect 118148 1226 118200 1232
rect 117792 870 117912 898
rect 117792 800 117820 870
rect 118252 800 118280 2246
rect 118344 1970 118372 2246
rect 118620 2106 118648 2887
rect 118988 2650 119016 4383
rect 119172 4264 119200 10200
rect 119436 9580 119488 9586
rect 119436 9522 119488 9528
rect 119342 4856 119398 4865
rect 119342 4791 119398 4800
rect 119356 4622 119384 4791
rect 119344 4616 119396 4622
rect 119344 4558 119396 4564
rect 119448 4434 119476 9522
rect 119540 5370 119568 10200
rect 119620 9580 119672 9586
rect 119620 9522 119672 9528
rect 119632 6225 119660 9522
rect 119724 9042 119752 10202
rect 119816 9518 119844 10338
rect 119986 10200 120042 11400
rect 120446 10200 120502 11400
rect 120814 10200 120870 11400
rect 121274 10200 121330 11400
rect 121734 10200 121790 11400
rect 122194 10200 122250 11400
rect 122562 10200 122618 11400
rect 123022 10200 123078 11400
rect 123482 10200 123538 11400
rect 123942 10200 123998 11400
rect 124310 10200 124366 11400
rect 124404 10532 124456 10538
rect 124404 10474 124456 10480
rect 119804 9512 119856 9518
rect 119804 9454 119856 9460
rect 119712 9036 119764 9042
rect 119712 8978 119764 8984
rect 119712 8900 119764 8906
rect 119712 8842 119764 8848
rect 119618 6216 119674 6225
rect 119618 6151 119674 6160
rect 119618 5672 119674 5681
rect 119618 5607 119674 5616
rect 119632 5574 119660 5607
rect 119620 5568 119672 5574
rect 119620 5510 119672 5516
rect 119528 5364 119580 5370
rect 119528 5306 119580 5312
rect 119618 4584 119674 4593
rect 119618 4519 119620 4528
rect 119672 4519 119674 4528
rect 119620 4490 119672 4496
rect 119448 4406 119660 4434
rect 119080 4236 119200 4264
rect 119080 3641 119108 4236
rect 119344 4072 119396 4078
rect 119396 4020 119568 4026
rect 119344 4014 119568 4020
rect 119356 3998 119568 4014
rect 119540 3942 119568 3998
rect 119528 3936 119580 3942
rect 119632 3913 119660 4406
rect 119528 3878 119580 3884
rect 119618 3904 119674 3913
rect 119618 3839 119674 3848
rect 119250 3768 119306 3777
rect 119250 3703 119306 3712
rect 119066 3632 119122 3641
rect 119066 3567 119122 3576
rect 118976 2644 119028 2650
rect 118976 2586 119028 2592
rect 118608 2100 118660 2106
rect 118608 2042 118660 2048
rect 118332 1964 118384 1970
rect 118332 1906 118384 1912
rect 118608 1896 118660 1902
rect 118660 1856 118740 1884
rect 118608 1838 118660 1844
rect 118712 800 118740 1856
rect 119158 1864 119214 1873
rect 119158 1799 119160 1808
rect 119212 1799 119214 1808
rect 119160 1770 119212 1776
rect 118804 1562 119200 1578
rect 118804 1556 119212 1562
rect 118804 1550 119160 1556
rect 118804 1426 118832 1550
rect 119160 1498 119212 1504
rect 118884 1488 118936 1494
rect 119264 1442 119292 3703
rect 119528 3392 119580 3398
rect 119528 3334 119580 3340
rect 119344 2984 119396 2990
rect 119344 2926 119396 2932
rect 118884 1430 118936 1436
rect 118792 1420 118844 1426
rect 118792 1362 118844 1368
rect 118896 950 118924 1430
rect 119172 1414 119292 1442
rect 118884 944 118936 950
rect 118884 886 118936 892
rect 119172 800 119200 1414
rect 119356 1358 119384 2926
rect 119344 1352 119396 1358
rect 119344 1294 119396 1300
rect 119540 800 119568 3334
rect 119724 814 119752 8842
rect 120000 8378 120028 10200
rect 120356 8968 120408 8974
rect 120356 8910 120408 8916
rect 119908 8350 120028 8378
rect 120264 8356 120316 8362
rect 119804 6860 119856 6866
rect 119804 6802 119856 6808
rect 119816 6458 119844 6802
rect 119804 6452 119856 6458
rect 119804 6394 119856 6400
rect 119804 4684 119856 4690
rect 119804 4626 119856 4632
rect 119816 3233 119844 4626
rect 119908 4282 119936 8350
rect 120264 8298 120316 8304
rect 119988 8288 120040 8294
rect 119988 8230 120040 8236
rect 120000 7818 120028 8230
rect 119988 7812 120040 7818
rect 119988 7754 120040 7760
rect 120172 7812 120224 7818
rect 120172 7754 120224 7760
rect 120080 7200 120132 7206
rect 120080 7142 120132 7148
rect 120092 6186 120120 7142
rect 120184 7002 120212 7754
rect 120172 6996 120224 7002
rect 120172 6938 120224 6944
rect 120276 6866 120304 8298
rect 120172 6860 120224 6866
rect 120172 6802 120224 6808
rect 120264 6860 120316 6866
rect 120264 6802 120316 6808
rect 120080 6180 120132 6186
rect 120080 6122 120132 6128
rect 120184 4690 120212 6802
rect 120368 6746 120396 8910
rect 120276 6718 120396 6746
rect 120172 4684 120224 4690
rect 120172 4626 120224 4632
rect 119896 4276 119948 4282
rect 119896 4218 119948 4224
rect 119988 4276 120040 4282
rect 119988 4218 120040 4224
rect 120000 4049 120028 4218
rect 119986 4040 120042 4049
rect 119986 3975 120042 3984
rect 120170 3632 120226 3641
rect 120170 3567 120226 3576
rect 119802 3224 119858 3233
rect 119802 3159 119858 3168
rect 120184 2922 120212 3567
rect 120172 2916 120224 2922
rect 120172 2858 120224 2864
rect 120172 2508 120224 2514
rect 120172 2450 120224 2456
rect 120184 2417 120212 2450
rect 120170 2408 120226 2417
rect 120170 2343 120226 2352
rect 120172 2304 120224 2310
rect 120172 2246 120224 2252
rect 119988 2032 120040 2038
rect 119988 1974 120040 1980
rect 119896 1896 119948 1902
rect 119896 1838 119948 1844
rect 119712 808 119764 814
rect 115296 604 115348 610
rect 115296 546 115348 552
rect 115662 -400 115718 800
rect 116030 -400 116086 800
rect 116490 -400 116546 800
rect 116950 -400 117006 800
rect 117410 -400 117466 800
rect 117778 -400 117834 800
rect 118238 -400 118294 800
rect 118698 -400 118754 800
rect 119158 -400 119214 800
rect 119526 -400 119582 800
rect 119712 750 119764 756
rect 119908 406 119936 1838
rect 120000 800 120028 1974
rect 120080 1828 120132 1834
rect 120080 1770 120132 1776
rect 120092 1737 120120 1770
rect 120078 1728 120134 1737
rect 120078 1663 120134 1672
rect 120184 1465 120212 2246
rect 120276 2106 120304 6718
rect 120460 5409 120488 10200
rect 120828 7206 120856 10200
rect 121288 10130 121316 10200
rect 121276 10124 121328 10130
rect 121276 10066 121328 10072
rect 121184 10056 121236 10062
rect 121184 9998 121236 10004
rect 121092 8492 121144 8498
rect 121092 8434 121144 8440
rect 121000 7268 121052 7274
rect 121000 7210 121052 7216
rect 120816 7200 120868 7206
rect 120816 7142 120868 7148
rect 120540 6316 120592 6322
rect 120540 6258 120592 6264
rect 120446 5400 120502 5409
rect 120446 5335 120502 5344
rect 120552 4690 120580 6258
rect 120632 6248 120684 6254
rect 120632 6190 120684 6196
rect 120816 6248 120868 6254
rect 120816 6190 120868 6196
rect 120644 5914 120672 6190
rect 120828 6118 120856 6190
rect 120816 6112 120868 6118
rect 120816 6054 120868 6060
rect 120632 5908 120684 5914
rect 120632 5850 120684 5856
rect 120540 4684 120592 4690
rect 120540 4626 120592 4632
rect 120356 3392 120408 3398
rect 120356 3334 120408 3340
rect 120368 3058 120396 3334
rect 120356 3052 120408 3058
rect 120356 2994 120408 3000
rect 120540 2984 120592 2990
rect 120540 2926 120592 2932
rect 120264 2100 120316 2106
rect 120264 2042 120316 2048
rect 120448 1556 120500 1562
rect 120448 1498 120500 1504
rect 120170 1456 120226 1465
rect 120170 1391 120226 1400
rect 120460 800 120488 1498
rect 120552 1222 120580 2926
rect 121012 2553 121040 7210
rect 120998 2544 121054 2553
rect 120998 2479 121054 2488
rect 120814 2272 120870 2281
rect 120814 2207 120870 2216
rect 120540 1216 120592 1222
rect 120540 1158 120592 1164
rect 120828 800 120856 2207
rect 121104 1562 121132 8434
rect 121196 4321 121224 9998
rect 121460 8424 121512 8430
rect 121460 8366 121512 8372
rect 121472 6322 121500 8366
rect 121552 7336 121604 7342
rect 121552 7278 121604 7284
rect 121460 6316 121512 6322
rect 121460 6258 121512 6264
rect 121368 5772 121420 5778
rect 121368 5714 121420 5720
rect 121274 5400 121330 5409
rect 121274 5335 121330 5344
rect 121288 5030 121316 5335
rect 121380 5030 121408 5714
rect 121276 5024 121328 5030
rect 121276 4966 121328 4972
rect 121368 5024 121420 5030
rect 121368 4966 121420 4972
rect 121182 4312 121238 4321
rect 121182 4247 121238 4256
rect 121564 4146 121592 7278
rect 121748 5545 121776 10200
rect 122208 9217 122236 10200
rect 122194 9208 122250 9217
rect 122194 9143 122250 9152
rect 122196 9036 122248 9042
rect 122196 8978 122248 8984
rect 122104 6792 122156 6798
rect 122104 6734 122156 6740
rect 122116 6458 122144 6734
rect 122012 6452 122064 6458
rect 122012 6394 122064 6400
rect 122104 6452 122156 6458
rect 122104 6394 122156 6400
rect 122024 5930 122052 6394
rect 122024 5902 122144 5930
rect 121828 5840 121880 5846
rect 121828 5782 121880 5788
rect 121734 5536 121790 5545
rect 121734 5471 121790 5480
rect 121644 4548 121696 4554
rect 121644 4490 121696 4496
rect 121552 4140 121604 4146
rect 121552 4082 121604 4088
rect 121656 3126 121684 4490
rect 121644 3120 121696 3126
rect 121644 3062 121696 3068
rect 121552 2848 121604 2854
rect 121552 2790 121604 2796
rect 121092 1556 121144 1562
rect 121092 1498 121144 1504
rect 121564 1442 121592 2790
rect 121840 1562 121868 5782
rect 122012 5704 122064 5710
rect 122012 5646 122064 5652
rect 122024 5302 122052 5646
rect 122012 5296 122064 5302
rect 122012 5238 122064 5244
rect 122116 4842 122144 5902
rect 121932 4814 122144 4842
rect 121932 1766 121960 4814
rect 122012 4140 122064 4146
rect 122012 4082 122064 4088
rect 122024 3602 122052 4082
rect 122208 3738 122236 8978
rect 122288 8016 122340 8022
rect 122288 7958 122340 7964
rect 122196 3732 122248 3738
rect 122196 3674 122248 3680
rect 122012 3596 122064 3602
rect 122012 3538 122064 3544
rect 122104 3596 122156 3602
rect 122104 3538 122156 3544
rect 122116 2689 122144 3538
rect 122102 2680 122158 2689
rect 122102 2615 122158 2624
rect 121920 1760 121972 1766
rect 121920 1702 121972 1708
rect 121828 1556 121880 1562
rect 121828 1498 121880 1504
rect 122300 1494 122328 7958
rect 122576 6338 122604 10200
rect 122656 7880 122708 7886
rect 122656 7822 122708 7828
rect 122484 6310 122604 6338
rect 122484 4282 122512 6310
rect 122668 5778 122696 7822
rect 122746 6760 122802 6769
rect 122746 6695 122802 6704
rect 122760 6458 122788 6695
rect 122748 6452 122800 6458
rect 122748 6394 122800 6400
rect 122840 6248 122892 6254
rect 122840 6190 122892 6196
rect 122656 5772 122708 5778
rect 122656 5714 122708 5720
rect 122472 4276 122524 4282
rect 122472 4218 122524 4224
rect 122562 2816 122618 2825
rect 122562 2751 122618 2760
rect 122196 1488 122248 1494
rect 121368 1420 121420 1426
rect 121564 1414 121776 1442
rect 122196 1430 122248 1436
rect 122288 1488 122340 1494
rect 122288 1430 122340 1436
rect 121368 1362 121420 1368
rect 121274 1184 121330 1193
rect 121274 1119 121330 1128
rect 121288 800 121316 1119
rect 119896 400 119948 406
rect 119896 342 119948 348
rect 119986 -400 120042 800
rect 120446 -400 120502 800
rect 120814 -400 120870 800
rect 121274 -400 121330 800
rect 121380 746 121408 1362
rect 121748 800 121776 1414
rect 122208 800 122236 1430
rect 122576 800 122604 2751
rect 122852 2038 122880 6190
rect 123036 5930 123064 10200
rect 123300 8356 123352 8362
rect 123300 8298 123352 8304
rect 123208 8016 123260 8022
rect 123208 7958 123260 7964
rect 123220 7546 123248 7958
rect 123312 7954 123340 8298
rect 123300 7948 123352 7954
rect 123300 7890 123352 7896
rect 123208 7540 123260 7546
rect 123208 7482 123260 7488
rect 123116 6452 123168 6458
rect 123116 6394 123168 6400
rect 122944 5902 123064 5930
rect 122944 5273 122972 5902
rect 123024 5704 123076 5710
rect 123024 5646 123076 5652
rect 122930 5264 122986 5273
rect 122930 5199 122986 5208
rect 123036 3602 123064 5646
rect 123128 4214 123156 6394
rect 123496 5794 123524 10200
rect 123850 7712 123906 7721
rect 123850 7647 123906 7656
rect 123668 6860 123720 6866
rect 123668 6802 123720 6808
rect 123404 5766 123524 5794
rect 123300 5160 123352 5166
rect 123300 5102 123352 5108
rect 123312 4214 123340 5102
rect 123404 4486 123432 5766
rect 123484 5704 123536 5710
rect 123484 5646 123536 5652
rect 123496 5370 123524 5646
rect 123574 5400 123630 5409
rect 123484 5364 123536 5370
rect 123574 5335 123576 5344
rect 123484 5306 123536 5312
rect 123628 5335 123630 5344
rect 123576 5306 123628 5312
rect 123484 5092 123536 5098
rect 123484 5034 123536 5040
rect 123392 4480 123444 4486
rect 123392 4422 123444 4428
rect 123496 4282 123524 5034
rect 123680 4434 123708 6802
rect 123758 6488 123814 6497
rect 123758 6423 123814 6432
rect 123772 6254 123800 6423
rect 123760 6248 123812 6254
rect 123760 6190 123812 6196
rect 123864 5352 123892 7647
rect 123956 5642 123984 10200
rect 124076 9820 124132 9840
rect 124076 9744 124132 9764
rect 124076 8732 124132 8752
rect 124076 8656 124132 8676
rect 124076 7644 124132 7664
rect 124076 7568 124132 7588
rect 124220 7268 124272 7274
rect 124220 7210 124272 7216
rect 124232 6798 124260 7210
rect 124324 6798 124352 10200
rect 124416 9042 124444 10474
rect 124770 10200 124826 11400
rect 125230 10200 125286 11400
rect 125690 10200 125746 11400
rect 126058 10200 126114 11400
rect 126518 10200 126574 11400
rect 126978 10200 127034 11400
rect 127438 10200 127494 11400
rect 127806 10200 127862 11400
rect 128266 10200 128322 11400
rect 128544 10260 128596 10266
rect 128544 10202 128596 10208
rect 124680 9580 124732 9586
rect 124680 9522 124732 9528
rect 124496 9512 124548 9518
rect 124496 9454 124548 9460
rect 124404 9036 124456 9042
rect 124404 8978 124456 8984
rect 124404 7812 124456 7818
rect 124404 7754 124456 7760
rect 124220 6792 124272 6798
rect 124220 6734 124272 6740
rect 124312 6792 124364 6798
rect 124312 6734 124364 6740
rect 124076 6556 124132 6576
rect 124076 6480 124132 6500
rect 124416 6390 124444 7754
rect 124404 6384 124456 6390
rect 124404 6326 124456 6332
rect 124404 6248 124456 6254
rect 124402 6216 124404 6225
rect 124456 6216 124458 6225
rect 124402 6151 124458 6160
rect 123944 5636 123996 5642
rect 123944 5578 123996 5584
rect 124076 5468 124132 5488
rect 124076 5392 124132 5412
rect 123864 5324 124260 5352
rect 123760 5024 123812 5030
rect 123760 4966 123812 4972
rect 123772 4593 123800 4966
rect 123852 4684 123904 4690
rect 123852 4626 123904 4632
rect 123758 4584 123814 4593
rect 123758 4519 123814 4528
rect 123680 4406 123800 4434
rect 123484 4276 123536 4282
rect 123484 4218 123536 4224
rect 123116 4208 123168 4214
rect 123116 4150 123168 4156
rect 123300 4208 123352 4214
rect 123300 4150 123352 4156
rect 123392 4072 123444 4078
rect 123392 4014 123444 4020
rect 123024 3596 123076 3602
rect 123024 3538 123076 3544
rect 123404 3448 123432 4014
rect 123404 3420 123708 3448
rect 123574 3224 123630 3233
rect 123300 3188 123352 3194
rect 123574 3159 123630 3168
rect 123300 3130 123352 3136
rect 123312 2854 123340 3130
rect 123588 3058 123616 3159
rect 123576 3052 123628 3058
rect 123576 2994 123628 3000
rect 123300 2848 123352 2854
rect 123300 2790 123352 2796
rect 123680 2650 123708 3420
rect 123668 2644 123720 2650
rect 123668 2586 123720 2592
rect 122840 2032 122892 2038
rect 123772 2009 123800 4406
rect 122840 1974 122892 1980
rect 123758 2000 123814 2009
rect 123758 1935 123814 1944
rect 123024 1828 123076 1834
rect 123024 1770 123076 1776
rect 123036 800 123064 1770
rect 123760 1556 123812 1562
rect 123760 1498 123812 1504
rect 123772 1426 123800 1498
rect 123760 1420 123812 1426
rect 123760 1362 123812 1368
rect 123392 1352 123444 1358
rect 123392 1294 123444 1300
rect 123404 898 123432 1294
rect 123864 921 123892 4626
rect 124128 4616 124180 4622
rect 124126 4584 124128 4593
rect 124180 4584 124182 4593
rect 124126 4519 124182 4528
rect 124232 4457 124260 5324
rect 124218 4448 124274 4457
rect 124076 4380 124132 4400
rect 124218 4383 124274 4392
rect 123942 4312 123998 4321
rect 124076 4304 124132 4324
rect 124218 4312 124274 4321
rect 123998 4256 124218 4264
rect 123942 4247 124274 4256
rect 123956 4236 124260 4247
rect 123942 3768 123998 3777
rect 123942 3703 123998 3712
rect 123956 3194 123984 3703
rect 124076 3292 124132 3312
rect 124076 3216 124132 3236
rect 123944 3188 123996 3194
rect 123944 3130 123996 3136
rect 123942 2816 123998 2825
rect 123942 2751 123998 2760
rect 123956 1902 123984 2751
rect 124312 2576 124364 2582
rect 124312 2518 124364 2524
rect 124076 2204 124132 2224
rect 124076 2128 124132 2148
rect 124218 2136 124274 2145
rect 124218 2071 124274 2080
rect 123944 1896 123996 1902
rect 123944 1838 123996 1844
rect 124232 1601 124260 2071
rect 124218 1592 124274 1601
rect 124218 1527 124274 1536
rect 124076 1116 124132 1136
rect 124076 1040 124132 1060
rect 123944 944 123996 950
rect 123850 912 123906 921
rect 123404 870 123524 898
rect 123496 800 123524 870
rect 123944 886 123996 892
rect 123850 847 123906 856
rect 123956 800 123984 886
rect 124324 800 124352 2518
rect 124508 2106 124536 9454
rect 124588 8492 124640 8498
rect 124588 8434 124640 8440
rect 124600 6866 124628 8434
rect 124588 6860 124640 6866
rect 124588 6802 124640 6808
rect 124692 6254 124720 9522
rect 124784 8090 124812 10200
rect 125140 10056 125192 10062
rect 125140 9998 125192 10004
rect 125152 8498 125180 9998
rect 125244 8838 125272 10200
rect 125508 9580 125560 9586
rect 125508 9522 125560 9528
rect 125232 8832 125284 8838
rect 125232 8774 125284 8780
rect 125140 8492 125192 8498
rect 125140 8434 125192 8440
rect 124772 8084 124824 8090
rect 124772 8026 124824 8032
rect 124864 7948 124916 7954
rect 124864 7890 124916 7896
rect 124772 7472 124824 7478
rect 124772 7414 124824 7420
rect 124784 7177 124812 7414
rect 124770 7168 124826 7177
rect 124770 7103 124826 7112
rect 124680 6248 124732 6254
rect 124680 6190 124732 6196
rect 124772 5772 124824 5778
rect 124772 5714 124824 5720
rect 124784 5370 124812 5714
rect 124772 5364 124824 5370
rect 124772 5306 124824 5312
rect 124680 5296 124732 5302
rect 124680 5238 124732 5244
rect 124692 5166 124720 5238
rect 124680 5160 124732 5166
rect 124680 5102 124732 5108
rect 124588 3392 124640 3398
rect 124588 3334 124640 3340
rect 124600 3210 124628 3334
rect 124600 3182 124812 3210
rect 124680 2508 124732 2514
rect 124680 2450 124732 2456
rect 124692 2417 124720 2450
rect 124678 2408 124734 2417
rect 124678 2343 124734 2352
rect 124496 2100 124548 2106
rect 124496 2042 124548 2048
rect 124680 1760 124732 1766
rect 124680 1702 124732 1708
rect 124692 1494 124720 1702
rect 124680 1488 124732 1494
rect 124680 1430 124732 1436
rect 124784 800 124812 3182
rect 124876 2106 124904 7890
rect 125048 7200 125100 7206
rect 125048 7142 125100 7148
rect 125232 7200 125284 7206
rect 125232 7142 125284 7148
rect 124956 6792 125008 6798
rect 124956 6734 125008 6740
rect 124968 4826 124996 6734
rect 124956 4820 125008 4826
rect 124956 4762 125008 4768
rect 125060 4690 125088 7142
rect 125048 4684 125100 4690
rect 125048 4626 125100 4632
rect 125244 4486 125272 7142
rect 125520 6866 125548 9522
rect 125704 7970 125732 10200
rect 125782 9072 125838 9081
rect 125782 9007 125838 9016
rect 125612 7942 125732 7970
rect 125508 6860 125560 6866
rect 125508 6802 125560 6808
rect 125612 6202 125640 7942
rect 125692 7880 125744 7886
rect 125692 7822 125744 7828
rect 125520 6174 125640 6202
rect 125520 6118 125548 6174
rect 125704 6118 125732 7822
rect 125796 6662 125824 9007
rect 125876 8900 125928 8906
rect 125876 8842 125928 8848
rect 125888 7721 125916 8842
rect 125874 7712 125930 7721
rect 125874 7647 125930 7656
rect 126072 7478 126100 10200
rect 126152 8356 126204 8362
rect 126152 8298 126204 8304
rect 126060 7472 126112 7478
rect 126060 7414 126112 7420
rect 126164 7342 126192 8298
rect 126152 7336 126204 7342
rect 126152 7278 126204 7284
rect 126152 7200 126204 7206
rect 126152 7142 126204 7148
rect 125968 6860 126020 6866
rect 125968 6802 126020 6808
rect 125980 6769 126008 6802
rect 125966 6760 126022 6769
rect 125966 6695 126022 6704
rect 125784 6656 125836 6662
rect 125784 6598 125836 6604
rect 125968 6656 126020 6662
rect 126164 6610 126192 7142
rect 125968 6598 126020 6604
rect 125980 6322 126008 6598
rect 126072 6582 126192 6610
rect 126072 6458 126100 6582
rect 126060 6452 126112 6458
rect 126060 6394 126112 6400
rect 125968 6316 126020 6322
rect 125968 6258 126020 6264
rect 125784 6248 125836 6254
rect 125784 6190 125836 6196
rect 125508 6112 125560 6118
rect 125508 6054 125560 6060
rect 125692 6112 125744 6118
rect 125692 6054 125744 6060
rect 125690 5264 125746 5273
rect 125690 5199 125746 5208
rect 125232 4480 125284 4486
rect 125232 4422 125284 4428
rect 125704 4010 125732 5199
rect 125692 4004 125744 4010
rect 125692 3946 125744 3952
rect 125506 3632 125562 3641
rect 125506 3567 125562 3576
rect 125600 3596 125652 3602
rect 125520 3398 125548 3567
rect 125600 3538 125652 3544
rect 125508 3392 125560 3398
rect 125508 3334 125560 3340
rect 125612 3058 125640 3538
rect 125600 3052 125652 3058
rect 125600 2994 125652 3000
rect 125138 2952 125194 2961
rect 125138 2887 125194 2896
rect 125324 2916 125376 2922
rect 125152 2854 125180 2887
rect 125324 2858 125376 2864
rect 125140 2848 125192 2854
rect 125140 2790 125192 2796
rect 125230 2544 125286 2553
rect 125230 2479 125286 2488
rect 125140 2372 125192 2378
rect 125140 2314 125192 2320
rect 124864 2100 124916 2106
rect 124864 2042 124916 2048
rect 124956 1828 125008 1834
rect 124956 1770 125008 1776
rect 124862 1456 124918 1465
rect 124968 1442 124996 1770
rect 125048 1760 125100 1766
rect 125048 1702 125100 1708
rect 125060 1601 125088 1702
rect 125046 1592 125102 1601
rect 125046 1527 125102 1536
rect 124968 1426 125088 1442
rect 124968 1420 125100 1426
rect 124968 1414 125048 1420
rect 124862 1391 124864 1400
rect 124916 1391 124918 1400
rect 124864 1362 124916 1368
rect 125048 1362 125100 1368
rect 125152 1358 125180 2314
rect 125244 1494 125272 2479
rect 125336 2106 125364 2858
rect 125416 2848 125468 2854
rect 125416 2790 125468 2796
rect 125428 2689 125456 2790
rect 125414 2680 125470 2689
rect 125796 2650 125824 6190
rect 126532 5930 126560 10200
rect 126794 9208 126850 9217
rect 126794 9143 126850 9152
rect 126612 8492 126664 8498
rect 126612 8434 126664 8440
rect 126624 8265 126652 8434
rect 126704 8424 126756 8430
rect 126704 8366 126756 8372
rect 126610 8256 126666 8265
rect 126610 8191 126666 8200
rect 126072 5902 126560 5930
rect 126612 5908 126664 5914
rect 126072 5030 126100 5902
rect 126612 5850 126664 5856
rect 126624 5794 126652 5850
rect 126348 5778 126652 5794
rect 126336 5772 126652 5778
rect 126388 5766 126652 5772
rect 126336 5714 126388 5720
rect 126244 5296 126296 5302
rect 126164 5256 126244 5284
rect 126060 5024 126112 5030
rect 126060 4966 126112 4972
rect 126164 4690 126192 5256
rect 126244 5238 126296 5244
rect 126244 5160 126296 5166
rect 126244 5102 126296 5108
rect 126256 4826 126284 5102
rect 126716 5030 126744 8366
rect 126808 5273 126836 9143
rect 126886 8392 126942 8401
rect 126886 8327 126942 8336
rect 126794 5264 126850 5273
rect 126794 5199 126850 5208
rect 126704 5024 126756 5030
rect 126704 4966 126756 4972
rect 126244 4820 126296 4826
rect 126244 4762 126296 4768
rect 126336 4752 126388 4758
rect 126336 4694 126388 4700
rect 126152 4684 126204 4690
rect 126152 4626 126204 4632
rect 126348 4554 126376 4694
rect 126796 4616 126848 4622
rect 126796 4558 126848 4564
rect 126336 4548 126388 4554
rect 126336 4490 126388 4496
rect 126520 4548 126572 4554
rect 126520 4490 126572 4496
rect 126532 4282 126560 4490
rect 126808 4486 126836 4558
rect 126796 4480 126848 4486
rect 126796 4422 126848 4428
rect 126520 4276 126572 4282
rect 126520 4218 126572 4224
rect 126900 4214 126928 8327
rect 126992 7290 127020 10200
rect 127254 7304 127310 7313
rect 126992 7262 127112 7290
rect 127084 5914 127112 7262
rect 127254 7239 127310 7248
rect 127268 6497 127296 7239
rect 127452 7206 127480 10200
rect 127820 8922 127848 10200
rect 128280 9738 128308 10200
rect 127544 8894 127848 8922
rect 128004 9710 128308 9738
rect 127440 7200 127492 7206
rect 127440 7142 127492 7148
rect 127544 6882 127572 8894
rect 127808 8832 127860 8838
rect 127808 8774 127860 8780
rect 127820 8498 127848 8774
rect 127808 8492 127860 8498
rect 127808 8434 127860 8440
rect 127900 8356 127952 8362
rect 127900 8298 127952 8304
rect 127716 7404 127768 7410
rect 127716 7346 127768 7352
rect 127622 7304 127678 7313
rect 127622 7239 127678 7248
rect 127360 6854 127572 6882
rect 127254 6488 127310 6497
rect 127254 6423 127310 6432
rect 127072 5908 127124 5914
rect 127072 5850 127124 5856
rect 127360 4865 127388 6854
rect 127636 6798 127664 7239
rect 127728 6934 127756 7346
rect 127808 7336 127860 7342
rect 127808 7278 127860 7284
rect 127716 6928 127768 6934
rect 127716 6870 127768 6876
rect 127624 6792 127676 6798
rect 127530 6760 127586 6769
rect 127624 6734 127676 6740
rect 127714 6760 127770 6769
rect 127530 6695 127586 6704
rect 127714 6695 127770 6704
rect 127544 5846 127572 6695
rect 127728 6225 127756 6695
rect 127714 6216 127770 6225
rect 127714 6151 127770 6160
rect 127624 6112 127676 6118
rect 127624 6054 127676 6060
rect 127440 5840 127492 5846
rect 127440 5782 127492 5788
rect 127532 5840 127584 5846
rect 127532 5782 127584 5788
rect 127346 4856 127402 4865
rect 127346 4791 127402 4800
rect 126336 4208 126388 4214
rect 126336 4150 126388 4156
rect 126428 4208 126480 4214
rect 126428 4150 126480 4156
rect 126888 4208 126940 4214
rect 126888 4150 126940 4156
rect 125876 4072 125928 4078
rect 125876 4014 125928 4020
rect 126242 4040 126298 4049
rect 125888 3482 125916 4014
rect 126242 3975 126298 3984
rect 125968 3936 126020 3942
rect 125968 3878 126020 3884
rect 126058 3904 126114 3913
rect 125980 3777 126008 3878
rect 126058 3839 126114 3848
rect 125966 3768 126022 3777
rect 125966 3703 126022 3712
rect 125966 3632 126022 3641
rect 126072 3602 126100 3839
rect 126256 3670 126284 3975
rect 126244 3664 126296 3670
rect 126244 3606 126296 3612
rect 125966 3567 125968 3576
rect 126020 3567 126022 3576
rect 126060 3596 126112 3602
rect 125968 3538 126020 3544
rect 126060 3538 126112 3544
rect 125888 3454 126192 3482
rect 126164 3398 126192 3454
rect 125968 3392 126020 3398
rect 125968 3334 126020 3340
rect 126152 3392 126204 3398
rect 126152 3334 126204 3340
rect 125414 2615 125470 2624
rect 125600 2644 125652 2650
rect 125600 2586 125652 2592
rect 125784 2644 125836 2650
rect 125784 2586 125836 2592
rect 125324 2100 125376 2106
rect 125324 2042 125376 2048
rect 125322 2000 125378 2009
rect 125322 1935 125378 1944
rect 125336 1834 125364 1935
rect 125324 1828 125376 1834
rect 125324 1770 125376 1776
rect 125232 1488 125284 1494
rect 125232 1430 125284 1436
rect 125140 1352 125192 1358
rect 125140 1294 125192 1300
rect 125612 1306 125640 2586
rect 125690 2544 125746 2553
rect 125690 2479 125692 2488
rect 125744 2479 125746 2488
rect 125692 2450 125744 2456
rect 125782 2000 125838 2009
rect 125782 1935 125838 1944
rect 125796 1902 125824 1935
rect 125784 1896 125836 1902
rect 125784 1838 125836 1844
rect 125612 1278 125732 1306
rect 125232 1216 125284 1222
rect 125232 1158 125284 1164
rect 125244 800 125272 1158
rect 125704 800 125732 1278
rect 125980 1222 126008 3334
rect 126348 3194 126376 4150
rect 126244 3188 126296 3194
rect 126244 3130 126296 3136
rect 126336 3188 126388 3194
rect 126336 3130 126388 3136
rect 126060 3120 126112 3126
rect 126060 3062 126112 3068
rect 125968 1216 126020 1222
rect 125968 1158 126020 1164
rect 126072 800 126100 3062
rect 126256 950 126284 3130
rect 126440 3058 126468 4150
rect 127164 4072 127216 4078
rect 127164 4014 127216 4020
rect 126794 3904 126850 3913
rect 126794 3839 126850 3848
rect 126428 3052 126480 3058
rect 126428 2994 126480 3000
rect 126808 2106 126836 3839
rect 126980 2984 127032 2990
rect 126980 2926 127032 2932
rect 126888 2916 126940 2922
rect 126888 2858 126940 2864
rect 126520 2100 126572 2106
rect 126520 2042 126572 2048
rect 126796 2100 126848 2106
rect 126796 2042 126848 2048
rect 126244 944 126296 950
rect 126244 886 126296 892
rect 126532 800 126560 2042
rect 126808 1902 126836 2042
rect 126900 1986 126928 2858
rect 126992 2650 127020 2926
rect 126980 2644 127032 2650
rect 126980 2586 127032 2592
rect 126900 1958 127020 1986
rect 126796 1896 126848 1902
rect 126888 1896 126940 1902
rect 126796 1838 126848 1844
rect 126886 1864 126888 1873
rect 126940 1864 126942 1873
rect 126886 1799 126942 1808
rect 126992 800 127020 1958
rect 121368 740 121420 746
rect 121368 682 121420 688
rect 121734 -400 121790 800
rect 122194 -400 122250 800
rect 122562 -400 122618 800
rect 123022 -400 123078 800
rect 123482 -400 123538 800
rect 123942 -400 123998 800
rect 124310 -400 124366 800
rect 124770 -400 124826 800
rect 125230 -400 125286 800
rect 125690 -400 125746 800
rect 126058 -400 126114 800
rect 126518 -400 126574 800
rect 126978 -400 127034 800
rect 127176 377 127204 4014
rect 127452 3602 127480 5782
rect 127636 5710 127664 6054
rect 127532 5704 127584 5710
rect 127532 5646 127584 5652
rect 127624 5704 127676 5710
rect 127624 5646 127676 5652
rect 127544 5545 127572 5646
rect 127530 5536 127586 5545
rect 127530 5471 127586 5480
rect 127440 3596 127492 3602
rect 127440 3538 127492 3544
rect 127348 2372 127400 2378
rect 127348 2314 127400 2320
rect 127440 2372 127492 2378
rect 127440 2314 127492 2320
rect 127360 1873 127388 2314
rect 127452 2145 127480 2314
rect 127438 2136 127494 2145
rect 127622 2136 127678 2145
rect 127438 2071 127494 2080
rect 127544 2094 127622 2122
rect 127346 1864 127402 1873
rect 127346 1799 127402 1808
rect 127544 1290 127572 2094
rect 127820 2106 127848 7278
rect 127912 6798 127940 8298
rect 127900 6792 127952 6798
rect 127900 6734 127952 6740
rect 128004 5681 128032 9710
rect 128360 9376 128412 9382
rect 128360 9318 128412 9324
rect 128452 9376 128504 9382
rect 128452 9318 128504 9324
rect 128084 9036 128136 9042
rect 128084 8978 128136 8984
rect 127990 5672 128046 5681
rect 127990 5607 128046 5616
rect 128096 5114 128124 8978
rect 128372 8922 128400 9318
rect 128464 9042 128492 9318
rect 128452 9036 128504 9042
rect 128452 8978 128504 8984
rect 128372 8894 128492 8922
rect 128360 7880 128412 7886
rect 128360 7822 128412 7828
rect 128268 6316 128320 6322
rect 128268 6258 128320 6264
rect 128280 5914 128308 6258
rect 128268 5908 128320 5914
rect 128268 5850 128320 5856
rect 128176 5772 128228 5778
rect 128176 5714 128228 5720
rect 128188 5681 128216 5714
rect 128174 5672 128230 5681
rect 128174 5607 128230 5616
rect 128174 5400 128230 5409
rect 128174 5335 128230 5344
rect 128188 5234 128216 5335
rect 128176 5228 128228 5234
rect 128176 5170 128228 5176
rect 128096 5086 128308 5114
rect 128084 5024 128136 5030
rect 128084 4966 128136 4972
rect 127992 4684 128044 4690
rect 127992 4626 128044 4632
rect 127900 4548 127952 4554
rect 127900 4490 127952 4496
rect 127912 3126 127940 4490
rect 127900 3120 127952 3126
rect 127900 3062 127952 3068
rect 127622 2071 127678 2080
rect 127808 2100 127860 2106
rect 127808 2042 127860 2048
rect 127900 1556 127952 1562
rect 127900 1498 127952 1504
rect 127808 1352 127860 1358
rect 127808 1294 127860 1300
rect 127532 1284 127584 1290
rect 127532 1226 127584 1232
rect 127440 1216 127492 1222
rect 127440 1158 127492 1164
rect 127624 1216 127676 1222
rect 127624 1158 127676 1164
rect 127452 800 127480 1158
rect 127636 882 127664 1158
rect 127624 876 127676 882
rect 127624 818 127676 824
rect 127820 800 127848 1294
rect 127912 1290 127940 1498
rect 127900 1284 127952 1290
rect 127900 1226 127952 1232
rect 128004 882 128032 4626
rect 128096 2446 128124 4966
rect 128176 4072 128228 4078
rect 128176 4014 128228 4020
rect 128188 2582 128216 4014
rect 128280 3738 128308 5086
rect 128268 3732 128320 3738
rect 128268 3674 128320 3680
rect 128268 3528 128320 3534
rect 128266 3496 128268 3505
rect 128320 3496 128322 3505
rect 128266 3431 128322 3440
rect 128268 3188 128320 3194
rect 128268 3130 128320 3136
rect 128176 2576 128228 2582
rect 128176 2518 128228 2524
rect 128084 2440 128136 2446
rect 128084 2382 128136 2388
rect 128176 1964 128228 1970
rect 128176 1906 128228 1912
rect 128188 1766 128216 1906
rect 128176 1760 128228 1766
rect 128176 1702 128228 1708
rect 128084 1556 128136 1562
rect 128084 1498 128136 1504
rect 128096 1426 128124 1498
rect 128084 1420 128136 1426
rect 128084 1362 128136 1368
rect 127992 876 128044 882
rect 127992 818 128044 824
rect 128280 800 128308 3130
rect 127162 368 127218 377
rect 127162 303 127218 312
rect 127438 -400 127494 800
rect 127806 -400 127862 800
rect 128266 -400 128322 800
rect 128372 105 128400 7822
rect 128464 7177 128492 8894
rect 128450 7168 128506 7177
rect 128450 7103 128506 7112
rect 128556 7018 128584 10202
rect 128726 10200 128782 11400
rect 128912 10396 128964 10402
rect 128912 10338 128964 10344
rect 128636 7200 128688 7206
rect 128636 7142 128688 7148
rect 128464 6990 128584 7018
rect 128464 4214 128492 6990
rect 128544 5568 128596 5574
rect 128544 5510 128596 5516
rect 128556 4865 128584 5510
rect 128648 5166 128676 7142
rect 128636 5160 128688 5166
rect 128636 5102 128688 5108
rect 128542 4856 128598 4865
rect 128542 4791 128598 4800
rect 128636 4480 128688 4486
rect 128636 4422 128688 4428
rect 128648 4214 128676 4422
rect 128452 4208 128504 4214
rect 128452 4150 128504 4156
rect 128636 4208 128688 4214
rect 128636 4150 128688 4156
rect 128740 4049 128768 10200
rect 128818 8936 128874 8945
rect 128818 8871 128874 8880
rect 128832 6730 128860 8871
rect 128820 6724 128872 6730
rect 128820 6666 128872 6672
rect 128924 6474 128952 10338
rect 129094 10200 129150 11400
rect 129554 10200 129610 11400
rect 130014 10200 130070 11400
rect 130384 10260 130436 10266
rect 130384 10202 130436 10208
rect 129108 10146 129136 10200
rect 129004 10124 129056 10130
rect 129108 10118 129228 10146
rect 129004 10066 129056 10072
rect 129016 8566 129044 10066
rect 129004 8560 129056 8566
rect 129004 8502 129056 8508
rect 129096 6860 129148 6866
rect 129096 6802 129148 6808
rect 128924 6446 129044 6474
rect 128820 5772 128872 5778
rect 128820 5714 128872 5720
rect 128726 4040 128782 4049
rect 128726 3975 128782 3984
rect 128634 3768 128690 3777
rect 128634 3703 128636 3712
rect 128688 3703 128690 3712
rect 128636 3674 128688 3680
rect 128450 3496 128506 3505
rect 128450 3431 128452 3440
rect 128504 3431 128506 3440
rect 128452 3402 128504 3408
rect 128726 3224 128782 3233
rect 128726 3159 128728 3168
rect 128780 3159 128782 3168
rect 128728 3130 128780 3136
rect 128636 2984 128688 2990
rect 128450 2952 128506 2961
rect 128688 2932 128768 2938
rect 128636 2926 128768 2932
rect 128648 2910 128768 2926
rect 128450 2887 128452 2896
rect 128504 2887 128506 2896
rect 128452 2858 128504 2864
rect 128544 2848 128596 2854
rect 128464 2796 128544 2802
rect 128464 2790 128596 2796
rect 128464 2774 128584 2790
rect 128464 2514 128492 2774
rect 128452 2508 128504 2514
rect 128452 2450 128504 2456
rect 128452 1420 128504 1426
rect 128452 1362 128504 1368
rect 128464 474 128492 1362
rect 128740 800 128768 2910
rect 128832 2689 128860 5714
rect 128912 5636 128964 5642
rect 128912 5578 128964 5584
rect 128818 2680 128874 2689
rect 128818 2615 128874 2624
rect 128924 1057 128952 5578
rect 129016 3890 129044 6446
rect 129108 4060 129136 6802
rect 129200 6118 129228 10118
rect 129280 9580 129332 9586
rect 129280 9522 129332 9528
rect 129292 8809 129320 9522
rect 129464 9512 129516 9518
rect 129464 9454 129516 9460
rect 129372 8900 129424 8906
rect 129372 8842 129424 8848
rect 129278 8800 129334 8809
rect 129278 8735 129334 8744
rect 129384 7585 129412 8842
rect 129370 7576 129426 7585
rect 129370 7511 129426 7520
rect 129280 6860 129332 6866
rect 129280 6802 129332 6808
rect 129188 6112 129240 6118
rect 129188 6054 129240 6060
rect 129292 5778 129320 6802
rect 129280 5772 129332 5778
rect 129280 5714 129332 5720
rect 129372 5636 129424 5642
rect 129372 5578 129424 5584
rect 129384 5370 129412 5578
rect 129372 5364 129424 5370
rect 129372 5306 129424 5312
rect 129108 4032 129228 4060
rect 129016 3862 129136 3890
rect 129004 3596 129056 3602
rect 129004 3538 129056 3544
rect 128910 1048 128966 1057
rect 128910 983 128966 992
rect 128452 468 128504 474
rect 128452 410 128504 416
rect 128358 96 128414 105
rect 128358 31 128414 40
rect 128726 -400 128782 800
rect 129016 134 129044 3538
rect 129108 3194 129136 3862
rect 129096 3188 129148 3194
rect 129096 3130 129148 3136
rect 129200 1986 129228 4032
rect 129278 3360 129334 3369
rect 129278 3295 129334 3304
rect 129292 3194 129320 3295
rect 129280 3188 129332 3194
rect 129280 3130 129332 3136
rect 129280 3052 129332 3058
rect 129280 2994 129332 3000
rect 129292 2378 129320 2994
rect 129372 2508 129424 2514
rect 129372 2450 129424 2456
rect 129280 2372 129332 2378
rect 129280 2314 129332 2320
rect 129200 1958 129320 1986
rect 129188 1828 129240 1834
rect 129188 1770 129240 1776
rect 129200 1494 129228 1770
rect 129188 1488 129240 1494
rect 129188 1430 129240 1436
rect 129292 1290 129320 1958
rect 129096 1284 129148 1290
rect 129096 1226 129148 1232
rect 129280 1284 129332 1290
rect 129280 1226 129332 1232
rect 129108 800 129136 1226
rect 129004 128 129056 134
rect 129004 70 129056 76
rect 129094 -400 129150 800
rect 129384 338 129412 2450
rect 129476 1494 129504 9454
rect 129568 9217 129596 10200
rect 129554 9208 129610 9217
rect 129554 9143 129610 9152
rect 129556 9036 129608 9042
rect 129556 8978 129608 8984
rect 129568 2650 129596 8978
rect 129648 8424 129700 8430
rect 129648 8366 129700 8372
rect 129660 2990 129688 8366
rect 129832 7744 129884 7750
rect 129832 7686 129884 7692
rect 129738 5400 129794 5409
rect 129738 5335 129740 5344
rect 129792 5335 129794 5344
rect 129740 5306 129792 5312
rect 129738 3360 129794 3369
rect 129738 3295 129794 3304
rect 129648 2984 129700 2990
rect 129648 2926 129700 2932
rect 129752 2836 129780 3295
rect 129660 2808 129780 2836
rect 129556 2644 129608 2650
rect 129556 2586 129608 2592
rect 129556 2508 129608 2514
rect 129556 2450 129608 2456
rect 129568 2310 129596 2450
rect 129556 2304 129608 2310
rect 129556 2246 129608 2252
rect 129556 1760 129608 1766
rect 129556 1702 129608 1708
rect 129464 1488 129516 1494
rect 129464 1430 129516 1436
rect 129568 800 129596 1702
rect 129660 1426 129688 2808
rect 129844 2310 129872 7686
rect 130028 5545 130056 10200
rect 130396 9586 130424 10202
rect 130474 10200 130530 11400
rect 130842 10200 130898 11400
rect 131302 10200 131358 11400
rect 131762 10200 131818 11400
rect 132222 10200 132278 11400
rect 132590 10200 132646 11400
rect 132960 10464 133012 10470
rect 132960 10406 133012 10412
rect 130384 9580 130436 9586
rect 130384 9522 130436 9528
rect 130384 9036 130436 9042
rect 130384 8978 130436 8984
rect 130292 7200 130344 7206
rect 130292 7142 130344 7148
rect 130200 6656 130252 6662
rect 130200 6598 130252 6604
rect 130212 6186 130240 6598
rect 130200 6180 130252 6186
rect 130200 6122 130252 6128
rect 130014 5536 130070 5545
rect 130014 5471 130070 5480
rect 130200 5160 130252 5166
rect 130200 5102 130252 5108
rect 129924 4684 129976 4690
rect 129924 4626 129976 4632
rect 129936 3505 129964 4626
rect 129922 3496 129978 3505
rect 129922 3431 129978 3440
rect 130108 3188 130160 3194
rect 130108 3130 130160 3136
rect 129924 2984 129976 2990
rect 129924 2926 129976 2932
rect 129936 2650 129964 2926
rect 129924 2644 129976 2650
rect 129924 2586 129976 2592
rect 129740 2304 129792 2310
rect 129740 2246 129792 2252
rect 129832 2304 129884 2310
rect 129832 2246 129884 2252
rect 129648 1420 129700 1426
rect 129648 1362 129700 1368
rect 129752 1306 129780 2246
rect 129660 1278 129780 1306
rect 129372 332 129424 338
rect 129372 274 129424 280
rect 129554 -400 129610 800
rect 129660 270 129688 1278
rect 130120 950 130148 3130
rect 130212 2446 130240 5102
rect 130304 3602 130332 7142
rect 130396 4214 130424 8978
rect 130488 8974 130516 10200
rect 130568 9580 130620 9586
rect 130568 9522 130620 9528
rect 130476 8968 130528 8974
rect 130476 8910 130528 8916
rect 130474 7304 130530 7313
rect 130474 7239 130530 7248
rect 130488 6662 130516 7239
rect 130476 6656 130528 6662
rect 130476 6598 130528 6604
rect 130476 5160 130528 5166
rect 130476 5102 130528 5108
rect 130384 4208 130436 4214
rect 130384 4150 130436 4156
rect 130292 3596 130344 3602
rect 130292 3538 130344 3544
rect 130488 3482 130516 5102
rect 130396 3454 130516 3482
rect 130200 2440 130252 2446
rect 130200 2382 130252 2388
rect 130396 2378 130424 3454
rect 130476 3392 130528 3398
rect 130476 3334 130528 3340
rect 130384 2372 130436 2378
rect 130384 2314 130436 2320
rect 130292 1896 130344 1902
rect 130292 1838 130344 1844
rect 130016 944 130068 950
rect 130016 886 130068 892
rect 130108 944 130160 950
rect 130108 886 130160 892
rect 130028 800 130056 886
rect 129648 264 129700 270
rect 129648 206 129700 212
rect 130014 -400 130070 800
rect 130304 202 130332 1838
rect 130488 800 130516 3334
rect 130292 196 130344 202
rect 130292 138 130344 144
rect 130474 -400 130530 800
rect 130580 649 130608 9522
rect 130856 9081 130884 10200
rect 130842 9072 130898 9081
rect 130842 9007 130898 9016
rect 130844 8968 130896 8974
rect 130844 8910 130896 8916
rect 130856 8362 130884 8910
rect 131316 8566 131344 10200
rect 131776 9994 131804 10200
rect 131764 9988 131816 9994
rect 131764 9930 131816 9936
rect 132236 8922 132264 10200
rect 132316 9512 132368 9518
rect 132316 9454 132368 9460
rect 132052 8894 132264 8922
rect 131670 8664 131726 8673
rect 131670 8599 131726 8608
rect 131304 8560 131356 8566
rect 131304 8502 131356 8508
rect 130844 8356 130896 8362
rect 130844 8298 130896 8304
rect 131396 7948 131448 7954
rect 131396 7890 131448 7896
rect 130844 7880 130896 7886
rect 130844 7822 130896 7828
rect 130660 5704 130712 5710
rect 130660 5646 130712 5652
rect 130672 3126 130700 5646
rect 130856 3194 130884 7822
rect 131304 6860 131356 6866
rect 131304 6802 131356 6808
rect 131212 6724 131264 6730
rect 131212 6666 131264 6672
rect 131026 6624 131082 6633
rect 131026 6559 131082 6568
rect 130936 6248 130988 6254
rect 130936 6190 130988 6196
rect 130948 4826 130976 6190
rect 131040 5302 131068 6559
rect 131120 6112 131172 6118
rect 131120 6054 131172 6060
rect 131028 5296 131080 5302
rect 131028 5238 131080 5244
rect 131132 5234 131160 6054
rect 131224 5370 131252 6666
rect 131316 5370 131344 6802
rect 131212 5364 131264 5370
rect 131212 5306 131264 5312
rect 131304 5364 131356 5370
rect 131304 5306 131356 5312
rect 131302 5264 131358 5273
rect 131120 5228 131172 5234
rect 131302 5199 131358 5208
rect 131120 5170 131172 5176
rect 131120 5092 131172 5098
rect 131120 5034 131172 5040
rect 131212 5092 131264 5098
rect 131212 5034 131264 5040
rect 130936 4820 130988 4826
rect 130936 4762 130988 4768
rect 131132 4282 131160 5034
rect 131120 4276 131172 4282
rect 131120 4218 131172 4224
rect 131028 4140 131080 4146
rect 131028 4082 131080 4088
rect 131040 4049 131068 4082
rect 131026 4040 131082 4049
rect 131026 3975 131082 3984
rect 131120 3596 131172 3602
rect 131120 3538 131172 3544
rect 130844 3188 130896 3194
rect 130844 3130 130896 3136
rect 130660 3120 130712 3126
rect 130660 3062 130712 3068
rect 131132 3058 131160 3538
rect 131224 3466 131252 5034
rect 131316 4622 131344 5199
rect 131304 4616 131356 4622
rect 131304 4558 131356 4564
rect 131304 3732 131356 3738
rect 131304 3674 131356 3680
rect 131212 3460 131264 3466
rect 131212 3402 131264 3408
rect 131120 3052 131172 3058
rect 131120 2994 131172 3000
rect 131212 2984 131264 2990
rect 131212 2926 131264 2932
rect 130844 2916 130896 2922
rect 130844 2858 130896 2864
rect 130752 2304 130804 2310
rect 130752 2246 130804 2252
rect 130764 1834 130792 2246
rect 130752 1828 130804 1834
rect 130752 1770 130804 1776
rect 130856 800 130884 2858
rect 130936 2508 130988 2514
rect 130936 2450 130988 2456
rect 130566 640 130622 649
rect 130566 575 130622 584
rect 130842 -400 130898 800
rect 130948 542 130976 2450
rect 131028 2304 131080 2310
rect 131028 2246 131080 2252
rect 131040 2038 131068 2246
rect 131028 2032 131080 2038
rect 131224 1986 131252 2926
rect 131316 2038 131344 3674
rect 131028 1974 131080 1980
rect 131132 1958 131252 1986
rect 131304 2032 131356 2038
rect 131304 1974 131356 1980
rect 130936 536 130988 542
rect 130936 478 130988 484
rect 131132 66 131160 1958
rect 131212 1896 131264 1902
rect 131408 1884 131436 7890
rect 131488 6860 131540 6866
rect 131488 6802 131540 6808
rect 131500 5234 131528 6802
rect 131580 6180 131632 6186
rect 131580 6122 131632 6128
rect 131592 5642 131620 6122
rect 131580 5636 131632 5642
rect 131580 5578 131632 5584
rect 131488 5228 131540 5234
rect 131488 5170 131540 5176
rect 131684 5114 131712 8599
rect 131762 7304 131818 7313
rect 131762 7239 131818 7248
rect 131776 6798 131804 7239
rect 131764 6792 131816 6798
rect 131764 6734 131816 6740
rect 132052 6730 132080 8894
rect 132224 8832 132276 8838
rect 132224 8774 132276 8780
rect 132236 8498 132264 8774
rect 132224 8492 132276 8498
rect 132224 8434 132276 8440
rect 132132 8424 132184 8430
rect 132132 8366 132184 8372
rect 132040 6724 132092 6730
rect 132040 6666 132092 6672
rect 131948 6452 132000 6458
rect 131868 6412 131948 6440
rect 131764 6384 131816 6390
rect 131868 6372 131896 6412
rect 131948 6394 132000 6400
rect 131816 6344 131896 6372
rect 131764 6326 131816 6332
rect 131764 5772 131816 5778
rect 131764 5714 131816 5720
rect 131592 5086 131712 5114
rect 131592 4214 131620 5086
rect 131672 4684 131724 4690
rect 131672 4626 131724 4632
rect 131580 4208 131632 4214
rect 131580 4150 131632 4156
rect 131684 3942 131712 4626
rect 131580 3936 131632 3942
rect 131580 3878 131632 3884
rect 131672 3936 131724 3942
rect 131672 3878 131724 3884
rect 131592 3482 131620 3878
rect 131488 3460 131540 3466
rect 131592 3454 131712 3482
rect 131488 3402 131540 3408
rect 131500 2145 131528 3402
rect 131684 3398 131712 3454
rect 131580 3392 131632 3398
rect 131580 3334 131632 3340
rect 131672 3392 131724 3398
rect 131672 3334 131724 3340
rect 131486 2136 131542 2145
rect 131486 2071 131542 2080
rect 131264 1856 131436 1884
rect 131212 1838 131264 1844
rect 131592 1442 131620 3334
rect 131672 2644 131724 2650
rect 131672 2586 131724 2592
rect 131684 1834 131712 2586
rect 131776 2145 131804 5714
rect 131948 5636 132000 5642
rect 131948 5578 132000 5584
rect 131854 3768 131910 3777
rect 131854 3703 131910 3712
rect 131868 2514 131896 3703
rect 131856 2508 131908 2514
rect 131856 2450 131908 2456
rect 131762 2136 131818 2145
rect 131762 2071 131818 2080
rect 131764 2032 131816 2038
rect 131764 1974 131816 1980
rect 131672 1828 131724 1834
rect 131672 1770 131724 1776
rect 131316 1414 131620 1442
rect 131316 800 131344 1414
rect 131776 800 131804 1974
rect 131120 60 131172 66
rect 131120 2 131172 8
rect 131302 -400 131358 800
rect 131762 -400 131818 800
rect 131960 513 131988 5578
rect 132040 4480 132092 4486
rect 132040 4422 132092 4428
rect 132052 4078 132080 4422
rect 132040 4072 132092 4078
rect 132040 4014 132092 4020
rect 132038 2680 132094 2689
rect 132144 2650 132172 8366
rect 132224 6248 132276 6254
rect 132224 6190 132276 6196
rect 132236 5710 132264 6190
rect 132224 5704 132276 5710
rect 132224 5646 132276 5652
rect 132224 5160 132276 5166
rect 132224 5102 132276 5108
rect 132236 2689 132264 5102
rect 132328 3738 132356 9454
rect 132406 8528 132462 8537
rect 132406 8463 132408 8472
rect 132460 8463 132462 8472
rect 132408 8434 132460 8440
rect 132604 7546 132632 10200
rect 132972 10146 133000 10406
rect 133050 10200 133106 11400
rect 133510 10200 133566 11400
rect 133604 10532 133656 10538
rect 133604 10474 133656 10480
rect 133064 10146 133092 10200
rect 132972 10118 133092 10146
rect 133420 9376 133472 9382
rect 133420 9318 133472 9324
rect 133328 8968 133380 8974
rect 133328 8910 133380 8916
rect 132960 8424 133012 8430
rect 132960 8366 133012 8372
rect 132774 8120 132830 8129
rect 132774 8055 132830 8064
rect 132592 7540 132644 7546
rect 132592 7482 132644 7488
rect 132500 6792 132552 6798
rect 132500 6734 132552 6740
rect 132406 5400 132462 5409
rect 132406 5335 132462 5344
rect 132420 5234 132448 5335
rect 132408 5228 132460 5234
rect 132408 5170 132460 5176
rect 132512 4146 132540 6734
rect 132592 6724 132644 6730
rect 132592 6666 132644 6672
rect 132604 6322 132632 6666
rect 132788 6322 132816 8055
rect 132592 6316 132644 6322
rect 132592 6258 132644 6264
rect 132776 6316 132828 6322
rect 132776 6258 132828 6264
rect 132590 5672 132646 5681
rect 132590 5607 132646 5616
rect 132604 5234 132632 5607
rect 132972 5556 133000 8366
rect 133236 7948 133288 7954
rect 133236 7890 133288 7896
rect 133052 7336 133104 7342
rect 133052 7278 133104 7284
rect 133144 7336 133196 7342
rect 133144 7278 133196 7284
rect 132880 5528 133000 5556
rect 133064 5545 133092 7278
rect 133156 7206 133184 7278
rect 133144 7200 133196 7206
rect 133144 7142 133196 7148
rect 133144 5772 133196 5778
rect 133144 5714 133196 5720
rect 133050 5536 133106 5545
rect 132592 5228 132644 5234
rect 132592 5170 132644 5176
rect 132592 5024 132644 5030
rect 132592 4966 132644 4972
rect 132684 5024 132736 5030
rect 132684 4966 132736 4972
rect 132500 4140 132552 4146
rect 132500 4082 132552 4088
rect 132408 4072 132460 4078
rect 132408 4014 132460 4020
rect 132316 3732 132368 3738
rect 132316 3674 132368 3680
rect 132420 3670 132448 4014
rect 132408 3664 132460 3670
rect 132408 3606 132460 3612
rect 132498 3496 132554 3505
rect 132498 3431 132554 3440
rect 132512 3126 132540 3431
rect 132500 3120 132552 3126
rect 132500 3062 132552 3068
rect 132222 2680 132278 2689
rect 132038 2615 132094 2624
rect 132132 2644 132184 2650
rect 132052 1193 132080 2615
rect 132604 2650 132632 4966
rect 132696 4865 132724 4966
rect 132682 4856 132738 4865
rect 132682 4791 132738 4800
rect 132222 2615 132278 2624
rect 132592 2644 132644 2650
rect 132132 2586 132184 2592
rect 132592 2586 132644 2592
rect 132224 2576 132276 2582
rect 132224 2518 132276 2524
rect 132316 2576 132368 2582
rect 132316 2518 132368 2524
rect 132038 1184 132094 1193
rect 132038 1119 132094 1128
rect 132236 800 132264 2518
rect 132328 1873 132356 2518
rect 132880 2106 132908 5528
rect 133050 5471 133106 5480
rect 132958 4856 133014 4865
rect 132958 4791 133014 4800
rect 132972 4321 133000 4791
rect 132958 4312 133014 4321
rect 132958 4247 133014 4256
rect 133156 3754 133184 5714
rect 133064 3726 133184 3754
rect 133064 3670 133092 3726
rect 133052 3664 133104 3670
rect 133052 3606 133104 3612
rect 133144 3596 133196 3602
rect 133144 3538 133196 3544
rect 132868 2100 132920 2106
rect 132868 2042 132920 2048
rect 132314 1864 132370 1873
rect 132314 1799 132370 1808
rect 132408 1420 132460 1426
rect 132408 1362 132460 1368
rect 132420 814 132448 1362
rect 133052 944 133104 950
rect 133052 886 133104 892
rect 132500 876 132552 882
rect 132552 836 132632 864
rect 132500 818 132552 824
rect 132408 808 132460 814
rect 131946 504 132002 513
rect 131946 439 132002 448
rect 132222 -400 132278 800
rect 132604 800 132632 836
rect 133064 800 133092 886
rect 132408 750 132460 756
rect 132590 -400 132646 800
rect 132868 128 132920 134
rect 132866 96 132868 105
rect 132920 96 132922 105
rect 132866 31 132922 40
rect 133050 -400 133106 800
rect 133156 134 133184 3538
rect 133248 1426 133276 7890
rect 133340 6882 133368 8910
rect 133432 8401 133460 9318
rect 133418 8392 133474 8401
rect 133418 8327 133474 8336
rect 133524 7818 133552 10200
rect 133616 9382 133644 10474
rect 133970 10200 134026 11400
rect 134338 10200 134394 11400
rect 134798 10200 134854 11400
rect 135258 10200 135314 11400
rect 135718 10200 135774 11400
rect 136086 10200 136142 11400
rect 136546 10200 136602 11400
rect 137006 10200 137062 11400
rect 137374 10200 137430 11400
rect 137834 10200 137890 11400
rect 138294 10200 138350 11400
rect 138754 10200 138810 11400
rect 139122 10200 139178 11400
rect 139582 10200 139638 11400
rect 140042 10200 140098 11400
rect 140502 10200 140558 11400
rect 140870 10200 140926 11400
rect 140964 10260 141016 10266
rect 140964 10202 141016 10208
rect 133604 9376 133656 9382
rect 133604 9318 133656 9324
rect 133984 8378 134012 10200
rect 134352 8945 134380 10200
rect 134812 9722 134840 10200
rect 134800 9716 134852 9722
rect 134800 9658 134852 9664
rect 134524 9580 134576 9586
rect 134524 9522 134576 9528
rect 134536 9042 134564 9522
rect 134524 9036 134576 9042
rect 134524 8978 134576 8984
rect 135076 9036 135128 9042
rect 135076 8978 135128 8984
rect 134338 8936 134394 8945
rect 134338 8871 134394 8880
rect 134522 8800 134578 8809
rect 134522 8735 134578 8744
rect 133800 8350 134012 8378
rect 133800 8294 133828 8350
rect 133788 8288 133840 8294
rect 133880 8288 133932 8294
rect 133788 8230 133840 8236
rect 133878 8256 133880 8265
rect 133932 8256 133934 8265
rect 133878 8191 133934 8200
rect 134062 8256 134118 8265
rect 134062 8191 134118 8200
rect 134076 7857 134104 8191
rect 134340 7948 134392 7954
rect 134536 7936 134564 8735
rect 134982 8392 135038 8401
rect 134982 8327 135038 8336
rect 134996 8129 135024 8327
rect 134982 8120 135038 8129
rect 134982 8055 135038 8064
rect 134536 7908 134840 7936
rect 134340 7890 134392 7896
rect 134062 7848 134118 7857
rect 133512 7812 133564 7818
rect 133512 7754 133564 7760
rect 133604 7812 133656 7818
rect 134062 7783 134118 7792
rect 133604 7754 133656 7760
rect 133340 6854 133460 6882
rect 133328 6792 133380 6798
rect 133328 6734 133380 6740
rect 133340 6633 133368 6734
rect 133326 6624 133382 6633
rect 133326 6559 133382 6568
rect 133432 6202 133460 6854
rect 133510 6624 133566 6633
rect 133510 6559 133566 6568
rect 133524 6254 133552 6559
rect 133616 6322 133644 7754
rect 133970 7576 134026 7585
rect 134154 7576 134210 7585
rect 133970 7511 133972 7520
rect 134024 7511 134026 7520
rect 134076 7534 134154 7562
rect 133972 7482 134024 7488
rect 134076 7426 134104 7534
rect 134154 7511 134210 7520
rect 133984 7398 134104 7426
rect 133880 7268 133932 7274
rect 133880 7210 133932 7216
rect 133696 7200 133748 7206
rect 133696 7142 133748 7148
rect 133788 7200 133840 7206
rect 133788 7142 133840 7148
rect 133604 6316 133656 6322
rect 133604 6258 133656 6264
rect 133340 6174 133460 6202
rect 133512 6248 133564 6254
rect 133512 6190 133564 6196
rect 133340 5352 133368 6174
rect 133604 6112 133656 6118
rect 133604 6054 133656 6060
rect 133616 5914 133644 6054
rect 133512 5908 133564 5914
rect 133512 5850 133564 5856
rect 133604 5908 133656 5914
rect 133604 5850 133656 5856
rect 133340 5324 133460 5352
rect 133328 5228 133380 5234
rect 133328 5170 133380 5176
rect 133340 4457 133368 5170
rect 133326 4448 133382 4457
rect 133326 4383 133382 4392
rect 133326 3904 133382 3913
rect 133326 3839 133382 3848
rect 133340 3641 133368 3839
rect 133326 3632 133382 3641
rect 133326 3567 133382 3576
rect 133432 2446 133460 5324
rect 133524 5234 133552 5850
rect 133604 5772 133656 5778
rect 133604 5714 133656 5720
rect 133512 5228 133564 5234
rect 133512 5170 133564 5176
rect 133616 5030 133644 5714
rect 133604 5024 133656 5030
rect 133604 4966 133656 4972
rect 133512 4684 133564 4690
rect 133512 4626 133564 4632
rect 133524 4554 133552 4626
rect 133512 4548 133564 4554
rect 133512 4490 133564 4496
rect 133708 4146 133736 7142
rect 133800 7041 133828 7142
rect 133786 7032 133842 7041
rect 133786 6967 133842 6976
rect 133892 6304 133920 7210
rect 133984 7177 134012 7398
rect 133970 7168 134026 7177
rect 133970 7103 134026 7112
rect 134154 7168 134210 7177
rect 134154 7103 134210 7112
rect 134064 6860 134116 6866
rect 134064 6802 134116 6808
rect 133972 6316 134024 6322
rect 133892 6276 133972 6304
rect 133972 6258 134024 6264
rect 133972 6180 134024 6186
rect 133892 6140 133972 6168
rect 133788 5908 133840 5914
rect 133788 5850 133840 5856
rect 133800 5030 133828 5850
rect 133788 5024 133840 5030
rect 133788 4966 133840 4972
rect 133696 4140 133748 4146
rect 133696 4082 133748 4088
rect 133696 4004 133748 4010
rect 133696 3946 133748 3952
rect 133602 3904 133658 3913
rect 133602 3839 133658 3848
rect 133510 3088 133566 3097
rect 133616 3058 133644 3839
rect 133708 3670 133736 3946
rect 133696 3664 133748 3670
rect 133696 3606 133748 3612
rect 133788 3596 133840 3602
rect 133788 3538 133840 3544
rect 133800 3398 133828 3538
rect 133696 3392 133748 3398
rect 133696 3334 133748 3340
rect 133788 3392 133840 3398
rect 133788 3334 133840 3340
rect 133708 3097 133736 3334
rect 133694 3088 133750 3097
rect 133510 3023 133566 3032
rect 133604 3052 133656 3058
rect 133524 2825 133552 3023
rect 133694 3023 133750 3032
rect 133604 2994 133656 3000
rect 133892 2990 133920 6140
rect 133972 6122 134024 6128
rect 134076 5914 134104 6802
rect 134064 5908 134116 5914
rect 134064 5850 134116 5856
rect 134168 5760 134196 7103
rect 134352 6866 134380 7890
rect 134614 7848 134670 7857
rect 134432 7812 134484 7818
rect 134614 7783 134616 7792
rect 134432 7754 134484 7760
rect 134668 7783 134670 7792
rect 134708 7812 134760 7818
rect 134616 7754 134668 7760
rect 134708 7754 134760 7760
rect 134444 6866 134472 7754
rect 134720 7478 134748 7754
rect 134708 7472 134760 7478
rect 134708 7414 134760 7420
rect 134616 7336 134668 7342
rect 134616 7278 134668 7284
rect 134628 7041 134656 7278
rect 134614 7032 134670 7041
rect 134614 6967 134670 6976
rect 134340 6860 134392 6866
rect 134340 6802 134392 6808
rect 134432 6860 134484 6866
rect 134432 6802 134484 6808
rect 134430 6352 134486 6361
rect 134430 6287 134486 6296
rect 134444 6254 134472 6287
rect 134432 6248 134484 6254
rect 134432 6190 134484 6196
rect 134708 6112 134760 6118
rect 134708 6054 134760 6060
rect 134614 5944 134670 5953
rect 134614 5879 134670 5888
rect 134628 5778 134656 5879
rect 134076 5732 134196 5760
rect 134616 5772 134668 5778
rect 133970 5264 134026 5273
rect 133970 5199 133972 5208
rect 134024 5199 134026 5208
rect 133972 5170 134024 5176
rect 133972 4276 134024 4282
rect 133972 4218 134024 4224
rect 133880 2984 133932 2990
rect 133880 2926 133932 2932
rect 133510 2816 133566 2825
rect 133510 2751 133566 2760
rect 133788 2644 133840 2650
rect 133788 2586 133840 2592
rect 133512 2508 133564 2514
rect 133512 2450 133564 2456
rect 133420 2440 133472 2446
rect 133420 2382 133472 2388
rect 133236 1420 133288 1426
rect 133236 1362 133288 1368
rect 133420 1420 133472 1426
rect 133420 1362 133472 1368
rect 133432 1290 133460 1362
rect 133420 1284 133472 1290
rect 133420 1226 133472 1232
rect 133524 800 133552 2450
rect 133696 1896 133748 1902
rect 133696 1838 133748 1844
rect 133708 1222 133736 1838
rect 133696 1216 133748 1222
rect 133696 1158 133748 1164
rect 133800 1018 133828 2586
rect 133984 2106 134012 4218
rect 134076 3720 134104 5732
rect 134616 5714 134668 5720
rect 134156 5636 134208 5642
rect 134156 5578 134208 5584
rect 134616 5636 134668 5642
rect 134616 5578 134668 5584
rect 134168 3890 134196 5578
rect 134628 5030 134656 5578
rect 134340 5024 134392 5030
rect 134340 4966 134392 4972
rect 134524 5024 134576 5030
rect 134524 4966 134576 4972
rect 134616 5024 134668 5030
rect 134616 4966 134668 4972
rect 134352 4690 134380 4966
rect 134340 4684 134392 4690
rect 134340 4626 134392 4632
rect 134248 4140 134300 4146
rect 134248 4082 134300 4088
rect 134260 4010 134288 4082
rect 134248 4004 134300 4010
rect 134248 3946 134300 3952
rect 134340 3936 134392 3942
rect 134168 3862 134288 3890
rect 134340 3878 134392 3884
rect 134076 3692 134196 3720
rect 134064 3596 134116 3602
rect 134064 3538 134116 3544
rect 134076 3466 134104 3538
rect 134064 3460 134116 3466
rect 134064 3402 134116 3408
rect 134064 3052 134116 3058
rect 134064 2994 134116 3000
rect 134076 2514 134104 2994
rect 134064 2508 134116 2514
rect 134064 2450 134116 2456
rect 133972 2100 134024 2106
rect 133972 2042 134024 2048
rect 134064 2100 134116 2106
rect 134064 2042 134116 2048
rect 133880 1896 133932 1902
rect 133932 1856 134012 1884
rect 133880 1838 133932 1844
rect 133788 1012 133840 1018
rect 133788 954 133840 960
rect 133984 800 134012 1856
rect 134076 1426 134104 2042
rect 134168 1766 134196 3692
rect 134260 1834 134288 3862
rect 134248 1828 134300 1834
rect 134248 1770 134300 1776
rect 134156 1760 134208 1766
rect 134156 1702 134208 1708
rect 134064 1420 134116 1426
rect 134064 1362 134116 1368
rect 134352 800 134380 3878
rect 134536 3602 134564 4966
rect 134720 4486 134748 6054
rect 134812 5710 134840 7908
rect 135088 7154 135116 8978
rect 135168 8492 135220 8498
rect 135168 8434 135220 8440
rect 135180 8129 135208 8434
rect 135166 8120 135222 8129
rect 135166 8055 135222 8064
rect 135168 7472 135220 7478
rect 135168 7414 135220 7420
rect 134904 7126 135116 7154
rect 134904 6372 134932 7126
rect 134982 7032 135038 7041
rect 135180 7018 135208 7414
rect 135038 6990 135208 7018
rect 134982 6967 135038 6976
rect 135272 6798 135300 10200
rect 135444 9988 135496 9994
rect 135444 9930 135496 9936
rect 135352 7268 135404 7274
rect 135352 7210 135404 7216
rect 135260 6792 135312 6798
rect 134982 6760 135038 6769
rect 135260 6734 135312 6740
rect 134982 6695 135038 6704
rect 134996 6497 135024 6695
rect 134982 6488 135038 6497
rect 134982 6423 135038 6432
rect 134904 6344 135116 6372
rect 134984 6248 135036 6254
rect 134984 6190 135036 6196
rect 134996 5953 135024 6190
rect 134982 5944 135038 5953
rect 134982 5879 135038 5888
rect 134892 5772 134944 5778
rect 134892 5714 134944 5720
rect 134800 5704 134852 5710
rect 134800 5646 134852 5652
rect 134708 4480 134760 4486
rect 134708 4422 134760 4428
rect 134616 4072 134668 4078
rect 134616 4014 134668 4020
rect 134524 3596 134576 3602
rect 134524 3538 134576 3544
rect 134432 2984 134484 2990
rect 134432 2926 134484 2932
rect 134444 1873 134472 2926
rect 134628 2446 134656 4014
rect 134708 3936 134760 3942
rect 134708 3878 134760 3884
rect 134798 3904 134854 3913
rect 134720 3194 134748 3878
rect 134798 3839 134854 3848
rect 134812 3398 134840 3839
rect 134800 3392 134852 3398
rect 134800 3334 134852 3340
rect 134708 3188 134760 3194
rect 134708 3130 134760 3136
rect 134800 2644 134852 2650
rect 134800 2586 134852 2592
rect 134616 2440 134668 2446
rect 134616 2382 134668 2388
rect 134812 1902 134840 2586
rect 134616 1896 134668 1902
rect 134430 1864 134486 1873
rect 134616 1838 134668 1844
rect 134800 1896 134852 1902
rect 134800 1838 134852 1844
rect 134430 1799 134486 1808
rect 134628 1766 134656 1838
rect 134616 1760 134668 1766
rect 134616 1702 134668 1708
rect 134904 1018 134932 5714
rect 135088 5352 135116 6344
rect 134996 5324 135116 5352
rect 134996 4298 135024 5324
rect 135166 5264 135222 5273
rect 135088 5234 135166 5250
rect 135076 5228 135166 5234
rect 135128 5222 135166 5228
rect 135364 5234 135392 7210
rect 135166 5199 135222 5208
rect 135352 5228 135404 5234
rect 135076 5170 135128 5176
rect 135352 5170 135404 5176
rect 135350 4448 135406 4457
rect 135350 4383 135406 4392
rect 134996 4270 135116 4298
rect 134984 4072 135036 4078
rect 134984 4014 135036 4020
rect 134996 1358 135024 4014
rect 135088 3194 135116 4270
rect 135076 3188 135128 3194
rect 135076 3130 135128 3136
rect 135364 1902 135392 4383
rect 135456 4010 135484 9930
rect 135732 9466 135760 10200
rect 135640 9438 135760 9466
rect 135640 8673 135668 9438
rect 135720 9376 135772 9382
rect 135720 9318 135772 9324
rect 135626 8664 135682 8673
rect 135626 8599 135682 8608
rect 135732 8566 135760 9318
rect 135720 8560 135772 8566
rect 135720 8502 135772 8508
rect 136100 8498 136128 10200
rect 136180 9716 136232 9722
rect 136180 9658 136232 9664
rect 135536 8492 135588 8498
rect 135536 8434 135588 8440
rect 136088 8492 136140 8498
rect 136088 8434 136140 8440
rect 135548 6866 135576 8434
rect 135996 8424 136048 8430
rect 135996 8366 136048 8372
rect 135812 7336 135864 7342
rect 135812 7278 135864 7284
rect 135626 7032 135682 7041
rect 135626 6967 135682 6976
rect 135536 6860 135588 6866
rect 135536 6802 135588 6808
rect 135640 6798 135668 6967
rect 135720 6860 135772 6866
rect 135720 6802 135772 6808
rect 135628 6792 135680 6798
rect 135628 6734 135680 6740
rect 135536 6180 135588 6186
rect 135536 6122 135588 6128
rect 135548 5642 135576 6122
rect 135536 5636 135588 5642
rect 135536 5578 135588 5584
rect 135732 4264 135760 6802
rect 135824 5681 135852 7278
rect 135904 6316 135956 6322
rect 135904 6258 135956 6264
rect 135810 5672 135866 5681
rect 135916 5642 135944 6258
rect 135810 5607 135866 5616
rect 135904 5636 135956 5642
rect 135904 5578 135956 5584
rect 135548 4236 135760 4264
rect 135444 4004 135496 4010
rect 135444 3946 135496 3952
rect 135444 3392 135496 3398
rect 135444 3334 135496 3340
rect 135352 1896 135404 1902
rect 135352 1838 135404 1844
rect 135456 1494 135484 3334
rect 135548 2378 135576 4236
rect 135720 4140 135772 4146
rect 135720 4082 135772 4088
rect 135628 3188 135680 3194
rect 135628 3130 135680 3136
rect 135640 2961 135668 3130
rect 135626 2952 135682 2961
rect 135626 2887 135682 2896
rect 135628 2440 135680 2446
rect 135628 2382 135680 2388
rect 135536 2372 135588 2378
rect 135536 2314 135588 2320
rect 135640 1494 135668 2382
rect 135444 1488 135496 1494
rect 135444 1430 135496 1436
rect 135628 1488 135680 1494
rect 135628 1430 135680 1436
rect 135260 1420 135312 1426
rect 135260 1362 135312 1368
rect 134984 1352 135036 1358
rect 134984 1294 135036 1300
rect 134800 1012 134852 1018
rect 134800 954 134852 960
rect 134892 1012 134944 1018
rect 134892 954 134944 960
rect 134812 800 134840 954
rect 135272 800 135300 1362
rect 135732 800 135760 4082
rect 136008 2990 136036 8366
rect 136192 5574 136220 9658
rect 136272 9648 136324 9654
rect 136272 9590 136324 9596
rect 136180 5568 136232 5574
rect 136180 5510 136232 5516
rect 136180 5228 136232 5234
rect 136180 5170 136232 5176
rect 136088 4684 136140 4690
rect 136088 4626 136140 4632
rect 136100 4282 136128 4626
rect 136192 4486 136220 5170
rect 136180 4480 136232 4486
rect 136180 4422 136232 4428
rect 136088 4276 136140 4282
rect 136088 4218 136140 4224
rect 136284 3126 136312 9590
rect 136364 9444 136416 9450
rect 136364 9386 136416 9392
rect 136376 8634 136404 9386
rect 136364 8628 136416 8634
rect 136364 8570 136416 8576
rect 136560 6254 136588 10200
rect 136916 10056 136968 10062
rect 136916 9998 136968 10004
rect 136928 9042 136956 9998
rect 136916 9036 136968 9042
rect 136916 8978 136968 8984
rect 136730 7712 136786 7721
rect 136730 7647 136786 7656
rect 136744 7410 136772 7647
rect 137020 7426 137048 10200
rect 137388 7834 137416 10200
rect 137848 8974 137876 10200
rect 137926 10160 137982 10169
rect 137926 10095 137982 10104
rect 137836 8968 137888 8974
rect 137836 8910 137888 8916
rect 137940 8498 137968 10095
rect 138204 8628 138256 8634
rect 138204 8570 138256 8576
rect 137928 8492 137980 8498
rect 137928 8434 137980 8440
rect 138018 8256 138074 8265
rect 138074 8214 138152 8242
rect 138018 8191 138074 8200
rect 137836 8016 137888 8022
rect 137834 7984 137836 7993
rect 137888 7984 137890 7993
rect 138018 7984 138074 7993
rect 137834 7919 137890 7928
rect 137940 7942 138018 7970
rect 137940 7857 137968 7942
rect 138018 7919 138074 7928
rect 138124 7857 138152 8214
rect 137204 7806 137416 7834
rect 137926 7848 137982 7857
rect 137204 7478 137232 7806
rect 137926 7783 137982 7792
rect 138110 7848 138166 7857
rect 138110 7783 138166 7792
rect 137374 7712 137430 7721
rect 137374 7647 137430 7656
rect 137388 7478 137416 7647
rect 136732 7404 136784 7410
rect 136732 7346 136784 7352
rect 136836 7398 137048 7426
rect 137192 7472 137244 7478
rect 137192 7414 137244 7420
rect 137376 7472 137428 7478
rect 137376 7414 137428 7420
rect 137468 7472 137520 7478
rect 137468 7414 137520 7420
rect 136640 6792 136692 6798
rect 136640 6734 136692 6740
rect 136548 6248 136600 6254
rect 136548 6190 136600 6196
rect 136652 5778 136680 6734
rect 136732 6248 136784 6254
rect 136732 6190 136784 6196
rect 136640 5772 136692 5778
rect 136640 5714 136692 5720
rect 136638 4584 136694 4593
rect 136364 4548 136416 4554
rect 136416 4508 136496 4536
rect 136638 4519 136640 4528
rect 136364 4490 136416 4496
rect 136364 3596 136416 3602
rect 136364 3538 136416 3544
rect 136272 3120 136324 3126
rect 136272 3062 136324 3068
rect 135904 2984 135956 2990
rect 135902 2952 135904 2961
rect 135996 2984 136048 2990
rect 135956 2952 135958 2961
rect 135996 2926 136048 2932
rect 135902 2887 135958 2896
rect 135812 2508 135864 2514
rect 136180 2508 136232 2514
rect 135864 2468 136180 2496
rect 135812 2450 135864 2456
rect 136180 2450 136232 2456
rect 135812 2372 135864 2378
rect 135864 2332 136036 2360
rect 135812 2314 135864 2320
rect 136008 1902 136036 2332
rect 135812 1896 135864 1902
rect 135812 1838 135864 1844
rect 135996 1896 136048 1902
rect 135996 1838 136048 1844
rect 135824 1748 135852 1838
rect 136180 1760 136232 1766
rect 135824 1720 136128 1748
rect 136100 800 136128 1720
rect 136180 1702 136232 1708
rect 136192 1494 136220 1702
rect 136376 1494 136404 3538
rect 136180 1488 136232 1494
rect 136180 1430 136232 1436
rect 136364 1488 136416 1494
rect 136364 1430 136416 1436
rect 136468 898 136496 4508
rect 136692 4519 136694 4528
rect 136640 4490 136692 4496
rect 136548 4276 136600 4282
rect 136548 4218 136600 4224
rect 136560 4146 136588 4218
rect 136548 4140 136600 4146
rect 136548 4082 136600 4088
rect 136640 4140 136692 4146
rect 136640 4082 136692 4088
rect 136652 4049 136680 4082
rect 136638 4040 136694 4049
rect 136548 4004 136600 4010
rect 136638 3975 136694 3984
rect 136548 3946 136600 3952
rect 136560 3534 136588 3946
rect 136548 3528 136600 3534
rect 136548 3470 136600 3476
rect 136640 2372 136692 2378
rect 136640 2314 136692 2320
rect 136652 1766 136680 2314
rect 136744 2106 136772 6190
rect 136836 5098 136864 7398
rect 137008 7336 137060 7342
rect 137008 7278 137060 7284
rect 137100 7336 137152 7342
rect 137100 7278 137152 7284
rect 137020 7177 137048 7278
rect 137006 7168 137062 7177
rect 137006 7103 137062 7112
rect 136914 5536 136970 5545
rect 136914 5471 136970 5480
rect 136824 5092 136876 5098
rect 136824 5034 136876 5040
rect 136928 4729 136956 5471
rect 137008 5160 137060 5166
rect 137008 5102 137060 5108
rect 136914 4720 136970 4729
rect 136914 4655 136970 4664
rect 136824 4072 136876 4078
rect 136824 4014 136876 4020
rect 136732 2100 136784 2106
rect 136732 2042 136784 2048
rect 136640 1760 136692 1766
rect 136640 1702 136692 1708
rect 136836 1494 136864 4014
rect 136914 3904 136970 3913
rect 136914 3839 136970 3848
rect 136928 3369 136956 3839
rect 137020 3777 137048 5102
rect 137006 3768 137062 3777
rect 137006 3703 137062 3712
rect 137112 3534 137140 7278
rect 137480 7002 137508 7414
rect 137558 7168 137614 7177
rect 137558 7103 137614 7112
rect 137468 6996 137520 7002
rect 137468 6938 137520 6944
rect 137572 6322 137600 7103
rect 137928 6996 137980 7002
rect 137928 6938 137980 6944
rect 137652 6792 137704 6798
rect 137652 6734 137704 6740
rect 137560 6316 137612 6322
rect 137560 6258 137612 6264
rect 137664 5760 137692 6734
rect 137572 5732 137692 5760
rect 137572 5574 137600 5732
rect 137652 5636 137704 5642
rect 137940 5624 137968 6938
rect 137652 5578 137704 5584
rect 137756 5596 137968 5624
rect 137560 5568 137612 5574
rect 137664 5545 137692 5578
rect 137560 5510 137612 5516
rect 137650 5536 137706 5545
rect 137650 5471 137706 5480
rect 137204 5358 137508 5386
rect 137204 5234 137232 5358
rect 137284 5296 137336 5302
rect 137284 5238 137336 5244
rect 137192 5228 137244 5234
rect 137192 5170 137244 5176
rect 137190 4584 137246 4593
rect 137190 4519 137246 4528
rect 137204 4214 137232 4519
rect 137296 4214 137324 5238
rect 137480 5216 137508 5358
rect 137652 5228 137704 5234
rect 137480 5188 137652 5216
rect 137652 5170 137704 5176
rect 137376 5160 137428 5166
rect 137376 5102 137428 5108
rect 137388 4622 137416 5102
rect 137560 4820 137612 4826
rect 137560 4762 137612 4768
rect 137652 4820 137704 4826
rect 137652 4762 137704 4768
rect 137572 4690 137600 4762
rect 137560 4684 137612 4690
rect 137560 4626 137612 4632
rect 137376 4616 137428 4622
rect 137664 4593 137692 4762
rect 137376 4558 137428 4564
rect 137650 4584 137706 4593
rect 137650 4519 137706 4528
rect 137756 4486 137784 5596
rect 137926 5536 137982 5545
rect 137926 5471 137982 5480
rect 137940 5386 137968 5471
rect 137940 5358 138152 5386
rect 138216 5370 138244 8570
rect 138308 6458 138336 10200
rect 138388 9036 138440 9042
rect 138388 8978 138440 8984
rect 138296 6452 138348 6458
rect 138296 6394 138348 6400
rect 138294 5400 138350 5409
rect 138124 5250 138152 5358
rect 138204 5364 138256 5370
rect 138294 5335 138350 5344
rect 138204 5306 138256 5312
rect 138308 5250 138336 5335
rect 138124 5222 138336 5250
rect 138296 4752 138348 4758
rect 138296 4694 138348 4700
rect 137940 4644 138152 4672
rect 137744 4480 137796 4486
rect 137744 4422 137796 4428
rect 137836 4480 137888 4486
rect 137836 4422 137888 4428
rect 137848 4282 137876 4422
rect 137836 4276 137888 4282
rect 137836 4218 137888 4224
rect 137192 4208 137244 4214
rect 137192 4150 137244 4156
rect 137284 4208 137336 4214
rect 137284 4150 137336 4156
rect 137940 4128 137968 4644
rect 138018 4584 138074 4593
rect 138018 4519 138074 4528
rect 137848 4100 137968 4128
rect 137744 4004 137796 4010
rect 137744 3946 137796 3952
rect 137376 3936 137428 3942
rect 137376 3878 137428 3884
rect 137100 3528 137152 3534
rect 137100 3470 137152 3476
rect 137388 3466 137416 3878
rect 137756 3720 137784 3946
rect 137848 3738 137876 4100
rect 138032 3992 138060 4519
rect 138124 4078 138152 4644
rect 138204 4208 138256 4214
rect 138204 4150 138256 4156
rect 138112 4072 138164 4078
rect 138112 4014 138164 4020
rect 137940 3964 138060 3992
rect 137572 3692 137784 3720
rect 137836 3732 137888 3738
rect 137468 3596 137520 3602
rect 137468 3538 137520 3544
rect 137284 3460 137336 3466
rect 137284 3402 137336 3408
rect 137376 3460 137428 3466
rect 137376 3402 137428 3408
rect 136914 3360 136970 3369
rect 136914 3295 136970 3304
rect 137190 3360 137246 3369
rect 137190 3295 137246 3304
rect 137008 3120 137060 3126
rect 137008 3062 137060 3068
rect 137020 2922 137048 3062
rect 137204 3058 137232 3295
rect 137192 3052 137244 3058
rect 137192 2994 137244 3000
rect 137008 2916 137060 2922
rect 137008 2858 137060 2864
rect 137296 2836 137324 3402
rect 137480 3398 137508 3538
rect 137468 3392 137520 3398
rect 137466 3360 137468 3369
rect 137520 3360 137522 3369
rect 137466 3295 137522 3304
rect 137466 3088 137522 3097
rect 137466 3023 137522 3032
rect 137296 2808 137416 2836
rect 137192 2304 137244 2310
rect 137192 2246 137244 2252
rect 137098 1864 137154 1873
rect 137098 1799 137154 1808
rect 137112 1766 137140 1799
rect 137100 1760 137152 1766
rect 137100 1702 137152 1708
rect 136824 1488 136876 1494
rect 136824 1430 136876 1436
rect 137204 1426 137232 2246
rect 137284 1896 137336 1902
rect 137282 1864 137284 1873
rect 137336 1864 137338 1873
rect 137282 1799 137338 1808
rect 137008 1420 137060 1426
rect 137008 1362 137060 1368
rect 137192 1420 137244 1426
rect 137192 1362 137244 1368
rect 136468 870 136588 898
rect 136560 800 136588 870
rect 137020 800 137048 1362
rect 137100 1352 137152 1358
rect 137100 1294 137152 1300
rect 137284 1352 137336 1358
rect 137284 1294 137336 1300
rect 137112 814 137140 1294
rect 137296 1018 137324 1294
rect 137284 1012 137336 1018
rect 137284 954 137336 960
rect 137100 808 137152 814
rect 133144 128 133196 134
rect 133144 70 133196 76
rect 133510 -400 133566 800
rect 133970 -400 134026 800
rect 134338 -400 134394 800
rect 134798 -400 134854 800
rect 135258 -400 135314 800
rect 135718 -400 135774 800
rect 136086 -400 136142 800
rect 136546 -400 136602 800
rect 137006 -400 137062 800
rect 137388 800 137416 2808
rect 137480 1544 137508 3023
rect 137572 2106 137600 3692
rect 137836 3674 137888 3680
rect 137940 3670 137968 3964
rect 138216 3890 138244 4150
rect 138032 3862 138244 3890
rect 137928 3664 137980 3670
rect 137928 3606 137980 3612
rect 137836 3528 137888 3534
rect 137836 3470 137888 3476
rect 137848 2514 137876 3470
rect 137928 3120 137980 3126
rect 137928 3062 137980 3068
rect 137940 2854 137968 3062
rect 138032 3058 138060 3862
rect 138110 3768 138166 3777
rect 138110 3703 138166 3712
rect 138204 3732 138256 3738
rect 138124 3194 138152 3703
rect 138204 3674 138256 3680
rect 138112 3188 138164 3194
rect 138112 3130 138164 3136
rect 138020 3052 138072 3058
rect 138020 2994 138072 3000
rect 138216 2990 138244 3674
rect 138204 2984 138256 2990
rect 138204 2926 138256 2932
rect 137928 2848 137980 2854
rect 137928 2790 137980 2796
rect 138202 2680 138258 2689
rect 138202 2615 138258 2624
rect 137836 2508 137888 2514
rect 137836 2450 137888 2456
rect 138020 2508 138072 2514
rect 138020 2450 138072 2456
rect 137744 2440 137796 2446
rect 137796 2388 137968 2394
rect 137744 2382 137968 2388
rect 137756 2366 137968 2382
rect 137652 2304 137704 2310
rect 137652 2246 137704 2252
rect 137664 2106 137692 2246
rect 137742 2136 137798 2145
rect 137560 2100 137612 2106
rect 137560 2042 137612 2048
rect 137652 2100 137704 2106
rect 137798 2094 137876 2122
rect 137742 2071 137798 2080
rect 137652 2042 137704 2048
rect 137848 2038 137876 2094
rect 137744 2032 137796 2038
rect 137744 1974 137796 1980
rect 137836 2032 137888 2038
rect 137836 1974 137888 1980
rect 137756 1873 137784 1974
rect 137558 1864 137614 1873
rect 137742 1864 137798 1873
rect 137614 1822 137692 1850
rect 137558 1799 137614 1808
rect 137664 1578 137692 1822
rect 137742 1799 137798 1808
rect 137940 1714 137968 2366
rect 138032 1834 138060 2450
rect 138216 2378 138244 2615
rect 138308 2394 138336 4694
rect 138400 3670 138428 8978
rect 138768 7342 138796 10200
rect 139136 9722 139164 10200
rect 139124 9716 139176 9722
rect 139124 9658 139176 9664
rect 139124 9376 139176 9382
rect 139124 9318 139176 9324
rect 139136 8838 139164 9318
rect 139124 8832 139176 8838
rect 139124 8774 139176 8780
rect 139124 8424 139176 8430
rect 139124 8366 139176 8372
rect 138756 7336 138808 7342
rect 138756 7278 138808 7284
rect 139032 6792 139084 6798
rect 139032 6734 139084 6740
rect 138480 6724 138532 6730
rect 138480 6666 138532 6672
rect 138492 6254 138520 6666
rect 138662 6352 138718 6361
rect 138662 6287 138718 6296
rect 138480 6248 138532 6254
rect 138480 6190 138532 6196
rect 138676 5953 138704 6287
rect 138662 5944 138718 5953
rect 138662 5879 138718 5888
rect 138756 5704 138808 5710
rect 138756 5646 138808 5652
rect 138570 5128 138626 5137
rect 138570 5063 138626 5072
rect 138478 3768 138534 3777
rect 138478 3703 138534 3712
rect 138388 3664 138440 3670
rect 138388 3606 138440 3612
rect 138388 3392 138440 3398
rect 138388 3334 138440 3340
rect 138400 2514 138428 3334
rect 138492 2854 138520 3703
rect 138584 2854 138612 5063
rect 138768 4826 138796 5646
rect 138848 5092 138900 5098
rect 138848 5034 138900 5040
rect 138756 4820 138808 4826
rect 138756 4762 138808 4768
rect 138664 4004 138716 4010
rect 138664 3946 138716 3952
rect 138676 3670 138704 3946
rect 138664 3664 138716 3670
rect 138664 3606 138716 3612
rect 138756 3392 138808 3398
rect 138756 3334 138808 3340
rect 138768 3194 138796 3334
rect 138756 3188 138808 3194
rect 138756 3130 138808 3136
rect 138664 2916 138716 2922
rect 138664 2858 138716 2864
rect 138480 2848 138532 2854
rect 138480 2790 138532 2796
rect 138572 2848 138624 2854
rect 138572 2790 138624 2796
rect 138676 2650 138704 2858
rect 138664 2644 138716 2650
rect 138664 2586 138716 2592
rect 138756 2644 138808 2650
rect 138860 2632 138888 5034
rect 138940 3936 138992 3942
rect 138940 3878 138992 3884
rect 138952 3534 138980 3878
rect 138940 3528 138992 3534
rect 138940 3470 138992 3476
rect 138940 3392 138992 3398
rect 138940 3334 138992 3340
rect 138808 2604 138888 2632
rect 138756 2586 138808 2592
rect 138388 2508 138440 2514
rect 138388 2450 138440 2456
rect 138204 2372 138256 2378
rect 138308 2366 138704 2394
rect 138204 2314 138256 2320
rect 138124 2106 138612 2122
rect 138124 2100 138624 2106
rect 138124 2094 138572 2100
rect 138020 1828 138072 1834
rect 138020 1770 138072 1776
rect 138124 1766 138152 2094
rect 138572 2042 138624 2048
rect 138204 1964 138256 1970
rect 138676 1952 138704 2366
rect 138204 1906 138256 1912
rect 138492 1924 138704 1952
rect 138112 1760 138164 1766
rect 137940 1686 138060 1714
rect 138216 1737 138244 1906
rect 138296 1760 138348 1766
rect 138112 1702 138164 1708
rect 138202 1728 138258 1737
rect 138032 1578 138060 1686
rect 138296 1702 138348 1708
rect 138202 1663 138258 1672
rect 138308 1578 138336 1702
rect 137664 1550 137968 1578
rect 138032 1550 138336 1578
rect 137480 1516 137600 1544
rect 137572 1057 137600 1516
rect 137940 1494 137968 1550
rect 137836 1488 137888 1494
rect 137836 1430 137888 1436
rect 137928 1488 137980 1494
rect 138492 1476 138520 1924
rect 138848 1828 138900 1834
rect 138848 1770 138900 1776
rect 138860 1494 138888 1770
rect 137928 1430 137980 1436
rect 138308 1448 138520 1476
rect 138848 1488 138900 1494
rect 137558 1048 137614 1057
rect 137558 983 137614 992
rect 137848 800 137876 1430
rect 138308 800 138336 1448
rect 138848 1430 138900 1436
rect 138952 1426 138980 3334
rect 139044 1426 139072 6734
rect 139136 4214 139164 8366
rect 139492 7948 139544 7954
rect 139492 7890 139544 7896
rect 139124 4208 139176 4214
rect 139124 4150 139176 4156
rect 139124 4072 139176 4078
rect 139124 4014 139176 4020
rect 139216 4072 139268 4078
rect 139400 4072 139452 4078
rect 139216 4014 139268 4020
rect 139320 4032 139400 4060
rect 139136 3516 139164 4014
rect 139228 3670 139256 4014
rect 139216 3664 139268 3670
rect 139216 3606 139268 3612
rect 139320 3516 139348 4032
rect 139400 4014 139452 4020
rect 139136 3488 139348 3516
rect 139504 2310 139532 7890
rect 139596 7002 139624 10200
rect 139952 7948 140004 7954
rect 139952 7890 140004 7896
rect 139964 7818 139992 7890
rect 139952 7812 140004 7818
rect 139952 7754 140004 7760
rect 140056 7562 140084 10200
rect 140412 9988 140464 9994
rect 140412 9930 140464 9936
rect 140226 8936 140282 8945
rect 140226 8871 140228 8880
rect 140280 8871 140282 8880
rect 140228 8842 140280 8848
rect 140226 8664 140282 8673
rect 140226 8599 140282 8608
rect 140240 7818 140268 8599
rect 140424 8498 140452 9930
rect 140412 8492 140464 8498
rect 140412 8434 140464 8440
rect 140516 7954 140544 10200
rect 140780 9920 140832 9926
rect 140780 9862 140832 9868
rect 140792 8498 140820 9862
rect 140780 8492 140832 8498
rect 140780 8434 140832 8440
rect 140780 8288 140832 8294
rect 140780 8230 140832 8236
rect 140504 7948 140556 7954
rect 140504 7890 140556 7896
rect 140792 7886 140820 8230
rect 140780 7880 140832 7886
rect 140686 7848 140742 7857
rect 140228 7812 140280 7818
rect 140228 7754 140280 7760
rect 140320 7812 140372 7818
rect 140780 7822 140832 7828
rect 140686 7783 140742 7792
rect 140320 7754 140372 7760
rect 140332 7585 140360 7754
rect 139688 7534 140084 7562
rect 140318 7576 140374 7585
rect 139584 6996 139636 7002
rect 139584 6938 139636 6944
rect 139584 6248 139636 6254
rect 139584 6190 139636 6196
rect 139492 2304 139544 2310
rect 139492 2246 139544 2252
rect 139490 2136 139546 2145
rect 139596 2106 139624 6190
rect 139688 4758 139716 7534
rect 140318 7511 140374 7520
rect 140502 7576 140558 7585
rect 140502 7511 140558 7520
rect 140516 7478 140544 7511
rect 140320 7472 140372 7478
rect 140320 7414 140372 7420
rect 140504 7472 140556 7478
rect 140504 7414 140556 7420
rect 139768 7268 139820 7274
rect 139768 7210 139820 7216
rect 139780 7002 139808 7210
rect 140332 7002 140360 7414
rect 140504 7336 140556 7342
rect 140504 7278 140556 7284
rect 139768 6996 139820 7002
rect 139768 6938 139820 6944
rect 140320 6996 140372 7002
rect 140320 6938 140372 6944
rect 140226 6624 140282 6633
rect 140226 6559 140282 6568
rect 140410 6624 140466 6633
rect 140410 6559 140466 6568
rect 139860 5772 139912 5778
rect 139860 5714 139912 5720
rect 139676 4752 139728 4758
rect 139676 4694 139728 4700
rect 139766 4584 139822 4593
rect 139766 4519 139822 4528
rect 139780 3670 139808 4519
rect 139768 3664 139820 3670
rect 139768 3606 139820 3612
rect 139872 2650 139900 5714
rect 140044 4616 140096 4622
rect 140044 4558 140096 4564
rect 140056 4146 140084 4558
rect 140044 4140 140096 4146
rect 140044 4082 140096 4088
rect 140042 2680 140098 2689
rect 139676 2644 139728 2650
rect 139676 2586 139728 2592
rect 139860 2644 139912 2650
rect 139860 2586 139912 2592
rect 139952 2644 140004 2650
rect 140042 2615 140098 2624
rect 139952 2586 140004 2592
rect 139688 2530 139716 2586
rect 139964 2530 139992 2586
rect 139688 2502 139992 2530
rect 140056 2145 140084 2615
rect 140042 2136 140098 2145
rect 139490 2071 139546 2080
rect 139584 2100 139636 2106
rect 139216 1896 139268 1902
rect 139504 1873 139532 2071
rect 140042 2071 140098 2080
rect 139584 2042 139636 2048
rect 140044 1964 140096 1970
rect 140044 1906 140096 1912
rect 140136 1964 140188 1970
rect 140136 1906 140188 1912
rect 139216 1838 139268 1844
rect 139306 1864 139362 1873
rect 139228 1442 139256 1838
rect 139490 1864 139546 1873
rect 139362 1822 139440 1850
rect 139306 1799 139362 1808
rect 139412 1714 139440 1822
rect 139490 1799 139546 1808
rect 139676 1828 139728 1834
rect 139676 1770 139728 1776
rect 139412 1686 139624 1714
rect 138572 1420 138624 1426
rect 138572 1362 138624 1368
rect 138940 1420 138992 1426
rect 138940 1362 138992 1368
rect 139032 1420 139084 1426
rect 139228 1414 139348 1442
rect 139032 1362 139084 1368
rect 138584 1170 138612 1362
rect 138848 1216 138900 1222
rect 138584 1142 138796 1170
rect 139124 1216 139176 1222
rect 138900 1176 139124 1204
rect 138848 1158 138900 1164
rect 139124 1158 139176 1164
rect 138768 800 138796 1142
rect 139320 1000 139348 1414
rect 139136 972 139348 1000
rect 139136 800 139164 972
rect 139596 800 139624 1686
rect 139688 1426 139716 1770
rect 139676 1420 139728 1426
rect 139676 1362 139728 1368
rect 140056 800 140084 1906
rect 140148 1766 140176 1906
rect 140240 1766 140268 6559
rect 140424 6118 140452 6559
rect 140516 6322 140544 7278
rect 140700 6934 140728 7783
rect 140688 6928 140740 6934
rect 140688 6870 140740 6876
rect 140504 6316 140556 6322
rect 140504 6258 140556 6264
rect 140412 6112 140464 6118
rect 140412 6054 140464 6060
rect 140686 5128 140742 5137
rect 140686 5063 140742 5072
rect 140410 4992 140466 5001
rect 140410 4927 140466 4936
rect 140320 3936 140372 3942
rect 140320 3878 140372 3884
rect 140332 3738 140360 3878
rect 140320 3732 140372 3738
rect 140320 3674 140372 3680
rect 140424 2854 140452 4927
rect 140700 4554 140728 5063
rect 140780 5024 140832 5030
rect 140780 4966 140832 4972
rect 140688 4548 140740 4554
rect 140688 4490 140740 4496
rect 140596 4208 140648 4214
rect 140792 4185 140820 4966
rect 140596 4150 140648 4156
rect 140778 4176 140834 4185
rect 140412 2848 140464 2854
rect 140412 2790 140464 2796
rect 140320 2508 140372 2514
rect 140320 2450 140372 2456
rect 140136 1760 140188 1766
rect 140136 1702 140188 1708
rect 140228 1760 140280 1766
rect 140228 1702 140280 1708
rect 140332 1562 140360 2450
rect 140320 1556 140372 1562
rect 140320 1498 140372 1504
rect 140504 944 140556 950
rect 140504 886 140556 892
rect 140516 800 140544 886
rect 137100 750 137152 756
rect 137374 -400 137430 800
rect 137652 332 137704 338
rect 137652 274 137704 280
rect 137664 105 137692 274
rect 137650 96 137706 105
rect 137650 31 137706 40
rect 137834 -400 137890 800
rect 138294 -400 138350 800
rect 138754 -400 138810 800
rect 139122 -400 139178 800
rect 139582 -400 139638 800
rect 140042 -400 140098 800
rect 140502 -400 140558 800
rect 140608 610 140636 4150
rect 140884 4146 140912 10200
rect 140976 9450 141004 10202
rect 141330 10200 141386 11400
rect 141790 10200 141846 11400
rect 142250 10200 142306 11400
rect 142618 10200 142674 11400
rect 143078 10200 143134 11400
rect 143538 10200 143594 11400
rect 143998 10200 144054 11400
rect 144366 10200 144422 11400
rect 144826 10200 144882 11400
rect 145286 10200 145342 11400
rect 145564 10328 145616 10334
rect 145564 10270 145616 10276
rect 140964 9444 141016 9450
rect 140964 9386 141016 9392
rect 141148 8968 141200 8974
rect 141148 8910 141200 8916
rect 141160 8090 141188 8910
rect 141240 8832 141292 8838
rect 141240 8774 141292 8780
rect 141252 8090 141280 8774
rect 141148 8084 141200 8090
rect 141148 8026 141200 8032
rect 141240 8084 141292 8090
rect 141240 8026 141292 8032
rect 141344 7970 141372 10200
rect 141804 10062 141832 10200
rect 141792 10056 141844 10062
rect 141792 9998 141844 10004
rect 142068 9376 142120 9382
rect 142068 9318 142120 9324
rect 142080 9178 142108 9318
rect 142068 9172 142120 9178
rect 142068 9114 142120 9120
rect 142160 8968 142212 8974
rect 142160 8910 142212 8916
rect 142172 8566 142200 8910
rect 142160 8560 142212 8566
rect 142160 8502 142212 8508
rect 141068 7942 141372 7970
rect 141976 8016 142028 8022
rect 142264 7970 142292 10200
rect 142632 9654 142660 10200
rect 142988 10192 143040 10198
rect 143092 10146 143120 10200
rect 143040 10140 143120 10146
rect 142988 10134 143120 10140
rect 143000 10118 143120 10134
rect 142620 9648 142672 9654
rect 142620 9590 142672 9596
rect 142802 8120 142858 8129
rect 142802 8055 142858 8064
rect 141976 7958 142028 7964
rect 141068 6866 141096 7942
rect 141148 7880 141200 7886
rect 141148 7822 141200 7828
rect 141160 6866 141188 7822
rect 141988 7342 142016 7958
rect 142172 7942 142292 7970
rect 142172 7449 142200 7942
rect 142252 7880 142304 7886
rect 142816 7857 142844 8055
rect 142252 7822 142304 7828
rect 142802 7848 142858 7857
rect 142158 7440 142214 7449
rect 142264 7410 142292 7822
rect 142802 7783 142858 7792
rect 142528 7540 142580 7546
rect 142528 7482 142580 7488
rect 142540 7410 142568 7482
rect 143446 7440 143502 7449
rect 142158 7375 142214 7384
rect 142252 7404 142304 7410
rect 142252 7346 142304 7352
rect 142528 7404 142580 7410
rect 143446 7375 143448 7384
rect 142528 7346 142580 7352
rect 143500 7375 143502 7384
rect 143448 7346 143500 7352
rect 141976 7336 142028 7342
rect 141976 7278 142028 7284
rect 142710 7304 142766 7313
rect 141240 7268 141292 7274
rect 142710 7239 142712 7248
rect 141240 7210 141292 7216
rect 142764 7239 142766 7248
rect 142712 7210 142764 7216
rect 141056 6860 141108 6866
rect 141056 6802 141108 6808
rect 141148 6860 141200 6866
rect 141148 6802 141200 6808
rect 141148 6724 141200 6730
rect 141148 6666 141200 6672
rect 141160 5778 141188 6666
rect 141148 5772 141200 5778
rect 141148 5714 141200 5720
rect 140962 4856 141018 4865
rect 140962 4791 141018 4800
rect 141056 4820 141108 4826
rect 140778 4111 140834 4120
rect 140872 4140 140924 4146
rect 140872 4082 140924 4088
rect 140976 3738 141004 4791
rect 141056 4762 141108 4768
rect 140964 3732 141016 3738
rect 140964 3674 141016 3680
rect 141068 2854 141096 4762
rect 141148 3596 141200 3602
rect 141148 3538 141200 3544
rect 141056 2848 141108 2854
rect 141056 2790 141108 2796
rect 140872 1828 140924 1834
rect 140872 1770 140924 1776
rect 140688 1216 140740 1222
rect 140688 1158 140740 1164
rect 140700 950 140728 1158
rect 140688 944 140740 950
rect 140688 886 140740 892
rect 140884 800 140912 1770
rect 141160 1426 141188 3538
rect 141252 1562 141280 7210
rect 142620 6316 142672 6322
rect 142620 6258 142672 6264
rect 142158 6080 142214 6089
rect 142158 6015 142214 6024
rect 142172 5914 142200 6015
rect 142160 5908 142212 5914
rect 142160 5850 142212 5856
rect 142632 5234 142660 6258
rect 143264 5908 143316 5914
rect 143264 5850 143316 5856
rect 143276 5234 143304 5850
rect 142620 5228 142672 5234
rect 142620 5170 142672 5176
rect 143264 5228 143316 5234
rect 143264 5170 143316 5176
rect 143356 5160 143408 5166
rect 143356 5102 143408 5108
rect 141608 4684 141660 4690
rect 141608 4626 141660 4632
rect 141514 4584 141570 4593
rect 141514 4519 141516 4528
rect 141568 4519 141570 4528
rect 141516 4490 141568 4496
rect 141514 4312 141570 4321
rect 141514 4247 141570 4256
rect 141330 4176 141386 4185
rect 141528 4146 141556 4247
rect 141330 4111 141386 4120
rect 141516 4140 141568 4146
rect 141344 3670 141372 4111
rect 141516 4082 141568 4088
rect 141332 3664 141384 3670
rect 141332 3606 141384 3612
rect 141422 2816 141478 2825
rect 141422 2751 141478 2760
rect 141240 1556 141292 1562
rect 141240 1498 141292 1504
rect 141436 1442 141464 2751
rect 141620 2689 141648 4626
rect 142436 4616 142488 4622
rect 142436 4558 142488 4564
rect 142448 4457 142476 4558
rect 142434 4448 142490 4457
rect 142434 4383 142490 4392
rect 142250 3768 142306 3777
rect 142250 3703 142306 3712
rect 142264 3602 142292 3703
rect 142160 3596 142212 3602
rect 142160 3538 142212 3544
rect 142252 3596 142304 3602
rect 142252 3538 142304 3544
rect 142172 3194 142200 3538
rect 142986 3360 143042 3369
rect 142724 3318 142986 3346
rect 142724 3233 142752 3318
rect 142986 3295 143042 3304
rect 142710 3224 142766 3233
rect 141700 3188 141752 3194
rect 141700 3130 141752 3136
rect 142160 3188 142212 3194
rect 142710 3159 142766 3168
rect 142160 3130 142212 3136
rect 141606 2680 141662 2689
rect 141606 2615 141662 2624
rect 141712 1562 141740 3130
rect 141790 3088 141846 3097
rect 141790 3023 141846 3032
rect 141804 2854 141832 3023
rect 141792 2848 141844 2854
rect 141792 2790 141844 2796
rect 143368 2106 143396 5102
rect 143552 4214 143580 10200
rect 144012 7002 144040 10200
rect 144380 10130 144408 10200
rect 144368 10124 144420 10130
rect 144368 10066 144420 10072
rect 144076 9276 144132 9296
rect 144076 9200 144132 9220
rect 144736 8968 144788 8974
rect 144736 8910 144788 8916
rect 144458 8664 144514 8673
rect 144458 8599 144514 8608
rect 144472 8401 144500 8599
rect 144458 8392 144514 8401
rect 144458 8327 144514 8336
rect 144076 8188 144132 8208
rect 144076 8112 144132 8132
rect 144276 7268 144328 7274
rect 144276 7210 144328 7216
rect 144288 7177 144316 7210
rect 144274 7168 144330 7177
rect 144076 7100 144132 7120
rect 144274 7103 144330 7112
rect 144076 7024 144132 7044
rect 144000 6996 144052 7002
rect 144000 6938 144052 6944
rect 143630 6896 143686 6905
rect 143630 6831 143632 6840
rect 143684 6831 143686 6840
rect 143632 6802 143684 6808
rect 143908 6248 143960 6254
rect 143908 6190 143960 6196
rect 144458 6216 144514 6225
rect 143920 5914 143948 6190
rect 144458 6151 144514 6160
rect 144076 6012 144132 6032
rect 144076 5936 144132 5956
rect 143908 5908 143960 5914
rect 143908 5850 143960 5856
rect 144472 5817 144500 6151
rect 144458 5808 144514 5817
rect 144458 5743 144514 5752
rect 144458 5536 144514 5545
rect 144458 5471 144514 5480
rect 144642 5536 144698 5545
rect 144642 5471 144698 5480
rect 144368 5228 144420 5234
rect 144368 5170 144420 5176
rect 144076 4924 144132 4944
rect 144076 4848 144132 4868
rect 144380 4842 144408 5170
rect 144472 5137 144500 5471
rect 144458 5128 144514 5137
rect 144458 5063 144514 5072
rect 144656 4842 144684 5471
rect 144380 4814 144684 4842
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 143906 3904 143962 3913
rect 143906 3839 143962 3848
rect 143920 3618 143948 3839
rect 144076 3836 144132 3856
rect 144076 3760 144132 3780
rect 144550 3768 144606 3777
rect 144748 3720 144776 8910
rect 144840 8634 144868 10200
rect 144920 9376 144972 9382
rect 144920 9318 144972 9324
rect 144828 8628 144880 8634
rect 144828 8570 144880 8576
rect 144932 8498 144960 9318
rect 144920 8492 144972 8498
rect 144920 8434 144972 8440
rect 145012 7948 145064 7954
rect 145012 7890 145064 7896
rect 144920 6792 144972 6798
rect 144920 6734 144972 6740
rect 144932 6361 144960 6734
rect 144918 6352 144974 6361
rect 144918 6287 144974 6296
rect 144828 5364 144880 5370
rect 144828 5306 144880 5312
rect 144840 5234 144868 5306
rect 144828 5228 144880 5234
rect 144828 5170 144880 5176
rect 144828 5024 144880 5030
rect 144828 4966 144880 4972
rect 144550 3703 144606 3712
rect 144458 3632 144514 3641
rect 143920 3590 144458 3618
rect 144458 3567 144514 3576
rect 144000 3528 144052 3534
rect 144000 3470 144052 3476
rect 144276 3528 144328 3534
rect 144276 3470 144328 3476
rect 143724 2984 143776 2990
rect 143724 2926 143776 2932
rect 143356 2100 143408 2106
rect 143356 2042 143408 2048
rect 142250 1728 142306 1737
rect 142250 1663 142306 1672
rect 141700 1556 141752 1562
rect 141700 1498 141752 1504
rect 141148 1420 141200 1426
rect 141148 1362 141200 1368
rect 141344 1414 141464 1442
rect 141516 1420 141568 1426
rect 141344 800 141372 1414
rect 141516 1362 141568 1368
rect 141528 1290 141556 1362
rect 141516 1284 141568 1290
rect 141516 1226 141568 1232
rect 141790 1048 141846 1057
rect 141790 983 141846 992
rect 141804 800 141832 983
rect 142264 800 142292 1663
rect 143080 1556 143132 1562
rect 143080 1498 143132 1504
rect 142988 1488 143040 1494
rect 142988 1430 143040 1436
rect 142434 1320 142490 1329
rect 142434 1255 142490 1264
rect 142448 1057 142476 1255
rect 142896 1216 142948 1222
rect 142896 1158 142948 1164
rect 142434 1048 142490 1057
rect 142434 983 142490 992
rect 142540 870 142660 898
rect 140596 604 140648 610
rect 140596 546 140648 552
rect 140870 -400 140926 800
rect 141330 -400 141386 800
rect 141790 -400 141846 800
rect 142250 -400 142306 800
rect 142540 746 142568 870
rect 142632 800 142660 870
rect 142908 814 142936 1158
rect 143000 814 143028 1430
rect 142896 808 142948 814
rect 142528 740 142580 746
rect 142528 682 142580 688
rect 142618 -400 142674 800
rect 142896 750 142948 756
rect 142988 808 143040 814
rect 143092 800 143120 1498
rect 143552 870 143672 898
rect 143552 800 143580 870
rect 142988 750 143040 756
rect 143078 -400 143134 800
rect 143538 -400 143594 800
rect 143644 610 143672 870
rect 143736 746 143764 2926
rect 143906 1592 143962 1601
rect 143906 1527 143962 1536
rect 143816 1420 143868 1426
rect 143816 1362 143868 1368
rect 143828 882 143856 1362
rect 143920 1329 143948 1527
rect 143906 1320 143962 1329
rect 143906 1255 143962 1264
rect 143816 876 143868 882
rect 143816 818 143868 824
rect 144012 800 144040 3470
rect 144288 3398 144316 3470
rect 144276 3392 144328 3398
rect 144276 3334 144328 3340
rect 144460 3392 144512 3398
rect 144564 3369 144592 3703
rect 144656 3692 144776 3720
rect 144460 3334 144512 3340
rect 144550 3360 144606 3369
rect 144472 3210 144500 3334
rect 144550 3295 144606 3304
rect 144656 3210 144684 3692
rect 144736 3596 144788 3602
rect 144736 3538 144788 3544
rect 144748 3398 144776 3538
rect 144840 3516 144868 4966
rect 144920 3528 144972 3534
rect 144840 3488 144920 3516
rect 144920 3470 144972 3476
rect 144736 3392 144788 3398
rect 144734 3360 144736 3369
rect 144828 3392 144880 3398
rect 144788 3360 144790 3369
rect 144828 3334 144880 3340
rect 144734 3295 144790 3304
rect 144472 3182 144684 3210
rect 144840 3126 144868 3334
rect 144828 3120 144880 3126
rect 144828 3062 144880 3068
rect 144368 2916 144420 2922
rect 144368 2858 144420 2864
rect 144552 2916 144604 2922
rect 144552 2858 144604 2864
rect 144076 2748 144132 2768
rect 144076 2672 144132 2692
rect 144184 2644 144236 2650
rect 144184 2586 144236 2592
rect 144196 2038 144224 2586
rect 144184 2032 144236 2038
rect 144184 1974 144236 1980
rect 144276 1964 144328 1970
rect 144276 1906 144328 1912
rect 144288 1737 144316 1906
rect 144274 1728 144330 1737
rect 144076 1660 144132 1680
rect 144274 1663 144330 1672
rect 144076 1584 144132 1604
rect 144380 800 144408 2858
rect 144460 2848 144512 2854
rect 144458 2816 144460 2825
rect 144512 2816 144514 2825
rect 144458 2751 144514 2760
rect 144564 2650 144592 2858
rect 144552 2644 144604 2650
rect 144552 2586 144604 2592
rect 144552 2508 144604 2514
rect 144552 2450 144604 2456
rect 144460 2372 144512 2378
rect 144460 2314 144512 2320
rect 144472 2038 144500 2314
rect 144460 2032 144512 2038
rect 144460 1974 144512 1980
rect 144564 950 144592 2450
rect 145024 2378 145052 7890
rect 145104 6248 145156 6254
rect 145104 6190 145156 6196
rect 145116 6118 145144 6190
rect 145104 6112 145156 6118
rect 145104 6054 145156 6060
rect 145300 4321 145328 10200
rect 145576 10146 145604 10270
rect 145654 10200 145710 11400
rect 145840 10260 145892 10266
rect 145840 10202 145892 10208
rect 145668 10146 145696 10200
rect 145576 10118 145696 10146
rect 145472 9036 145524 9042
rect 145472 8978 145524 8984
rect 145380 6316 145432 6322
rect 145380 6258 145432 6264
rect 145392 5370 145420 6258
rect 145380 5364 145432 5370
rect 145380 5306 145432 5312
rect 145380 4480 145432 4486
rect 145380 4422 145432 4428
rect 145286 4312 145342 4321
rect 145286 4247 145342 4256
rect 145196 2984 145248 2990
rect 145194 2952 145196 2961
rect 145288 2984 145340 2990
rect 145248 2952 145250 2961
rect 145288 2926 145340 2932
rect 145194 2887 145250 2896
rect 144644 2372 144696 2378
rect 144644 2314 144696 2320
rect 145012 2372 145064 2378
rect 145012 2314 145064 2320
rect 144656 1426 144684 2314
rect 144736 1896 144788 1902
rect 144736 1838 144788 1844
rect 144644 1420 144696 1426
rect 144644 1362 144696 1368
rect 144642 1320 144698 1329
rect 144642 1255 144644 1264
rect 144696 1255 144698 1264
rect 144644 1226 144696 1232
rect 144552 944 144604 950
rect 144748 932 144776 1838
rect 144932 1822 145236 1850
rect 145300 1834 145328 2926
rect 144932 1494 144960 1822
rect 145208 1766 145236 1822
rect 145288 1828 145340 1834
rect 145288 1770 145340 1776
rect 145104 1760 145156 1766
rect 145104 1702 145156 1708
rect 145196 1760 145248 1766
rect 145196 1702 145248 1708
rect 145116 1494 145144 1702
rect 144920 1488 144972 1494
rect 144920 1430 144972 1436
rect 145104 1488 145156 1494
rect 145104 1430 145156 1436
rect 145012 1216 145064 1222
rect 145064 1176 145144 1204
rect 145012 1158 145064 1164
rect 144748 904 144960 932
rect 144552 886 144604 892
rect 144656 836 144868 864
rect 143724 740 143776 746
rect 143724 682 143776 688
rect 143632 604 143684 610
rect 143632 546 143684 552
rect 143998 -400 144054 800
rect 144366 -400 144422 800
rect 144656 746 144684 836
rect 144840 800 144868 836
rect 144644 740 144696 746
rect 144644 682 144696 688
rect 144826 -400 144882 800
rect 144932 746 144960 904
rect 144920 740 144972 746
rect 144920 682 144972 688
rect 145116 218 145144 1176
rect 145392 1034 145420 4422
rect 145484 3738 145512 8978
rect 145852 8974 145880 10202
rect 146114 10200 146170 11400
rect 146574 10200 146630 11400
rect 147034 10200 147090 11400
rect 147312 10600 147364 10606
rect 147312 10542 147364 10548
rect 146128 9450 146156 10200
rect 146116 9444 146168 9450
rect 146116 9386 146168 9392
rect 146114 9072 146170 9081
rect 146114 9007 146170 9016
rect 145840 8968 145892 8974
rect 145840 8910 145892 8916
rect 146128 8566 146156 9007
rect 146116 8560 146168 8566
rect 146116 8502 146168 8508
rect 146208 8424 146260 8430
rect 146208 8366 146260 8372
rect 145564 8356 145616 8362
rect 145564 8298 145616 8304
rect 145472 3732 145524 3738
rect 145472 3674 145524 3680
rect 145576 3126 145604 8298
rect 145932 7880 145984 7886
rect 145932 7822 145984 7828
rect 145944 7410 145972 7822
rect 145932 7404 145984 7410
rect 145932 7346 145984 7352
rect 145840 6112 145892 6118
rect 145840 6054 145892 6060
rect 145656 4276 145708 4282
rect 145656 4218 145708 4224
rect 145564 3120 145616 3126
rect 145564 3062 145616 3068
rect 145562 2136 145618 2145
rect 145562 2071 145618 2080
rect 145576 1902 145604 2071
rect 145472 1896 145524 1902
rect 145472 1838 145524 1844
rect 145564 1896 145616 1902
rect 145564 1838 145616 1844
rect 145484 1426 145512 1838
rect 145668 1442 145696 4218
rect 145748 3528 145800 3534
rect 145748 3470 145800 3476
rect 145760 2582 145788 3470
rect 145748 2576 145800 2582
rect 145748 2518 145800 2524
rect 145852 2145 145880 6054
rect 146116 5704 146168 5710
rect 146116 5646 146168 5652
rect 146024 3460 146076 3466
rect 146024 3402 146076 3408
rect 145838 2136 145894 2145
rect 145838 2071 145894 2080
rect 145472 1420 145524 1426
rect 145668 1414 145880 1442
rect 145472 1362 145524 1368
rect 145746 1320 145802 1329
rect 145746 1255 145748 1264
rect 145800 1255 145802 1264
rect 145748 1226 145800 1232
rect 145852 1034 145880 1414
rect 146036 1306 146064 3402
rect 146128 3126 146156 5646
rect 146116 3120 146168 3126
rect 146116 3062 146168 3068
rect 146116 2916 146168 2922
rect 146116 2858 146168 2864
rect 146128 2446 146156 2858
rect 146116 2440 146168 2446
rect 146116 2382 146168 2388
rect 146114 2272 146170 2281
rect 146114 2207 146170 2216
rect 146128 1442 146156 2207
rect 146220 1562 146248 8366
rect 146392 5704 146444 5710
rect 146392 5646 146444 5652
rect 146404 5234 146432 5646
rect 146392 5228 146444 5234
rect 146392 5170 146444 5176
rect 146392 2304 146444 2310
rect 146390 2272 146392 2281
rect 146444 2272 146446 2281
rect 146390 2207 146446 2216
rect 146208 1556 146260 1562
rect 146208 1498 146260 1504
rect 146128 1414 146248 1442
rect 146220 1306 146248 1414
rect 146036 1278 146156 1306
rect 146220 1278 146340 1306
rect 145300 1006 145420 1034
rect 145668 1006 145880 1034
rect 145300 800 145328 1006
rect 145668 800 145696 1006
rect 146128 800 146156 1278
rect 146312 1034 146340 1278
rect 146588 1170 146616 10200
rect 147048 6474 147076 10200
rect 147324 10146 147352 10542
rect 147402 10200 147458 11400
rect 147862 10200 147918 11400
rect 148322 10200 148378 11400
rect 148782 10200 148838 11400
rect 149150 10200 149206 11400
rect 149610 10200 149666 11400
rect 150070 10200 150126 11400
rect 150530 10200 150586 11400
rect 150898 10200 150954 11400
rect 151358 10200 151414 11400
rect 151818 10200 151874 11400
rect 152186 10200 152242 11400
rect 152646 10200 152702 11400
rect 153106 10200 153162 11400
rect 153566 10200 153622 11400
rect 153934 10200 153990 11400
rect 154394 10200 154450 11400
rect 154854 10200 154910 11400
rect 155314 10200 155370 11400
rect 155682 10200 155738 11400
rect 156142 10200 156198 11400
rect 156602 10200 156658 11400
rect 157062 10200 157118 11400
rect 157430 10200 157486 11400
rect 157890 10200 157946 11400
rect 158350 10200 158406 11400
rect 158810 10200 158866 11400
rect 159178 10200 159234 11400
rect 159638 10200 159694 11400
rect 160098 10200 160154 11400
rect 160466 10200 160522 11400
rect 160926 10200 160982 11400
rect 161386 10200 161442 11400
rect 161846 10200 161902 11400
rect 162214 10200 162270 11400
rect 162674 10200 162730 11400
rect 163134 10200 163190 11400
rect 163594 10200 163650 11400
rect 163962 10200 164018 11400
rect 164422 10200 164478 11400
rect 164882 10200 164938 11400
rect 165342 10200 165398 11400
rect 165710 10200 165766 11400
rect 166170 10200 166226 11400
rect 166630 10200 166686 11400
rect 167090 10200 167146 11400
rect 167458 10200 167514 11400
rect 167918 10200 167974 11400
rect 168378 10200 168434 11400
rect 168746 10200 168802 11400
rect 169206 10200 169262 11400
rect 169576 10260 169628 10266
rect 169576 10202 169628 10208
rect 147416 10146 147444 10200
rect 147324 10118 147444 10146
rect 147680 9376 147732 9382
rect 147680 9318 147732 9324
rect 147692 9110 147720 9318
rect 147680 9104 147732 9110
rect 147680 9046 147732 9052
rect 147220 8016 147272 8022
rect 147272 7976 147352 8004
rect 147220 7958 147272 7964
rect 146772 6446 147076 6474
rect 146668 2508 146720 2514
rect 146668 2450 146720 2456
rect 146680 1426 146708 2450
rect 146668 1420 146720 1426
rect 146668 1362 146720 1368
rect 146588 1142 146708 1170
rect 146312 1006 146616 1034
rect 146588 800 146616 1006
rect 145194 232 145250 241
rect 145116 190 145194 218
rect 145194 167 145250 176
rect 145286 -400 145342 800
rect 145654 -400 145710 800
rect 146114 -400 146170 800
rect 146574 -400 146630 800
rect 146680 785 146708 1142
rect 146772 1057 146800 6446
rect 147128 3120 147180 3126
rect 147128 3062 147180 3068
rect 147036 2848 147088 2854
rect 147036 2790 147088 2796
rect 146944 2032 146996 2038
rect 146944 1974 146996 1980
rect 146852 1828 146904 1834
rect 146852 1770 146904 1776
rect 146864 1562 146892 1770
rect 146852 1556 146904 1562
rect 146852 1498 146904 1504
rect 146956 1494 146984 1974
rect 146944 1488 146996 1494
rect 146944 1430 146996 1436
rect 146758 1048 146814 1057
rect 146758 983 146814 992
rect 147048 800 147076 2790
rect 147140 2106 147168 3062
rect 147324 2106 147352 7976
rect 147772 7880 147824 7886
rect 147772 7822 147824 7828
rect 147680 7336 147732 7342
rect 147680 7278 147732 7284
rect 147692 6322 147720 7278
rect 147784 6866 147812 7822
rect 147876 6934 147904 10200
rect 148230 9344 148286 9353
rect 148230 9279 148286 9288
rect 148244 8906 148272 9279
rect 148336 9178 148364 10200
rect 148416 9376 148468 9382
rect 148416 9318 148468 9324
rect 148324 9172 148376 9178
rect 148324 9114 148376 9120
rect 148232 8900 148284 8906
rect 148232 8842 148284 8848
rect 148428 8498 148456 9318
rect 148416 8492 148468 8498
rect 148416 8434 148468 8440
rect 148692 8492 148744 8498
rect 148692 8434 148744 8440
rect 147864 6928 147916 6934
rect 147864 6870 147916 6876
rect 147772 6860 147824 6866
rect 147772 6802 147824 6808
rect 147956 6860 148008 6866
rect 147956 6802 148008 6808
rect 147680 6316 147732 6322
rect 147680 6258 147732 6264
rect 147588 3596 147640 3602
rect 147588 3538 147640 3544
rect 147600 3126 147628 3538
rect 147588 3120 147640 3126
rect 147588 3062 147640 3068
rect 147968 2650 147996 6802
rect 148704 6769 148732 8434
rect 148690 6760 148746 6769
rect 148690 6695 148746 6704
rect 148796 5710 148824 10200
rect 148966 10024 149022 10033
rect 148966 9959 149022 9968
rect 148980 7410 149008 9959
rect 148968 7404 149020 7410
rect 148968 7346 149020 7352
rect 148876 7336 148928 7342
rect 148876 7278 148928 7284
rect 148784 5704 148836 5710
rect 148784 5646 148836 5652
rect 148324 4820 148376 4826
rect 148324 4762 148376 4768
rect 148336 4622 148364 4762
rect 148324 4616 148376 4622
rect 148324 4558 148376 4564
rect 148324 2984 148376 2990
rect 148324 2926 148376 2932
rect 147956 2644 148008 2650
rect 147956 2586 148008 2592
rect 147404 2440 147456 2446
rect 147404 2382 147456 2388
rect 147128 2100 147180 2106
rect 147128 2042 147180 2048
rect 147312 2100 147364 2106
rect 147312 2042 147364 2048
rect 147416 2038 147444 2382
rect 147404 2032 147456 2038
rect 147404 1974 147456 1980
rect 147404 1556 147456 1562
rect 147404 1498 147456 1504
rect 147416 800 147444 1498
rect 147864 1216 147916 1222
rect 147864 1158 147916 1164
rect 148232 1216 148284 1222
rect 148232 1158 148284 1164
rect 147876 800 147904 1158
rect 148244 882 148272 1158
rect 148232 876 148284 882
rect 148232 818 148284 824
rect 148336 800 148364 2926
rect 148888 2106 148916 7278
rect 149164 6905 149192 10200
rect 149150 6896 149206 6905
rect 149150 6831 149206 6840
rect 149624 5302 149652 10200
rect 149704 10124 149756 10130
rect 149704 10066 149756 10072
rect 149716 8498 149744 10066
rect 149704 8492 149756 8498
rect 149704 8434 149756 8440
rect 150084 7970 150112 10200
rect 150440 9036 150492 9042
rect 150440 8978 150492 8984
rect 149992 7942 150112 7970
rect 149992 6458 150020 7942
rect 150072 7880 150124 7886
rect 150072 7822 150124 7828
rect 150084 7478 150112 7822
rect 150072 7472 150124 7478
rect 150072 7414 150124 7420
rect 150348 7268 150400 7274
rect 150348 7210 150400 7216
rect 149980 6452 150032 6458
rect 149980 6394 150032 6400
rect 149612 5296 149664 5302
rect 149612 5238 149664 5244
rect 149704 3392 149756 3398
rect 149704 3334 149756 3340
rect 149244 2848 149296 2854
rect 149244 2790 149296 2796
rect 149060 2440 149112 2446
rect 149060 2382 149112 2388
rect 148876 2100 148928 2106
rect 148876 2042 148928 2048
rect 148784 1488 148836 1494
rect 148784 1430 148836 1436
rect 148796 800 148824 1430
rect 149072 1426 149100 2382
rect 149150 1592 149206 1601
rect 149150 1527 149206 1536
rect 149060 1420 149112 1426
rect 149060 1362 149112 1368
rect 149164 800 149192 1527
rect 146666 776 146722 785
rect 146666 711 146722 720
rect 147034 -400 147090 800
rect 147402 -400 147458 800
rect 147862 -400 147918 800
rect 148322 -400 148378 800
rect 148782 -400 148838 800
rect 149150 -400 149206 800
rect 149256 610 149284 2790
rect 149612 1828 149664 1834
rect 149612 1770 149664 1776
rect 149624 800 149652 1770
rect 149716 1018 149744 3334
rect 150256 2576 150308 2582
rect 150256 2518 150308 2524
rect 150072 2032 150124 2038
rect 150072 1974 150124 1980
rect 149704 1012 149756 1018
rect 149704 954 149756 960
rect 150084 800 150112 1974
rect 150268 1426 150296 2518
rect 150360 1562 150388 7210
rect 150452 3738 150480 8978
rect 150544 6633 150572 10200
rect 150624 9512 150676 9518
rect 150624 9454 150676 9460
rect 150530 6624 150586 6633
rect 150530 6559 150586 6568
rect 150636 6322 150664 9454
rect 150716 9104 150768 9110
rect 150716 9046 150768 9052
rect 150728 8498 150756 9046
rect 150716 8492 150768 8498
rect 150716 8434 150768 8440
rect 150716 7336 150768 7342
rect 150716 7278 150768 7284
rect 150728 6866 150756 7278
rect 150716 6860 150768 6866
rect 150716 6802 150768 6808
rect 150624 6316 150676 6322
rect 150624 6258 150676 6264
rect 150440 3732 150492 3738
rect 150440 3674 150492 3680
rect 150912 2088 150940 10200
rect 151268 10056 151320 10062
rect 151268 9998 151320 10004
rect 151280 9586 151308 9998
rect 151268 9580 151320 9586
rect 151268 9522 151320 9528
rect 151084 8968 151136 8974
rect 151084 8910 151136 8916
rect 151096 8634 151124 8910
rect 151084 8628 151136 8634
rect 151084 8570 151136 8576
rect 151084 7880 151136 7886
rect 151084 7822 151136 7828
rect 151096 6866 151124 7822
rect 151084 6860 151136 6866
rect 151084 6802 151136 6808
rect 151372 5642 151400 10200
rect 151636 9444 151688 9450
rect 151636 9386 151688 9392
rect 151648 8498 151676 9386
rect 151636 8492 151688 8498
rect 151636 8434 151688 8440
rect 151728 7404 151780 7410
rect 151728 7346 151780 7352
rect 151740 6633 151768 7346
rect 151726 6624 151782 6633
rect 151726 6559 151782 6568
rect 151634 6488 151690 6497
rect 151634 6423 151690 6432
rect 151648 6322 151676 6423
rect 151636 6316 151688 6322
rect 151636 6258 151688 6264
rect 151832 6089 151860 10200
rect 152096 9716 152148 9722
rect 152096 9658 152148 9664
rect 152108 9178 152136 9658
rect 152096 9172 152148 9178
rect 152096 9114 152148 9120
rect 152200 6186 152228 10200
rect 152370 7984 152426 7993
rect 152370 7919 152426 7928
rect 152384 7721 152412 7919
rect 152464 7812 152516 7818
rect 152464 7754 152516 7760
rect 152370 7712 152426 7721
rect 152370 7647 152426 7656
rect 152188 6180 152240 6186
rect 152188 6122 152240 6128
rect 151818 6080 151874 6089
rect 151818 6015 151874 6024
rect 151360 5636 151412 5642
rect 151360 5578 151412 5584
rect 152372 4072 152424 4078
rect 152372 4014 152424 4020
rect 151728 3936 151780 3942
rect 151266 3904 151322 3913
rect 151728 3878 151780 3884
rect 151266 3839 151322 3848
rect 151174 2408 151230 2417
rect 151174 2343 151230 2352
rect 150820 2060 150940 2088
rect 150348 1556 150400 1562
rect 150348 1498 150400 1504
rect 150530 1456 150586 1465
rect 150256 1420 150308 1426
rect 150530 1391 150586 1400
rect 150256 1362 150308 1368
rect 150544 800 150572 1391
rect 149244 604 149296 610
rect 149244 546 149296 552
rect 149610 -400 149666 800
rect 150070 -400 150126 800
rect 150530 -400 150586 800
rect 150820 406 150848 2060
rect 150900 1964 150952 1970
rect 150900 1906 150952 1912
rect 150912 800 150940 1906
rect 151188 1601 151216 2343
rect 151174 1592 151230 1601
rect 151174 1527 151230 1536
rect 151280 1442 151308 3839
rect 151634 3496 151690 3505
rect 151634 3431 151690 3440
rect 151360 3120 151412 3126
rect 151412 3080 151584 3108
rect 151360 3062 151412 3068
rect 151556 2990 151584 3080
rect 151452 2984 151504 2990
rect 151452 2926 151504 2932
rect 151544 2984 151596 2990
rect 151544 2926 151596 2932
rect 151648 2938 151676 3431
rect 151740 3074 151768 3878
rect 151820 3664 151872 3670
rect 151820 3606 151872 3612
rect 151832 3534 151860 3606
rect 151820 3528 151872 3534
rect 152384 3505 152412 4014
rect 151820 3470 151872 3476
rect 152370 3496 152426 3505
rect 152370 3431 152426 3440
rect 152002 3088 152058 3097
rect 151740 3046 152002 3074
rect 152002 3023 152058 3032
rect 151280 1414 151400 1442
rect 151372 800 151400 1414
rect 150808 400 150860 406
rect 150808 342 150860 348
rect 150898 -400 150954 800
rect 151358 -400 151414 800
rect 151464 610 151492 2926
rect 151648 2910 151860 2938
rect 151832 800 151860 2910
rect 152186 2000 152242 2009
rect 152186 1935 152242 1944
rect 152200 800 152228 1935
rect 152476 1562 152504 7754
rect 152554 7712 152610 7721
rect 152554 7647 152610 7656
rect 152568 6798 152596 7647
rect 152556 6792 152608 6798
rect 152556 6734 152608 6740
rect 152660 3584 152688 10200
rect 152832 8968 152884 8974
rect 152832 8910 152884 8916
rect 152844 8498 152872 8910
rect 152832 8492 152884 8498
rect 152832 8434 152884 8440
rect 153016 7880 153068 7886
rect 153120 7868 153148 10200
rect 153476 9512 153528 9518
rect 153476 9454 153528 9460
rect 153068 7840 153148 7868
rect 153292 7880 153344 7886
rect 153016 7822 153068 7828
rect 153292 7822 153344 7828
rect 153106 6896 153162 6905
rect 153016 6860 153068 6866
rect 153106 6831 153162 6840
rect 153016 6802 153068 6808
rect 152924 5636 152976 5642
rect 152924 5578 152976 5584
rect 152660 3556 152780 3584
rect 152648 3460 152700 3466
rect 152648 3402 152700 3408
rect 152464 1556 152516 1562
rect 152464 1498 152516 1504
rect 152660 800 152688 3402
rect 152752 882 152780 3556
rect 152936 1018 152964 5578
rect 153028 2310 153056 6802
rect 153120 6798 153148 6831
rect 153108 6792 153160 6798
rect 153108 6734 153160 6740
rect 153304 6322 153332 7822
rect 153292 6316 153344 6322
rect 153292 6258 153344 6264
rect 153292 5704 153344 5710
rect 153292 5646 153344 5652
rect 153304 5234 153332 5646
rect 153292 5228 153344 5234
rect 153292 5170 153344 5176
rect 153106 3632 153162 3641
rect 153106 3567 153162 3576
rect 153290 3632 153346 3641
rect 153290 3567 153346 3576
rect 153016 2304 153068 2310
rect 153016 2246 153068 2252
rect 152924 1012 152976 1018
rect 152924 954 152976 960
rect 152740 876 152792 882
rect 152740 818 152792 824
rect 153120 800 153148 3567
rect 153304 3233 153332 3567
rect 153290 3224 153346 3233
rect 153290 3159 153346 3168
rect 153488 2106 153516 9454
rect 153580 6361 153608 10200
rect 153844 9580 153896 9586
rect 153844 9522 153896 9528
rect 153856 9489 153884 9522
rect 153842 9480 153898 9489
rect 153842 9415 153898 9424
rect 153844 8424 153896 8430
rect 153844 8366 153896 8372
rect 153856 7410 153884 8366
rect 153844 7404 153896 7410
rect 153844 7346 153896 7352
rect 153566 6352 153622 6361
rect 153566 6287 153622 6296
rect 153948 6254 153976 10200
rect 154028 8356 154080 8362
rect 154028 8298 154080 8304
rect 153936 6248 153988 6254
rect 153936 6190 153988 6196
rect 153660 5772 153712 5778
rect 153660 5714 153712 5720
rect 153566 3496 153622 3505
rect 153566 3431 153622 3440
rect 153580 3233 153608 3431
rect 153566 3224 153622 3233
rect 153566 3159 153622 3168
rect 153566 2544 153622 2553
rect 153566 2479 153622 2488
rect 153476 2100 153528 2106
rect 153476 2042 153528 2048
rect 153580 800 153608 2479
rect 153672 2378 153700 5714
rect 153934 3768 153990 3777
rect 153934 3703 153990 3712
rect 153660 2372 153712 2378
rect 153660 2314 153712 2320
rect 153844 2032 153896 2038
rect 153844 1974 153896 1980
rect 153856 1426 153884 1974
rect 153844 1420 153896 1426
rect 153844 1362 153896 1368
rect 153948 800 153976 3703
rect 154040 1562 154068 8298
rect 154132 7954 154344 7970
rect 154120 7948 154356 7954
rect 154172 7942 154304 7948
rect 154120 7890 154172 7896
rect 154304 7890 154356 7896
rect 154408 5846 154436 10200
rect 154486 9208 154542 9217
rect 154486 9143 154542 9152
rect 154500 8974 154528 9143
rect 154488 8968 154540 8974
rect 154488 8910 154540 8916
rect 154868 6662 154896 10200
rect 154856 6656 154908 6662
rect 154856 6598 154908 6604
rect 155328 6390 155356 10200
rect 155592 9444 155644 9450
rect 155592 9386 155644 9392
rect 155500 9376 155552 9382
rect 155500 9318 155552 9324
rect 155408 8424 155460 8430
rect 155408 8366 155460 8372
rect 155316 6384 155368 6390
rect 155316 6326 155368 6332
rect 154396 5840 154448 5846
rect 154396 5782 154448 5788
rect 155420 2514 155448 8366
rect 155512 4826 155540 9318
rect 155604 7177 155632 9386
rect 155590 7168 155646 7177
rect 155590 7103 155646 7112
rect 155696 6225 155724 10200
rect 156052 9988 156104 9994
rect 156052 9930 156104 9936
rect 155776 9172 155828 9178
rect 155776 9114 155828 9120
rect 155788 7041 155816 9114
rect 155868 7948 155920 7954
rect 155868 7890 155920 7896
rect 155774 7032 155830 7041
rect 155774 6967 155830 6976
rect 155774 6760 155830 6769
rect 155774 6695 155830 6704
rect 155682 6216 155738 6225
rect 155682 6151 155738 6160
rect 155500 4820 155552 4826
rect 155500 4762 155552 4768
rect 155316 2508 155368 2514
rect 155316 2450 155368 2456
rect 155408 2508 155460 2514
rect 155408 2450 155460 2456
rect 155224 1964 155276 1970
rect 155224 1906 155276 1912
rect 154854 1592 154910 1601
rect 154028 1556 154080 1562
rect 154854 1527 154910 1536
rect 154028 1498 154080 1504
rect 154316 836 154436 864
rect 151452 604 151504 610
rect 151452 546 151504 552
rect 151818 -400 151874 800
rect 152186 -400 152242 800
rect 152646 -400 152702 800
rect 153106 -400 153162 800
rect 153566 -400 153622 800
rect 153934 -400 153990 800
rect 154316 241 154344 836
rect 154408 800 154436 836
rect 154868 800 154896 1527
rect 155040 1352 155092 1358
rect 155040 1294 155092 1300
rect 154302 232 154358 241
rect 154302 167 154358 176
rect 154394 -400 154450 800
rect 154854 -400 154910 800
rect 155052 406 155080 1294
rect 155040 400 155092 406
rect 155040 342 155092 348
rect 155236 241 155264 1906
rect 155328 1340 155356 2450
rect 155684 2032 155736 2038
rect 155788 2009 155816 6695
rect 155684 1974 155736 1980
rect 155774 2000 155830 2009
rect 155696 1562 155724 1974
rect 155774 1935 155830 1944
rect 155880 1952 155908 7890
rect 155960 7812 156012 7818
rect 155960 7754 156012 7760
rect 155972 5370 156000 7754
rect 156064 7342 156092 9930
rect 156156 9738 156184 10200
rect 156156 9710 156552 9738
rect 156328 9512 156380 9518
rect 156328 9454 156380 9460
rect 156236 8968 156288 8974
rect 156236 8910 156288 8916
rect 156248 8498 156276 8910
rect 156236 8492 156288 8498
rect 156236 8434 156288 8440
rect 156144 8424 156196 8430
rect 156144 8366 156196 8372
rect 156052 7336 156104 7342
rect 156052 7278 156104 7284
rect 155960 5364 156012 5370
rect 155960 5306 156012 5312
rect 156156 5273 156184 8366
rect 156142 5264 156198 5273
rect 156142 5199 156198 5208
rect 156234 4176 156290 4185
rect 156234 4111 156290 4120
rect 156144 2916 156196 2922
rect 156144 2858 156196 2864
rect 156052 2508 156104 2514
rect 156052 2450 156104 2456
rect 155960 1964 156012 1970
rect 155880 1924 155960 1952
rect 155960 1906 156012 1912
rect 156064 1766 156092 2450
rect 155960 1760 156012 1766
rect 155960 1702 156012 1708
rect 156052 1760 156104 1766
rect 156052 1702 156104 1708
rect 155684 1556 155736 1562
rect 155684 1498 155736 1504
rect 155500 1352 155552 1358
rect 155328 1312 155500 1340
rect 155500 1294 155552 1300
rect 155328 870 155448 898
rect 155328 800 155356 870
rect 155222 232 155278 241
rect 155222 167 155278 176
rect 155314 -400 155370 800
rect 155420 474 155448 870
rect 155604 870 155724 898
rect 155972 882 156000 1702
rect 156052 1352 156104 1358
rect 156052 1294 156104 1300
rect 155604 678 155632 870
rect 155696 800 155724 870
rect 155960 876 156012 882
rect 155960 818 156012 824
rect 155592 672 155644 678
rect 155592 614 155644 620
rect 155408 468 155460 474
rect 155408 410 155460 416
rect 155682 -400 155738 800
rect 156064 678 156092 1294
rect 156156 800 156184 2858
rect 156052 672 156104 678
rect 156052 614 156104 620
rect 156142 -400 156198 800
rect 156248 474 156276 4111
rect 156340 1426 156368 9454
rect 156418 8800 156474 8809
rect 156418 8735 156474 8744
rect 156432 7721 156460 8735
rect 156418 7712 156474 7721
rect 156418 7647 156474 7656
rect 156524 5574 156552 9710
rect 156616 9382 156644 10200
rect 156696 9648 156748 9654
rect 156694 9616 156696 9625
rect 156748 9616 156750 9625
rect 156694 9551 156750 9560
rect 156604 9376 156656 9382
rect 156604 9318 156656 9324
rect 157076 9194 157104 10200
rect 157444 9602 157472 10200
rect 157444 9574 157564 9602
rect 157432 9444 157484 9450
rect 157432 9386 157484 9392
rect 157340 9376 157392 9382
rect 157340 9318 157392 9324
rect 156616 9166 157104 9194
rect 156616 7886 156644 9166
rect 156696 9036 156748 9042
rect 156696 8978 156748 8984
rect 156880 9036 156932 9042
rect 156880 8978 156932 8984
rect 156604 7880 156656 7886
rect 156604 7822 156656 7828
rect 156602 7712 156658 7721
rect 156602 7647 156658 7656
rect 156616 6497 156644 7647
rect 156602 6488 156658 6497
rect 156602 6423 156658 6432
rect 156512 5568 156564 5574
rect 156512 5510 156564 5516
rect 156512 5092 156564 5098
rect 156512 5034 156564 5040
rect 156420 2984 156472 2990
rect 156420 2926 156472 2932
rect 156328 1420 156380 1426
rect 156328 1362 156380 1368
rect 156432 785 156460 2926
rect 156524 1329 156552 5034
rect 156602 4040 156658 4049
rect 156602 3975 156658 3984
rect 156616 1601 156644 3975
rect 156708 3126 156736 8978
rect 156788 7948 156840 7954
rect 156788 7890 156840 7896
rect 156800 7546 156828 7890
rect 156892 7857 156920 8978
rect 157156 8832 157208 8838
rect 157156 8774 157208 8780
rect 157062 8664 157118 8673
rect 157062 8599 157118 8608
rect 157076 7993 157104 8599
rect 157168 8265 157196 8774
rect 157154 8256 157210 8265
rect 157352 8242 157380 9318
rect 157444 8265 157472 9386
rect 157154 8191 157210 8200
rect 157260 8214 157380 8242
rect 157430 8256 157486 8265
rect 157062 7984 157118 7993
rect 157062 7919 157118 7928
rect 156878 7848 156934 7857
rect 156878 7783 156934 7792
rect 156788 7540 156840 7546
rect 156788 7482 156840 7488
rect 156878 7440 156934 7449
rect 157260 7426 157288 8214
rect 157430 8191 157486 8200
rect 157536 8129 157564 9574
rect 157614 8800 157670 8809
rect 157614 8735 157670 8744
rect 157522 8120 157578 8129
rect 157522 8055 157578 8064
rect 157628 7857 157656 8735
rect 157706 8392 157762 8401
rect 157706 8327 157762 8336
rect 157720 7886 157748 8327
rect 157708 7880 157760 7886
rect 157614 7848 157670 7857
rect 157708 7822 157760 7828
rect 157614 7783 157670 7792
rect 157430 7576 157486 7585
rect 157904 7562 157932 10200
rect 158076 9648 158128 9654
rect 158076 9590 158128 9596
rect 157984 8968 158036 8974
rect 157984 8910 158036 8916
rect 157996 7954 158024 8910
rect 157984 7948 158036 7954
rect 157984 7890 158036 7896
rect 157430 7511 157486 7520
rect 157536 7534 157932 7562
rect 156934 7398 157288 7426
rect 157340 7472 157392 7478
rect 157340 7414 157392 7420
rect 156878 7375 156934 7384
rect 157064 7336 157116 7342
rect 157352 7290 157380 7414
rect 157444 7324 157472 7511
rect 157536 7449 157564 7534
rect 157708 7472 157760 7478
rect 157522 7440 157578 7449
rect 157522 7375 157578 7384
rect 157706 7440 157708 7449
rect 157760 7440 157762 7449
rect 157706 7375 157762 7384
rect 158088 7324 158116 9590
rect 158364 7886 158392 10200
rect 158824 9178 158852 10200
rect 159088 10192 159140 10198
rect 159088 10134 159140 10140
rect 159100 9586 159128 10134
rect 159192 9994 159220 10200
rect 159180 9988 159232 9994
rect 159180 9930 159232 9936
rect 159088 9580 159140 9586
rect 159088 9522 159140 9528
rect 158812 9172 158864 9178
rect 158812 9114 158864 9120
rect 159548 8560 159600 8566
rect 159548 8502 159600 8508
rect 159560 8362 159588 8502
rect 159548 8356 159600 8362
rect 159548 8298 159600 8304
rect 159652 8294 159680 10200
rect 160112 9602 160140 10200
rect 160112 9574 160232 9602
rect 160100 9512 160152 9518
rect 160100 9454 160152 9460
rect 160112 9178 160140 9454
rect 160100 9172 160152 9178
rect 160100 9114 160152 9120
rect 160204 9042 160232 9574
rect 160284 9172 160336 9178
rect 160284 9114 160336 9120
rect 160192 9036 160244 9042
rect 160192 8978 160244 8984
rect 160008 8968 160060 8974
rect 160008 8910 160060 8916
rect 159824 8628 159876 8634
rect 159824 8570 159876 8576
rect 159916 8628 159968 8634
rect 159916 8570 159968 8576
rect 159640 8288 159692 8294
rect 159640 8230 159692 8236
rect 159836 7993 159864 8570
rect 159928 8498 159956 8570
rect 160020 8498 160048 8910
rect 159916 8492 159968 8498
rect 159916 8434 159968 8440
rect 160008 8492 160060 8498
rect 160008 8434 160060 8440
rect 159822 7984 159878 7993
rect 159822 7919 159878 7928
rect 159916 7948 159968 7954
rect 159916 7890 159968 7896
rect 158352 7880 158404 7886
rect 158352 7822 158404 7828
rect 158904 7540 158956 7546
rect 158904 7482 158956 7488
rect 158916 7449 158944 7482
rect 159928 7449 159956 7890
rect 160296 7478 160324 9114
rect 160480 8838 160508 10200
rect 160468 8832 160520 8838
rect 160468 8774 160520 8780
rect 160940 8673 160968 10200
rect 160926 8664 160982 8673
rect 160926 8599 160982 8608
rect 161400 8537 161428 10200
rect 161860 9761 161888 10200
rect 161846 9752 161902 9761
rect 161846 9687 161902 9696
rect 162228 9450 162256 10200
rect 162216 9444 162268 9450
rect 162216 9386 162268 9392
rect 162124 9104 162176 9110
rect 162124 9046 162176 9052
rect 161940 8968 161992 8974
rect 161940 8910 161992 8916
rect 161386 8528 161442 8537
rect 161386 8463 161442 8472
rect 161846 8528 161902 8537
rect 161846 8463 161902 8472
rect 160652 8288 160704 8294
rect 160652 8230 160704 8236
rect 160664 8022 160692 8230
rect 160652 8016 160704 8022
rect 160652 7958 160704 7964
rect 161204 7880 161256 7886
rect 161202 7848 161204 7857
rect 161256 7848 161258 7857
rect 161202 7783 161258 7792
rect 160284 7472 160336 7478
rect 158902 7440 158958 7449
rect 158902 7375 158958 7384
rect 159914 7440 159970 7449
rect 160284 7414 160336 7420
rect 161860 7410 161888 8463
rect 161952 7410 161980 8910
rect 162136 8129 162164 9046
rect 162584 8424 162636 8430
rect 162584 8366 162636 8372
rect 162122 8120 162178 8129
rect 162122 8055 162178 8064
rect 162308 7880 162360 7886
rect 162308 7822 162360 7828
rect 162320 7478 162348 7822
rect 162308 7472 162360 7478
rect 162596 7449 162624 8366
rect 162688 7721 162716 10200
rect 163148 8265 163176 10200
rect 163608 8809 163636 10200
rect 163594 8800 163650 8809
rect 163594 8735 163650 8744
rect 163976 8294 164004 10200
rect 164076 9820 164132 9840
rect 164076 9744 164132 9764
rect 164238 9752 164294 9761
rect 164160 9710 164238 9738
rect 164160 9654 164188 9710
rect 164238 9687 164294 9696
rect 164148 9648 164200 9654
rect 164148 9590 164200 9596
rect 164332 9376 164384 9382
rect 164332 9318 164384 9324
rect 164344 9042 164372 9318
rect 164332 9036 164384 9042
rect 164436 9024 164464 10200
rect 164896 9602 164924 10200
rect 165252 9988 165304 9994
rect 165252 9930 165304 9936
rect 165264 9654 165292 9930
rect 165356 9738 165384 10200
rect 165724 10169 165752 10200
rect 165710 10160 165766 10169
rect 165710 10095 165766 10104
rect 166184 9926 166212 10200
rect 166172 9920 166224 9926
rect 166172 9862 166224 9868
rect 166264 9920 166316 9926
rect 166264 9862 166316 9868
rect 165356 9710 165476 9738
rect 165252 9648 165304 9654
rect 164896 9574 165016 9602
rect 165252 9590 165304 9596
rect 165344 9648 165396 9654
rect 165344 9590 165396 9596
rect 164884 9512 164936 9518
rect 164884 9454 164936 9460
rect 164436 8996 164740 9024
rect 164332 8978 164384 8984
rect 164424 8900 164476 8906
rect 164424 8842 164476 8848
rect 164076 8732 164132 8752
rect 164076 8656 164132 8676
rect 164436 8634 164464 8842
rect 164332 8628 164384 8634
rect 164332 8570 164384 8576
rect 164424 8628 164476 8634
rect 164424 8570 164476 8576
rect 164344 8514 164372 8570
rect 164514 8528 164570 8537
rect 164344 8486 164514 8514
rect 164514 8463 164570 8472
rect 164240 8424 164292 8430
rect 164240 8366 164292 8372
rect 163964 8288 164016 8294
rect 163134 8256 163190 8265
rect 163134 8191 163190 8200
rect 163318 8256 163374 8265
rect 163964 8230 164016 8236
rect 163318 8191 163374 8200
rect 162674 7712 162730 7721
rect 162674 7647 162730 7656
rect 163332 7585 163360 8191
rect 164252 8090 164280 8366
rect 164516 8288 164568 8294
rect 164516 8230 164568 8236
rect 164608 8288 164660 8294
rect 164608 8230 164660 8236
rect 164240 8084 164292 8090
rect 164240 8026 164292 8032
rect 164332 8084 164384 8090
rect 164332 8026 164384 8032
rect 164344 7970 164372 8026
rect 164252 7954 164372 7970
rect 164528 7954 164556 8230
rect 164620 8022 164648 8230
rect 164608 8016 164660 8022
rect 164608 7958 164660 7964
rect 164240 7948 164372 7954
rect 164292 7942 164372 7948
rect 164516 7948 164568 7954
rect 164240 7890 164292 7896
rect 164516 7890 164568 7896
rect 164076 7644 164132 7664
rect 163318 7576 163374 7585
rect 164076 7568 164132 7588
rect 163318 7511 163374 7520
rect 164712 7449 164740 8996
rect 164792 8900 164844 8906
rect 164792 8842 164844 8848
rect 164804 8401 164832 8842
rect 164790 8392 164846 8401
rect 164790 8327 164846 8336
rect 164896 7449 164924 9454
rect 164988 7585 165016 9574
rect 165068 9580 165120 9586
rect 165068 9522 165120 9528
rect 165080 8090 165108 9522
rect 165356 8498 165384 9590
rect 165344 8492 165396 8498
rect 165344 8434 165396 8440
rect 165068 8084 165120 8090
rect 165068 8026 165120 8032
rect 165448 7857 165476 9710
rect 166276 9586 166304 9862
rect 166264 9580 166316 9586
rect 166264 9522 166316 9528
rect 166644 9178 166672 10200
rect 166998 9888 167054 9897
rect 166998 9823 167054 9832
rect 166632 9172 166684 9178
rect 166632 9114 166684 9120
rect 165620 9104 165672 9110
rect 165620 9046 165672 9052
rect 166448 9104 166500 9110
rect 166448 9046 166500 9052
rect 165434 7848 165490 7857
rect 165434 7783 165490 7792
rect 165632 7585 165660 9046
rect 166460 7750 166488 9046
rect 166816 8492 166868 8498
rect 166816 8434 166868 8440
rect 166540 8356 166592 8362
rect 166540 8298 166592 8304
rect 166448 7744 166500 7750
rect 166448 7686 166500 7692
rect 164974 7576 165030 7585
rect 164974 7511 165030 7520
rect 165618 7576 165674 7585
rect 165618 7511 165674 7520
rect 166552 7449 166580 8298
rect 166828 8129 166856 8434
rect 166814 8120 166870 8129
rect 166814 8055 166870 8064
rect 167012 7818 167040 9823
rect 167104 8294 167132 10200
rect 167472 9081 167500 10200
rect 167736 9512 167788 9518
rect 167736 9454 167788 9460
rect 167458 9072 167514 9081
rect 167458 9007 167514 9016
rect 167366 8664 167422 8673
rect 167366 8599 167422 8608
rect 167184 8424 167236 8430
rect 167184 8366 167236 8372
rect 167092 8288 167144 8294
rect 167196 8265 167224 8366
rect 167092 8230 167144 8236
rect 167182 8256 167238 8265
rect 167182 8191 167238 8200
rect 167276 8084 167328 8090
rect 167276 8026 167328 8032
rect 167288 7886 167316 8026
rect 167276 7880 167328 7886
rect 167276 7822 167328 7828
rect 167000 7812 167052 7818
rect 167000 7754 167052 7760
rect 167380 7585 167408 8599
rect 167748 8401 167776 9454
rect 167932 8945 167960 10200
rect 168392 9654 168420 10200
rect 168760 9761 168788 10200
rect 168746 9752 168802 9761
rect 168746 9687 168802 9696
rect 168380 9648 168432 9654
rect 168380 9590 168432 9596
rect 169116 9376 169168 9382
rect 169116 9318 169168 9324
rect 169024 9036 169076 9042
rect 169024 8978 169076 8984
rect 167918 8936 167974 8945
rect 167918 8871 167974 8880
rect 168472 8492 168524 8498
rect 168472 8434 168524 8440
rect 167734 8392 167790 8401
rect 167734 8327 167790 8336
rect 168484 8022 168512 8434
rect 169036 8401 169064 8978
rect 169022 8392 169078 8401
rect 169022 8327 169078 8336
rect 168472 8016 168524 8022
rect 168472 7958 168524 7964
rect 167736 7880 167788 7886
rect 167736 7822 167788 7828
rect 167366 7576 167422 7585
rect 167366 7511 167422 7520
rect 167748 7449 167776 7822
rect 169128 7449 169156 9318
rect 169220 8974 169248 10200
rect 169588 10146 169616 10202
rect 169666 10200 169722 11400
rect 170126 10200 170182 11400
rect 170494 10200 170550 11400
rect 170954 10200 171010 11400
rect 171414 10200 171470 11400
rect 171874 10200 171930 11400
rect 172242 10200 172298 11400
rect 172702 10200 172758 11400
rect 173162 10200 173218 11400
rect 173622 10200 173678 11400
rect 173990 10200 174046 11400
rect 174450 10200 174506 11400
rect 174910 10200 174966 11400
rect 175370 10200 175426 11400
rect 175738 10200 175794 11400
rect 176198 10200 176254 11400
rect 176658 10200 176714 11400
rect 177026 10200 177082 11400
rect 177486 10200 177542 11400
rect 177946 10200 178002 11400
rect 178406 10200 178462 11400
rect 178774 10200 178830 11400
rect 179234 10200 179290 11400
rect 179694 10200 179750 11400
rect 180154 10200 180210 11400
rect 180522 10200 180578 11400
rect 180982 10200 181038 11400
rect 181442 10200 181498 11400
rect 181902 10200 181958 11400
rect 182270 10200 182326 11400
rect 182730 10200 182786 11400
rect 183190 10200 183246 11400
rect 183650 10200 183706 11400
rect 184018 10200 184074 11400
rect 184478 10200 184534 11400
rect 184938 10200 184994 11400
rect 185306 10200 185362 11400
rect 185766 10200 185822 11400
rect 186226 10200 186282 11400
rect 186686 10200 186742 11400
rect 187054 10200 187110 11400
rect 187514 10200 187570 11400
rect 187974 10200 188030 11400
rect 188434 10200 188490 11400
rect 188802 10200 188858 11400
rect 189262 10200 189318 11400
rect 189722 10200 189778 11400
rect 190182 10200 190238 11400
rect 190550 10200 190606 11400
rect 191010 10200 191066 11400
rect 191470 10200 191526 11400
rect 191930 10200 191986 11400
rect 192298 10200 192354 11400
rect 192758 10200 192814 11400
rect 193218 10200 193274 11400
rect 193586 10200 193642 11400
rect 194046 10200 194102 11400
rect 194506 10200 194562 11400
rect 194966 10200 195022 11400
rect 195334 10200 195390 11400
rect 195794 10200 195850 11400
rect 196254 10200 196310 11400
rect 196714 10200 196770 11400
rect 197082 10200 197138 11400
rect 197542 10200 197598 11400
rect 198002 10200 198058 11400
rect 198462 10200 198518 11400
rect 198830 10200 198886 11400
rect 199290 10200 199346 11400
rect 199750 10200 199806 11400
rect 169680 10146 169708 10200
rect 169588 10118 169708 10146
rect 169944 10192 169996 10198
rect 169944 10134 169996 10140
rect 169760 9512 169812 9518
rect 169760 9454 169812 9460
rect 169208 8968 169260 8974
rect 169208 8910 169260 8916
rect 169390 8120 169446 8129
rect 169390 8055 169446 8064
rect 169404 7449 169432 8055
rect 169772 7449 169800 9454
rect 169956 9042 169984 10134
rect 170140 9353 170168 10200
rect 170126 9344 170182 9353
rect 170126 9279 170182 9288
rect 169944 9036 169996 9042
rect 169944 8978 169996 8984
rect 170036 8560 170088 8566
rect 170508 8537 170536 10200
rect 170968 9110 170996 10200
rect 171324 10192 171376 10198
rect 171324 10134 171376 10140
rect 171336 9654 171364 10134
rect 171324 9648 171376 9654
rect 171324 9590 171376 9596
rect 171428 9602 171456 10200
rect 171428 9574 171640 9602
rect 171416 9512 171468 9518
rect 171416 9454 171468 9460
rect 170956 9104 171008 9110
rect 170956 9046 171008 9052
rect 171232 9036 171284 9042
rect 171232 8978 171284 8984
rect 170036 8502 170088 8508
rect 170494 8528 170550 8537
rect 170048 8129 170076 8502
rect 170494 8463 170550 8472
rect 170772 8424 170824 8430
rect 170770 8392 170772 8401
rect 170824 8392 170826 8401
rect 170770 8327 170826 8336
rect 171048 8356 171100 8362
rect 171048 8298 171100 8304
rect 170034 8120 170090 8129
rect 170034 8055 170090 8064
rect 171060 7750 171088 8298
rect 171140 8288 171192 8294
rect 171140 8230 171192 8236
rect 171152 8090 171180 8230
rect 171140 8084 171192 8090
rect 171140 8026 171192 8032
rect 170036 7744 170088 7750
rect 170036 7686 170088 7692
rect 171048 7744 171100 7750
rect 171048 7686 171100 7692
rect 170048 7449 170076 7686
rect 171244 7449 171272 8978
rect 171428 7449 171456 9454
rect 171508 9104 171560 9110
rect 171508 9046 171560 9052
rect 171520 8566 171548 9046
rect 171612 8809 171640 9574
rect 171888 9217 171916 10200
rect 172256 9897 172284 10200
rect 172242 9888 172298 9897
rect 172242 9823 172298 9832
rect 172518 9752 172574 9761
rect 172518 9687 172574 9696
rect 172152 9580 172204 9586
rect 172152 9522 172204 9528
rect 171874 9208 171930 9217
rect 171874 9143 171930 9152
rect 171598 8800 171654 8809
rect 171598 8735 171654 8744
rect 171508 8560 171560 8566
rect 172164 8537 172192 9522
rect 172336 9512 172388 9518
rect 172336 9454 172388 9460
rect 171508 8502 171560 8508
rect 172150 8528 172206 8537
rect 172150 8463 172206 8472
rect 171784 8424 171836 8430
rect 171784 8366 171836 8372
rect 171796 7449 171824 8366
rect 172348 8090 172376 9454
rect 172532 8906 172560 9687
rect 172520 8900 172572 8906
rect 172520 8842 172572 8848
rect 172716 8242 172744 10200
rect 173176 8838 173204 10200
rect 173164 8832 173216 8838
rect 173164 8774 173216 8780
rect 172624 8214 172744 8242
rect 172336 8084 172388 8090
rect 172336 8026 172388 8032
rect 172624 7449 172652 8214
rect 172704 8084 172756 8090
rect 172704 8026 172756 8032
rect 172716 7818 172744 8026
rect 173532 7948 173584 7954
rect 173532 7890 173584 7896
rect 172704 7812 172756 7818
rect 172704 7754 172756 7760
rect 173544 7449 173572 7890
rect 173636 7857 173664 10200
rect 173716 9512 173768 9518
rect 173716 9454 173768 9460
rect 173728 9081 173756 9454
rect 174004 9217 174032 10200
rect 173990 9208 174046 9217
rect 173990 9143 174046 9152
rect 173714 9072 173770 9081
rect 173714 9007 173770 9016
rect 173716 8968 173768 8974
rect 173716 8910 173768 8916
rect 173728 7954 173756 8910
rect 174268 8832 174320 8838
rect 174268 8774 174320 8780
rect 173900 8288 173952 8294
rect 173900 8230 173952 8236
rect 173716 7948 173768 7954
rect 173716 7890 173768 7896
rect 173622 7848 173678 7857
rect 173912 7818 173940 8230
rect 173622 7783 173678 7792
rect 173900 7812 173952 7818
rect 173900 7754 173952 7760
rect 174280 7585 174308 8774
rect 174464 7585 174492 10200
rect 174924 9382 174952 10200
rect 175384 9489 175412 10200
rect 175464 9512 175516 9518
rect 175370 9480 175426 9489
rect 175464 9454 175516 9460
rect 175370 9415 175426 9424
rect 174912 9376 174964 9382
rect 174912 9318 174964 9324
rect 174912 9036 174964 9042
rect 174912 8978 174964 8984
rect 174266 7576 174322 7585
rect 174266 7511 174322 7520
rect 174450 7576 174506 7585
rect 174450 7511 174506 7520
rect 174924 7449 174952 8978
rect 175476 7449 175504 9454
rect 175752 8634 175780 10200
rect 176212 9761 176240 10200
rect 176198 9752 176254 9761
rect 176198 9687 176254 9696
rect 175924 9444 175976 9450
rect 175924 9386 175976 9392
rect 175936 9353 175964 9386
rect 175922 9344 175978 9353
rect 175922 9279 175978 9288
rect 175740 8628 175792 8634
rect 175740 8570 175792 8576
rect 176200 8628 176252 8634
rect 176200 8570 176252 8576
rect 176212 7818 176240 8570
rect 176672 8514 176700 10200
rect 177040 9994 177068 10200
rect 177028 9988 177080 9994
rect 177028 9930 177080 9936
rect 176752 8832 176804 8838
rect 176752 8774 176804 8780
rect 176844 8832 176896 8838
rect 176844 8774 176896 8780
rect 176488 8486 176700 8514
rect 176384 8424 176436 8430
rect 176382 8392 176384 8401
rect 176436 8392 176438 8401
rect 176488 8362 176516 8486
rect 176568 8424 176620 8430
rect 176568 8366 176620 8372
rect 176382 8327 176438 8336
rect 176476 8356 176528 8362
rect 176476 8298 176528 8304
rect 176382 8256 176438 8265
rect 176382 8191 176438 8200
rect 176396 7818 176424 8191
rect 176476 7948 176528 7954
rect 176476 7890 176528 7896
rect 176200 7812 176252 7818
rect 176200 7754 176252 7760
rect 176384 7812 176436 7818
rect 176384 7754 176436 7760
rect 176488 7585 176516 7890
rect 176580 7857 176608 8366
rect 176764 8265 176792 8774
rect 176856 8566 176884 8774
rect 176844 8560 176896 8566
rect 176844 8502 176896 8508
rect 177500 8294 177528 10200
rect 177856 9512 177908 9518
rect 177856 9454 177908 9460
rect 177488 8288 177540 8294
rect 176750 8256 176806 8265
rect 177488 8230 177540 8236
rect 176750 8191 176806 8200
rect 176566 7848 176622 7857
rect 176566 7783 176622 7792
rect 177486 7848 177542 7857
rect 177486 7783 177542 7792
rect 176568 7744 176620 7750
rect 176660 7744 176712 7750
rect 176620 7704 176660 7732
rect 176568 7686 176620 7692
rect 176660 7686 176712 7692
rect 176474 7576 176530 7585
rect 176474 7511 176530 7520
rect 162308 7414 162360 7420
rect 162582 7440 162638 7449
rect 159914 7375 159970 7384
rect 161848 7404 161900 7410
rect 161848 7346 161900 7352
rect 161940 7404 161992 7410
rect 162582 7375 162638 7384
rect 164698 7440 164754 7449
rect 164698 7375 164754 7384
rect 164882 7440 164938 7449
rect 164882 7375 164938 7384
rect 166538 7440 166594 7449
rect 166538 7375 166594 7384
rect 167734 7440 167790 7449
rect 167734 7375 167790 7384
rect 169114 7440 169170 7449
rect 169114 7375 169170 7384
rect 169390 7440 169446 7449
rect 169390 7375 169446 7384
rect 169758 7440 169814 7449
rect 169758 7375 169814 7384
rect 170034 7440 170090 7449
rect 170034 7375 170090 7384
rect 171230 7440 171286 7449
rect 171230 7375 171286 7384
rect 171414 7440 171470 7449
rect 171414 7375 171470 7384
rect 171782 7440 171838 7449
rect 171782 7375 171838 7384
rect 172610 7440 172666 7449
rect 172610 7375 172666 7384
rect 173530 7440 173586 7449
rect 173530 7375 173586 7384
rect 174910 7440 174966 7449
rect 174910 7375 174966 7384
rect 175462 7440 175518 7449
rect 175462 7375 175518 7384
rect 161940 7346 161992 7352
rect 157444 7296 158116 7324
rect 177500 7313 177528 7783
rect 177868 7313 177896 9454
rect 177960 7449 177988 10200
rect 178420 10033 178448 10200
rect 178406 10024 178462 10033
rect 178406 9959 178462 9968
rect 178040 8968 178092 8974
rect 178040 8910 178092 8916
rect 178052 7954 178080 8910
rect 178788 8537 178816 10200
rect 179248 9654 179276 10200
rect 179512 9920 179564 9926
rect 179512 9862 179564 9868
rect 179236 9648 179288 9654
rect 179236 9590 179288 9596
rect 179524 9178 179552 9862
rect 179708 9625 179736 10200
rect 179694 9616 179750 9625
rect 179694 9551 179750 9560
rect 179512 9172 179564 9178
rect 179512 9114 179564 9120
rect 178960 8628 179012 8634
rect 178960 8570 179012 8576
rect 178972 8537 179000 8570
rect 178774 8528 178830 8537
rect 178774 8463 178830 8472
rect 178958 8528 179014 8537
rect 178958 8463 179014 8472
rect 179512 8288 179564 8294
rect 180168 8265 180196 10200
rect 180536 8673 180564 10200
rect 180522 8664 180578 8673
rect 180522 8599 180578 8608
rect 180996 8362 181024 10200
rect 181260 10056 181312 10062
rect 181260 9998 181312 10004
rect 181272 9586 181300 9998
rect 181260 9580 181312 9586
rect 181260 9522 181312 9528
rect 181456 8514 181484 10200
rect 181536 9988 181588 9994
rect 181536 9930 181588 9936
rect 181548 9722 181576 9930
rect 181536 9716 181588 9722
rect 181536 9658 181588 9664
rect 181628 9648 181680 9654
rect 181628 9590 181680 9596
rect 181640 9042 181668 9590
rect 181628 9036 181680 9042
rect 181628 8978 181680 8984
rect 181916 8809 181944 10200
rect 182088 10056 182140 10062
rect 182088 9998 182140 10004
rect 181996 9036 182048 9042
rect 181996 8978 182048 8984
rect 181902 8800 181958 8809
rect 181902 8735 181958 8744
rect 181272 8486 181484 8514
rect 180984 8356 181036 8362
rect 180984 8298 181036 8304
rect 179512 8230 179564 8236
rect 180154 8256 180210 8265
rect 178040 7948 178092 7954
rect 178040 7890 178092 7896
rect 179524 7886 179552 8230
rect 180154 8191 180210 8200
rect 180614 8256 180670 8265
rect 180614 8191 180670 8200
rect 179512 7880 179564 7886
rect 180628 7857 180656 8191
rect 181272 8129 181300 8486
rect 181444 8424 181496 8430
rect 181442 8392 181444 8401
rect 181496 8392 181498 8401
rect 181442 8327 181498 8336
rect 181258 8120 181314 8129
rect 181258 8055 181314 8064
rect 181352 8084 181404 8090
rect 181352 8026 181404 8032
rect 181536 8084 181588 8090
rect 181536 8026 181588 8032
rect 181168 7880 181220 7886
rect 179512 7822 179564 7828
rect 180614 7848 180670 7857
rect 178408 7812 178460 7818
rect 181168 7822 181220 7828
rect 180614 7783 180670 7792
rect 178408 7754 178460 7760
rect 178420 7449 178448 7754
rect 180890 7712 180946 7721
rect 180890 7647 180946 7656
rect 180904 7478 180932 7647
rect 180892 7472 180944 7478
rect 177946 7440 178002 7449
rect 177946 7375 178002 7384
rect 178406 7440 178462 7449
rect 181180 7449 181208 7822
rect 181364 7546 181392 8026
rect 181352 7540 181404 7546
rect 181352 7482 181404 7488
rect 180892 7414 180944 7420
rect 181166 7440 181222 7449
rect 178406 7375 178462 7384
rect 181548 7410 181576 8026
rect 181812 7744 181864 7750
rect 181812 7686 181864 7692
rect 181824 7410 181852 7686
rect 182008 7449 182036 8978
rect 182100 8906 182128 9998
rect 182088 8900 182140 8906
rect 182088 8842 182140 8848
rect 182088 7948 182140 7954
rect 182088 7890 182140 7896
rect 182100 7585 182128 7890
rect 182086 7576 182142 7585
rect 182086 7511 182142 7520
rect 182284 7449 182312 10200
rect 182744 10146 182772 10200
rect 182560 10118 182772 10146
rect 182560 9654 182588 10118
rect 182732 9988 182784 9994
rect 182732 9930 182784 9936
rect 182744 9654 182772 9930
rect 183204 9926 183232 10200
rect 183192 9920 183244 9926
rect 183192 9862 183244 9868
rect 182548 9648 182600 9654
rect 182548 9590 182600 9596
rect 182732 9648 182784 9654
rect 182732 9590 182784 9596
rect 182640 9512 182692 9518
rect 182640 9454 182692 9460
rect 182824 9512 182876 9518
rect 182824 9454 182876 9460
rect 182652 9042 182680 9454
rect 182640 9036 182692 9042
rect 182640 8978 182692 8984
rect 182836 8838 182864 9454
rect 183006 9344 183062 9353
rect 183006 9279 183062 9288
rect 182824 8832 182876 8838
rect 182824 8774 182876 8780
rect 183020 8430 183048 9279
rect 183664 8922 183692 10200
rect 183928 9716 183980 9722
rect 183928 9658 183980 9664
rect 183744 9512 183796 9518
rect 183744 9454 183796 9460
rect 183572 8906 183692 8922
rect 183560 8900 183692 8906
rect 183612 8894 183692 8900
rect 183560 8842 183612 8848
rect 183008 8424 183060 8430
rect 183008 8366 183060 8372
rect 182454 8120 182510 8129
rect 182454 8055 182510 8064
rect 183282 8120 183338 8129
rect 183756 8090 183784 9454
rect 183940 8498 183968 9658
rect 184032 9450 184060 10200
rect 184020 9444 184072 9450
rect 184020 9386 184072 9392
rect 184492 9330 184520 10200
rect 184308 9302 184520 9330
rect 184076 9276 184132 9296
rect 184076 9200 184132 9220
rect 183836 8492 183888 8498
rect 183836 8434 183888 8440
rect 183928 8492 183980 8498
rect 183928 8434 183980 8440
rect 184112 8492 184164 8498
rect 184112 8434 184164 8440
rect 183848 8378 183876 8434
rect 184124 8378 184152 8434
rect 183848 8350 184152 8378
rect 184076 8188 184132 8208
rect 184076 8112 184132 8132
rect 183282 8055 183338 8064
rect 183744 8084 183796 8090
rect 182468 7954 182496 8055
rect 182456 7948 182508 7954
rect 183296 7936 183324 8055
rect 183744 8026 183796 8032
rect 183560 7948 183612 7954
rect 183296 7908 183560 7936
rect 182456 7890 182508 7896
rect 183560 7890 183612 7896
rect 182548 7880 182600 7886
rect 182824 7880 182876 7886
rect 182600 7840 182772 7868
rect 182548 7822 182600 7828
rect 182640 7744 182692 7750
rect 182640 7686 182692 7692
rect 181994 7440 182050 7449
rect 181166 7375 181222 7384
rect 181536 7404 181588 7410
rect 181536 7346 181588 7352
rect 181812 7404 181864 7410
rect 181994 7375 182050 7384
rect 182270 7440 182326 7449
rect 182652 7410 182680 7686
rect 182744 7410 182772 7840
rect 182824 7822 182876 7828
rect 182836 7721 182864 7822
rect 183560 7812 183612 7818
rect 183560 7754 183612 7760
rect 183572 7721 183600 7754
rect 182822 7712 182878 7721
rect 182822 7647 182878 7656
rect 183558 7712 183614 7721
rect 183558 7647 183614 7656
rect 184308 7449 184336 9302
rect 184480 9172 184532 9178
rect 184480 9114 184532 9120
rect 184294 7440 184350 7449
rect 182270 7375 182326 7384
rect 182640 7404 182692 7410
rect 181812 7346 181864 7352
rect 182640 7346 182692 7352
rect 182732 7404 182784 7410
rect 184294 7375 184350 7384
rect 182732 7346 182784 7352
rect 177486 7304 177542 7313
rect 157064 7278 157116 7284
rect 156970 7032 157026 7041
rect 156970 6967 157026 6976
rect 156984 5681 157012 6967
rect 157076 6633 157104 7278
rect 157260 7262 157380 7290
rect 157062 6624 157118 6633
rect 157062 6559 157118 6568
rect 157154 6352 157210 6361
rect 157154 6287 157210 6296
rect 156970 5672 157026 5681
rect 156970 5607 157026 5616
rect 157062 5128 157118 5137
rect 157062 5063 157118 5072
rect 156970 4720 157026 4729
rect 156970 4655 157026 4664
rect 156786 4040 156842 4049
rect 156786 3975 156842 3984
rect 156696 3120 156748 3126
rect 156696 3062 156748 3068
rect 156602 1592 156658 1601
rect 156602 1527 156658 1536
rect 156800 1465 156828 3975
rect 156880 3596 156932 3602
rect 156880 3538 156932 3544
rect 156786 1456 156842 1465
rect 156786 1391 156842 1400
rect 156510 1320 156566 1329
rect 156510 1255 156566 1264
rect 156892 950 156920 3538
rect 156984 3126 157012 4655
rect 156972 3120 157024 3126
rect 156972 3062 157024 3068
rect 157076 2689 157104 5063
rect 157168 4842 157196 6287
rect 157260 5545 157288 7262
rect 177486 7239 177542 7248
rect 177854 7304 177910 7313
rect 177854 7239 177910 7248
rect 157246 5536 157302 5545
rect 157246 5471 157302 5480
rect 157168 4814 157288 4842
rect 157156 3528 157208 3534
rect 157156 3470 157208 3476
rect 157062 2680 157118 2689
rect 157062 2615 157118 2624
rect 157062 2544 157118 2553
rect 157168 2514 157196 3470
rect 157062 2479 157064 2488
rect 157116 2479 157118 2488
rect 157156 2508 157208 2514
rect 157064 2450 157116 2456
rect 157156 2450 157208 2456
rect 157260 1426 157288 4814
rect 161204 2984 161256 2990
rect 162676 2984 162728 2990
rect 161256 2944 161428 2972
rect 161204 2926 161256 2932
rect 157432 2848 157484 2854
rect 157432 2790 157484 2796
rect 158352 2848 158404 2854
rect 158352 2790 158404 2796
rect 158536 2848 158588 2854
rect 158536 2790 158588 2796
rect 157248 1420 157300 1426
rect 157248 1362 157300 1368
rect 156880 944 156932 950
rect 156524 870 156644 898
rect 156880 886 156932 892
rect 156418 776 156474 785
rect 156418 711 156474 720
rect 156236 468 156288 474
rect 156236 410 156288 416
rect 156524 338 156552 870
rect 156616 800 156644 870
rect 156984 870 157104 898
rect 156512 332 156564 338
rect 156512 274 156564 280
rect 156602 -400 156658 800
rect 156984 542 157012 870
rect 157076 800 157104 870
rect 157444 800 157472 2790
rect 157904 2638 158116 2666
rect 157904 2582 157932 2638
rect 157892 2576 157944 2582
rect 157892 2518 157944 2524
rect 157984 2576 158036 2582
rect 157984 2518 158036 2524
rect 157524 2508 157576 2514
rect 157524 2450 157576 2456
rect 156972 536 157024 542
rect 156972 478 157024 484
rect 157062 -400 157118 800
rect 157430 -400 157486 800
rect 157536 338 157564 2450
rect 157996 2378 158024 2518
rect 158088 2496 158116 2638
rect 158260 2508 158312 2514
rect 158088 2468 158260 2496
rect 158260 2450 158312 2456
rect 157984 2372 158036 2378
rect 157984 2314 158036 2320
rect 157812 836 157932 864
rect 157524 332 157576 338
rect 157524 274 157576 280
rect 157812 270 157840 836
rect 157904 800 157932 836
rect 158364 800 158392 2790
rect 158548 2009 158576 2790
rect 161032 2514 161244 2530
rect 161020 2508 161244 2514
rect 161072 2502 161244 2508
rect 161216 2496 161244 2502
rect 161296 2508 161348 2514
rect 161216 2468 161296 2496
rect 161020 2450 161072 2456
rect 161296 2450 161348 2456
rect 158812 2440 158864 2446
rect 158812 2382 158864 2388
rect 159088 2440 159140 2446
rect 159088 2382 159140 2388
rect 161112 2440 161164 2446
rect 161112 2382 161164 2388
rect 158534 2000 158590 2009
rect 158534 1935 158590 1944
rect 158718 2000 158774 2009
rect 158718 1935 158720 1944
rect 158772 1935 158774 1944
rect 158720 1906 158772 1912
rect 158824 800 158852 2382
rect 159100 1358 159128 2382
rect 160928 2304 160980 2310
rect 159454 2272 159510 2281
rect 159454 2207 159510 2216
rect 159730 2272 159786 2281
rect 160928 2246 160980 2252
rect 159730 2207 159786 2216
rect 159468 2106 159496 2207
rect 159364 2100 159416 2106
rect 159364 2042 159416 2048
rect 159456 2100 159508 2106
rect 159456 2042 159508 2048
rect 159376 1834 159404 2042
rect 159548 2032 159600 2038
rect 159548 1974 159600 1980
rect 159364 1828 159416 1834
rect 159364 1770 159416 1776
rect 159088 1352 159140 1358
rect 159088 1294 159140 1300
rect 159100 836 159220 864
rect 157800 264 157852 270
rect 157800 206 157852 212
rect 157890 -400 157946 800
rect 158350 -400 158406 800
rect 158810 -400 158866 800
rect 159100 202 159128 836
rect 159192 800 159220 836
rect 159088 196 159140 202
rect 159088 138 159140 144
rect 159178 -400 159234 800
rect 159272 332 159324 338
rect 159272 274 159324 280
rect 159284 241 159312 274
rect 159560 270 159588 1974
rect 159744 1970 159772 2207
rect 160834 2136 160890 2145
rect 160940 2106 160968 2246
rect 160834 2071 160836 2080
rect 160888 2071 160890 2080
rect 160928 2100 160980 2106
rect 160836 2042 160888 2048
rect 160928 2042 160980 2048
rect 159732 1964 159784 1970
rect 159732 1906 159784 1912
rect 159824 1964 159876 1970
rect 159824 1906 159876 1912
rect 159638 1592 159694 1601
rect 159638 1527 159694 1536
rect 159652 800 159680 1527
rect 159836 1494 159864 1906
rect 161124 1902 161152 2382
rect 160560 1896 160612 1902
rect 160560 1838 160612 1844
rect 160744 1896 160796 1902
rect 160744 1838 160796 1844
rect 161112 1896 161164 1902
rect 161112 1838 161164 1844
rect 161202 1864 161258 1873
rect 159824 1488 159876 1494
rect 159824 1430 159876 1436
rect 160100 1216 160152 1222
rect 160100 1158 160152 1164
rect 160112 800 160140 1158
rect 160572 950 160600 1838
rect 160652 1420 160704 1426
rect 160652 1362 160704 1368
rect 160468 944 160520 950
rect 160468 886 160520 892
rect 160560 944 160612 950
rect 160560 886 160612 892
rect 160480 800 160508 886
rect 159548 264 159600 270
rect 159270 232 159326 241
rect 159548 206 159600 212
rect 159270 167 159326 176
rect 159638 -400 159694 800
rect 160098 -400 160154 800
rect 160466 -400 160522 800
rect 160664 542 160692 1362
rect 160652 536 160704 542
rect 160652 478 160704 484
rect 160650 232 160706 241
rect 160756 202 160784 1838
rect 161202 1799 161258 1808
rect 161018 1592 161074 1601
rect 161216 1562 161244 1799
rect 161018 1527 161020 1536
rect 161072 1527 161074 1536
rect 161204 1556 161256 1562
rect 161020 1498 161072 1504
rect 161204 1498 161256 1504
rect 160848 836 160968 864
rect 160848 785 160876 836
rect 160940 800 160968 836
rect 161400 800 161428 2944
rect 162214 2952 162270 2961
rect 162596 2944 162676 2972
rect 162270 2910 162348 2938
rect 162214 2887 162270 2896
rect 161480 2848 161532 2854
rect 161480 2790 161532 2796
rect 161492 2446 161520 2790
rect 162214 2680 162270 2689
rect 162214 2615 162270 2624
rect 162032 2576 162084 2582
rect 162032 2518 162084 2524
rect 161480 2440 161532 2446
rect 161480 2382 161532 2388
rect 161572 2440 161624 2446
rect 161572 2382 161624 2388
rect 161584 1902 161612 2382
rect 161754 2272 161810 2281
rect 161754 2207 161810 2216
rect 161768 1902 161796 2207
rect 161572 1896 161624 1902
rect 161478 1864 161534 1873
rect 161572 1838 161624 1844
rect 161756 1896 161808 1902
rect 161756 1838 161808 1844
rect 161478 1799 161480 1808
rect 161532 1799 161534 1808
rect 161480 1770 161532 1776
rect 162044 1766 162072 2518
rect 162228 1970 162256 2615
rect 162216 1964 162268 1970
rect 162216 1906 162268 1912
rect 161940 1760 161992 1766
rect 161940 1702 161992 1708
rect 162032 1760 162084 1766
rect 162032 1702 162084 1708
rect 161768 836 161888 864
rect 160834 776 160890 785
rect 160834 711 160890 720
rect 160650 167 160652 176
rect 160704 167 160706 176
rect 160744 196 160796 202
rect 160652 138 160704 144
rect 160744 138 160796 144
rect 160926 -400 160982 800
rect 161386 -400 161442 800
rect 161768 474 161796 836
rect 161860 800 161888 836
rect 161756 468 161808 474
rect 161756 410 161808 416
rect 161846 -400 161902 800
rect 161952 796 161980 1702
rect 162124 1488 162176 1494
rect 162124 1430 162176 1436
rect 162032 1352 162084 1358
rect 162032 1294 162084 1300
rect 162044 950 162072 1294
rect 162136 1034 162164 1430
rect 162320 1222 162348 2910
rect 162490 2816 162546 2825
rect 162490 2751 162546 2760
rect 162504 2650 162532 2751
rect 162492 2644 162544 2650
rect 162492 2586 162544 2592
rect 162400 2508 162452 2514
rect 162400 2450 162452 2456
rect 162412 2258 162440 2450
rect 162412 2230 162532 2258
rect 162400 2100 162452 2106
rect 162400 2042 162452 2048
rect 162412 1358 162440 2042
rect 162504 1748 162532 2230
rect 162596 1884 162624 2944
rect 162676 2926 162728 2932
rect 162768 2984 162820 2990
rect 166724 2984 166776 2990
rect 162768 2926 162820 2932
rect 165342 2952 165398 2961
rect 162780 2514 162808 2926
rect 165342 2887 165398 2896
rect 165526 2952 165582 2961
rect 173808 2984 173860 2990
rect 167274 2952 167330 2961
rect 166724 2926 166776 2932
rect 165526 2887 165582 2896
rect 166264 2916 166316 2922
rect 165356 2854 165384 2887
rect 165068 2848 165120 2854
rect 163778 2816 163834 2825
rect 163778 2751 163834 2760
rect 164330 2816 164386 2825
rect 165068 2790 165120 2796
rect 165344 2848 165396 2854
rect 165344 2790 165396 2796
rect 164330 2751 164386 2760
rect 163044 2576 163096 2582
rect 163096 2524 163176 2530
rect 163044 2518 163176 2524
rect 162768 2508 162820 2514
rect 163056 2502 163176 2518
rect 163148 2496 163176 2502
rect 163228 2508 163280 2514
rect 163148 2468 163228 2496
rect 162768 2450 162820 2456
rect 163228 2450 163280 2456
rect 163688 2508 163740 2514
rect 163688 2450 163740 2456
rect 163700 2417 163728 2450
rect 162950 2408 163006 2417
rect 162950 2343 163006 2352
rect 163134 2408 163190 2417
rect 163134 2343 163190 2352
rect 163686 2408 163742 2417
rect 163686 2343 163742 2352
rect 162964 2020 162992 2343
rect 163148 2310 163176 2343
rect 163136 2304 163188 2310
rect 163136 2246 163188 2252
rect 163320 2304 163372 2310
rect 163320 2246 163372 2252
rect 163228 2032 163280 2038
rect 162964 1992 163228 2020
rect 163228 1974 163280 1980
rect 163044 1896 163096 1902
rect 162596 1856 163044 1884
rect 163044 1838 163096 1844
rect 162504 1720 162992 1748
rect 162492 1556 162544 1562
rect 162492 1498 162544 1504
rect 162504 1408 162532 1498
rect 162768 1420 162820 1426
rect 162504 1380 162768 1408
rect 162768 1362 162820 1368
rect 162400 1352 162452 1358
rect 162400 1294 162452 1300
rect 162308 1216 162360 1222
rect 162308 1158 162360 1164
rect 162768 1216 162820 1222
rect 162768 1158 162820 1164
rect 162860 1216 162912 1222
rect 162860 1158 162912 1164
rect 162136 1006 162440 1034
rect 162032 944 162084 950
rect 162032 886 162084 892
rect 162136 836 162256 864
rect 162136 796 162164 836
rect 162228 800 162256 836
rect 161952 768 162164 796
rect 162122 504 162178 513
rect 162122 439 162178 448
rect 162136 105 162164 439
rect 162122 96 162178 105
rect 162122 31 162178 40
rect 162214 -400 162270 800
rect 162306 776 162362 785
rect 162412 762 162440 1006
rect 162596 836 162716 864
rect 162490 776 162546 785
rect 162412 734 162490 762
rect 162306 711 162362 720
rect 162490 711 162546 720
rect 162320 241 162348 711
rect 162306 232 162362 241
rect 162306 167 162362 176
rect 162596 66 162624 836
rect 162688 800 162716 836
rect 162584 60 162636 66
rect 162584 2 162636 8
rect 162674 -400 162730 800
rect 162780 66 162808 1158
rect 162872 1018 162900 1158
rect 162964 1018 162992 1720
rect 162860 1012 162912 1018
rect 162860 954 162912 960
rect 162952 1012 163004 1018
rect 162952 954 163004 960
rect 163056 836 163176 864
rect 163056 134 163084 836
rect 163148 800 163176 836
rect 163044 128 163096 134
rect 163044 70 163096 76
rect 162768 60 162820 66
rect 162768 2 162820 8
rect 163134 -400 163190 800
rect 163226 504 163282 513
rect 163226 439 163282 448
rect 163240 134 163268 439
rect 163332 377 163360 2246
rect 163686 1864 163742 1873
rect 163596 1828 163648 1834
rect 163686 1799 163688 1808
rect 163596 1770 163648 1776
rect 163740 1799 163742 1808
rect 163688 1770 163740 1776
rect 163608 1426 163636 1770
rect 163688 1556 163740 1562
rect 163688 1498 163740 1504
rect 163596 1420 163648 1426
rect 163596 1362 163648 1368
rect 163424 870 163636 898
rect 163424 814 163452 870
rect 163412 808 163464 814
rect 163608 800 163636 870
rect 163412 750 163464 756
rect 163318 368 163374 377
rect 163318 303 163374 312
rect 163228 128 163280 134
rect 163228 70 163280 76
rect 163594 -400 163650 800
rect 163700 377 163728 1498
rect 163792 814 163820 2751
rect 164344 2650 164372 2751
rect 164332 2644 164384 2650
rect 164332 2586 164384 2592
rect 164436 2502 164924 2530
rect 164436 2446 164464 2502
rect 164424 2440 164476 2446
rect 164424 2382 164476 2388
rect 164896 2310 164924 2502
rect 164884 2304 164936 2310
rect 163884 2264 164188 2292
rect 163884 2145 163912 2264
rect 164160 2258 164188 2264
rect 164238 2272 164294 2281
rect 164160 2230 164238 2258
rect 164076 2204 164132 2224
rect 164238 2207 164294 2216
rect 164344 2230 164556 2258
rect 164884 2246 164936 2252
rect 163870 2136 163926 2145
rect 164076 2128 164132 2148
rect 164238 2136 164294 2145
rect 163870 2071 163926 2080
rect 164238 2071 164294 2080
rect 164252 1902 164280 2071
rect 164344 2038 164372 2230
rect 164528 2106 164556 2230
rect 164516 2100 164568 2106
rect 164516 2042 164568 2048
rect 164620 2060 164924 2088
rect 164332 2032 164384 2038
rect 164620 1986 164648 2060
rect 164332 1974 164384 1980
rect 164436 1958 164648 1986
rect 164712 1970 164832 1986
rect 164700 1964 164832 1970
rect 164240 1896 164292 1902
rect 163870 1864 163926 1873
rect 164240 1838 164292 1844
rect 163870 1799 163926 1808
rect 163884 1193 163912 1799
rect 164436 1714 164464 1958
rect 164752 1958 164832 1964
rect 164700 1906 164752 1912
rect 164344 1686 164464 1714
rect 164238 1592 164294 1601
rect 164238 1527 164294 1536
rect 163870 1184 163926 1193
rect 163870 1119 163926 1128
rect 164076 1116 164132 1136
rect 163870 1048 163926 1057
rect 164076 1040 164132 1060
rect 164252 1057 164280 1527
rect 164344 1358 164372 1686
rect 164514 1592 164570 1601
rect 164514 1527 164570 1536
rect 164528 1494 164556 1527
rect 164516 1488 164568 1494
rect 164516 1430 164568 1436
rect 164698 1456 164754 1465
rect 164698 1391 164754 1400
rect 164332 1352 164384 1358
rect 164712 1340 164740 1391
rect 164332 1294 164384 1300
rect 164436 1312 164740 1340
rect 164238 1048 164294 1057
rect 163870 983 163926 992
rect 164238 983 164294 992
rect 163884 898 163912 983
rect 163884 870 164004 898
rect 163780 808 163832 814
rect 163976 800 164004 870
rect 164436 800 164464 1312
rect 164804 932 164832 1958
rect 164896 1358 164924 2060
rect 164976 1556 165028 1562
rect 164976 1498 165028 1504
rect 164988 1426 165016 1498
rect 165080 1426 165108 2790
rect 165250 2680 165306 2689
rect 165434 2680 165490 2689
rect 165306 2638 165384 2666
rect 165250 2615 165306 2624
rect 165252 2032 165304 2038
rect 165252 1974 165304 1980
rect 165264 1494 165292 1974
rect 165252 1488 165304 1494
rect 165252 1430 165304 1436
rect 164976 1420 165028 1426
rect 164976 1362 165028 1368
rect 165068 1420 165120 1426
rect 165068 1362 165120 1368
rect 164884 1352 164936 1358
rect 164884 1294 164936 1300
rect 164804 921 165016 932
rect 164804 912 165030 921
rect 164804 904 164974 912
rect 164804 836 164924 864
rect 164974 847 165030 856
rect 163780 750 163832 756
rect 163686 368 163742 377
rect 163686 303 163742 312
rect 163962 -400 164018 800
rect 164422 -400 164478 800
rect 164804 746 164832 836
rect 164896 800 164924 836
rect 165356 800 165384 2638
rect 165540 2650 165568 2887
rect 166264 2858 166316 2864
rect 165434 2615 165490 2624
rect 165528 2644 165580 2650
rect 165448 2446 165476 2615
rect 165528 2586 165580 2592
rect 165436 2440 165488 2446
rect 165436 2382 165488 2388
rect 165894 2408 165950 2417
rect 165894 2343 165950 2352
rect 165620 2032 165672 2038
rect 165620 1974 165672 1980
rect 165712 2032 165764 2038
rect 165712 1974 165764 1980
rect 165436 1896 165488 1902
rect 165436 1838 165488 1844
rect 165526 1864 165582 1873
rect 165448 921 165476 1838
rect 165526 1799 165582 1808
rect 165540 1494 165568 1799
rect 165528 1488 165580 1494
rect 165528 1430 165580 1436
rect 165632 1000 165660 1974
rect 165724 1737 165752 1974
rect 165908 1737 165936 2343
rect 165710 1728 165766 1737
rect 165710 1663 165766 1672
rect 165894 1728 165950 1737
rect 165894 1663 165950 1672
rect 166080 1012 166132 1018
rect 165632 972 166080 1000
rect 166080 954 166132 960
rect 165434 912 165490 921
rect 165434 847 165490 856
rect 165632 836 165752 864
rect 164792 740 164844 746
rect 164792 682 164844 688
rect 164882 -400 164938 800
rect 165342 -400 165398 800
rect 165632 678 165660 836
rect 165724 800 165752 836
rect 166092 836 166212 864
rect 165620 672 165672 678
rect 165620 614 165672 620
rect 165710 -400 165766 800
rect 166092 649 166120 836
rect 166184 800 166212 836
rect 166078 640 166134 649
rect 166078 575 166134 584
rect 166170 -400 166226 800
rect 166276 678 166304 2858
rect 166736 2825 166764 2926
rect 167104 2910 167274 2938
rect 167104 2854 167132 2910
rect 167274 2887 167330 2896
rect 169482 2952 169538 2961
rect 169482 2887 169538 2896
rect 169758 2952 169814 2961
rect 169758 2887 169814 2896
rect 170034 2952 170090 2961
rect 170034 2887 170090 2896
rect 171690 2952 171746 2961
rect 180156 2984 180208 2990
rect 173808 2926 173860 2932
rect 174910 2952 174966 2961
rect 171690 2887 171746 2896
rect 171784 2916 171836 2922
rect 167092 2848 167144 2854
rect 166722 2816 166778 2825
rect 167092 2790 167144 2796
rect 168562 2816 168618 2825
rect 166722 2751 166778 2760
rect 168562 2751 168618 2760
rect 167274 2680 167330 2689
rect 167274 2615 167330 2624
rect 167734 2680 167790 2689
rect 167734 2615 167790 2624
rect 167288 2514 167316 2615
rect 167460 2576 167512 2582
rect 167460 2518 167512 2524
rect 167276 2508 167328 2514
rect 167276 2450 167328 2456
rect 167092 2304 167144 2310
rect 166998 2272 167054 2281
rect 167092 2246 167144 2252
rect 167184 2304 167236 2310
rect 167184 2246 167236 2252
rect 166998 2207 167054 2216
rect 166906 2136 166962 2145
rect 166906 2071 166962 2080
rect 166920 1358 166948 2071
rect 167012 1970 167040 2207
rect 167104 2106 167132 2246
rect 167092 2100 167144 2106
rect 167092 2042 167144 2048
rect 167196 2038 167224 2246
rect 167184 2032 167236 2038
rect 167184 1974 167236 1980
rect 167000 1964 167052 1970
rect 167000 1906 167052 1912
rect 167366 1456 167422 1465
rect 167366 1391 167422 1400
rect 167380 1358 167408 1391
rect 167472 1358 167500 2518
rect 167748 2514 167776 2615
rect 167736 2508 167788 2514
rect 167736 2450 167788 2456
rect 167552 2440 167604 2446
rect 167552 2382 167604 2388
rect 167564 2038 167592 2382
rect 168576 2106 168604 2751
rect 169116 2508 169168 2514
rect 169116 2450 169168 2456
rect 169300 2508 169352 2514
rect 169300 2450 169352 2456
rect 168654 2272 168710 2281
rect 168654 2207 168710 2216
rect 168668 2106 168696 2207
rect 168564 2100 168616 2106
rect 168564 2042 168616 2048
rect 168656 2100 168708 2106
rect 168656 2042 168708 2048
rect 167552 2032 167604 2038
rect 167552 1974 167604 1980
rect 168380 1896 168432 1902
rect 168432 1856 168788 1884
rect 168380 1838 168432 1844
rect 168104 1488 168156 1494
rect 168104 1430 168156 1436
rect 167920 1420 167972 1426
rect 167920 1362 167972 1368
rect 166908 1352 166960 1358
rect 166908 1294 166960 1300
rect 167368 1352 167420 1358
rect 167368 1294 167420 1300
rect 167460 1352 167512 1358
rect 167460 1294 167512 1300
rect 167012 882 167132 898
rect 167000 876 167132 882
rect 166552 836 166672 864
rect 166264 672 166316 678
rect 166264 614 166316 620
rect 166552 542 166580 836
rect 166644 800 166672 836
rect 167052 870 167132 876
rect 167000 818 167052 824
rect 167104 800 167132 870
rect 167380 870 167500 898
rect 166540 536 166592 542
rect 166540 478 166592 484
rect 166630 -400 166686 800
rect 166906 504 166962 513
rect 166906 439 166962 448
rect 166920 270 166948 439
rect 166908 264 166960 270
rect 166908 206 166960 212
rect 167090 -400 167146 800
rect 167380 542 167408 870
rect 167472 800 167500 870
rect 167932 800 167960 1362
rect 168116 1057 168144 1430
rect 168102 1048 168158 1057
rect 168102 983 168158 992
rect 168286 1048 168342 1057
rect 168286 983 168342 992
rect 168300 950 168328 983
rect 168288 944 168340 950
rect 168288 886 168340 892
rect 168392 870 168512 898
rect 168392 800 168420 870
rect 167368 536 167420 542
rect 167368 478 167420 484
rect 167458 -400 167514 800
rect 167918 -400 167974 800
rect 168378 -400 168434 800
rect 168484 134 168512 870
rect 168760 800 168788 1856
rect 169022 1728 169078 1737
rect 169022 1663 169078 1672
rect 169036 882 169064 1663
rect 169128 1018 169156 2450
rect 169312 1562 169340 2450
rect 169496 1902 169524 2887
rect 169666 2816 169722 2825
rect 169666 2751 169722 2760
rect 169680 1902 169708 2751
rect 169772 2582 169800 2887
rect 169760 2576 169812 2582
rect 169760 2518 169812 2524
rect 169758 2272 169814 2281
rect 169758 2207 169814 2216
rect 169484 1896 169536 1902
rect 169390 1864 169446 1873
rect 169484 1838 169536 1844
rect 169668 1896 169720 1902
rect 169668 1838 169720 1844
rect 169390 1799 169446 1808
rect 169300 1556 169352 1562
rect 169300 1498 169352 1504
rect 169404 1426 169432 1799
rect 169772 1766 169800 2207
rect 169944 1896 169996 1902
rect 169944 1838 169996 1844
rect 169760 1760 169812 1766
rect 169760 1702 169812 1708
rect 169956 1494 169984 1838
rect 170048 1562 170076 2887
rect 171138 2680 171194 2689
rect 171138 2615 171140 2624
rect 171192 2615 171194 2624
rect 171322 2680 171378 2689
rect 171704 2650 171732 2887
rect 171784 2858 171836 2864
rect 171322 2615 171378 2624
rect 171692 2644 171744 2650
rect 171140 2586 171192 2592
rect 171336 2417 171364 2615
rect 171692 2586 171744 2592
rect 171322 2408 171378 2417
rect 171322 2343 171378 2352
rect 171322 2136 171378 2145
rect 171322 2071 171378 2080
rect 171232 2032 171284 2038
rect 171232 1974 171284 1980
rect 170036 1556 170088 1562
rect 170036 1498 170088 1504
rect 169944 1488 169996 1494
rect 169944 1430 169996 1436
rect 171138 1456 171194 1465
rect 169392 1420 169444 1426
rect 171244 1426 171272 1974
rect 171336 1494 171364 2071
rect 171324 1488 171376 1494
rect 171324 1430 171376 1436
rect 171138 1391 171194 1400
rect 171232 1420 171284 1426
rect 169392 1362 169444 1368
rect 169116 1012 169168 1018
rect 169116 954 169168 960
rect 170954 912 171010 921
rect 169024 876 169076 882
rect 169024 818 169076 824
rect 169128 870 169248 898
rect 168472 128 168524 134
rect 168472 70 168524 76
rect 168746 -400 168802 800
rect 169128 785 169156 870
rect 169220 800 169248 870
rect 169588 870 169708 898
rect 169114 776 169170 785
rect 169114 711 169170 720
rect 169206 -400 169262 800
rect 169588 746 169616 870
rect 169680 800 169708 870
rect 170048 870 170168 898
rect 169576 740 169628 746
rect 169576 682 169628 688
rect 169666 -400 169722 800
rect 170048 270 170076 870
rect 170140 800 170168 870
rect 170416 870 170536 898
rect 170036 264 170088 270
rect 170036 206 170088 212
rect 170126 -400 170182 800
rect 170416 377 170444 870
rect 170508 800 170536 870
rect 170954 847 171010 856
rect 170968 800 170996 847
rect 171152 814 171180 1391
rect 171232 1362 171284 1368
rect 171796 1306 171824 2858
rect 173348 2848 173400 2854
rect 173254 2816 173310 2825
rect 173348 2790 173400 2796
rect 173254 2751 173310 2760
rect 171874 2000 171930 2009
rect 171874 1935 171930 1944
rect 171888 1902 171916 1935
rect 171876 1896 171928 1902
rect 171876 1838 171928 1844
rect 172980 1896 173032 1902
rect 172980 1838 173032 1844
rect 173072 1896 173124 1902
rect 173072 1838 173124 1844
rect 173162 1864 173218 1873
rect 172992 1766 173020 1838
rect 172428 1760 172480 1766
rect 172428 1702 172480 1708
rect 172980 1760 173032 1766
rect 172980 1702 173032 1708
rect 172440 1426 172468 1702
rect 173084 1494 173112 1838
rect 173162 1799 173218 1808
rect 173072 1488 173124 1494
rect 173072 1430 173124 1436
rect 172428 1420 172480 1426
rect 172428 1362 172480 1368
rect 171796 1278 171916 1306
rect 171336 870 171456 898
rect 171140 808 171192 814
rect 170402 368 170458 377
rect 170402 303 170458 312
rect 170494 -400 170550 800
rect 170954 -400 171010 800
rect 171140 750 171192 756
rect 171336 610 171364 870
rect 171428 800 171456 870
rect 171888 800 171916 1278
rect 172704 944 172756 950
rect 172164 870 172284 898
rect 172704 886 172756 892
rect 171324 604 171376 610
rect 171324 546 171376 552
rect 171414 -400 171470 800
rect 171874 -400 171930 800
rect 172164 66 172192 870
rect 172256 800 172284 870
rect 172716 800 172744 886
rect 173176 800 173204 1799
rect 173268 1426 173296 2751
rect 173360 2514 173388 2790
rect 173348 2508 173400 2514
rect 173348 2450 173400 2456
rect 173820 1902 173848 2926
rect 174910 2887 174966 2896
rect 175922 2952 175978 2961
rect 175922 2887 175978 2896
rect 176474 2952 176530 2961
rect 176750 2952 176806 2961
rect 176474 2887 176476 2896
rect 174924 2514 174952 2887
rect 175278 2816 175334 2825
rect 175278 2751 175334 2760
rect 173992 2508 174044 2514
rect 173992 2450 174044 2456
rect 174912 2508 174964 2514
rect 174912 2450 174964 2456
rect 174004 2106 174032 2450
rect 173992 2100 174044 2106
rect 173992 2042 174044 2048
rect 173624 1896 173676 1902
rect 173624 1838 173676 1844
rect 173808 1896 173860 1902
rect 173808 1838 173860 1844
rect 173636 1494 173664 1838
rect 174912 1556 174964 1562
rect 174912 1498 174964 1504
rect 173624 1488 173676 1494
rect 173624 1430 173676 1436
rect 174452 1488 174504 1494
rect 174452 1430 174504 1436
rect 173256 1420 173308 1426
rect 173256 1362 173308 1368
rect 173348 1420 173400 1426
rect 173532 1420 173584 1426
rect 173400 1380 173532 1408
rect 173348 1362 173400 1368
rect 173532 1362 173584 1368
rect 173544 870 173664 898
rect 172152 60 172204 66
rect 172152 2 172204 8
rect 172242 -400 172298 800
rect 172702 -400 172758 800
rect 173162 -400 173218 800
rect 173544 474 173572 870
rect 173636 800 173664 870
rect 173912 870 174032 898
rect 173532 468 173584 474
rect 173532 410 173584 416
rect 173622 -400 173678 800
rect 173912 678 173940 870
rect 174004 800 174032 870
rect 174464 800 174492 1430
rect 174924 800 174952 1498
rect 175292 1442 175320 2751
rect 175936 2650 175964 2887
rect 176528 2887 176530 2896
rect 176660 2916 176712 2922
rect 176476 2858 176528 2864
rect 176750 2887 176806 2896
rect 177854 2952 177910 2961
rect 180156 2926 180208 2932
rect 180340 2984 180392 2990
rect 180340 2926 180392 2932
rect 180430 2952 180486 2961
rect 177854 2887 177910 2896
rect 176660 2858 176712 2864
rect 176566 2816 176622 2825
rect 176566 2751 176622 2760
rect 175740 2644 175792 2650
rect 175740 2586 175792 2592
rect 175924 2644 175976 2650
rect 175924 2586 175976 2592
rect 175752 2106 175780 2586
rect 175832 2508 175884 2514
rect 175832 2450 175884 2456
rect 175740 2100 175792 2106
rect 175740 2042 175792 2048
rect 175740 1556 175792 1562
rect 175740 1498 175792 1504
rect 175292 1414 175412 1442
rect 175384 1358 175412 1414
rect 175372 1352 175424 1358
rect 175372 1294 175424 1300
rect 175188 1284 175240 1290
rect 175188 1226 175240 1232
rect 175464 1284 175516 1290
rect 175464 1226 175516 1232
rect 175200 1170 175228 1226
rect 175476 1170 175504 1226
rect 175200 1142 175504 1170
rect 175292 882 175412 898
rect 175280 876 175412 882
rect 175332 870 175412 876
rect 175280 818 175332 824
rect 175384 800 175412 870
rect 175752 800 175780 1498
rect 175844 882 175872 2450
rect 176292 2440 176344 2446
rect 176290 2408 176292 2417
rect 176344 2408 176346 2417
rect 176290 2343 176346 2352
rect 176198 2272 176254 2281
rect 176254 2230 176332 2258
rect 176198 2207 176254 2216
rect 176304 1902 176332 2230
rect 176476 2032 176528 2038
rect 176476 1974 176528 1980
rect 176200 1896 176252 1902
rect 176200 1838 176252 1844
rect 176292 1896 176344 1902
rect 176292 1838 176344 1844
rect 176016 1760 176068 1766
rect 176014 1728 176016 1737
rect 176108 1760 176160 1766
rect 176068 1728 176070 1737
rect 176108 1702 176160 1708
rect 176014 1663 176070 1672
rect 176120 1426 176148 1702
rect 176108 1420 176160 1426
rect 176108 1362 176160 1368
rect 175832 876 175884 882
rect 175832 818 175884 824
rect 176212 800 176240 1838
rect 176488 1222 176516 1974
rect 176580 1562 176608 2751
rect 176568 1556 176620 1562
rect 176568 1498 176620 1504
rect 176476 1216 176528 1222
rect 176476 1158 176528 1164
rect 176672 800 176700 2858
rect 176764 2582 176792 2887
rect 176752 2576 176804 2582
rect 176752 2518 176804 2524
rect 177028 2508 177080 2514
rect 177080 2468 177160 2496
rect 177028 2450 177080 2456
rect 177026 2272 177082 2281
rect 177026 2207 177082 2216
rect 176844 1964 176896 1970
rect 176844 1906 176896 1912
rect 176856 1494 176884 1906
rect 176844 1488 176896 1494
rect 176844 1430 176896 1436
rect 177040 800 177068 2207
rect 177132 1873 177160 2468
rect 177764 2304 177816 2310
rect 177764 2246 177816 2252
rect 177776 2106 177804 2246
rect 177868 2106 177896 2887
rect 179236 2848 179288 2854
rect 179236 2790 179288 2796
rect 178132 2644 178184 2650
rect 178132 2586 178184 2592
rect 177764 2100 177816 2106
rect 177764 2042 177816 2048
rect 177856 2100 177908 2106
rect 177856 2042 177908 2048
rect 177118 1864 177174 1873
rect 177118 1799 177174 1808
rect 178144 1426 178172 2586
rect 178314 2136 178370 2145
rect 178314 2071 178370 2080
rect 178224 2032 178276 2038
rect 178224 1974 178276 1980
rect 178236 1902 178264 1974
rect 178224 1896 178276 1902
rect 178224 1838 178276 1844
rect 178328 1562 178356 2071
rect 178316 1556 178368 1562
rect 178316 1498 178368 1504
rect 177488 1420 177540 1426
rect 177488 1362 177540 1368
rect 178132 1420 178184 1426
rect 178132 1362 178184 1368
rect 177500 800 177528 1362
rect 178776 1216 178828 1222
rect 178776 1158 178828 1164
rect 177868 870 177988 898
rect 173900 672 173952 678
rect 173900 614 173952 620
rect 173990 -400 174046 800
rect 174450 -400 174506 800
rect 174910 -400 174966 800
rect 175370 -400 175426 800
rect 175738 -400 175794 800
rect 176198 -400 176254 800
rect 176658 -400 176714 800
rect 177026 -400 177082 800
rect 177486 -400 177542 800
rect 177868 406 177896 870
rect 177960 800 177988 870
rect 178328 870 178448 898
rect 177856 400 177908 406
rect 177856 342 177908 348
rect 177946 -400 178002 800
rect 178328 338 178356 870
rect 178420 800 178448 870
rect 178788 800 178816 1158
rect 179248 800 179276 2790
rect 179510 2408 179566 2417
rect 179510 2343 179566 2352
rect 179524 1902 179552 2343
rect 179604 2304 179656 2310
rect 179604 2246 179656 2252
rect 179616 2106 179644 2246
rect 179604 2100 179656 2106
rect 179604 2042 179656 2048
rect 179328 1896 179380 1902
rect 179328 1838 179380 1844
rect 179512 1896 179564 1902
rect 179512 1838 179564 1844
rect 179340 1562 179368 1838
rect 179328 1556 179380 1562
rect 179328 1498 179380 1504
rect 179616 870 179736 898
rect 178316 332 178368 338
rect 178316 274 178368 280
rect 178406 -400 178462 800
rect 178774 -400 178830 800
rect 179234 -400 179290 800
rect 179616 202 179644 870
rect 179708 800 179736 870
rect 180168 800 180196 2926
rect 180352 2038 180380 2926
rect 180430 2887 180432 2896
rect 180484 2887 180486 2896
rect 184204 2916 184256 2922
rect 180432 2858 180484 2864
rect 184204 2858 184256 2864
rect 184076 2748 184132 2768
rect 184076 2672 184132 2692
rect 181076 2508 181128 2514
rect 181076 2450 181128 2456
rect 180340 2032 180392 2038
rect 180340 1974 180392 1980
rect 181088 1970 181116 2450
rect 182546 2408 182602 2417
rect 181260 2372 181312 2378
rect 182546 2343 182548 2352
rect 181260 2314 181312 2320
rect 182600 2343 182602 2352
rect 182548 2314 182600 2320
rect 181076 1964 181128 1970
rect 181076 1906 181128 1912
rect 180708 1896 180760 1902
rect 180708 1838 180760 1844
rect 180720 1442 180748 1838
rect 180720 1414 181024 1442
rect 181272 1426 181300 2314
rect 181994 2136 182050 2145
rect 181994 2071 181996 2080
rect 182048 2071 182050 2080
rect 181996 2042 182048 2048
rect 183744 1896 183796 1902
rect 183374 1864 183430 1873
rect 181628 1828 181680 1834
rect 183374 1799 183430 1808
rect 183480 1844 183744 1850
rect 183480 1838 183796 1844
rect 183480 1822 183784 1838
rect 181628 1770 181680 1776
rect 181350 1728 181406 1737
rect 181350 1663 181406 1672
rect 180524 1352 180576 1358
rect 180524 1294 180576 1300
rect 180536 800 180564 1294
rect 180996 800 181024 1414
rect 181260 1420 181312 1426
rect 181260 1362 181312 1368
rect 181364 1222 181392 1663
rect 181640 1222 181668 1770
rect 182272 1556 182324 1562
rect 182324 1516 182772 1544
rect 182272 1498 182324 1504
rect 181352 1216 181404 1222
rect 181352 1158 181404 1164
rect 181628 1216 181680 1222
rect 181628 1158 181680 1164
rect 182272 1216 182324 1222
rect 182272 1158 182324 1164
rect 181534 1048 181590 1057
rect 181534 983 181590 992
rect 181548 950 181576 983
rect 181444 944 181496 950
rect 181444 886 181496 892
rect 181536 944 181588 950
rect 181536 886 181588 892
rect 181456 800 181484 886
rect 181812 876 181864 882
rect 181864 836 181944 864
rect 181812 818 181864 824
rect 181916 800 181944 836
rect 182284 800 182312 1158
rect 182744 800 182772 1516
rect 183388 1442 183416 1799
rect 183480 1766 183508 1822
rect 183468 1760 183520 1766
rect 183468 1702 183520 1708
rect 184076 1660 184132 1680
rect 183558 1592 183614 1601
rect 184076 1584 184132 1604
rect 183558 1527 183560 1536
rect 183612 1527 183614 1536
rect 183560 1498 183612 1504
rect 184216 1442 184244 2858
rect 184388 2644 184440 2650
rect 184388 2586 184440 2592
rect 183388 1414 183692 1442
rect 183192 1352 183244 1358
rect 183192 1294 183244 1300
rect 183204 800 183232 1294
rect 183664 800 183692 1414
rect 184032 1414 184244 1442
rect 184032 800 184060 1414
rect 184400 898 184428 2586
rect 184492 2446 184520 9114
rect 184952 9058 184980 10200
rect 184572 9036 184624 9042
rect 184952 9030 185072 9058
rect 184572 8978 184624 8984
rect 184584 2514 184612 8978
rect 184848 8968 184900 8974
rect 184848 8910 184900 8916
rect 184940 8968 184992 8974
rect 184940 8910 184992 8916
rect 184664 8628 184716 8634
rect 184664 8570 184716 8576
rect 184676 7818 184704 8570
rect 184756 8492 184808 8498
rect 184756 8434 184808 8440
rect 184664 7812 184716 7818
rect 184664 7754 184716 7760
rect 184572 2508 184624 2514
rect 184572 2450 184624 2456
rect 184480 2440 184532 2446
rect 184480 2382 184532 2388
rect 184768 1562 184796 8434
rect 184860 8090 184888 8910
rect 184952 8566 184980 8910
rect 184940 8560 184992 8566
rect 184940 8502 184992 8508
rect 184848 8084 184900 8090
rect 184848 8026 184900 8032
rect 184940 8084 184992 8090
rect 184940 8026 184992 8032
rect 184848 7812 184900 7818
rect 184848 7754 184900 7760
rect 184860 2106 184888 7754
rect 184952 7478 184980 8026
rect 185044 7857 185072 9030
rect 185320 8265 185348 10200
rect 185676 10192 185728 10198
rect 185780 10146 185808 10200
rect 185728 10140 185808 10146
rect 185676 10134 185808 10140
rect 185688 10118 185808 10134
rect 186240 9194 186268 10200
rect 186148 9166 186268 9194
rect 186148 8537 186176 9166
rect 186228 9036 186280 9042
rect 186228 8978 186280 8984
rect 186134 8528 186190 8537
rect 186134 8463 186190 8472
rect 185492 8424 185544 8430
rect 185492 8366 185544 8372
rect 185306 8256 185362 8265
rect 185306 8191 185362 8200
rect 185030 7848 185086 7857
rect 185030 7783 185086 7792
rect 185398 7576 185454 7585
rect 185398 7511 185454 7520
rect 184940 7472 184992 7478
rect 184940 7414 184992 7420
rect 185124 2644 185176 2650
rect 185124 2586 185176 2592
rect 185136 2378 185164 2586
rect 184940 2372 184992 2378
rect 184940 2314 184992 2320
rect 185124 2372 185176 2378
rect 185124 2314 185176 2320
rect 184952 2281 184980 2314
rect 184938 2272 184994 2281
rect 184938 2207 184994 2216
rect 185412 2106 185440 7511
rect 184848 2100 184900 2106
rect 184848 2042 184900 2048
rect 185400 2100 185452 2106
rect 185400 2042 185452 2048
rect 184940 1896 184992 1902
rect 184940 1838 184992 1844
rect 184756 1556 184808 1562
rect 184756 1498 184808 1504
rect 184400 870 184520 898
rect 184492 800 184520 870
rect 184952 800 184980 1838
rect 185308 1760 185360 1766
rect 185308 1702 185360 1708
rect 185320 800 185348 1702
rect 185504 1562 185532 8366
rect 185676 2576 185728 2582
rect 185676 2518 185728 2524
rect 186042 2544 186098 2553
rect 185688 2417 185716 2518
rect 185952 2508 186004 2514
rect 186042 2479 186098 2488
rect 185952 2450 186004 2456
rect 185674 2408 185730 2417
rect 185674 2343 185730 2352
rect 185768 1828 185820 1834
rect 185768 1770 185820 1776
rect 185492 1556 185544 1562
rect 185492 1498 185544 1504
rect 185780 800 185808 1770
rect 185964 1766 185992 2450
rect 186056 2446 186084 2479
rect 186044 2440 186096 2446
rect 186044 2382 186096 2388
rect 186134 2136 186190 2145
rect 186134 2071 186190 2080
rect 186044 1964 186096 1970
rect 186044 1906 186096 1912
rect 186056 1873 186084 1906
rect 186042 1864 186098 1873
rect 186042 1799 186098 1808
rect 185952 1760 186004 1766
rect 185952 1702 186004 1708
rect 186148 1494 186176 2071
rect 186240 2038 186268 8978
rect 186596 2372 186648 2378
rect 186596 2314 186648 2320
rect 186318 2272 186374 2281
rect 186318 2207 186374 2216
rect 186332 2106 186360 2207
rect 186410 2136 186466 2145
rect 186320 2100 186372 2106
rect 186410 2071 186412 2080
rect 186320 2042 186372 2048
rect 186464 2071 186466 2080
rect 186412 2042 186464 2048
rect 186608 2038 186636 2314
rect 186228 2032 186280 2038
rect 186228 1974 186280 1980
rect 186596 2032 186648 2038
rect 186596 1974 186648 1980
rect 186320 1828 186372 1834
rect 186320 1770 186372 1776
rect 186332 1494 186360 1770
rect 186700 1578 186728 10200
rect 187068 10062 187096 10200
rect 187056 10056 187108 10062
rect 187056 9998 187108 10004
rect 187424 9716 187476 9722
rect 187424 9658 187476 9664
rect 187056 2984 187108 2990
rect 187056 2926 187108 2932
rect 186872 2576 186924 2582
rect 186872 2518 186924 2524
rect 186608 1550 186728 1578
rect 186136 1488 186188 1494
rect 186136 1430 186188 1436
rect 186320 1488 186372 1494
rect 186320 1430 186372 1436
rect 186228 1352 186280 1358
rect 186228 1294 186280 1300
rect 186240 800 186268 1294
rect 186608 1290 186636 1550
rect 186884 1426 186912 2518
rect 186688 1420 186740 1426
rect 186688 1362 186740 1368
rect 186872 1420 186924 1426
rect 186872 1362 186924 1368
rect 186596 1284 186648 1290
rect 186596 1226 186648 1232
rect 186700 800 186728 1362
rect 187068 800 187096 2926
rect 187436 2446 187464 9658
rect 187528 8974 187556 10200
rect 187884 9104 187936 9110
rect 187884 9046 187936 9052
rect 187516 8968 187568 8974
rect 187516 8910 187568 8916
rect 187896 8566 187924 9046
rect 187884 8560 187936 8566
rect 187884 8502 187936 8508
rect 187884 7948 187936 7954
rect 187884 7890 187936 7896
rect 187424 2440 187476 2446
rect 187424 2382 187476 2388
rect 187514 2408 187570 2417
rect 187514 2343 187570 2352
rect 187528 2310 187556 2343
rect 187332 2304 187384 2310
rect 187332 2246 187384 2252
rect 187516 2304 187568 2310
rect 187516 2246 187568 2252
rect 187344 2145 187372 2246
rect 187330 2136 187386 2145
rect 187330 2071 187386 2080
rect 187700 1964 187752 1970
rect 187700 1906 187752 1912
rect 187148 1420 187200 1426
rect 187148 1362 187200 1368
rect 187160 1306 187188 1362
rect 187160 1278 187556 1306
rect 187528 800 187556 1278
rect 187712 1034 187740 1906
rect 187896 1562 187924 7890
rect 187988 7546 188016 10200
rect 188448 8498 188476 10200
rect 188436 8492 188488 8498
rect 188436 8434 188488 8440
rect 188068 8424 188120 8430
rect 188068 8366 188120 8372
rect 187976 7540 188028 7546
rect 187976 7482 188028 7488
rect 187884 1556 187936 1562
rect 187884 1498 187936 1504
rect 187712 1006 188016 1034
rect 187988 800 188016 1006
rect 188080 814 188108 8366
rect 188816 7478 188844 10200
rect 188988 9512 189040 9518
rect 188988 9454 189040 9460
rect 188896 8356 188948 8362
rect 188896 8298 188948 8304
rect 188804 7472 188856 7478
rect 188804 7414 188856 7420
rect 188908 1494 188936 8298
rect 189000 1562 189028 9454
rect 189172 7812 189224 7818
rect 189172 7754 189224 7760
rect 189184 7478 189212 7754
rect 189172 7472 189224 7478
rect 189172 7414 189224 7420
rect 189276 2106 189304 10200
rect 189448 9512 189500 9518
rect 189448 9454 189500 9460
rect 189356 9036 189408 9042
rect 189356 8978 189408 8984
rect 189368 2582 189396 8978
rect 189460 8090 189488 9454
rect 189736 8906 189764 10200
rect 190196 9586 190224 10200
rect 190184 9580 190236 9586
rect 190184 9522 190236 9528
rect 189724 8900 189776 8906
rect 189724 8842 189776 8848
rect 190564 8294 190592 10200
rect 190736 8900 190788 8906
rect 190736 8842 190788 8848
rect 190644 8424 190696 8430
rect 190644 8366 190696 8372
rect 190552 8288 190604 8294
rect 190552 8230 190604 8236
rect 189448 8084 189500 8090
rect 189448 8026 189500 8032
rect 190552 8084 190604 8090
rect 190552 8026 190604 8032
rect 190564 7954 190592 8026
rect 190552 7948 190604 7954
rect 190552 7890 190604 7896
rect 190460 2848 190512 2854
rect 190460 2790 190512 2796
rect 189356 2576 189408 2582
rect 189356 2518 189408 2524
rect 190184 2576 190236 2582
rect 190184 2518 190236 2524
rect 189724 2508 189776 2514
rect 189724 2450 189776 2456
rect 189264 2100 189316 2106
rect 189264 2042 189316 2048
rect 189448 2032 189500 2038
rect 189448 1974 189500 1980
rect 189460 1873 189488 1974
rect 189446 1864 189502 1873
rect 189264 1828 189316 1834
rect 189446 1799 189502 1808
rect 189264 1770 189316 1776
rect 188988 1556 189040 1562
rect 188988 1498 189040 1504
rect 188804 1488 188856 1494
rect 188804 1430 188856 1436
rect 188896 1488 188948 1494
rect 188896 1430 188948 1436
rect 188436 1420 188488 1426
rect 188436 1362 188488 1368
rect 188068 808 188120 814
rect 179604 196 179656 202
rect 179604 138 179656 144
rect 179694 -400 179750 800
rect 180154 -400 180210 800
rect 180522 -400 180578 800
rect 180982 -400 181038 800
rect 181442 -400 181498 800
rect 181902 -400 181958 800
rect 182270 -400 182326 800
rect 182730 -400 182786 800
rect 183190 -400 183246 800
rect 183650 -400 183706 800
rect 184018 -400 184074 800
rect 184478 -400 184534 800
rect 184938 -400 184994 800
rect 185306 -400 185362 800
rect 185766 -400 185822 800
rect 186226 -400 186282 800
rect 186686 -400 186742 800
rect 187054 -400 187110 800
rect 187514 -400 187570 800
rect 187974 -400 188030 800
rect 188448 800 188476 1362
rect 188816 800 188844 1430
rect 189276 800 189304 1770
rect 189736 800 189764 2450
rect 189814 2272 189870 2281
rect 189814 2207 189870 2216
rect 189828 1766 189856 2207
rect 189816 1760 189868 1766
rect 189816 1702 189868 1708
rect 190196 800 190224 2518
rect 190472 1902 190500 2790
rect 190552 2508 190604 2514
rect 190552 2450 190604 2456
rect 190460 1896 190512 1902
rect 190460 1838 190512 1844
rect 190564 800 190592 2450
rect 190656 1902 190684 8366
rect 190748 2514 190776 8842
rect 191024 8566 191052 10200
rect 191104 9920 191156 9926
rect 191104 9862 191156 9868
rect 191116 9654 191144 9862
rect 191104 9648 191156 9654
rect 191104 9590 191156 9596
rect 191196 9444 191248 9450
rect 191196 9386 191248 9392
rect 191208 8634 191236 9386
rect 191484 8974 191512 10200
rect 191944 9722 191972 10200
rect 191932 9716 191984 9722
rect 191932 9658 191984 9664
rect 191932 9376 191984 9382
rect 191932 9318 191984 9324
rect 191944 9042 191972 9318
rect 192116 9172 192168 9178
rect 192116 9114 192168 9120
rect 191932 9036 191984 9042
rect 191932 8978 191984 8984
rect 191472 8968 191524 8974
rect 191472 8910 191524 8916
rect 191196 8628 191248 8634
rect 191196 8570 191248 8576
rect 191012 8560 191064 8566
rect 191012 8502 191064 8508
rect 192128 8498 192156 9114
rect 192312 8974 192340 10200
rect 192668 9512 192720 9518
rect 192668 9454 192720 9460
rect 192300 8968 192352 8974
rect 192300 8910 192352 8916
rect 192116 8492 192168 8498
rect 192116 8434 192168 8440
rect 191654 7984 191710 7993
rect 191654 7919 191656 7928
rect 191708 7919 191710 7928
rect 191656 7890 191708 7896
rect 192680 7177 192708 9454
rect 192772 8922 192800 10200
rect 193232 10146 193260 10200
rect 193232 10118 193352 10146
rect 192772 8894 192892 8922
rect 192760 7948 192812 7954
rect 192760 7890 192812 7896
rect 192666 7168 192722 7177
rect 192666 7103 192722 7112
rect 192300 2848 192352 2854
rect 192300 2790 192352 2796
rect 190736 2508 190788 2514
rect 190736 2450 190788 2456
rect 191012 2372 191064 2378
rect 191012 2314 191064 2320
rect 190644 1896 190696 1902
rect 190644 1838 190696 1844
rect 191024 800 191052 2314
rect 191472 1964 191524 1970
rect 191472 1906 191524 1912
rect 191932 1964 191984 1970
rect 191932 1906 191984 1912
rect 191380 1556 191432 1562
rect 191380 1498 191432 1504
rect 191392 1358 191420 1498
rect 191380 1352 191432 1358
rect 191380 1294 191432 1300
rect 191484 800 191512 1906
rect 191944 800 191972 1906
rect 192312 800 192340 2790
rect 192772 2650 192800 7890
rect 192864 7886 192892 8894
rect 192852 7880 192904 7886
rect 192852 7822 192904 7828
rect 192944 7812 192996 7818
rect 192944 7754 192996 7760
rect 192760 2644 192812 2650
rect 192760 2586 192812 2592
rect 192760 2440 192812 2446
rect 192760 2382 192812 2388
rect 192668 2372 192720 2378
rect 192668 2314 192720 2320
rect 192680 2145 192708 2314
rect 192666 2136 192722 2145
rect 192666 2071 192722 2080
rect 192772 800 192800 2382
rect 192956 2106 192984 7754
rect 193220 2508 193272 2514
rect 193220 2450 193272 2456
rect 192944 2100 192996 2106
rect 192944 2042 192996 2048
rect 193232 800 193260 2450
rect 193324 2310 193352 10118
rect 193600 3754 193628 10200
rect 193864 8424 193916 8430
rect 193864 8366 193916 8372
rect 193508 3726 193628 3754
rect 193508 2378 193536 3726
rect 193588 2984 193640 2990
rect 193588 2926 193640 2932
rect 193496 2372 193548 2378
rect 193496 2314 193548 2320
rect 193312 2304 193364 2310
rect 193312 2246 193364 2252
rect 193310 2000 193366 2009
rect 193310 1935 193366 1944
rect 193324 1902 193352 1935
rect 193312 1896 193364 1902
rect 193312 1838 193364 1844
rect 193324 1426 193352 1838
rect 193312 1420 193364 1426
rect 193312 1362 193364 1368
rect 193600 800 193628 2926
rect 193876 2650 193904 8366
rect 194060 2650 194088 10200
rect 194520 9586 194548 10200
rect 194508 9580 194560 9586
rect 194508 9522 194560 9528
rect 194232 9512 194284 9518
rect 194232 9454 194284 9460
rect 194244 8634 194272 9454
rect 194876 8968 194928 8974
rect 194876 8910 194928 8916
rect 194232 8628 194284 8634
rect 194232 8570 194284 8576
rect 194508 8288 194560 8294
rect 194508 8230 194560 8236
rect 193864 2644 193916 2650
rect 193864 2586 193916 2592
rect 194048 2644 194100 2650
rect 194048 2586 194100 2592
rect 194048 2508 194100 2514
rect 194048 2450 194100 2456
rect 194060 800 194088 2450
rect 194520 800 194548 8230
rect 194888 7313 194916 8910
rect 194980 8498 195008 10200
rect 195152 10124 195204 10130
rect 195152 10066 195204 10072
rect 195164 9586 195192 10066
rect 195152 9580 195204 9586
rect 195152 9522 195204 9528
rect 195060 9444 195112 9450
rect 195060 9386 195112 9392
rect 194968 8492 195020 8498
rect 194968 8434 195020 8440
rect 194968 7948 195020 7954
rect 194968 7890 195020 7896
rect 194874 7304 194930 7313
rect 194874 7239 194930 7248
rect 194692 2848 194744 2854
rect 194692 2790 194744 2796
rect 194704 1970 194732 2790
rect 194980 2650 195008 7890
rect 195072 2650 195100 9386
rect 195348 8974 195376 10200
rect 195336 8968 195388 8974
rect 195336 8910 195388 8916
rect 195336 8084 195388 8090
rect 195336 8026 195388 8032
rect 194968 2644 195020 2650
rect 194968 2586 195020 2592
rect 195060 2644 195112 2650
rect 195060 2586 195112 2592
rect 195060 2100 195112 2106
rect 195060 2042 195112 2048
rect 194692 1964 194744 1970
rect 194692 1906 194744 1912
rect 194968 1556 195020 1562
rect 194968 1498 195020 1504
rect 194980 800 195008 1498
rect 195072 1426 195100 2042
rect 195152 1760 195204 1766
rect 195152 1702 195204 1708
rect 195164 1426 195192 1702
rect 195060 1420 195112 1426
rect 195060 1362 195112 1368
rect 195152 1420 195204 1426
rect 195152 1362 195204 1368
rect 195348 800 195376 8026
rect 195808 7886 195836 10200
rect 196268 9654 196296 10200
rect 196256 9648 196308 9654
rect 196256 9590 196308 9596
rect 196440 9036 196492 9042
rect 196440 8978 196492 8984
rect 196256 8560 196308 8566
rect 196256 8502 196308 8508
rect 195796 7880 195848 7886
rect 195796 7822 195848 7828
rect 195888 2916 195940 2922
rect 195888 2858 195940 2864
rect 195900 2106 195928 2858
rect 195888 2100 195940 2106
rect 195888 2042 195940 2048
rect 195796 1284 195848 1290
rect 195796 1226 195848 1232
rect 195808 800 195836 1226
rect 196268 800 196296 8502
rect 196452 2650 196480 8978
rect 196728 7478 196756 10200
rect 197096 8106 197124 10200
rect 197360 9512 197412 9518
rect 197360 9454 197412 9460
rect 197372 9178 197400 9454
rect 197360 9172 197412 9178
rect 197360 9114 197412 9120
rect 197268 9036 197320 9042
rect 197268 8978 197320 8984
rect 197004 8078 197124 8106
rect 196716 7472 196768 7478
rect 196716 7414 196768 7420
rect 197004 7410 197032 8078
rect 197084 7948 197136 7954
rect 197084 7890 197136 7896
rect 196992 7404 197044 7410
rect 196992 7346 197044 7352
rect 196900 2984 196952 2990
rect 196900 2926 196952 2932
rect 196440 2644 196492 2650
rect 196440 2586 196492 2592
rect 196912 2514 196940 2926
rect 196900 2508 196952 2514
rect 196900 2450 196952 2456
rect 196716 1352 196768 1358
rect 196716 1294 196768 1300
rect 196728 800 196756 1294
rect 197096 800 197124 7890
rect 197280 3534 197308 8978
rect 197360 8832 197412 8838
rect 197360 8774 197412 8780
rect 197372 8090 197400 8774
rect 197556 8498 197584 10200
rect 198016 9926 198044 10200
rect 198004 9920 198056 9926
rect 198004 9862 198056 9868
rect 198476 9110 198504 10200
rect 198844 9994 198872 10200
rect 198832 9988 198884 9994
rect 198832 9930 198884 9936
rect 198464 9104 198516 9110
rect 198464 9046 198516 9052
rect 197544 8492 197596 8498
rect 197544 8434 197596 8440
rect 197360 8084 197412 8090
rect 197360 8026 197412 8032
rect 199304 7750 199332 10200
rect 199764 9654 199792 10200
rect 199752 9648 199804 9654
rect 199752 9590 199804 9596
rect 199292 7744 199344 7750
rect 199292 7686 199344 7692
rect 197268 3528 197320 3534
rect 197268 3470 197320 3476
rect 198004 3528 198056 3534
rect 198004 3470 198056 3476
rect 197268 1828 197320 1834
rect 197268 1770 197320 1776
rect 197280 1714 197308 1770
rect 197280 1686 197400 1714
rect 197372 1170 197400 1686
rect 197372 1142 197584 1170
rect 197556 800 197584 1142
rect 198016 800 198044 3470
rect 199752 2916 199804 2922
rect 199752 2858 199804 2864
rect 199292 2848 199344 2854
rect 199292 2790 199344 2796
rect 198830 1456 198886 1465
rect 198464 1420 198516 1426
rect 198830 1391 198886 1400
rect 198464 1362 198516 1368
rect 198476 800 198504 1362
rect 198844 800 198872 1391
rect 199304 800 199332 2790
rect 199764 800 199792 2858
rect 188068 750 188120 756
rect 188434 -400 188490 800
rect 188802 -400 188858 800
rect 189262 -400 189318 800
rect 189722 -400 189778 800
rect 190182 -400 190238 800
rect 190550 -400 190606 800
rect 191010 -400 191066 800
rect 191470 -400 191526 800
rect 191930 -400 191986 800
rect 192298 -400 192354 800
rect 192758 -400 192814 800
rect 193218 -400 193274 800
rect 193586 -400 193642 800
rect 194046 -400 194102 800
rect 194506 -400 194562 800
rect 194966 -400 195022 800
rect 195334 -400 195390 800
rect 195794 -400 195850 800
rect 196254 -400 196310 800
rect 196714 -400 196770 800
rect 197082 -400 197138 800
rect 197542 -400 197598 800
rect 198002 -400 198058 800
rect 198462 -400 198518 800
rect 198830 -400 198886 800
rect 199290 -400 199346 800
rect 199750 -400 199806 800
<< via2 >>
rect 4076 9818 4132 9820
rect 4076 9766 4078 9818
rect 4078 9766 4130 9818
rect 4130 9766 4132 9818
rect 4076 9764 4132 9766
rect 4066 9152 4122 9208
rect 4076 8730 4132 8732
rect 4076 8678 4078 8730
rect 4078 8678 4130 8730
rect 4130 8678 4132 8730
rect 4076 8676 4132 8678
rect 4076 7642 4132 7644
rect 4076 7590 4078 7642
rect 4078 7590 4130 7642
rect 4130 7590 4132 7642
rect 4076 7588 4132 7590
rect 4076 6554 4132 6556
rect 4076 6502 4078 6554
rect 4078 6502 4130 6554
rect 4130 6502 4132 6554
rect 4076 6500 4132 6502
rect 2962 5480 3018 5536
rect 4076 5466 4132 5468
rect 4076 5414 4078 5466
rect 4078 5414 4130 5466
rect 4130 5414 4132 5466
rect 4076 5412 4132 5414
rect 4076 4378 4132 4380
rect 4076 4326 4078 4378
rect 4078 4326 4130 4378
rect 4130 4326 4132 4378
rect 4076 4324 4132 4326
rect 4076 3290 4132 3292
rect 4076 3238 4078 3290
rect 4078 3238 4130 3290
rect 4130 3238 4132 3290
rect 4076 3236 4132 3238
rect 4076 2202 4132 2204
rect 4076 2150 4078 2202
rect 4078 2150 4130 2202
rect 4130 2150 4132 2202
rect 4076 2148 4132 2150
rect 4066 1808 4122 1864
rect 4076 1114 4132 1116
rect 4076 1062 4078 1114
rect 4078 1062 4130 1114
rect 4130 1062 4132 1114
rect 4076 1060 4132 1062
rect 24076 9274 24132 9276
rect 24076 9222 24078 9274
rect 24078 9222 24130 9274
rect 24130 9222 24132 9274
rect 24076 9220 24132 9222
rect 24076 8186 24132 8188
rect 24076 8134 24078 8186
rect 24078 8134 24130 8186
rect 24130 8134 24132 8186
rect 24076 8132 24132 8134
rect 24076 7098 24132 7100
rect 24076 7046 24078 7098
rect 24078 7046 24130 7098
rect 24130 7046 24132 7098
rect 24076 7044 24132 7046
rect 24076 6010 24132 6012
rect 24076 5958 24078 6010
rect 24078 5958 24130 6010
rect 24130 5958 24132 6010
rect 24076 5956 24132 5958
rect 24076 4922 24132 4924
rect 24076 4870 24078 4922
rect 24078 4870 24130 4922
rect 24130 4870 24132 4922
rect 24076 4868 24132 4870
rect 24076 3834 24132 3836
rect 24076 3782 24078 3834
rect 24078 3782 24130 3834
rect 24130 3782 24132 3834
rect 24076 3780 24132 3782
rect 24076 2746 24132 2748
rect 24076 2694 24078 2746
rect 24078 2694 24130 2746
rect 24130 2694 24132 2746
rect 24076 2692 24132 2694
rect 24076 1658 24132 1660
rect 24076 1606 24078 1658
rect 24078 1606 24130 1658
rect 24130 1606 24132 1658
rect 24076 1604 24132 1606
rect 44076 9818 44132 9820
rect 44076 9766 44078 9818
rect 44078 9766 44130 9818
rect 44130 9766 44132 9818
rect 44076 9764 44132 9766
rect 44076 8730 44132 8732
rect 44076 8678 44078 8730
rect 44078 8678 44130 8730
rect 44130 8678 44132 8730
rect 44076 8676 44132 8678
rect 44076 7642 44132 7644
rect 44076 7590 44078 7642
rect 44078 7590 44130 7642
rect 44130 7590 44132 7642
rect 44076 7588 44132 7590
rect 44076 6554 44132 6556
rect 44076 6502 44078 6554
rect 44078 6502 44130 6554
rect 44130 6502 44132 6554
rect 44076 6500 44132 6502
rect 44076 5466 44132 5468
rect 44076 5414 44078 5466
rect 44078 5414 44130 5466
rect 44130 5414 44132 5466
rect 44076 5412 44132 5414
rect 44076 4378 44132 4380
rect 44076 4326 44078 4378
rect 44078 4326 44130 4378
rect 44130 4326 44132 4378
rect 44076 4324 44132 4326
rect 44076 3290 44132 3292
rect 44076 3238 44078 3290
rect 44078 3238 44130 3290
rect 44130 3238 44132 3290
rect 44076 3236 44132 3238
rect 44076 2202 44132 2204
rect 44076 2150 44078 2202
rect 44078 2150 44130 2202
rect 44130 2150 44132 2202
rect 44076 2148 44132 2150
rect 44076 1114 44132 1116
rect 44076 1062 44078 1114
rect 44078 1062 44130 1114
rect 44130 1062 44132 1114
rect 44076 1060 44132 1062
rect 60646 3984 60702 4040
rect 64076 9274 64132 9276
rect 64076 9222 64078 9274
rect 64078 9222 64130 9274
rect 64130 9222 64132 9274
rect 64076 9220 64132 9222
rect 64076 8186 64132 8188
rect 64076 8134 64078 8186
rect 64078 8134 64130 8186
rect 64130 8134 64132 8186
rect 64076 8132 64132 8134
rect 64076 7098 64132 7100
rect 64076 7046 64078 7098
rect 64078 7046 64130 7098
rect 64130 7046 64132 7098
rect 64076 7044 64132 7046
rect 64076 6010 64132 6012
rect 64076 5958 64078 6010
rect 64078 5958 64130 6010
rect 64130 5958 64132 6010
rect 64076 5956 64132 5958
rect 64076 4922 64132 4924
rect 64076 4870 64078 4922
rect 64078 4870 64130 4922
rect 64130 4870 64132 4922
rect 64076 4868 64132 4870
rect 64076 3834 64132 3836
rect 64076 3782 64078 3834
rect 64078 3782 64130 3834
rect 64130 3782 64132 3834
rect 64076 3780 64132 3782
rect 64076 2746 64132 2748
rect 64076 2694 64078 2746
rect 64078 2694 64130 2746
rect 64130 2694 64132 2746
rect 64076 2692 64132 2694
rect 64076 1658 64132 1660
rect 64076 1606 64078 1658
rect 64078 1606 64130 1658
rect 64130 1606 64132 1658
rect 64076 1604 64132 1606
rect 68742 7248 68798 7304
rect 70306 4564 70308 4584
rect 70308 4564 70360 4584
rect 70360 4564 70362 4584
rect 70306 4528 70362 4564
rect 79046 3576 79102 3632
rect 79138 2352 79194 2408
rect 80978 1400 81034 1456
rect 81254 2896 81310 2952
rect 81806 6180 81862 6216
rect 81806 6160 81808 6180
rect 81808 6160 81860 6180
rect 81860 6160 81862 6180
rect 82174 6180 82230 6216
rect 82174 6160 82176 6180
rect 82176 6160 82228 6180
rect 82228 6160 82230 6180
rect 84076 9818 84132 9820
rect 84076 9766 84078 9818
rect 84078 9766 84130 9818
rect 84130 9766 84132 9818
rect 84076 9764 84132 9766
rect 84076 8730 84132 8732
rect 84076 8678 84078 8730
rect 84078 8678 84130 8730
rect 84130 8678 84132 8730
rect 84076 8676 84132 8678
rect 84076 7642 84132 7644
rect 84076 7590 84078 7642
rect 84078 7590 84130 7642
rect 84130 7590 84132 7642
rect 84076 7588 84132 7590
rect 84076 6554 84132 6556
rect 84076 6502 84078 6554
rect 84078 6502 84130 6554
rect 84130 6502 84132 6554
rect 84076 6500 84132 6502
rect 84076 5466 84132 5468
rect 84076 5414 84078 5466
rect 84078 5414 84130 5466
rect 84130 5414 84132 5466
rect 84076 5412 84132 5414
rect 84076 4378 84132 4380
rect 84076 4326 84078 4378
rect 84078 4326 84130 4378
rect 84130 4326 84132 4378
rect 84076 4324 84132 4326
rect 84076 3290 84132 3292
rect 84076 3238 84078 3290
rect 84078 3238 84130 3290
rect 84130 3238 84132 3290
rect 84076 3236 84132 3238
rect 84076 2202 84132 2204
rect 84076 2150 84078 2202
rect 84078 2150 84130 2202
rect 84130 2150 84132 2202
rect 84076 2148 84132 2150
rect 84076 1114 84132 1116
rect 84076 1062 84078 1114
rect 84078 1062 84130 1114
rect 84130 1062 84132 1114
rect 84076 1060 84132 1062
rect 86774 1808 86830 1864
rect 89626 3304 89682 3360
rect 89994 5244 89996 5264
rect 89996 5244 90048 5264
rect 90048 5244 90050 5264
rect 89994 5208 90050 5244
rect 90270 2488 90326 2544
rect 91926 5480 91982 5536
rect 93306 7384 93362 7440
rect 92018 1944 92074 2000
rect 93766 7520 93822 7576
rect 93674 1264 93730 1320
rect 96158 7384 96214 7440
rect 97078 8880 97134 8936
rect 96894 6024 96950 6080
rect 97630 6296 97686 6352
rect 97538 6160 97594 6216
rect 97630 3440 97686 3496
rect 98274 6704 98330 6760
rect 98458 7420 98460 7440
rect 98460 7420 98512 7440
rect 98512 7420 98514 7440
rect 98458 7384 98514 7420
rect 99194 6840 99250 6896
rect 99286 6332 99288 6352
rect 99288 6332 99340 6352
rect 99340 6332 99342 6352
rect 99286 6296 99342 6332
rect 99286 6160 99342 6216
rect 99470 6196 99472 6216
rect 99472 6196 99524 6216
rect 99524 6196 99526 6216
rect 99470 6160 99526 6196
rect 99470 5908 99526 5944
rect 99746 6860 99802 6896
rect 99746 6840 99748 6860
rect 99748 6840 99800 6860
rect 99800 6840 99802 6860
rect 99746 6704 99802 6760
rect 99470 5888 99472 5908
rect 99472 5888 99524 5908
rect 99524 5888 99526 5908
rect 99286 5752 99342 5808
rect 100114 6024 100170 6080
rect 101218 5364 101274 5400
rect 101218 5344 101220 5364
rect 101220 5344 101272 5364
rect 101272 5344 101274 5364
rect 101126 2080 101182 2136
rect 102690 5888 102746 5944
rect 102966 6160 103022 6216
rect 102874 4664 102930 4720
rect 104076 9274 104132 9276
rect 104076 9222 104078 9274
rect 104078 9222 104130 9274
rect 104130 9222 104132 9274
rect 104076 9220 104132 9222
rect 104076 8186 104132 8188
rect 104076 8134 104078 8186
rect 104078 8134 104130 8186
rect 104130 8134 104132 8186
rect 104076 8132 104132 8134
rect 103886 7812 103942 7848
rect 103886 7792 103888 7812
rect 103888 7792 103940 7812
rect 103940 7792 103942 7812
rect 104076 7098 104132 7100
rect 104076 7046 104078 7098
rect 104078 7046 104130 7098
rect 104130 7046 104132 7098
rect 104076 7044 104132 7046
rect 104076 6010 104132 6012
rect 104076 5958 104078 6010
rect 104078 5958 104130 6010
rect 104130 5958 104132 6010
rect 104076 5956 104132 5958
rect 104622 8880 104678 8936
rect 104346 5772 104402 5808
rect 104346 5752 104348 5772
rect 104348 5752 104400 5772
rect 104400 5752 104402 5772
rect 104076 4922 104132 4924
rect 104076 4870 104078 4922
rect 104078 4870 104130 4922
rect 104130 4870 104132 4922
rect 104076 4868 104132 4870
rect 104076 3834 104132 3836
rect 104076 3782 104078 3834
rect 104078 3782 104130 3834
rect 104130 3782 104132 3834
rect 104076 3780 104132 3782
rect 104076 2746 104132 2748
rect 104076 2694 104078 2746
rect 104078 2694 104130 2746
rect 104130 2694 104132 2746
rect 104076 2692 104132 2694
rect 105266 8064 105322 8120
rect 105358 7656 105414 7712
rect 105174 5344 105230 5400
rect 105082 5108 105084 5128
rect 105084 5108 105136 5128
rect 105136 5108 105138 5128
rect 105082 5072 105138 5108
rect 105358 4256 105414 4312
rect 105450 4120 105506 4176
rect 106370 4972 106372 4992
rect 106372 4972 106424 4992
rect 106424 4972 106426 4992
rect 106370 4936 106426 4972
rect 106278 4800 106334 4856
rect 105910 4256 105966 4312
rect 104622 2624 104678 2680
rect 104076 1658 104132 1660
rect 104076 1606 104078 1658
rect 104078 1606 104130 1658
rect 104130 1606 104132 1658
rect 104076 1604 104132 1606
rect 105450 2080 105506 2136
rect 105818 3440 105874 3496
rect 106646 5344 106702 5400
rect 106646 4936 106702 4992
rect 106646 4800 106702 4856
rect 106554 4392 106610 4448
rect 106646 3440 106702 3496
rect 106646 2216 106702 2272
rect 107014 5072 107070 5128
rect 106922 4936 106978 4992
rect 107566 7948 107622 7984
rect 108302 8336 108358 8392
rect 107566 7928 107568 7948
rect 107568 7928 107620 7948
rect 107620 7928 107622 7948
rect 107474 7112 107530 7168
rect 107566 4800 107622 4856
rect 107658 3848 107714 3904
rect 107014 2760 107070 2816
rect 107290 1672 107346 1728
rect 108118 6840 108174 6896
rect 108118 5108 108120 5128
rect 108120 5108 108172 5128
rect 108172 5108 108174 5128
rect 108118 5072 108174 5108
rect 107934 4664 107990 4720
rect 108762 6432 108818 6488
rect 108394 5616 108450 5672
rect 108394 4936 108450 4992
rect 108394 2100 108450 2136
rect 108394 2080 108396 2100
rect 108396 2080 108448 2100
rect 108448 2080 108450 2100
rect 108762 5772 108818 5808
rect 108762 5752 108764 5772
rect 108764 5752 108816 5772
rect 108816 5752 108818 5772
rect 109130 6432 109186 6488
rect 109222 5888 109278 5944
rect 109590 6976 109646 7032
rect 109590 6024 109646 6080
rect 109682 4120 109738 4176
rect 109590 3984 109646 4040
rect 109590 3712 109646 3768
rect 109222 3168 109278 3224
rect 108762 2216 108818 2272
rect 109038 2216 109094 2272
rect 109038 1556 109094 1592
rect 109038 1536 109040 1556
rect 109040 1536 109092 1556
rect 109092 1536 109094 1556
rect 109222 2080 109278 2136
rect 109498 2080 109554 2136
rect 109682 1672 109738 1728
rect 109774 1556 109830 1592
rect 109774 1536 109776 1556
rect 109776 1536 109828 1556
rect 109828 1536 109830 1556
rect 98366 176 98422 232
rect 110418 4936 110474 4992
rect 110510 4800 110566 4856
rect 110418 4392 110474 4448
rect 110326 3984 110382 4040
rect 110510 2760 110566 2816
rect 110878 4800 110934 4856
rect 111062 4120 111118 4176
rect 111062 3848 111118 3904
rect 111246 6024 111302 6080
rect 111246 4392 111302 4448
rect 110970 2216 111026 2272
rect 110142 1536 110198 1592
rect 110694 1420 110750 1456
rect 110694 1400 110696 1420
rect 110696 1400 110748 1420
rect 110748 1400 110750 1420
rect 111614 4664 111670 4720
rect 111706 3848 111762 3904
rect 111522 2080 111578 2136
rect 112074 3168 112130 3224
rect 112074 1844 112076 1864
rect 112076 1844 112128 1864
rect 112128 1844 112130 1864
rect 112074 1808 112130 1844
rect 111982 1400 112038 1456
rect 113454 8336 113510 8392
rect 113638 4392 113694 4448
rect 113454 3984 113510 4040
rect 114006 7520 114062 7576
rect 113730 3712 113786 3768
rect 112442 3304 112498 3360
rect 112350 2388 112352 2408
rect 112352 2388 112404 2408
rect 112404 2388 112406 2408
rect 112350 2352 112406 2388
rect 112258 1808 112314 1864
rect 113822 3052 113878 3088
rect 113822 3032 113824 3052
rect 113824 3032 113876 3052
rect 113876 3032 113878 3052
rect 113546 2916 113602 2952
rect 113546 2896 113548 2916
rect 113548 2896 113600 2916
rect 113600 2896 113602 2916
rect 113546 1964 113602 2000
rect 114466 8064 114522 8120
rect 114282 7112 114338 7168
rect 114466 6432 114522 6488
rect 114466 6296 114522 6352
rect 114834 6160 114890 6216
rect 114742 5652 114744 5672
rect 114744 5652 114796 5672
rect 114796 5652 114798 5672
rect 114742 5616 114798 5652
rect 115386 3848 115442 3904
rect 114190 3440 114246 3496
rect 115202 2524 115204 2544
rect 115204 2524 115256 2544
rect 115256 2524 115258 2544
rect 115202 2488 115258 2524
rect 113546 1944 113548 1964
rect 113548 1944 113600 1964
rect 113600 1944 113602 1964
rect 115938 3440 115994 3496
rect 115846 3168 115902 3224
rect 116950 5344 117006 5400
rect 116950 4428 116952 4448
rect 116952 4428 117004 4448
rect 117004 4428 117006 4448
rect 116950 4392 117006 4428
rect 116490 3340 116492 3360
rect 116492 3340 116544 3360
rect 116544 3340 116546 3360
rect 116490 3304 116546 3340
rect 116858 3848 116914 3904
rect 116674 2896 116730 2952
rect 116858 2760 116914 2816
rect 116306 2252 116308 2272
rect 116308 2252 116360 2272
rect 116360 2252 116362 2272
rect 116306 2216 116362 2252
rect 110050 720 110106 776
rect 116858 1128 116914 1184
rect 117502 9152 117558 9208
rect 118054 6024 118110 6080
rect 117594 4800 117650 4856
rect 117410 4528 117466 4584
rect 117318 3304 117374 3360
rect 117502 3304 117558 3360
rect 117134 2216 117190 2272
rect 118790 7248 118846 7304
rect 118606 7112 118662 7168
rect 118882 6160 118938 6216
rect 118514 5364 118570 5400
rect 118514 5344 118516 5364
rect 118516 5344 118568 5364
rect 118568 5344 118570 5364
rect 118514 3984 118570 4040
rect 118514 3712 118570 3768
rect 118698 3340 118700 3360
rect 118700 3340 118752 3360
rect 118752 3340 118754 3360
rect 118698 3304 118754 3340
rect 118330 3168 118386 3224
rect 118974 4392 119030 4448
rect 118606 2896 118662 2952
rect 118238 2644 118294 2680
rect 118238 2624 118240 2644
rect 118240 2624 118292 2644
rect 118292 2624 118294 2644
rect 119342 4800 119398 4856
rect 119618 6160 119674 6216
rect 119618 5616 119674 5672
rect 119618 4548 119674 4584
rect 119618 4528 119620 4548
rect 119620 4528 119672 4548
rect 119672 4528 119674 4548
rect 119618 3848 119674 3904
rect 119250 3712 119306 3768
rect 119066 3576 119122 3632
rect 119158 1828 119214 1864
rect 119158 1808 119160 1828
rect 119160 1808 119212 1828
rect 119212 1808 119214 1828
rect 119986 3984 120042 4040
rect 120170 3576 120226 3632
rect 119802 3168 119858 3224
rect 120170 2352 120226 2408
rect 120078 1672 120134 1728
rect 120446 5344 120502 5400
rect 120170 1400 120226 1456
rect 120998 2488 121054 2544
rect 120814 2216 120870 2272
rect 121274 5344 121330 5400
rect 121182 4256 121238 4312
rect 122194 9152 122250 9208
rect 121734 5480 121790 5536
rect 122102 2624 122158 2680
rect 122746 6704 122802 6760
rect 122562 2760 122618 2816
rect 121274 1128 121330 1184
rect 122930 5208 122986 5264
rect 123850 7656 123906 7712
rect 123574 5364 123630 5400
rect 123574 5344 123576 5364
rect 123576 5344 123628 5364
rect 123628 5344 123630 5364
rect 123758 6432 123814 6488
rect 124076 9818 124132 9820
rect 124076 9766 124078 9818
rect 124078 9766 124130 9818
rect 124130 9766 124132 9818
rect 124076 9764 124132 9766
rect 124076 8730 124132 8732
rect 124076 8678 124078 8730
rect 124078 8678 124130 8730
rect 124130 8678 124132 8730
rect 124076 8676 124132 8678
rect 124076 7642 124132 7644
rect 124076 7590 124078 7642
rect 124078 7590 124130 7642
rect 124130 7590 124132 7642
rect 124076 7588 124132 7590
rect 124076 6554 124132 6556
rect 124076 6502 124078 6554
rect 124078 6502 124130 6554
rect 124130 6502 124132 6554
rect 124076 6500 124132 6502
rect 124402 6196 124404 6216
rect 124404 6196 124456 6216
rect 124456 6196 124458 6216
rect 124402 6160 124458 6196
rect 124076 5466 124132 5468
rect 124076 5414 124078 5466
rect 124078 5414 124130 5466
rect 124130 5414 124132 5466
rect 124076 5412 124132 5414
rect 123758 4528 123814 4584
rect 123574 3168 123630 3224
rect 123758 1944 123814 2000
rect 124126 4564 124128 4584
rect 124128 4564 124180 4584
rect 124180 4564 124182 4584
rect 124126 4528 124182 4564
rect 124218 4392 124274 4448
rect 124076 4378 124132 4380
rect 124076 4326 124078 4378
rect 124078 4326 124130 4378
rect 124130 4326 124132 4378
rect 124076 4324 124132 4326
rect 123942 4256 123998 4312
rect 124218 4256 124274 4312
rect 123942 3712 123998 3768
rect 124076 3290 124132 3292
rect 124076 3238 124078 3290
rect 124078 3238 124130 3290
rect 124130 3238 124132 3290
rect 124076 3236 124132 3238
rect 123942 2760 123998 2816
rect 124076 2202 124132 2204
rect 124076 2150 124078 2202
rect 124078 2150 124130 2202
rect 124130 2150 124132 2202
rect 124076 2148 124132 2150
rect 124218 2080 124274 2136
rect 124218 1536 124274 1592
rect 124076 1114 124132 1116
rect 124076 1062 124078 1114
rect 124078 1062 124130 1114
rect 124130 1062 124132 1114
rect 124076 1060 124132 1062
rect 123850 856 123906 912
rect 124770 7112 124826 7168
rect 124678 2352 124734 2408
rect 125782 9016 125838 9072
rect 125874 7656 125930 7712
rect 125966 6704 126022 6760
rect 125690 5208 125746 5264
rect 125506 3576 125562 3632
rect 125138 2896 125194 2952
rect 125230 2488 125286 2544
rect 124862 1420 124918 1456
rect 124862 1400 124864 1420
rect 124864 1400 124916 1420
rect 124916 1400 124918 1420
rect 125046 1536 125102 1592
rect 125414 2624 125470 2680
rect 126794 9152 126850 9208
rect 126610 8200 126666 8256
rect 126886 8336 126942 8392
rect 126794 5208 126850 5264
rect 127254 7248 127310 7304
rect 127622 7248 127678 7304
rect 127254 6432 127310 6488
rect 127530 6704 127586 6760
rect 127714 6704 127770 6760
rect 127714 6160 127770 6216
rect 127346 4800 127402 4856
rect 126242 3984 126298 4040
rect 126058 3848 126114 3904
rect 125966 3712 126022 3768
rect 125966 3596 126022 3632
rect 125966 3576 125968 3596
rect 125968 3576 126020 3596
rect 126020 3576 126022 3596
rect 125322 1944 125378 2000
rect 125690 2508 125746 2544
rect 125690 2488 125692 2508
rect 125692 2488 125744 2508
rect 125744 2488 125746 2508
rect 125782 1944 125838 2000
rect 126794 3848 126850 3904
rect 126886 1844 126888 1864
rect 126888 1844 126940 1864
rect 126940 1844 126942 1864
rect 126886 1808 126942 1844
rect 127530 5480 127586 5536
rect 127438 2080 127494 2136
rect 127346 1808 127402 1864
rect 127622 2080 127678 2136
rect 127990 5616 128046 5672
rect 128174 5616 128230 5672
rect 128174 5344 128230 5400
rect 128266 3476 128268 3496
rect 128268 3476 128320 3496
rect 128320 3476 128322 3496
rect 128266 3440 128322 3476
rect 127162 312 127218 368
rect 128450 7112 128506 7168
rect 128542 4800 128598 4856
rect 128818 8880 128874 8936
rect 128726 3984 128782 4040
rect 128634 3732 128690 3768
rect 128634 3712 128636 3732
rect 128636 3712 128688 3732
rect 128688 3712 128690 3732
rect 128450 3460 128506 3496
rect 128450 3440 128452 3460
rect 128452 3440 128504 3460
rect 128504 3440 128506 3460
rect 128726 3188 128782 3224
rect 128726 3168 128728 3188
rect 128728 3168 128780 3188
rect 128780 3168 128782 3188
rect 128450 2916 128506 2952
rect 128450 2896 128452 2916
rect 128452 2896 128504 2916
rect 128504 2896 128506 2916
rect 128818 2624 128874 2680
rect 129278 8744 129334 8800
rect 129370 7520 129426 7576
rect 128910 992 128966 1048
rect 128358 40 128414 96
rect 129278 3304 129334 3360
rect 129554 9152 129610 9208
rect 129738 5364 129794 5400
rect 129738 5344 129740 5364
rect 129740 5344 129792 5364
rect 129792 5344 129794 5364
rect 129738 3304 129794 3360
rect 130014 5480 130070 5536
rect 129922 3440 129978 3496
rect 130474 7248 130530 7304
rect 130842 9016 130898 9072
rect 131670 8608 131726 8664
rect 131026 6568 131082 6624
rect 131302 5208 131358 5264
rect 131026 3984 131082 4040
rect 130566 584 130622 640
rect 131762 7248 131818 7304
rect 131486 2080 131542 2136
rect 131854 3712 131910 3768
rect 131762 2080 131818 2136
rect 132038 2624 132094 2680
rect 132406 8492 132462 8528
rect 132406 8472 132408 8492
rect 132408 8472 132460 8492
rect 132460 8472 132462 8492
rect 132774 8064 132830 8120
rect 132406 5344 132462 5400
rect 132590 5616 132646 5672
rect 132498 3440 132554 3496
rect 132222 2624 132278 2680
rect 132682 4800 132738 4856
rect 132038 1128 132094 1184
rect 133050 5480 133106 5536
rect 132958 4800 133014 4856
rect 132958 4256 133014 4312
rect 132314 1808 132370 1864
rect 131946 448 132002 504
rect 132866 76 132868 96
rect 132868 76 132920 96
rect 132920 76 132922 96
rect 132866 40 132922 76
rect 133418 8336 133474 8392
rect 134338 8880 134394 8936
rect 134522 8744 134578 8800
rect 133878 8236 133880 8256
rect 133880 8236 133932 8256
rect 133932 8236 133934 8256
rect 133878 8200 133934 8236
rect 134062 8200 134118 8256
rect 134982 8336 135038 8392
rect 134982 8064 135038 8120
rect 134062 7792 134118 7848
rect 133326 6568 133382 6624
rect 133510 6568 133566 6624
rect 133970 7540 134026 7576
rect 133970 7520 133972 7540
rect 133972 7520 134024 7540
rect 134024 7520 134026 7540
rect 134154 7520 134210 7576
rect 133326 4392 133382 4448
rect 133326 3848 133382 3904
rect 133326 3576 133382 3632
rect 133786 6976 133842 7032
rect 133970 7112 134026 7168
rect 134154 7112 134210 7168
rect 133602 3848 133658 3904
rect 133510 3032 133566 3088
rect 133694 3032 133750 3088
rect 134614 7812 134670 7848
rect 134614 7792 134616 7812
rect 134616 7792 134668 7812
rect 134668 7792 134670 7812
rect 134614 6976 134670 7032
rect 134430 6296 134486 6352
rect 134614 5888 134670 5944
rect 133970 5228 134026 5264
rect 133970 5208 133972 5228
rect 133972 5208 134024 5228
rect 134024 5208 134026 5228
rect 133510 2760 133566 2816
rect 135166 8064 135222 8120
rect 134982 6976 135038 7032
rect 134982 6704 135038 6760
rect 134982 6432 135038 6488
rect 134982 5888 135038 5944
rect 134798 3848 134854 3904
rect 134430 1808 134486 1864
rect 135166 5208 135222 5264
rect 135350 4392 135406 4448
rect 135626 8608 135682 8664
rect 135626 6976 135682 7032
rect 135810 5616 135866 5672
rect 135626 2896 135682 2952
rect 136730 7656 136786 7712
rect 137926 10104 137982 10160
rect 138018 8200 138074 8256
rect 137834 7964 137836 7984
rect 137836 7964 137888 7984
rect 137888 7964 137890 7984
rect 137834 7928 137890 7964
rect 138018 7928 138074 7984
rect 137926 7792 137982 7848
rect 138110 7792 138166 7848
rect 137374 7656 137430 7712
rect 136638 4548 136694 4584
rect 136638 4528 136640 4548
rect 136640 4528 136692 4548
rect 136692 4528 136694 4548
rect 135902 2932 135904 2952
rect 135904 2932 135956 2952
rect 135956 2932 135958 2952
rect 135902 2896 135958 2932
rect 136638 3984 136694 4040
rect 137006 7112 137062 7168
rect 136914 5480 136970 5536
rect 136914 4664 136970 4720
rect 136914 3848 136970 3904
rect 137006 3712 137062 3768
rect 137558 7112 137614 7168
rect 137650 5480 137706 5536
rect 137190 4528 137246 4584
rect 137650 4528 137706 4584
rect 137926 5480 137982 5536
rect 138294 5344 138350 5400
rect 138018 4528 138074 4584
rect 136914 3304 136970 3360
rect 137190 3304 137246 3360
rect 137466 3340 137468 3360
rect 137468 3340 137520 3360
rect 137520 3340 137522 3360
rect 137466 3304 137522 3340
rect 137466 3032 137522 3088
rect 137098 1808 137154 1864
rect 137282 1844 137284 1864
rect 137284 1844 137336 1864
rect 137336 1844 137338 1864
rect 137282 1808 137338 1844
rect 138110 3712 138166 3768
rect 138202 2624 138258 2680
rect 137742 2080 137798 2136
rect 137558 1808 137614 1864
rect 137742 1808 137798 1864
rect 138662 6296 138718 6352
rect 138662 5888 138718 5944
rect 138570 5072 138626 5128
rect 138478 3712 138534 3768
rect 138202 1672 138258 1728
rect 137558 992 137614 1048
rect 140226 8900 140282 8936
rect 140226 8880 140228 8900
rect 140228 8880 140280 8900
rect 140280 8880 140282 8900
rect 140226 8608 140282 8664
rect 140686 7792 140742 7848
rect 139490 2080 139546 2136
rect 140318 7520 140374 7576
rect 140502 7520 140558 7576
rect 140226 6568 140282 6624
rect 140410 6568 140466 6624
rect 139766 4528 139822 4584
rect 140042 2624 140098 2680
rect 140042 2080 140098 2136
rect 139306 1808 139362 1864
rect 139490 1808 139546 1864
rect 140686 5072 140742 5128
rect 140410 4936 140466 4992
rect 137650 40 137706 96
rect 140778 4120 140834 4176
rect 142802 8064 142858 8120
rect 142158 7384 142214 7440
rect 142802 7792 142858 7848
rect 143446 7404 143502 7440
rect 143446 7384 143448 7404
rect 143448 7384 143500 7404
rect 143500 7384 143502 7404
rect 142710 7268 142766 7304
rect 142710 7248 142712 7268
rect 142712 7248 142764 7268
rect 142764 7248 142766 7268
rect 140962 4800 141018 4856
rect 142158 6024 142214 6080
rect 141514 4548 141570 4584
rect 141514 4528 141516 4548
rect 141516 4528 141568 4548
rect 141568 4528 141570 4548
rect 141514 4256 141570 4312
rect 141330 4120 141386 4176
rect 141422 2760 141478 2816
rect 142434 4392 142490 4448
rect 142250 3712 142306 3768
rect 142986 3304 143042 3360
rect 142710 3168 142766 3224
rect 141606 2624 141662 2680
rect 141790 3032 141846 3088
rect 144076 9274 144132 9276
rect 144076 9222 144078 9274
rect 144078 9222 144130 9274
rect 144130 9222 144132 9274
rect 144076 9220 144132 9222
rect 144458 8608 144514 8664
rect 144458 8336 144514 8392
rect 144076 8186 144132 8188
rect 144076 8134 144078 8186
rect 144078 8134 144130 8186
rect 144130 8134 144132 8186
rect 144076 8132 144132 8134
rect 144274 7112 144330 7168
rect 144076 7098 144132 7100
rect 144076 7046 144078 7098
rect 144078 7046 144130 7098
rect 144130 7046 144132 7098
rect 144076 7044 144132 7046
rect 143630 6860 143686 6896
rect 143630 6840 143632 6860
rect 143632 6840 143684 6860
rect 143684 6840 143686 6860
rect 144458 6160 144514 6216
rect 144076 6010 144132 6012
rect 144076 5958 144078 6010
rect 144078 5958 144130 6010
rect 144130 5958 144132 6010
rect 144076 5956 144132 5958
rect 144458 5752 144514 5808
rect 144458 5480 144514 5536
rect 144642 5480 144698 5536
rect 144076 4922 144132 4924
rect 144076 4870 144078 4922
rect 144078 4870 144130 4922
rect 144130 4870 144132 4922
rect 144076 4868 144132 4870
rect 144458 5072 144514 5128
rect 143906 3848 143962 3904
rect 144076 3834 144132 3836
rect 144076 3782 144078 3834
rect 144078 3782 144130 3834
rect 144130 3782 144132 3834
rect 144076 3780 144132 3782
rect 144550 3712 144606 3768
rect 144918 6296 144974 6352
rect 144458 3576 144514 3632
rect 142250 1672 142306 1728
rect 141790 992 141846 1048
rect 142434 1264 142490 1320
rect 142434 992 142490 1048
rect 143906 1536 143962 1592
rect 143906 1264 143962 1320
rect 144550 3304 144606 3360
rect 144734 3340 144736 3360
rect 144736 3340 144788 3360
rect 144788 3340 144790 3360
rect 144734 3304 144790 3340
rect 144076 2746 144132 2748
rect 144076 2694 144078 2746
rect 144078 2694 144130 2746
rect 144130 2694 144132 2746
rect 144076 2692 144132 2694
rect 144274 1672 144330 1728
rect 144076 1658 144132 1660
rect 144076 1606 144078 1658
rect 144078 1606 144130 1658
rect 144130 1606 144132 1658
rect 144076 1604 144132 1606
rect 144458 2796 144460 2816
rect 144460 2796 144512 2816
rect 144512 2796 144514 2816
rect 144458 2760 144514 2796
rect 145286 4256 145342 4312
rect 145194 2932 145196 2952
rect 145196 2932 145248 2952
rect 145248 2932 145250 2952
rect 145194 2896 145250 2932
rect 144642 1284 144698 1320
rect 144642 1264 144644 1284
rect 144644 1264 144696 1284
rect 144696 1264 144698 1284
rect 146114 9016 146170 9072
rect 145562 2080 145618 2136
rect 145838 2080 145894 2136
rect 145746 1284 145802 1320
rect 145746 1264 145748 1284
rect 145748 1264 145800 1284
rect 145800 1264 145802 1284
rect 146114 2216 146170 2272
rect 146390 2252 146392 2272
rect 146392 2252 146444 2272
rect 146444 2252 146446 2272
rect 146390 2216 146446 2252
rect 145194 176 145250 232
rect 146758 992 146814 1048
rect 148230 9288 148286 9344
rect 148690 6704 148746 6760
rect 148966 9968 149022 10024
rect 149150 6840 149206 6896
rect 149150 1536 149206 1592
rect 146666 720 146722 776
rect 150530 6568 150586 6624
rect 151726 6568 151782 6624
rect 151634 6432 151690 6488
rect 152370 7928 152426 7984
rect 152370 7656 152426 7712
rect 151818 6024 151874 6080
rect 151266 3848 151322 3904
rect 151174 2352 151230 2408
rect 150530 1400 150586 1456
rect 151174 1536 151230 1592
rect 151634 3440 151690 3496
rect 152370 3440 152426 3496
rect 152002 3032 152058 3088
rect 152186 1944 152242 2000
rect 152554 7656 152610 7712
rect 153106 6840 153162 6896
rect 153106 3576 153162 3632
rect 153290 3576 153346 3632
rect 153290 3168 153346 3224
rect 153842 9424 153898 9480
rect 153566 6296 153622 6352
rect 153566 3440 153622 3496
rect 153566 3168 153622 3224
rect 153566 2488 153622 2544
rect 153934 3712 153990 3768
rect 154486 9152 154542 9208
rect 155590 7112 155646 7168
rect 155774 6976 155830 7032
rect 155774 6704 155830 6760
rect 155682 6160 155738 6216
rect 154854 1536 154910 1592
rect 154302 176 154358 232
rect 155774 1944 155830 2000
rect 156142 5208 156198 5264
rect 156234 4120 156290 4176
rect 155222 176 155278 232
rect 156418 8744 156474 8800
rect 156418 7656 156474 7712
rect 156694 9596 156696 9616
rect 156696 9596 156748 9616
rect 156748 9596 156750 9616
rect 156694 9560 156750 9596
rect 156602 7656 156658 7712
rect 156602 6432 156658 6488
rect 156602 3984 156658 4040
rect 157062 8608 157118 8664
rect 157154 8200 157210 8256
rect 157062 7928 157118 7984
rect 156878 7792 156934 7848
rect 156878 7384 156934 7440
rect 157430 8200 157486 8256
rect 157614 8744 157670 8800
rect 157522 8064 157578 8120
rect 157706 8336 157762 8392
rect 157614 7792 157670 7848
rect 157430 7520 157486 7576
rect 157522 7384 157578 7440
rect 157706 7420 157708 7440
rect 157708 7420 157760 7440
rect 157760 7420 157762 7440
rect 157706 7384 157762 7420
rect 159822 7928 159878 7984
rect 160926 8608 160982 8664
rect 161846 9696 161902 9752
rect 161386 8472 161442 8528
rect 161846 8472 161902 8528
rect 161202 7828 161204 7848
rect 161204 7828 161256 7848
rect 161256 7828 161258 7848
rect 161202 7792 161258 7828
rect 158902 7384 158958 7440
rect 159914 7384 159970 7440
rect 162122 8064 162178 8120
rect 163594 8744 163650 8800
rect 164076 9818 164132 9820
rect 164076 9766 164078 9818
rect 164078 9766 164130 9818
rect 164130 9766 164132 9818
rect 164076 9764 164132 9766
rect 164238 9696 164294 9752
rect 165710 10104 165766 10160
rect 164076 8730 164132 8732
rect 164076 8678 164078 8730
rect 164078 8678 164130 8730
rect 164130 8678 164132 8730
rect 164076 8676 164132 8678
rect 164514 8472 164570 8528
rect 163134 8200 163190 8256
rect 163318 8200 163374 8256
rect 162674 7656 162730 7712
rect 164076 7642 164132 7644
rect 164076 7590 164078 7642
rect 164078 7590 164130 7642
rect 164130 7590 164132 7642
rect 164076 7588 164132 7590
rect 163318 7520 163374 7576
rect 164790 8336 164846 8392
rect 166998 9832 167054 9888
rect 165434 7792 165490 7848
rect 164974 7520 165030 7576
rect 165618 7520 165674 7576
rect 166814 8064 166870 8120
rect 167458 9016 167514 9072
rect 167366 8608 167422 8664
rect 167182 8200 167238 8256
rect 168746 9696 168802 9752
rect 167918 8880 167974 8936
rect 167734 8336 167790 8392
rect 169022 8336 169078 8392
rect 167366 7520 167422 7576
rect 169390 8064 169446 8120
rect 170126 9288 170182 9344
rect 170494 8472 170550 8528
rect 170770 8372 170772 8392
rect 170772 8372 170824 8392
rect 170824 8372 170826 8392
rect 170770 8336 170826 8372
rect 170034 8064 170090 8120
rect 172242 9832 172298 9888
rect 172518 9696 172574 9752
rect 171874 9152 171930 9208
rect 171598 8744 171654 8800
rect 172150 8472 172206 8528
rect 173990 9152 174046 9208
rect 173714 9016 173770 9072
rect 173622 7792 173678 7848
rect 175370 9424 175426 9480
rect 174266 7520 174322 7576
rect 174450 7520 174506 7576
rect 176198 9696 176254 9752
rect 175922 9288 175978 9344
rect 176382 8372 176384 8392
rect 176384 8372 176436 8392
rect 176436 8372 176438 8392
rect 176382 8336 176438 8372
rect 176382 8200 176438 8256
rect 176750 8200 176806 8256
rect 176566 7792 176622 7848
rect 177486 7792 177542 7848
rect 176474 7520 176530 7576
rect 162582 7384 162638 7440
rect 164698 7384 164754 7440
rect 164882 7384 164938 7440
rect 166538 7384 166594 7440
rect 167734 7384 167790 7440
rect 169114 7384 169170 7440
rect 169390 7384 169446 7440
rect 169758 7384 169814 7440
rect 170034 7384 170090 7440
rect 171230 7384 171286 7440
rect 171414 7384 171470 7440
rect 171782 7384 171838 7440
rect 172610 7384 172666 7440
rect 173530 7384 173586 7440
rect 174910 7384 174966 7440
rect 175462 7384 175518 7440
rect 178406 9968 178462 10024
rect 179694 9560 179750 9616
rect 178774 8472 178830 8528
rect 178958 8472 179014 8528
rect 180522 8608 180578 8664
rect 181902 8744 181958 8800
rect 180154 8200 180210 8256
rect 180614 8200 180670 8256
rect 181442 8372 181444 8392
rect 181444 8372 181496 8392
rect 181496 8372 181498 8392
rect 181442 8336 181498 8372
rect 181258 8064 181314 8120
rect 180614 7792 180670 7848
rect 180890 7656 180946 7712
rect 177946 7384 178002 7440
rect 178406 7384 178462 7440
rect 181166 7384 181222 7440
rect 182086 7520 182142 7576
rect 183006 9288 183062 9344
rect 182454 8064 182510 8120
rect 183282 8064 183338 8120
rect 184076 9274 184132 9276
rect 184076 9222 184078 9274
rect 184078 9222 184130 9274
rect 184130 9222 184132 9274
rect 184076 9220 184132 9222
rect 184076 8186 184132 8188
rect 184076 8134 184078 8186
rect 184078 8134 184130 8186
rect 184130 8134 184132 8186
rect 184076 8132 184132 8134
rect 181994 7384 182050 7440
rect 182270 7384 182326 7440
rect 182822 7656 182878 7712
rect 183558 7656 183614 7712
rect 184294 7384 184350 7440
rect 156970 6976 157026 7032
rect 157062 6568 157118 6624
rect 157154 6296 157210 6352
rect 156970 5616 157026 5672
rect 157062 5072 157118 5128
rect 156970 4664 157026 4720
rect 156786 3984 156842 4040
rect 156602 1536 156658 1592
rect 156786 1400 156842 1456
rect 156510 1264 156566 1320
rect 177486 7248 177542 7304
rect 177854 7248 177910 7304
rect 157246 5480 157302 5536
rect 157062 2624 157118 2680
rect 157062 2508 157118 2544
rect 157062 2488 157064 2508
rect 157064 2488 157116 2508
rect 157116 2488 157118 2508
rect 156418 720 156474 776
rect 158534 1944 158590 2000
rect 158718 1964 158774 2000
rect 158718 1944 158720 1964
rect 158720 1944 158772 1964
rect 158772 1944 158774 1964
rect 159454 2216 159510 2272
rect 159730 2216 159786 2272
rect 160834 2100 160890 2136
rect 160834 2080 160836 2100
rect 160836 2080 160888 2100
rect 160888 2080 160890 2100
rect 159638 1536 159694 1592
rect 159270 176 159326 232
rect 160650 196 160706 232
rect 161202 1808 161258 1864
rect 161018 1556 161074 1592
rect 161018 1536 161020 1556
rect 161020 1536 161072 1556
rect 161072 1536 161074 1556
rect 162214 2896 162270 2952
rect 162214 2624 162270 2680
rect 161754 2216 161810 2272
rect 161478 1828 161534 1864
rect 161478 1808 161480 1828
rect 161480 1808 161532 1828
rect 161532 1808 161534 1828
rect 160834 720 160890 776
rect 160650 176 160652 196
rect 160652 176 160704 196
rect 160704 176 160706 196
rect 162490 2760 162546 2816
rect 165342 2896 165398 2952
rect 165526 2896 165582 2952
rect 163778 2760 163834 2816
rect 164330 2760 164386 2816
rect 162950 2352 163006 2408
rect 163134 2352 163190 2408
rect 163686 2352 163742 2408
rect 162122 448 162178 504
rect 162122 40 162178 96
rect 162306 720 162362 776
rect 162490 720 162546 776
rect 162306 176 162362 232
rect 163226 448 163282 504
rect 163686 1828 163742 1864
rect 163686 1808 163688 1828
rect 163688 1808 163740 1828
rect 163740 1808 163742 1828
rect 163318 312 163374 368
rect 164238 2216 164294 2272
rect 164076 2202 164132 2204
rect 164076 2150 164078 2202
rect 164078 2150 164130 2202
rect 164130 2150 164132 2202
rect 164076 2148 164132 2150
rect 163870 2080 163926 2136
rect 164238 2080 164294 2136
rect 163870 1808 163926 1864
rect 164238 1536 164294 1592
rect 163870 1128 163926 1184
rect 164076 1114 164132 1116
rect 164076 1062 164078 1114
rect 164078 1062 164130 1114
rect 164130 1062 164132 1114
rect 164076 1060 164132 1062
rect 163870 992 163926 1048
rect 164514 1536 164570 1592
rect 164698 1400 164754 1456
rect 164238 992 164294 1048
rect 165250 2624 165306 2680
rect 164974 856 165030 912
rect 163686 312 163742 368
rect 165434 2624 165490 2680
rect 165894 2352 165950 2408
rect 165526 1808 165582 1864
rect 165710 1672 165766 1728
rect 165894 1672 165950 1728
rect 165434 856 165490 912
rect 166078 584 166134 640
rect 167274 2896 167330 2952
rect 169482 2896 169538 2952
rect 169758 2896 169814 2952
rect 170034 2896 170090 2952
rect 171690 2896 171746 2952
rect 166722 2760 166778 2816
rect 168562 2760 168618 2816
rect 167274 2624 167330 2680
rect 167734 2624 167790 2680
rect 166998 2216 167054 2272
rect 166906 2080 166962 2136
rect 167366 1400 167422 1456
rect 168654 2216 168710 2272
rect 166906 448 166962 504
rect 168102 992 168158 1048
rect 168286 992 168342 1048
rect 169022 1672 169078 1728
rect 169666 2760 169722 2816
rect 169758 2216 169814 2272
rect 169390 1808 169446 1864
rect 171138 2644 171194 2680
rect 171138 2624 171140 2644
rect 171140 2624 171192 2644
rect 171192 2624 171194 2644
rect 171322 2624 171378 2680
rect 171322 2352 171378 2408
rect 171322 2080 171378 2136
rect 171138 1400 171194 1456
rect 169114 720 169170 776
rect 170954 856 171010 912
rect 173254 2760 173310 2816
rect 171874 1944 171930 2000
rect 173162 1808 173218 1864
rect 170402 312 170458 368
rect 174910 2896 174966 2952
rect 175922 2896 175978 2952
rect 176474 2916 176530 2952
rect 176474 2896 176476 2916
rect 176476 2896 176528 2916
rect 176528 2896 176530 2916
rect 175278 2760 175334 2816
rect 176750 2896 176806 2952
rect 177854 2896 177910 2952
rect 176566 2760 176622 2816
rect 176290 2388 176292 2408
rect 176292 2388 176344 2408
rect 176344 2388 176346 2408
rect 176290 2352 176346 2388
rect 176198 2216 176254 2272
rect 176014 1708 176016 1728
rect 176016 1708 176068 1728
rect 176068 1708 176070 1728
rect 176014 1672 176070 1708
rect 177026 2216 177082 2272
rect 177118 1808 177174 1864
rect 178314 2080 178370 2136
rect 179510 2352 179566 2408
rect 180430 2916 180486 2952
rect 180430 2896 180432 2916
rect 180432 2896 180484 2916
rect 180484 2896 180486 2916
rect 184076 2746 184132 2748
rect 184076 2694 184078 2746
rect 184078 2694 184130 2746
rect 184130 2694 184132 2746
rect 184076 2692 184132 2694
rect 182546 2372 182602 2408
rect 182546 2352 182548 2372
rect 182548 2352 182600 2372
rect 182600 2352 182602 2372
rect 181994 2100 182050 2136
rect 181994 2080 181996 2100
rect 181996 2080 182048 2100
rect 182048 2080 182050 2100
rect 183374 1808 183430 1864
rect 181350 1672 181406 1728
rect 181534 992 181590 1048
rect 184076 1658 184132 1660
rect 184076 1606 184078 1658
rect 184078 1606 184130 1658
rect 184130 1606 184132 1658
rect 184076 1604 184132 1606
rect 183558 1556 183614 1592
rect 183558 1536 183560 1556
rect 183560 1536 183612 1556
rect 183612 1536 183614 1556
rect 186134 8472 186190 8528
rect 185306 8200 185362 8256
rect 185030 7792 185086 7848
rect 185398 7520 185454 7576
rect 184938 2216 184994 2272
rect 186042 2488 186098 2544
rect 185674 2352 185730 2408
rect 186134 2080 186190 2136
rect 186042 1808 186098 1864
rect 186318 2216 186374 2272
rect 186410 2100 186466 2136
rect 186410 2080 186412 2100
rect 186412 2080 186464 2100
rect 186464 2080 186466 2100
rect 187514 2352 187570 2408
rect 187330 2080 187386 2136
rect 189446 1808 189502 1864
rect 189814 2216 189870 2272
rect 191654 7948 191710 7984
rect 191654 7928 191656 7948
rect 191656 7928 191708 7948
rect 191708 7928 191710 7948
rect 192666 7112 192722 7168
rect 192666 2080 192722 2136
rect 193310 1944 193366 2000
rect 194874 7248 194930 7304
rect 198830 1400 198886 1456
<< metal3 >>
rect -1594 12420 -1588 12484
rect -1524 12482 -1518 12484
rect 25666 12482 25672 12484
rect -1524 12422 25672 12482
rect -1524 12420 -1518 12422
rect 25666 12420 25672 12422
rect 25736 12482 25742 12484
rect 65666 12482 65672 12484
rect 25736 12422 65672 12482
rect 25736 12420 25742 12422
rect 65666 12420 65672 12422
rect 65736 12482 65742 12484
rect 105666 12482 105672 12484
rect 65736 12422 105672 12482
rect 65736 12420 65742 12422
rect 105666 12420 105672 12422
rect 105736 12482 105742 12484
rect 145666 12482 145672 12484
rect 105736 12422 145672 12482
rect 105736 12420 105742 12422
rect 145666 12420 145672 12422
rect 145736 12482 145742 12484
rect 185666 12482 185672 12484
rect 145736 12422 185672 12482
rect 145736 12420 145742 12422
rect 185666 12420 185672 12422
rect 185736 12482 185742 12484
rect 201434 12482 201440 12484
rect 185736 12422 201440 12482
rect 185736 12420 185742 12422
rect 201434 12420 201440 12422
rect 201504 12420 201510 12484
rect -1454 12280 -1448 12344
rect -1384 12342 -1378 12344
rect 5666 12342 5672 12344
rect -1384 12282 5672 12342
rect -1384 12280 -1378 12282
rect 5666 12280 5672 12282
rect 5736 12342 5742 12344
rect 45666 12342 45672 12344
rect 5736 12282 45672 12342
rect 5736 12280 5742 12282
rect 45666 12280 45672 12282
rect 45736 12342 45742 12344
rect 85666 12342 85672 12344
rect 45736 12282 85672 12342
rect 45736 12280 45742 12282
rect 85666 12280 85672 12282
rect 85736 12342 85742 12344
rect 125666 12342 125672 12344
rect 85736 12282 125672 12342
rect 85736 12280 85742 12282
rect 125666 12280 125672 12282
rect 125736 12342 125742 12344
rect 165666 12342 165672 12344
rect 125736 12282 165672 12342
rect 125736 12280 125742 12282
rect 165666 12280 165672 12282
rect 165736 12342 165742 12344
rect 201294 12342 201300 12344
rect 165736 12282 201300 12342
rect 165736 12280 165742 12282
rect 201294 12280 201300 12282
rect 201364 12280 201370 12344
rect -1314 12140 -1308 12204
rect -1244 12202 -1238 12204
rect 25266 12202 25272 12204
rect -1244 12142 25272 12202
rect -1244 12140 -1238 12142
rect 25266 12140 25272 12142
rect 25336 12202 25342 12204
rect 65266 12202 65272 12204
rect 25336 12142 65272 12202
rect 25336 12140 25342 12142
rect 65266 12140 65272 12142
rect 65336 12202 65342 12204
rect 105266 12202 105272 12204
rect 65336 12142 105272 12202
rect 65336 12140 65342 12142
rect 105266 12140 105272 12142
rect 105336 12202 105342 12204
rect 145266 12202 145272 12204
rect 105336 12142 145272 12202
rect 105336 12140 105342 12142
rect 145266 12140 145272 12142
rect 145336 12202 145342 12204
rect 185266 12202 185272 12204
rect 145336 12142 185272 12202
rect 145336 12140 145342 12142
rect 185266 12140 185272 12142
rect 185336 12202 185342 12204
rect 201154 12202 201160 12204
rect 185336 12142 201160 12202
rect 185336 12140 185342 12142
rect 201154 12140 201160 12142
rect 201224 12140 201230 12204
rect -1174 12000 -1168 12064
rect -1104 12062 -1098 12064
rect 5266 12062 5272 12064
rect -1104 12002 5272 12062
rect -1104 12000 -1098 12002
rect 5266 12000 5272 12002
rect 5336 12062 5342 12064
rect 45266 12062 45272 12064
rect 5336 12002 45272 12062
rect 5336 12000 5342 12002
rect 45266 12000 45272 12002
rect 45336 12062 45342 12064
rect 85266 12062 85272 12064
rect 45336 12002 85272 12062
rect 45336 12000 45342 12002
rect 85266 12000 85272 12002
rect 85336 12062 85342 12064
rect 125266 12062 125272 12064
rect 85336 12002 125272 12062
rect 85336 12000 85342 12002
rect 125266 12000 125272 12002
rect 125336 12062 125342 12064
rect 165266 12062 165272 12064
rect 125336 12002 165272 12062
rect 125336 12000 125342 12002
rect 165266 12000 165272 12002
rect 165336 12062 165342 12064
rect 201014 12062 201020 12064
rect 165336 12002 201020 12062
rect 165336 12000 165342 12002
rect 201014 12000 201020 12002
rect 201084 12000 201090 12064
rect -1034 11860 -1028 11924
rect -964 11922 -958 11924
rect 24866 11922 24872 11924
rect -964 11862 24872 11922
rect -964 11860 -958 11862
rect 24866 11860 24872 11862
rect 24936 11922 24942 11924
rect 64866 11922 64872 11924
rect 24936 11862 64872 11922
rect 24936 11860 24942 11862
rect 64866 11860 64872 11862
rect 64936 11922 64942 11924
rect 104866 11922 104872 11924
rect 64936 11862 104872 11922
rect 64936 11860 64942 11862
rect 104866 11860 104872 11862
rect 104936 11922 104942 11924
rect 144866 11922 144872 11924
rect 104936 11862 144872 11922
rect 104936 11860 104942 11862
rect 144866 11860 144872 11862
rect 144936 11922 144942 11924
rect 184866 11922 184872 11924
rect 144936 11862 184872 11922
rect 144936 11860 144942 11862
rect 184866 11860 184872 11862
rect 184936 11922 184942 11924
rect 200874 11922 200880 11924
rect 184936 11862 200880 11922
rect 184936 11860 184942 11862
rect 200874 11860 200880 11862
rect 200944 11860 200950 11924
rect -894 11720 -888 11784
rect -824 11782 -818 11784
rect 4866 11782 4872 11784
rect -824 11722 4872 11782
rect -824 11720 -818 11722
rect 4866 11720 4872 11722
rect 4936 11782 4942 11784
rect 44866 11782 44872 11784
rect 4936 11722 44872 11782
rect 4936 11720 4942 11722
rect 44866 11720 44872 11722
rect 44936 11782 44942 11784
rect 84866 11782 84872 11784
rect 44936 11722 84872 11782
rect 44936 11720 44942 11722
rect 84866 11720 84872 11722
rect 84936 11782 84942 11784
rect 124866 11782 124872 11784
rect 84936 11722 124872 11782
rect 84936 11720 84942 11722
rect 124866 11720 124872 11722
rect 124936 11782 124942 11784
rect 164866 11782 164872 11784
rect 124936 11722 164872 11782
rect 124936 11720 124942 11722
rect 164866 11720 164872 11722
rect 164936 11782 164942 11784
rect 200734 11782 200740 11784
rect 164936 11722 200740 11782
rect 164936 11720 164942 11722
rect 200734 11720 200740 11722
rect 200804 11720 200810 11784
rect -754 11580 -748 11644
rect -684 11642 -678 11644
rect 24466 11642 24472 11644
rect -684 11582 24472 11642
rect -684 11580 -678 11582
rect 24466 11580 24472 11582
rect 24536 11642 24542 11644
rect 64466 11642 64472 11644
rect 24536 11582 64472 11642
rect 24536 11580 24542 11582
rect 64466 11580 64472 11582
rect 64536 11642 64542 11644
rect 104466 11642 104472 11644
rect 64536 11582 104472 11642
rect 64536 11580 64542 11582
rect 104466 11580 104472 11582
rect 104536 11642 104542 11644
rect 144466 11642 144472 11644
rect 104536 11582 144472 11642
rect 104536 11580 104542 11582
rect 144466 11580 144472 11582
rect 144536 11642 144542 11644
rect 184466 11642 184472 11644
rect 144536 11582 184472 11642
rect 144536 11580 144542 11582
rect 184466 11580 184472 11582
rect 184536 11642 184542 11644
rect 200594 11642 200600 11644
rect 184536 11582 200600 11642
rect 184536 11580 184542 11582
rect 200594 11580 200600 11582
rect 200664 11580 200670 11644
rect -614 11440 -608 11504
rect -544 11502 -538 11504
rect 4466 11502 4472 11504
rect -544 11442 4472 11502
rect -544 11440 -538 11442
rect 4466 11440 4472 11442
rect 4536 11502 4542 11504
rect 44466 11502 44472 11504
rect 4536 11442 44472 11502
rect 4536 11440 4542 11442
rect 44466 11440 44472 11442
rect 44536 11502 44542 11504
rect 84466 11502 84472 11504
rect 44536 11442 84472 11502
rect 44536 11440 44542 11442
rect 84466 11440 84472 11442
rect 84536 11502 84542 11504
rect 124466 11502 124472 11504
rect 84536 11442 124472 11502
rect 84536 11440 84542 11442
rect 124466 11440 124472 11442
rect 124536 11502 124542 11504
rect 164466 11502 164472 11504
rect 124536 11442 164472 11502
rect 124536 11440 124542 11442
rect 164466 11440 164472 11442
rect 164536 11502 164542 11504
rect 200454 11502 200460 11504
rect 164536 11442 200460 11502
rect 164536 11440 164542 11442
rect 200454 11440 200460 11442
rect 200524 11440 200530 11504
rect -474 11300 -468 11364
rect -404 11362 -398 11364
rect 24066 11362 24072 11364
rect -404 11302 24072 11362
rect -404 11300 -398 11302
rect 24066 11300 24072 11302
rect 24136 11362 24142 11364
rect 64066 11362 64072 11364
rect 24136 11302 64072 11362
rect 24136 11300 24142 11302
rect 64066 11300 64072 11302
rect 64136 11362 64142 11364
rect 104066 11362 104072 11364
rect 64136 11302 104072 11362
rect 64136 11300 64142 11302
rect 104066 11300 104072 11302
rect 104136 11362 104142 11364
rect 144066 11362 144072 11364
rect 104136 11302 144072 11362
rect 104136 11300 104142 11302
rect 144066 11300 144072 11302
rect 144136 11362 144142 11364
rect 184066 11362 184072 11364
rect 144136 11302 184072 11362
rect 144136 11300 144142 11302
rect 184066 11300 184072 11302
rect 184136 11362 184142 11364
rect 200314 11362 200320 11364
rect 184136 11302 200320 11362
rect 184136 11300 184142 11302
rect 200314 11300 200320 11302
rect 200384 11300 200390 11364
rect -334 11160 -328 11224
rect -264 11222 -258 11224
rect 4066 11222 4072 11224
rect -264 11162 4072 11222
rect -264 11160 -258 11162
rect 4066 11160 4072 11162
rect 4136 11222 4142 11224
rect 44066 11222 44072 11224
rect 4136 11162 44072 11222
rect 4136 11160 4142 11162
rect 44066 11160 44072 11162
rect 44136 11222 44142 11224
rect 84066 11222 84072 11224
rect 44136 11162 84072 11222
rect 44136 11160 44142 11162
rect 84066 11160 84072 11162
rect 84136 11222 84142 11224
rect 124066 11222 124072 11224
rect 84136 11162 124072 11222
rect 84136 11160 84142 11162
rect 124066 11160 124072 11162
rect 124136 11222 124142 11224
rect 164066 11222 164072 11224
rect 124136 11162 164072 11222
rect 124136 11160 124142 11162
rect 164066 11160 164072 11162
rect 164136 11222 164142 11224
rect 200174 11222 200180 11224
rect 164136 11162 200180 11222
rect 164136 11160 164142 11162
rect 200174 11160 200180 11162
rect 200244 11160 200250 11224
rect 137921 10162 137987 10165
rect 165705 10162 165771 10165
rect 137921 10160 165771 10162
rect 137921 10104 137926 10160
rect 137982 10104 165710 10160
rect 165766 10104 165771 10160
rect 137921 10102 165771 10104
rect 137921 10099 137987 10102
rect 165705 10099 165771 10102
rect 148961 10026 149027 10029
rect 178401 10026 178467 10029
rect 148961 10024 178467 10026
rect 148961 9968 148966 10024
rect 149022 9968 178406 10024
rect 178462 9968 178467 10024
rect 148961 9966 178467 9968
rect 148961 9963 149027 9966
rect 178401 9963 178467 9966
rect 166993 9890 167059 9893
rect 172237 9890 172303 9893
rect 166993 9888 172303 9890
rect 166993 9832 166998 9888
rect 167054 9832 172242 9888
rect 172298 9832 172303 9888
rect 166993 9830 172303 9832
rect 166993 9827 167059 9830
rect 172237 9827 172303 9830
rect 4071 9824 4137 9825
rect 44071 9824 44137 9825
rect 84071 9824 84137 9825
rect 124071 9824 124137 9825
rect 164071 9824 164137 9825
rect 4066 9760 4072 9824
rect 4136 9760 4142 9824
rect 44066 9760 44072 9824
rect 44136 9760 44142 9824
rect 84066 9760 84072 9824
rect 84136 9760 84142 9824
rect 124066 9760 124072 9824
rect 124136 9760 124142 9824
rect 164066 9760 164072 9824
rect 164136 9760 164142 9824
rect 4071 9759 4137 9760
rect 44071 9759 44137 9760
rect 84071 9759 84137 9760
rect 124071 9759 124137 9760
rect 164071 9759 164137 9760
rect 157374 9692 157380 9756
rect 157444 9754 157450 9756
rect 161841 9754 161907 9757
rect 157444 9752 161907 9754
rect 157444 9696 161846 9752
rect 161902 9696 161907 9752
rect 157444 9694 161907 9696
rect 157444 9692 157450 9694
rect 161841 9691 161907 9694
rect 164233 9754 164299 9757
rect 168741 9754 168807 9757
rect 164233 9752 168807 9754
rect 164233 9696 164238 9752
rect 164294 9696 168746 9752
rect 168802 9696 168807 9752
rect 164233 9694 168807 9696
rect 164233 9691 164299 9694
rect 168741 9691 168807 9694
rect 172513 9754 172579 9757
rect 176193 9754 176259 9757
rect 172513 9752 176259 9754
rect 172513 9696 172518 9752
rect 172574 9696 176198 9752
rect 176254 9696 176259 9752
rect 172513 9694 176259 9696
rect 172513 9691 172579 9694
rect 176193 9691 176259 9694
rect 156689 9618 156755 9621
rect 179689 9618 179755 9621
rect 156689 9616 179755 9618
rect 156689 9560 156694 9616
rect 156750 9560 179694 9616
rect 179750 9560 179755 9616
rect 156689 9558 179755 9560
rect 156689 9555 156755 9558
rect 179689 9555 179755 9558
rect 153837 9482 153903 9485
rect 175365 9482 175431 9485
rect 153837 9480 175431 9482
rect 153837 9424 153842 9480
rect 153898 9424 175370 9480
rect 175426 9424 175431 9480
rect 153837 9422 175431 9424
rect 153837 9419 153903 9422
rect 175365 9419 175431 9422
rect 148225 9346 148291 9349
rect 170121 9346 170187 9349
rect 148225 9344 170187 9346
rect 148225 9288 148230 9344
rect 148286 9288 170126 9344
rect 170182 9288 170187 9344
rect 148225 9286 170187 9288
rect 148225 9283 148291 9286
rect 170121 9283 170187 9286
rect 175917 9346 175983 9349
rect 183001 9346 183067 9349
rect 175917 9344 183067 9346
rect 175917 9288 175922 9344
rect 175978 9288 183006 9344
rect 183062 9288 183067 9344
rect 175917 9286 183067 9288
rect 175917 9283 175983 9286
rect 183001 9283 183067 9286
rect 24071 9280 24137 9281
rect 64071 9280 64137 9281
rect 104071 9280 104137 9281
rect 144071 9280 144137 9281
rect 184071 9280 184137 9281
rect -400 9210 800 9240
rect 24066 9216 24072 9280
rect 24136 9216 24142 9280
rect 64066 9216 64072 9280
rect 64136 9216 64142 9280
rect 104066 9216 104072 9280
rect 104136 9216 104142 9280
rect 144066 9216 144072 9280
rect 144136 9216 144142 9280
rect 184066 9216 184072 9280
rect 184136 9216 184142 9280
rect 24071 9215 24137 9216
rect 64071 9215 64137 9216
rect 104071 9215 104137 9216
rect 144071 9215 144137 9216
rect 184071 9215 184137 9216
rect 4061 9210 4127 9213
rect -400 9208 4127 9210
rect -400 9152 4066 9208
rect 4122 9152 4127 9208
rect -400 9150 4127 9152
rect -400 9120 800 9150
rect 4061 9147 4127 9150
rect 117497 9210 117563 9213
rect 122189 9210 122255 9213
rect 117497 9208 122255 9210
rect 117497 9152 117502 9208
rect 117558 9152 122194 9208
rect 122250 9152 122255 9208
rect 117497 9150 122255 9152
rect 117497 9147 117563 9150
rect 122189 9147 122255 9150
rect 126789 9210 126855 9213
rect 129549 9210 129615 9213
rect 126789 9208 129615 9210
rect 126789 9152 126794 9208
rect 126850 9152 129554 9208
rect 129610 9152 129615 9208
rect 126789 9150 129615 9152
rect 126789 9147 126855 9150
rect 129549 9147 129615 9150
rect 154481 9210 154547 9213
rect 171869 9210 171935 9213
rect 173985 9210 174051 9213
rect 154481 9208 171935 9210
rect 154481 9152 154486 9208
rect 154542 9152 171874 9208
rect 171930 9152 171935 9208
rect 154481 9150 171935 9152
rect 154481 9147 154547 9150
rect 171869 9147 171935 9150
rect 172470 9208 174051 9210
rect 172470 9152 173990 9208
rect 174046 9152 174051 9208
rect 172470 9150 174051 9152
rect 125777 9074 125843 9077
rect 130837 9074 130903 9077
rect 125777 9072 130903 9074
rect 125777 9016 125782 9072
rect 125838 9016 130842 9072
rect 130898 9016 130903 9072
rect 125777 9014 130903 9016
rect 125777 9011 125843 9014
rect 130837 9011 130903 9014
rect 146109 9074 146175 9077
rect 167453 9074 167519 9077
rect 146109 9072 167519 9074
rect 146109 9016 146114 9072
rect 146170 9016 167458 9072
rect 167514 9016 167519 9072
rect 146109 9014 167519 9016
rect 146109 9011 146175 9014
rect 167453 9011 167519 9014
rect 167862 9012 167868 9076
rect 167932 9074 167938 9076
rect 172470 9074 172530 9150
rect 173985 9147 174051 9150
rect 167932 9014 172530 9074
rect 173709 9076 173775 9077
rect 173709 9072 173756 9076
rect 173820 9074 173826 9076
rect 173709 9016 173714 9072
rect 167932 9012 167938 9014
rect 173709 9012 173756 9016
rect 173820 9014 173866 9074
rect 173820 9012 173826 9014
rect 173709 9011 173775 9012
rect 97073 8938 97139 8941
rect 104617 8938 104683 8941
rect 97073 8936 104683 8938
rect 97073 8880 97078 8936
rect 97134 8880 104622 8936
rect 104678 8880 104683 8936
rect 97073 8878 104683 8880
rect 97073 8875 97139 8878
rect 104617 8875 104683 8878
rect 128813 8938 128879 8941
rect 134333 8938 134399 8941
rect 128813 8936 134399 8938
rect 128813 8880 128818 8936
rect 128874 8880 134338 8936
rect 134394 8880 134399 8936
rect 128813 8878 134399 8880
rect 128813 8875 128879 8878
rect 134333 8875 134399 8878
rect 140221 8938 140287 8941
rect 167913 8938 167979 8941
rect 140221 8936 167979 8938
rect 140221 8880 140226 8936
rect 140282 8880 167918 8936
rect 167974 8880 167979 8936
rect 140221 8878 167979 8880
rect 140221 8875 140287 8878
rect 167913 8875 167979 8878
rect 168966 8876 168972 8940
rect 169036 8938 169042 8940
rect 169036 8878 171794 8938
rect 169036 8876 169042 8878
rect 129273 8802 129339 8805
rect 134517 8802 134583 8805
rect 129273 8800 134583 8802
rect 129273 8744 129278 8800
rect 129334 8744 134522 8800
rect 134578 8744 134583 8800
rect 129273 8742 134583 8744
rect 129273 8739 129339 8742
rect 134517 8739 134583 8742
rect 156413 8802 156479 8805
rect 157609 8802 157675 8805
rect 156413 8800 157675 8802
rect 156413 8744 156418 8800
rect 156474 8744 157614 8800
rect 157670 8744 157675 8800
rect 156413 8742 157675 8744
rect 156413 8739 156479 8742
rect 157609 8739 157675 8742
rect 157742 8740 157748 8804
rect 157812 8802 157818 8804
rect 163589 8802 163655 8805
rect 171593 8802 171659 8805
rect 157812 8800 163655 8802
rect 157812 8744 163594 8800
rect 163650 8744 163655 8800
rect 157812 8742 163655 8744
rect 157812 8740 157818 8742
rect 163589 8739 163655 8742
rect 164374 8800 171659 8802
rect 164374 8744 171598 8800
rect 171654 8744 171659 8800
rect 164374 8742 171659 8744
rect 171734 8802 171794 8878
rect 181897 8802 181963 8805
rect 171734 8800 181963 8802
rect 171734 8744 181902 8800
rect 181958 8744 181963 8800
rect 171734 8742 181963 8744
rect 4071 8736 4137 8737
rect 44071 8736 44137 8737
rect 84071 8736 84137 8737
rect 124071 8736 124137 8737
rect 164071 8736 164137 8737
rect 4066 8672 4072 8736
rect 4136 8672 4142 8736
rect 44066 8672 44072 8736
rect 44136 8672 44142 8736
rect 84066 8672 84072 8736
rect 84136 8672 84142 8736
rect 124066 8672 124072 8736
rect 124136 8672 124142 8736
rect 164066 8672 164072 8736
rect 164136 8672 164142 8736
rect 4071 8671 4137 8672
rect 44071 8671 44137 8672
rect 84071 8671 84137 8672
rect 124071 8671 124137 8672
rect 164071 8671 164137 8672
rect 131665 8666 131731 8669
rect 135621 8666 135687 8669
rect 131665 8664 135687 8666
rect 131665 8608 131670 8664
rect 131726 8608 135626 8664
rect 135682 8608 135687 8664
rect 131665 8606 135687 8608
rect 131665 8603 131731 8606
rect 135621 8603 135687 8606
rect 140221 8666 140287 8669
rect 144453 8666 144519 8669
rect 140221 8664 144519 8666
rect 140221 8608 140226 8664
rect 140282 8608 144458 8664
rect 144514 8608 144519 8664
rect 140221 8606 144519 8608
rect 140221 8603 140287 8606
rect 144453 8603 144519 8606
rect 157057 8666 157123 8669
rect 160921 8666 160987 8669
rect 157057 8664 160987 8666
rect 157057 8608 157062 8664
rect 157118 8608 160926 8664
rect 160982 8608 160987 8664
rect 157057 8606 160987 8608
rect 157057 8603 157123 8606
rect 160921 8603 160987 8606
rect 132401 8530 132467 8533
rect 161381 8530 161447 8533
rect 132401 8528 161447 8530
rect 132401 8472 132406 8528
rect 132462 8472 161386 8528
rect 161442 8472 161447 8528
rect 132401 8470 161447 8472
rect 132401 8467 132467 8470
rect 161381 8467 161447 8470
rect 161841 8530 161907 8533
rect 164374 8530 164434 8742
rect 171593 8739 171659 8742
rect 181897 8739 181963 8742
rect 167361 8666 167427 8669
rect 180517 8666 180583 8669
rect 167361 8664 180583 8666
rect 167361 8608 167366 8664
rect 167422 8608 180522 8664
rect 180578 8608 180583 8664
rect 167361 8606 180583 8608
rect 167361 8603 167427 8606
rect 180517 8603 180583 8606
rect 161841 8528 164434 8530
rect 161841 8472 161846 8528
rect 161902 8472 164434 8528
rect 161841 8470 164434 8472
rect 164509 8530 164575 8533
rect 170489 8530 170555 8533
rect 164509 8528 170555 8530
rect 164509 8472 164514 8528
rect 164570 8472 170494 8528
rect 170550 8472 170555 8528
rect 164509 8470 170555 8472
rect 161841 8467 161907 8470
rect 164509 8467 164575 8470
rect 170489 8467 170555 8470
rect 172145 8530 172211 8533
rect 178769 8530 178835 8533
rect 172145 8528 178835 8530
rect 172145 8472 172150 8528
rect 172206 8472 178774 8528
rect 178830 8472 178835 8528
rect 172145 8470 178835 8472
rect 172145 8467 172211 8470
rect 178769 8467 178835 8470
rect 178953 8530 179019 8533
rect 186129 8530 186195 8533
rect 178953 8528 186195 8530
rect 178953 8472 178958 8528
rect 179014 8472 186134 8528
rect 186190 8472 186195 8528
rect 178953 8470 186195 8472
rect 178953 8467 179019 8470
rect 186129 8467 186195 8470
rect 108297 8394 108363 8397
rect 113449 8394 113515 8397
rect 108297 8392 113515 8394
rect 108297 8336 108302 8392
rect 108358 8336 113454 8392
rect 113510 8336 113515 8392
rect 108297 8334 113515 8336
rect 108297 8331 108363 8334
rect 113449 8331 113515 8334
rect 126881 8394 126947 8397
rect 133413 8394 133479 8397
rect 126881 8392 133479 8394
rect 126881 8336 126886 8392
rect 126942 8336 133418 8392
rect 133474 8336 133479 8392
rect 126881 8334 133479 8336
rect 126881 8331 126947 8334
rect 133413 8331 133479 8334
rect 134977 8394 135043 8397
rect 144453 8394 144519 8397
rect 157558 8394 157564 8396
rect 134977 8392 138260 8394
rect 134977 8336 134982 8392
rect 135038 8336 138260 8392
rect 134977 8334 138260 8336
rect 134977 8331 135043 8334
rect 126605 8258 126671 8261
rect 133873 8258 133939 8261
rect 126605 8256 133939 8258
rect 126605 8200 126610 8256
rect 126666 8200 133878 8256
rect 133934 8200 133939 8256
rect 126605 8198 133939 8200
rect 126605 8195 126671 8198
rect 133873 8195 133939 8198
rect 134057 8258 134123 8261
rect 138013 8258 138079 8261
rect 134057 8256 138079 8258
rect 134057 8200 134062 8256
rect 134118 8200 138018 8256
rect 138074 8200 138079 8256
rect 134057 8198 138079 8200
rect 138200 8258 138260 8334
rect 143904 8334 144378 8394
rect 143904 8258 143964 8334
rect 138200 8198 143964 8258
rect 144318 8258 144378 8334
rect 144453 8392 157564 8394
rect 144453 8336 144458 8392
rect 144514 8336 157564 8392
rect 144453 8334 157564 8336
rect 144453 8331 144519 8334
rect 157558 8332 157564 8334
rect 157628 8332 157634 8396
rect 157701 8394 157767 8397
rect 164785 8394 164851 8397
rect 157701 8392 164851 8394
rect 157701 8336 157706 8392
rect 157762 8336 164790 8392
rect 164846 8336 164851 8392
rect 157701 8334 164851 8336
rect 157701 8331 157767 8334
rect 164785 8331 164851 8334
rect 165470 8332 165476 8396
rect 165540 8394 165546 8396
rect 167729 8394 167795 8397
rect 165540 8392 167795 8394
rect 165540 8336 167734 8392
rect 167790 8336 167795 8392
rect 165540 8334 167795 8336
rect 165540 8332 165546 8334
rect 167729 8331 167795 8334
rect 169017 8394 169083 8397
rect 170765 8396 170831 8397
rect 169518 8394 169524 8396
rect 169017 8392 169524 8394
rect 169017 8336 169022 8392
rect 169078 8336 169524 8392
rect 169017 8334 169524 8336
rect 169017 8331 169083 8334
rect 169518 8332 169524 8334
rect 169588 8332 169594 8396
rect 170765 8392 170812 8396
rect 170876 8394 170882 8396
rect 170765 8336 170770 8392
rect 170765 8332 170812 8336
rect 170876 8334 170922 8394
rect 170876 8332 170882 8334
rect 175958 8332 175964 8396
rect 176028 8394 176034 8396
rect 176377 8394 176443 8397
rect 176028 8392 176443 8394
rect 176028 8336 176382 8392
rect 176438 8336 176443 8392
rect 176028 8334 176443 8336
rect 176028 8332 176034 8334
rect 170765 8331 170831 8332
rect 176377 8331 176443 8334
rect 177614 8332 177620 8396
rect 177684 8394 177690 8396
rect 181437 8394 181503 8397
rect 177684 8392 181503 8394
rect 177684 8336 181442 8392
rect 181498 8336 181503 8392
rect 177684 8334 181503 8336
rect 177684 8332 177690 8334
rect 181437 8331 181503 8334
rect 183878 8334 184306 8394
rect 157149 8258 157215 8261
rect 144318 8256 157215 8258
rect 144318 8200 157154 8256
rect 157210 8200 157215 8256
rect 144318 8198 157215 8200
rect 134057 8195 134123 8198
rect 138013 8195 138079 8198
rect 157149 8195 157215 8198
rect 157425 8258 157491 8261
rect 163129 8258 163195 8261
rect 157425 8256 163195 8258
rect 157425 8200 157430 8256
rect 157486 8200 163134 8256
rect 163190 8200 163195 8256
rect 157425 8198 163195 8200
rect 157425 8195 157491 8198
rect 163129 8195 163195 8198
rect 163313 8258 163379 8261
rect 167177 8258 167243 8261
rect 176377 8258 176443 8261
rect 163313 8256 167010 8258
rect 163313 8200 163318 8256
rect 163374 8200 167010 8256
rect 163313 8198 167010 8200
rect 163313 8195 163379 8198
rect 24071 8192 24137 8193
rect 64071 8192 64137 8193
rect 104071 8192 104137 8193
rect 144071 8192 144137 8193
rect 24066 8128 24072 8192
rect 24136 8128 24142 8192
rect 64066 8128 64072 8192
rect 64136 8128 64142 8192
rect 104066 8128 104072 8192
rect 104136 8128 104142 8192
rect 144066 8128 144072 8192
rect 144136 8128 144142 8192
rect 24071 8127 24137 8128
rect 64071 8127 64137 8128
rect 104071 8127 104137 8128
rect 144071 8127 144137 8128
rect 105261 8122 105327 8125
rect 114461 8122 114527 8125
rect 105261 8120 114527 8122
rect 105261 8064 105266 8120
rect 105322 8064 114466 8120
rect 114522 8064 114527 8120
rect 105261 8062 114527 8064
rect 105261 8059 105327 8062
rect 114461 8059 114527 8062
rect 132769 8122 132835 8125
rect 134977 8122 135043 8125
rect 132769 8120 135043 8122
rect 132769 8064 132774 8120
rect 132830 8064 134982 8120
rect 135038 8064 135043 8120
rect 132769 8062 135043 8064
rect 132769 8059 132835 8062
rect 134977 8059 135043 8062
rect 135161 8122 135227 8125
rect 142797 8122 142863 8125
rect 157517 8122 157583 8125
rect 161974 8122 161980 8124
rect 135161 8120 142863 8122
rect 135161 8064 135166 8120
rect 135222 8064 142802 8120
rect 142858 8064 142863 8120
rect 135161 8062 142863 8064
rect 135161 8059 135227 8062
rect 142797 8059 142863 8062
rect 149654 8120 157583 8122
rect 149654 8064 157522 8120
rect 157578 8064 157583 8120
rect 149654 8062 157583 8064
rect 107561 7986 107627 7989
rect 137829 7986 137895 7989
rect 107561 7984 137895 7986
rect 107561 7928 107566 7984
rect 107622 7928 137834 7984
rect 137890 7928 137895 7984
rect 107561 7926 137895 7928
rect 107561 7923 107627 7926
rect 137829 7923 137895 7926
rect 138013 7986 138079 7989
rect 149654 7986 149714 8062
rect 157517 8059 157583 8062
rect 157704 8062 161980 8122
rect 138013 7984 149714 7986
rect 138013 7928 138018 7984
rect 138074 7928 149714 7984
rect 138013 7926 149714 7928
rect 152365 7986 152431 7989
rect 157057 7986 157123 7989
rect 157704 7986 157764 8062
rect 161974 8060 161980 8062
rect 162044 8060 162050 8124
rect 162117 8122 162183 8125
rect 166809 8122 166875 8125
rect 162117 8120 166875 8122
rect 162117 8064 162122 8120
rect 162178 8064 166814 8120
rect 166870 8064 166875 8120
rect 162117 8062 166875 8064
rect 166950 8122 167010 8198
rect 167177 8256 176443 8258
rect 167177 8200 167182 8256
rect 167238 8200 176382 8256
rect 176438 8200 176443 8256
rect 167177 8198 176443 8200
rect 167177 8195 167243 8198
rect 176377 8195 176443 8198
rect 176745 8258 176811 8261
rect 180149 8258 180215 8261
rect 176745 8256 180215 8258
rect 176745 8200 176750 8256
rect 176806 8200 180154 8256
rect 180210 8200 180215 8256
rect 176745 8198 180215 8200
rect 176745 8195 176811 8198
rect 180149 8195 180215 8198
rect 180609 8258 180675 8261
rect 183878 8258 183938 8334
rect 180609 8256 183938 8258
rect 180609 8200 180614 8256
rect 180670 8200 183938 8256
rect 180609 8198 183938 8200
rect 184246 8258 184306 8334
rect 185301 8258 185367 8261
rect 184246 8256 185367 8258
rect 184246 8200 185306 8256
rect 185362 8200 185367 8256
rect 184246 8198 185367 8200
rect 180609 8195 180675 8198
rect 185301 8195 185367 8198
rect 184071 8192 184137 8193
rect 184066 8128 184072 8192
rect 184136 8128 184142 8192
rect 184071 8127 184137 8128
rect 169385 8122 169451 8125
rect 166950 8120 169451 8122
rect 166950 8064 169390 8120
rect 169446 8064 169451 8120
rect 166950 8062 169451 8064
rect 162117 8059 162183 8062
rect 166809 8059 166875 8062
rect 169385 8059 169451 8062
rect 170029 8122 170095 8125
rect 181253 8122 181319 8125
rect 170029 8120 181319 8122
rect 170029 8064 170034 8120
rect 170090 8064 181258 8120
rect 181314 8064 181319 8120
rect 170029 8062 181319 8064
rect 170029 8059 170095 8062
rect 181253 8059 181319 8062
rect 182449 8122 182515 8125
rect 183277 8122 183343 8125
rect 182449 8120 183343 8122
rect 182449 8064 182454 8120
rect 182510 8064 183282 8120
rect 183338 8064 183343 8120
rect 182449 8062 183343 8064
rect 182449 8059 182515 8062
rect 183277 8059 183343 8062
rect 152365 7984 157123 7986
rect 152365 7928 152370 7984
rect 152426 7928 157062 7984
rect 157118 7928 157123 7984
rect 152365 7926 157123 7928
rect 138013 7923 138079 7926
rect 152365 7923 152431 7926
rect 157057 7923 157123 7926
rect 157198 7926 157764 7986
rect 159817 7986 159883 7989
rect 191649 7986 191715 7989
rect 159817 7984 191715 7986
rect 159817 7928 159822 7984
rect 159878 7928 191654 7984
rect 191710 7928 191715 7984
rect 159817 7926 191715 7928
rect 103881 7850 103947 7853
rect 134057 7850 134123 7853
rect 103881 7848 134123 7850
rect 103881 7792 103886 7848
rect 103942 7792 134062 7848
rect 134118 7792 134123 7848
rect 103881 7790 134123 7792
rect 103881 7787 103947 7790
rect 134057 7787 134123 7790
rect 134609 7850 134675 7853
rect 137921 7850 137987 7853
rect 134609 7848 137987 7850
rect 134609 7792 134614 7848
rect 134670 7792 137926 7848
rect 137982 7792 137987 7848
rect 134609 7790 137987 7792
rect 134609 7787 134675 7790
rect 137921 7787 137987 7790
rect 138105 7850 138171 7853
rect 140681 7850 140747 7853
rect 138105 7848 140747 7850
rect 138105 7792 138110 7848
rect 138166 7792 140686 7848
rect 140742 7792 140747 7848
rect 138105 7790 140747 7792
rect 138105 7787 138171 7790
rect 140681 7787 140747 7790
rect 142797 7850 142863 7853
rect 156873 7850 156939 7853
rect 157198 7850 157258 7926
rect 159817 7923 159883 7926
rect 191649 7923 191715 7926
rect 142797 7848 156939 7850
rect 142797 7792 142802 7848
rect 142858 7792 156878 7848
rect 156934 7792 156939 7848
rect 142797 7790 156939 7792
rect 142797 7787 142863 7790
rect 156873 7787 156939 7790
rect 157014 7790 157258 7850
rect 157609 7850 157675 7853
rect 161197 7850 161263 7853
rect 165429 7850 165495 7853
rect 167126 7850 167132 7852
rect 157609 7848 157994 7850
rect 157609 7792 157614 7848
rect 157670 7792 157994 7848
rect 157609 7790 157994 7792
rect 105353 7714 105419 7717
rect 123845 7714 123911 7717
rect 105353 7712 123911 7714
rect 105353 7656 105358 7712
rect 105414 7656 123850 7712
rect 123906 7656 123911 7712
rect 105353 7654 123911 7656
rect 105353 7651 105419 7654
rect 123845 7651 123911 7654
rect 125869 7714 125935 7717
rect 136725 7714 136791 7717
rect 125869 7712 136791 7714
rect 125869 7656 125874 7712
rect 125930 7656 136730 7712
rect 136786 7656 136791 7712
rect 125869 7654 136791 7656
rect 125869 7651 125935 7654
rect 136725 7651 136791 7654
rect 137369 7714 137435 7717
rect 152365 7714 152431 7717
rect 137369 7712 152431 7714
rect 137369 7656 137374 7712
rect 137430 7656 152370 7712
rect 152426 7656 152431 7712
rect 137369 7654 152431 7656
rect 137369 7651 137435 7654
rect 152365 7651 152431 7654
rect 152549 7714 152615 7717
rect 156413 7714 156479 7717
rect 152549 7712 156479 7714
rect 152549 7656 152554 7712
rect 152610 7656 156418 7712
rect 156474 7656 156479 7712
rect 152549 7654 156479 7656
rect 152549 7651 152615 7654
rect 156413 7651 156479 7654
rect 156597 7714 156663 7717
rect 157014 7714 157074 7790
rect 157609 7787 157675 7790
rect 156597 7712 157074 7714
rect 156597 7656 156602 7712
rect 156658 7656 157074 7712
rect 156597 7654 157074 7656
rect 156597 7651 156663 7654
rect 157190 7652 157196 7716
rect 157260 7714 157266 7716
rect 157934 7714 157994 7790
rect 161197 7848 164434 7850
rect 161197 7792 161202 7848
rect 161258 7792 164434 7848
rect 161197 7790 164434 7792
rect 161197 7787 161263 7790
rect 162669 7714 162735 7717
rect 157260 7654 157626 7714
rect 157934 7712 162735 7714
rect 157934 7656 162674 7712
rect 162730 7656 162735 7712
rect 157934 7654 162735 7656
rect 164374 7714 164434 7790
rect 165429 7848 167132 7850
rect 165429 7792 165434 7848
rect 165490 7792 167132 7848
rect 165429 7790 167132 7792
rect 165429 7787 165495 7790
rect 167126 7788 167132 7790
rect 167196 7788 167202 7852
rect 167310 7788 167316 7852
rect 167380 7850 167386 7852
rect 173617 7850 173683 7853
rect 167380 7848 173683 7850
rect 167380 7792 173622 7848
rect 173678 7792 173683 7848
rect 167380 7790 173683 7792
rect 167380 7788 167386 7790
rect 173617 7787 173683 7790
rect 175590 7788 175596 7852
rect 175660 7850 175666 7852
rect 176561 7850 176627 7853
rect 175660 7848 176627 7850
rect 175660 7792 176566 7848
rect 176622 7792 176627 7848
rect 175660 7790 176627 7792
rect 175660 7788 175666 7790
rect 176561 7787 176627 7790
rect 177481 7850 177547 7853
rect 180609 7850 180675 7853
rect 185025 7850 185091 7853
rect 177481 7848 180675 7850
rect 177481 7792 177486 7848
rect 177542 7792 180614 7848
rect 180670 7792 180675 7848
rect 177481 7790 180675 7792
rect 177481 7787 177547 7790
rect 180609 7787 180675 7790
rect 180750 7848 185091 7850
rect 180750 7792 185030 7848
rect 185086 7792 185091 7848
rect 180750 7790 185091 7792
rect 180750 7714 180810 7790
rect 185025 7787 185091 7790
rect 164374 7654 180810 7714
rect 180885 7714 180951 7717
rect 182817 7714 182883 7717
rect 183553 7716 183619 7717
rect 180885 7712 182883 7714
rect 180885 7656 180890 7712
rect 180946 7656 182822 7712
rect 182878 7656 182883 7712
rect 180885 7654 182883 7656
rect 157260 7652 157266 7654
rect 4071 7648 4137 7649
rect 44071 7648 44137 7649
rect 84071 7648 84137 7649
rect 124071 7648 124137 7649
rect 4066 7584 4072 7648
rect 4136 7584 4142 7648
rect 44066 7584 44072 7648
rect 44136 7584 44142 7648
rect 84066 7584 84072 7648
rect 84136 7584 84142 7648
rect 124066 7584 124072 7648
rect 124136 7584 124142 7648
rect 4071 7583 4137 7584
rect 44071 7583 44137 7584
rect 84071 7583 84137 7584
rect 124071 7583 124137 7584
rect 93761 7578 93827 7581
rect 114001 7578 114067 7581
rect 93761 7576 114067 7578
rect 93761 7520 93766 7576
rect 93822 7520 114006 7576
rect 114062 7520 114067 7576
rect 93761 7518 114067 7520
rect 93761 7515 93827 7518
rect 114001 7515 114067 7518
rect 129365 7578 129431 7581
rect 133965 7578 134031 7581
rect 129365 7576 134031 7578
rect 129365 7520 129370 7576
rect 129426 7520 133970 7576
rect 134026 7520 134031 7576
rect 129365 7518 134031 7520
rect 129365 7515 129431 7518
rect 133965 7515 134031 7518
rect 134149 7578 134215 7581
rect 140313 7578 140379 7581
rect 134149 7576 140379 7578
rect 134149 7520 134154 7576
rect 134210 7520 140318 7576
rect 140374 7520 140379 7576
rect 134149 7518 140379 7520
rect 134149 7515 134215 7518
rect 140313 7515 140379 7518
rect 140497 7578 140563 7581
rect 157425 7578 157491 7581
rect 140497 7576 157491 7578
rect 140497 7520 140502 7576
rect 140558 7520 157430 7576
rect 157486 7520 157491 7576
rect 140497 7518 157491 7520
rect 157566 7578 157626 7654
rect 162669 7651 162735 7654
rect 180885 7651 180951 7654
rect 182817 7651 182883 7654
rect 183502 7652 183508 7716
rect 183572 7714 183619 7716
rect 183572 7712 183664 7714
rect 183614 7656 183664 7712
rect 183572 7654 183664 7656
rect 183572 7652 183619 7654
rect 183553 7651 183619 7652
rect 164071 7648 164137 7649
rect 164066 7584 164072 7648
rect 164136 7584 164142 7648
rect 164071 7583 164137 7584
rect 163313 7578 163379 7581
rect 157566 7576 163379 7578
rect 157566 7520 163318 7576
rect 163374 7520 163379 7576
rect 157566 7518 163379 7520
rect 140497 7515 140563 7518
rect 157425 7515 157491 7518
rect 163313 7515 163379 7518
rect 164969 7578 165035 7581
rect 165102 7578 165108 7580
rect 164969 7576 165108 7578
rect 164969 7520 164974 7576
rect 165030 7520 165108 7576
rect 164969 7518 165108 7520
rect 164969 7515 165035 7518
rect 165102 7516 165108 7518
rect 165172 7516 165178 7580
rect 165613 7578 165679 7581
rect 166022 7578 166028 7580
rect 165613 7576 166028 7578
rect 165613 7520 165618 7576
rect 165674 7520 166028 7576
rect 165613 7518 166028 7520
rect 165613 7515 165679 7518
rect 166022 7516 166028 7518
rect 166092 7516 166098 7580
rect 167361 7578 167427 7581
rect 174261 7578 174327 7581
rect 166398 7576 167427 7578
rect 166398 7520 167366 7576
rect 167422 7520 167427 7576
rect 166398 7518 167427 7520
rect 93301 7442 93367 7445
rect 96153 7442 96219 7445
rect 93301 7440 96219 7442
rect 93301 7384 93306 7440
rect 93362 7384 96158 7440
rect 96214 7384 96219 7440
rect 93301 7382 96219 7384
rect 93301 7379 93367 7382
rect 96153 7379 96219 7382
rect 98453 7442 98519 7445
rect 142153 7442 142219 7445
rect 98453 7440 142219 7442
rect 98453 7384 98458 7440
rect 98514 7384 142158 7440
rect 142214 7384 142219 7440
rect 98453 7382 142219 7384
rect 98453 7379 98519 7382
rect 142153 7379 142219 7382
rect 143441 7442 143507 7445
rect 156873 7442 156939 7445
rect 143441 7440 156939 7442
rect 143441 7384 143446 7440
rect 143502 7384 156878 7440
rect 156934 7384 156939 7440
rect 143441 7382 156939 7384
rect 143441 7379 143507 7382
rect 156873 7379 156939 7382
rect 157006 7380 157012 7444
rect 157076 7442 157082 7444
rect 157517 7442 157583 7445
rect 157076 7440 157583 7442
rect 157076 7384 157522 7440
rect 157578 7384 157583 7440
rect 157076 7382 157583 7384
rect 157076 7380 157082 7382
rect 157517 7379 157583 7382
rect 157701 7442 157767 7445
rect 158897 7444 158963 7445
rect 158662 7442 158668 7444
rect 157701 7440 158668 7442
rect 157701 7384 157706 7440
rect 157762 7384 158668 7440
rect 157701 7382 158668 7384
rect 157701 7379 157767 7382
rect 158662 7380 158668 7382
rect 158732 7380 158738 7444
rect 158846 7442 158852 7444
rect 158806 7382 158852 7442
rect 158916 7440 158963 7444
rect 158958 7384 158963 7440
rect 158846 7380 158852 7382
rect 158916 7380 158963 7384
rect 158897 7379 158963 7380
rect 159909 7444 159975 7445
rect 159909 7440 159956 7444
rect 160020 7442 160026 7444
rect 159909 7384 159914 7440
rect 159909 7380 159956 7384
rect 160020 7382 160066 7442
rect 160020 7380 160026 7382
rect 161422 7380 161428 7444
rect 161492 7442 161498 7444
rect 162577 7442 162643 7445
rect 164693 7444 164759 7445
rect 164693 7442 164740 7444
rect 161492 7440 162643 7442
rect 161492 7384 162582 7440
rect 162638 7384 162643 7440
rect 161492 7382 162643 7384
rect 164648 7440 164740 7442
rect 164648 7384 164698 7440
rect 164648 7382 164740 7384
rect 161492 7380 161498 7382
rect 159909 7379 159975 7380
rect 162577 7379 162643 7382
rect 164693 7380 164740 7382
rect 164804 7380 164810 7444
rect 164877 7442 164943 7445
rect 165838 7442 165844 7444
rect 164877 7440 165844 7442
rect 164877 7384 164882 7440
rect 164938 7384 165844 7440
rect 164877 7382 165844 7384
rect 164693 7379 164759 7380
rect 164877 7379 164943 7382
rect 165838 7380 165844 7382
rect 165908 7380 165914 7444
rect 68737 7306 68803 7309
rect 118785 7306 118851 7309
rect 68737 7304 118851 7306
rect 68737 7248 68742 7304
rect 68798 7248 118790 7304
rect 118846 7248 118851 7304
rect 68737 7246 118851 7248
rect 68737 7243 68803 7246
rect 118785 7243 118851 7246
rect 124254 7244 124260 7308
rect 124324 7306 124330 7308
rect 127249 7306 127315 7309
rect 124324 7304 127315 7306
rect 124324 7248 127254 7304
rect 127310 7248 127315 7304
rect 124324 7246 127315 7248
rect 124324 7244 124330 7246
rect 127249 7243 127315 7246
rect 127617 7306 127683 7309
rect 130469 7306 130535 7309
rect 127617 7304 130535 7306
rect 127617 7248 127622 7304
rect 127678 7248 130474 7304
rect 130530 7248 130535 7304
rect 127617 7246 130535 7248
rect 127617 7243 127683 7246
rect 130469 7243 130535 7246
rect 131757 7306 131823 7309
rect 142705 7306 142771 7309
rect 157374 7306 157380 7308
rect 131757 7304 142771 7306
rect 131757 7248 131762 7304
rect 131818 7248 142710 7304
rect 142766 7248 142771 7304
rect 131757 7246 142771 7248
rect 131757 7243 131823 7246
rect 142705 7243 142771 7246
rect 142846 7246 157380 7306
rect 107469 7170 107535 7173
rect 114277 7170 114343 7173
rect 107469 7168 114343 7170
rect 107469 7112 107474 7168
rect 107530 7112 114282 7168
rect 114338 7112 114343 7168
rect 107469 7110 114343 7112
rect 107469 7107 107535 7110
rect 114277 7107 114343 7110
rect 118601 7170 118667 7173
rect 124765 7170 124831 7173
rect 118601 7168 124831 7170
rect 118601 7112 118606 7168
rect 118662 7112 124770 7168
rect 124826 7112 124831 7168
rect 118601 7110 124831 7112
rect 118601 7107 118667 7110
rect 124765 7107 124831 7110
rect 128445 7170 128511 7173
rect 133965 7170 134031 7173
rect 128445 7168 134031 7170
rect 128445 7112 128450 7168
rect 128506 7112 133970 7168
rect 134026 7112 134031 7168
rect 128445 7110 134031 7112
rect 128445 7107 128511 7110
rect 133965 7107 134031 7110
rect 134149 7170 134215 7173
rect 137001 7170 137067 7173
rect 134149 7168 137067 7170
rect 134149 7112 134154 7168
rect 134210 7112 137006 7168
rect 137062 7112 137067 7168
rect 134149 7110 137067 7112
rect 134149 7107 134215 7110
rect 137001 7107 137067 7110
rect 137553 7170 137619 7173
rect 142846 7170 142906 7246
rect 157374 7244 157380 7246
rect 157444 7244 157450 7308
rect 166398 7306 166458 7518
rect 167361 7515 167427 7518
rect 167502 7576 174327 7578
rect 167502 7520 174266 7576
rect 174322 7520 174327 7576
rect 167502 7518 174327 7520
rect 166533 7442 166599 7445
rect 167502 7442 167562 7518
rect 174261 7515 174327 7518
rect 174445 7578 174511 7581
rect 176469 7580 176535 7581
rect 175038 7578 175044 7580
rect 174445 7576 175044 7578
rect 174445 7520 174450 7576
rect 174506 7520 175044 7576
rect 174445 7518 175044 7520
rect 174445 7515 174511 7518
rect 175038 7516 175044 7518
rect 175108 7516 175114 7580
rect 176469 7576 176516 7580
rect 176580 7578 176586 7580
rect 182081 7578 182147 7581
rect 185393 7578 185459 7581
rect 176469 7520 176474 7576
rect 176469 7516 176516 7520
rect 176580 7518 176626 7578
rect 182081 7576 185459 7578
rect 182081 7520 182086 7576
rect 182142 7520 185398 7576
rect 185454 7520 185459 7576
rect 182081 7518 185459 7520
rect 176580 7516 176586 7518
rect 176469 7515 176535 7516
rect 182081 7515 182147 7518
rect 185393 7515 185459 7518
rect 167729 7444 167795 7445
rect 167678 7442 167684 7444
rect 166533 7440 167562 7442
rect 166533 7384 166538 7440
rect 166594 7384 167562 7440
rect 166533 7382 167562 7384
rect 167638 7382 167684 7442
rect 167748 7440 167795 7444
rect 167790 7384 167795 7440
rect 166533 7379 166599 7382
rect 167678 7380 167684 7382
rect 167748 7380 167795 7384
rect 167729 7379 167795 7380
rect 169109 7440 169175 7445
rect 169109 7384 169114 7440
rect 169170 7384 169175 7440
rect 169109 7379 169175 7384
rect 169385 7440 169451 7445
rect 169753 7444 169819 7445
rect 169702 7442 169708 7444
rect 169385 7384 169390 7440
rect 169446 7384 169451 7440
rect 169385 7379 169451 7384
rect 169662 7382 169708 7442
rect 169772 7440 169819 7444
rect 170029 7444 170095 7445
rect 171225 7444 171291 7445
rect 171409 7444 171475 7445
rect 171777 7444 171843 7445
rect 170029 7442 170076 7444
rect 169814 7384 169819 7440
rect 169702 7380 169708 7382
rect 169772 7380 169819 7384
rect 169984 7440 170076 7442
rect 169984 7384 170034 7440
rect 169984 7382 170076 7384
rect 169753 7379 169819 7380
rect 170029 7380 170076 7382
rect 170140 7380 170146 7444
rect 171174 7442 171180 7444
rect 171134 7382 171180 7442
rect 171244 7440 171291 7444
rect 171286 7384 171291 7440
rect 171174 7380 171180 7382
rect 171244 7380 171291 7384
rect 171358 7380 171364 7444
rect 171428 7442 171475 7444
rect 171726 7442 171732 7444
rect 171428 7440 171520 7442
rect 171470 7384 171520 7440
rect 171428 7382 171520 7384
rect 171686 7382 171732 7442
rect 171796 7440 171843 7444
rect 171838 7384 171843 7440
rect 171428 7380 171475 7382
rect 171726 7380 171732 7382
rect 171796 7380 171843 7384
rect 172462 7380 172468 7444
rect 172532 7442 172538 7444
rect 172605 7442 172671 7445
rect 172532 7440 172671 7442
rect 172532 7384 172610 7440
rect 172666 7384 172671 7440
rect 172532 7382 172671 7384
rect 172532 7380 172538 7382
rect 170029 7379 170095 7380
rect 171225 7379 171291 7380
rect 171409 7379 171475 7380
rect 171777 7379 171843 7380
rect 172605 7379 172671 7382
rect 173382 7380 173388 7444
rect 173452 7442 173458 7444
rect 173525 7442 173591 7445
rect 174905 7444 174971 7445
rect 174854 7442 174860 7444
rect 173452 7440 173591 7442
rect 173452 7384 173530 7440
rect 173586 7384 173591 7440
rect 173452 7382 173591 7384
rect 174814 7382 174860 7442
rect 174924 7440 174971 7444
rect 174966 7384 174971 7440
rect 173452 7380 173458 7382
rect 173525 7379 173591 7382
rect 174854 7380 174860 7382
rect 174924 7380 174971 7384
rect 174905 7379 174971 7380
rect 175457 7442 175523 7445
rect 175774 7442 175780 7444
rect 175457 7440 175780 7442
rect 175457 7384 175462 7440
rect 175518 7384 175780 7440
rect 175457 7382 175780 7384
rect 175457 7379 175523 7382
rect 175774 7380 175780 7382
rect 175844 7380 175850 7444
rect 177062 7380 177068 7444
rect 177132 7442 177138 7444
rect 177941 7442 178007 7445
rect 177132 7440 178007 7442
rect 177132 7384 177946 7440
rect 178002 7384 178007 7440
rect 177132 7382 178007 7384
rect 177132 7380 177138 7382
rect 177941 7379 178007 7382
rect 178401 7440 178467 7445
rect 178401 7384 178406 7440
rect 178462 7384 178467 7440
rect 178401 7379 178467 7384
rect 180742 7380 180748 7444
rect 180812 7442 180818 7444
rect 181161 7442 181227 7445
rect 181989 7444 182055 7445
rect 182265 7444 182331 7445
rect 181989 7442 182036 7444
rect 180812 7440 181227 7442
rect 180812 7384 181166 7440
rect 181222 7384 181227 7440
rect 180812 7382 181227 7384
rect 181944 7440 182036 7442
rect 181944 7384 181994 7440
rect 181944 7382 182036 7384
rect 180812 7380 180818 7382
rect 181161 7379 181227 7382
rect 181989 7380 182036 7382
rect 182100 7380 182106 7444
rect 182214 7442 182220 7444
rect 182174 7382 182220 7442
rect 182284 7440 182331 7444
rect 182326 7384 182331 7440
rect 182214 7380 182220 7382
rect 182284 7380 182331 7384
rect 182398 7380 182404 7444
rect 182468 7442 182474 7444
rect 184289 7442 184355 7445
rect 182468 7440 184355 7442
rect 182468 7384 184294 7440
rect 184350 7384 184355 7440
rect 182468 7382 184355 7384
rect 182468 7380 182474 7382
rect 181989 7379 182055 7380
rect 182265 7379 182331 7380
rect 184289 7379 184355 7382
rect 169112 7306 169172 7379
rect 157934 7246 166458 7306
rect 167916 7246 169172 7306
rect 169388 7306 169448 7379
rect 177481 7306 177547 7309
rect 177849 7308 177915 7309
rect 177798 7306 177804 7308
rect 169388 7304 177547 7306
rect 169388 7248 177486 7304
rect 177542 7248 177547 7304
rect 169388 7246 177547 7248
rect 177758 7246 177804 7306
rect 177868 7304 177915 7308
rect 177910 7248 177915 7304
rect 137553 7168 142906 7170
rect 137553 7112 137558 7168
rect 137614 7112 142906 7168
rect 137553 7110 142906 7112
rect 144269 7170 144335 7173
rect 155585 7170 155651 7173
rect 157934 7170 157994 7246
rect 167916 7170 167976 7246
rect 177481 7243 177547 7246
rect 177798 7244 177804 7246
rect 177868 7244 177915 7248
rect 178404 7306 178464 7379
rect 194869 7306 194935 7309
rect 178404 7304 194935 7306
rect 178404 7248 194874 7304
rect 194930 7248 194935 7304
rect 178404 7246 194935 7248
rect 177849 7243 177915 7244
rect 194869 7243 194935 7246
rect 144269 7168 155651 7170
rect 144269 7112 144274 7168
rect 144330 7112 155590 7168
rect 155646 7112 155651 7168
rect 144269 7110 155651 7112
rect 137553 7107 137619 7110
rect 144269 7107 144335 7110
rect 155585 7107 155651 7110
rect 156462 7110 157994 7170
rect 158118 7110 167976 7170
rect 24071 7104 24137 7105
rect 64071 7104 64137 7105
rect 104071 7104 104137 7105
rect 144071 7104 144137 7105
rect 24066 7040 24072 7104
rect 24136 7040 24142 7104
rect 64066 7040 64072 7104
rect 64136 7040 64142 7104
rect 104066 7040 104072 7104
rect 104136 7040 104142 7104
rect 144066 7040 144072 7104
rect 144136 7040 144142 7104
rect 24071 7039 24137 7040
rect 64071 7039 64137 7040
rect 104071 7039 104137 7040
rect 144071 7039 144137 7040
rect 109585 7034 109651 7037
rect 133781 7034 133847 7037
rect 109585 7032 133847 7034
rect 109585 6976 109590 7032
rect 109646 6976 133786 7032
rect 133842 6976 133847 7032
rect 109585 6974 133847 6976
rect 109585 6971 109651 6974
rect 133781 6971 133847 6974
rect 134609 7034 134675 7037
rect 134977 7034 135043 7037
rect 134609 7032 135043 7034
rect 134609 6976 134614 7032
rect 134670 6976 134982 7032
rect 135038 6976 135043 7032
rect 134609 6974 135043 6976
rect 134609 6971 134675 6974
rect 134977 6971 135043 6974
rect 135621 7034 135687 7037
rect 155769 7034 155835 7037
rect 135621 7032 143964 7034
rect 135621 6976 135626 7032
rect 135682 6976 143964 7032
rect 135621 6974 143964 6976
rect 135621 6971 135687 6974
rect 99189 6898 99255 6901
rect 99741 6898 99807 6901
rect 99189 6896 99807 6898
rect 99189 6840 99194 6896
rect 99250 6840 99746 6896
rect 99802 6840 99807 6896
rect 99189 6838 99807 6840
rect 99189 6835 99255 6838
rect 99741 6835 99807 6838
rect 108113 6898 108179 6901
rect 135164 6898 135362 6932
rect 143625 6898 143691 6901
rect 108113 6896 143691 6898
rect 108113 6840 108118 6896
rect 108174 6872 143630 6896
rect 108174 6840 135224 6872
rect 108113 6838 135224 6840
rect 135302 6840 143630 6872
rect 143686 6840 143691 6896
rect 135302 6838 143691 6840
rect 143904 6898 143964 6974
rect 144318 7032 155835 7034
rect 144318 6976 155774 7032
rect 155830 6976 155835 7032
rect 144318 6974 155835 6976
rect 144318 6898 144378 6974
rect 155769 6971 155835 6974
rect 149145 6898 149211 6901
rect 143904 6838 144378 6898
rect 147078 6896 149211 6898
rect 147078 6840 149150 6896
rect 149206 6840 149211 6896
rect 147078 6838 149211 6840
rect 108113 6835 108179 6838
rect 143625 6835 143691 6838
rect 98269 6762 98335 6765
rect 99741 6762 99807 6765
rect 98269 6760 99807 6762
rect 98269 6704 98274 6760
rect 98330 6704 99746 6760
rect 99802 6704 99807 6760
rect 98269 6702 99807 6704
rect 98269 6699 98335 6702
rect 99741 6699 99807 6702
rect 122741 6762 122807 6765
rect 124208 6762 124214 6764
rect 122741 6760 124214 6762
rect 122741 6704 122746 6760
rect 122802 6704 124214 6760
rect 122741 6702 124214 6704
rect 122741 6699 122807 6702
rect 124208 6700 124214 6702
rect 124278 6700 124284 6764
rect 125961 6762 126027 6765
rect 127525 6762 127591 6765
rect 125961 6760 127591 6762
rect 125961 6704 125966 6760
rect 126022 6704 127530 6760
rect 127586 6704 127591 6760
rect 125961 6702 127591 6704
rect 125961 6699 126027 6702
rect 127525 6699 127591 6702
rect 127709 6762 127775 6765
rect 134742 6762 134748 6764
rect 127709 6760 134748 6762
rect 127709 6704 127714 6760
rect 127770 6704 134748 6760
rect 127709 6702 134748 6704
rect 127709 6699 127775 6702
rect 134742 6700 134748 6702
rect 134812 6700 134818 6764
rect 134977 6762 135043 6765
rect 147078 6762 147138 6838
rect 149145 6835 149211 6838
rect 153101 6898 153167 6901
rect 156462 6898 156522 7110
rect 156965 7034 157031 7037
rect 158118 7034 158178 7110
rect 168046 7108 168052 7172
rect 168116 7170 168122 7172
rect 192661 7170 192727 7173
rect 168116 7168 192727 7170
rect 168116 7112 192666 7168
rect 192722 7112 192727 7168
rect 168116 7110 192727 7112
rect 168116 7108 168122 7110
rect 192661 7107 192727 7110
rect 156965 7032 158178 7034
rect 156965 6976 156970 7032
rect 157026 6976 158178 7032
rect 156965 6974 158178 6976
rect 156965 6971 157031 6974
rect 158662 6972 158668 7036
rect 158732 7034 158738 7036
rect 182398 7034 182404 7036
rect 158732 6974 182404 7034
rect 158732 6972 158738 6974
rect 182398 6972 182404 6974
rect 182468 6972 182474 7036
rect 153101 6896 156522 6898
rect 153101 6840 153106 6896
rect 153162 6840 156522 6896
rect 153101 6838 156522 6840
rect 153101 6835 153167 6838
rect 134977 6760 147138 6762
rect 134977 6704 134982 6760
rect 135038 6704 147138 6760
rect 134977 6702 147138 6704
rect 148685 6762 148751 6765
rect 155769 6762 155835 6765
rect 148685 6760 155835 6762
rect 148685 6704 148690 6760
rect 148746 6704 155774 6760
rect 155830 6704 155835 6760
rect 148685 6702 155835 6704
rect 134977 6699 135043 6702
rect 148685 6699 148751 6702
rect 155769 6699 155835 6702
rect 131021 6626 131087 6629
rect 133321 6626 133387 6629
rect 131021 6624 133387 6626
rect 131021 6568 131026 6624
rect 131082 6568 133326 6624
rect 133382 6568 133387 6624
rect 131021 6566 133387 6568
rect 131021 6563 131087 6566
rect 133321 6563 133387 6566
rect 133505 6626 133571 6629
rect 140221 6626 140287 6629
rect 133505 6624 140287 6626
rect 133505 6568 133510 6624
rect 133566 6568 140226 6624
rect 140282 6568 140287 6624
rect 133505 6566 140287 6568
rect 133505 6563 133571 6566
rect 140221 6563 140287 6566
rect 140405 6626 140471 6629
rect 150525 6626 150591 6629
rect 140405 6624 150591 6626
rect 140405 6568 140410 6624
rect 140466 6568 150530 6624
rect 150586 6568 150591 6624
rect 140405 6566 150591 6568
rect 140405 6563 140471 6566
rect 150525 6563 150591 6566
rect 151721 6626 151787 6629
rect 157057 6626 157123 6629
rect 151721 6624 157123 6626
rect 151721 6568 151726 6624
rect 151782 6568 157062 6624
rect 157118 6568 157123 6624
rect 151721 6566 157123 6568
rect 151721 6563 151787 6566
rect 157057 6563 157123 6566
rect 4071 6560 4137 6561
rect 44071 6560 44137 6561
rect 84071 6560 84137 6561
rect 124071 6560 124137 6561
rect 4066 6496 4072 6560
rect 4136 6496 4142 6560
rect 44066 6496 44072 6560
rect 44136 6496 44142 6560
rect 84066 6496 84072 6560
rect 84136 6496 84142 6560
rect 124066 6496 124072 6560
rect 124136 6496 124142 6560
rect 4071 6495 4137 6496
rect 44071 6495 44137 6496
rect 84071 6495 84137 6496
rect 124071 6495 124137 6496
rect 108757 6490 108823 6493
rect 109125 6490 109191 6493
rect 108757 6488 109191 6490
rect 108757 6432 108762 6488
rect 108818 6432 109130 6488
rect 109186 6432 109191 6488
rect 108757 6430 109191 6432
rect 108757 6427 108823 6430
rect 109125 6427 109191 6430
rect 114461 6490 114527 6493
rect 123753 6490 123819 6493
rect 114461 6488 123819 6490
rect 114461 6432 114466 6488
rect 114522 6432 123758 6488
rect 123814 6432 123819 6488
rect 114461 6430 123819 6432
rect 114461 6427 114527 6430
rect 123753 6427 123819 6430
rect 127249 6490 127315 6493
rect 134977 6490 135043 6493
rect 127249 6488 135043 6490
rect 127249 6432 127254 6488
rect 127310 6432 134982 6488
rect 135038 6432 135043 6488
rect 127249 6430 135043 6432
rect 127249 6427 127315 6430
rect 134977 6427 135043 6430
rect 135110 6428 135116 6492
rect 135180 6490 135186 6492
rect 151629 6490 151695 6493
rect 156597 6490 156663 6493
rect 135180 6430 149024 6490
rect 135180 6428 135186 6430
rect 97625 6354 97691 6357
rect 99281 6354 99347 6357
rect 97625 6352 99347 6354
rect 97625 6296 97630 6352
rect 97686 6296 99286 6352
rect 99342 6296 99347 6352
rect 97625 6294 99347 6296
rect 97625 6291 97691 6294
rect 99281 6291 99347 6294
rect 114461 6354 114527 6357
rect 134425 6354 134491 6357
rect 138657 6354 138723 6357
rect 144913 6354 144979 6357
rect 114461 6352 134491 6354
rect 114461 6296 114466 6352
rect 114522 6296 134430 6352
rect 134486 6296 134491 6352
rect 114461 6294 134491 6296
rect 114461 6291 114527 6294
rect 134425 6291 134491 6294
rect 134612 6294 135408 6354
rect 81801 6218 81867 6221
rect 82169 6218 82235 6221
rect 81801 6216 82235 6218
rect 81801 6160 81806 6216
rect 81862 6160 82174 6216
rect 82230 6160 82235 6216
rect 81801 6158 82235 6160
rect 81801 6155 81867 6158
rect 82169 6155 82235 6158
rect 97533 6218 97599 6221
rect 99281 6218 99347 6221
rect 97533 6216 99347 6218
rect 97533 6160 97538 6216
rect 97594 6160 99286 6216
rect 99342 6160 99347 6216
rect 97533 6158 99347 6160
rect 97533 6155 97599 6158
rect 99281 6155 99347 6158
rect 99465 6218 99531 6221
rect 102961 6218 103027 6221
rect 99465 6216 103027 6218
rect 99465 6160 99470 6216
rect 99526 6160 102966 6216
rect 103022 6160 103027 6216
rect 99465 6158 103027 6160
rect 99465 6155 99531 6158
rect 102961 6155 103027 6158
rect 114829 6218 114895 6221
rect 118877 6218 118943 6221
rect 114829 6216 118943 6218
rect 114829 6160 114834 6216
rect 114890 6160 118882 6216
rect 118938 6160 118943 6216
rect 114829 6158 118943 6160
rect 114829 6155 114895 6158
rect 118877 6155 118943 6158
rect 119613 6218 119679 6221
rect 124254 6218 124260 6220
rect 119613 6216 124260 6218
rect 119613 6160 119618 6216
rect 119674 6160 124260 6216
rect 119613 6158 124260 6160
rect 119613 6155 119679 6158
rect 124254 6156 124260 6158
rect 124324 6156 124330 6220
rect 124397 6218 124463 6221
rect 127709 6218 127775 6221
rect 134612 6218 134672 6294
rect 135348 6218 135408 6294
rect 138657 6352 144979 6354
rect 138657 6296 138662 6352
rect 138718 6296 144918 6352
rect 144974 6296 144979 6352
rect 138657 6294 144979 6296
rect 148964 6354 149024 6430
rect 151629 6488 156663 6490
rect 151629 6432 151634 6488
rect 151690 6432 156602 6488
rect 156658 6432 156663 6488
rect 151629 6430 156663 6432
rect 151629 6427 151695 6430
rect 156597 6427 156663 6430
rect 157198 6357 157258 6868
rect 185666 6803 185672 6867
rect 185736 6803 185742 6867
rect 164466 6680 164472 6744
rect 164536 6680 164542 6744
rect 185266 6403 185272 6467
rect 185336 6403 185342 6467
rect 153561 6354 153627 6357
rect 148964 6352 153627 6354
rect 148964 6296 153566 6352
rect 153622 6296 153627 6352
rect 148964 6294 153627 6296
rect 138657 6291 138723 6294
rect 144913 6291 144979 6294
rect 153561 6291 153627 6294
rect 157149 6352 157258 6357
rect 157149 6296 157154 6352
rect 157210 6296 157258 6352
rect 157149 6294 157258 6296
rect 157149 6291 157215 6294
rect 144453 6218 144519 6221
rect 155677 6218 155743 6221
rect 124397 6216 127775 6218
rect 124397 6160 124402 6216
rect 124458 6160 127714 6216
rect 127770 6160 127775 6216
rect 124397 6158 127775 6160
rect 124397 6155 124463 6158
rect 127709 6155 127775 6158
rect 129046 6158 134672 6218
rect 134750 6158 135178 6218
rect 135348 6158 144378 6218
rect 96889 6082 96955 6085
rect 100109 6082 100175 6085
rect 96889 6080 100175 6082
rect 96889 6024 96894 6080
rect 96950 6024 100114 6080
rect 100170 6024 100175 6080
rect 96889 6022 100175 6024
rect 96889 6019 96955 6022
rect 100109 6019 100175 6022
rect 109585 6082 109651 6085
rect 111241 6082 111307 6085
rect 109585 6080 111307 6082
rect 109585 6024 109590 6080
rect 109646 6024 111246 6080
rect 111302 6024 111307 6080
rect 109585 6022 111307 6024
rect 109585 6019 109651 6022
rect 111241 6019 111307 6022
rect 118049 6082 118115 6085
rect 129046 6082 129106 6158
rect 134750 6082 134810 6158
rect 118049 6080 129106 6082
rect 118049 6024 118054 6080
rect 118110 6024 129106 6080
rect 118049 6022 129106 6024
rect 133048 6022 134810 6082
rect 135118 6082 135178 6158
rect 142153 6082 142219 6085
rect 135118 6080 142219 6082
rect 135118 6024 142158 6080
rect 142214 6024 142219 6080
rect 135118 6022 142219 6024
rect 144318 6082 144378 6158
rect 144453 6216 155743 6218
rect 144453 6160 144458 6216
rect 144514 6160 155682 6216
rect 155738 6160 155743 6216
rect 144453 6158 155743 6160
rect 144453 6155 144519 6158
rect 155677 6155 155743 6158
rect 151813 6082 151879 6085
rect 144318 6080 151879 6082
rect 144318 6024 151818 6080
rect 151874 6024 151879 6080
rect 165666 6074 165672 6138
rect 165736 6074 165742 6138
rect 144318 6022 151879 6024
rect 118049 6019 118115 6022
rect 24071 6016 24137 6017
rect 64071 6016 64137 6017
rect 104071 6016 104137 6017
rect 24066 5952 24072 6016
rect 24136 5952 24142 6016
rect 64066 5952 64072 6016
rect 64136 5952 64142 6016
rect 104066 5952 104072 6016
rect 104136 5952 104142 6016
rect 24071 5951 24137 5952
rect 64071 5951 64137 5952
rect 104071 5951 104137 5952
rect 99465 5946 99531 5949
rect 102685 5946 102751 5949
rect 99465 5944 102751 5946
rect 99465 5888 99470 5944
rect 99526 5888 102690 5944
rect 102746 5888 102751 5944
rect 99465 5886 102751 5888
rect 99465 5883 99531 5886
rect 102685 5883 102751 5886
rect 109217 5946 109283 5949
rect 133048 5946 133108 6022
rect 142153 6019 142219 6022
rect 151813 6019 151879 6022
rect 144071 6016 144137 6017
rect 144066 5952 144072 6016
rect 144136 5952 144142 6016
rect 184466 5952 184472 6016
rect 184536 5952 184542 6016
rect 144071 5951 144137 5952
rect 109217 5944 133108 5946
rect 109217 5888 109222 5944
rect 109278 5888 133108 5944
rect 109217 5886 133108 5888
rect 134609 5946 134675 5949
rect 134977 5946 135043 5949
rect 138657 5946 138723 5949
rect 134609 5944 135043 5946
rect 134609 5888 134614 5944
rect 134670 5888 134982 5944
rect 135038 5888 135043 5944
rect 135302 5944 138723 5946
rect 135302 5912 138662 5944
rect 134609 5886 135043 5888
rect 109217 5883 109283 5886
rect 134609 5883 134675 5886
rect 134977 5883 135043 5886
rect 135118 5888 138662 5912
rect 138718 5888 138723 5944
rect 135118 5886 138723 5888
rect 135118 5852 135362 5886
rect 138657 5883 138723 5886
rect 99281 5810 99347 5813
rect 104341 5810 104407 5813
rect 99281 5808 104407 5810
rect 99281 5752 99286 5808
rect 99342 5752 104346 5808
rect 104402 5752 104407 5808
rect 99281 5750 104407 5752
rect 99281 5747 99347 5750
rect 104341 5747 104407 5750
rect 108757 5810 108823 5813
rect 135118 5810 135178 5852
rect 144453 5810 144519 5813
rect 108757 5808 135178 5810
rect 108757 5752 108762 5808
rect 108818 5752 135178 5808
rect 135486 5808 144519 5810
rect 135486 5776 144458 5808
rect 108757 5750 135178 5752
rect 135348 5752 144458 5776
rect 144514 5752 144519 5808
rect 135348 5750 144519 5752
rect 108757 5747 108823 5750
rect 135348 5716 135546 5750
rect 144453 5747 144519 5750
rect 108389 5674 108455 5677
rect 114737 5674 114803 5677
rect 108389 5672 114803 5674
rect 108389 5616 108394 5672
rect 108450 5616 114742 5672
rect 114798 5616 114803 5672
rect 108389 5614 114803 5616
rect 108389 5611 108455 5614
rect 114737 5611 114803 5614
rect 119613 5674 119679 5677
rect 127985 5674 128051 5677
rect 119613 5672 128051 5674
rect 119613 5616 119618 5672
rect 119674 5616 127990 5672
rect 128046 5616 128051 5672
rect 119613 5614 128051 5616
rect 119613 5611 119679 5614
rect 127985 5611 128051 5614
rect 128169 5674 128235 5677
rect 132585 5674 132651 5677
rect 135348 5674 135408 5716
rect 128169 5672 132651 5674
rect 128169 5616 128174 5672
rect 128230 5616 132590 5672
rect 132646 5616 132651 5672
rect 128169 5614 132651 5616
rect 128169 5611 128235 5614
rect 132585 5611 132651 5614
rect 132726 5614 135408 5674
rect 135805 5674 135871 5677
rect 156965 5674 157031 5677
rect 165266 5674 165272 5738
rect 165336 5674 165342 5738
rect 135805 5672 157031 5674
rect 135805 5616 135810 5672
rect 135866 5616 156970 5672
rect 157026 5616 157031 5672
rect 135805 5614 157031 5616
rect -400 5538 800 5568
rect 2957 5538 3023 5541
rect -400 5536 3023 5538
rect -400 5480 2962 5536
rect 3018 5480 3023 5536
rect -400 5478 3023 5480
rect -400 5448 800 5478
rect 2957 5475 3023 5478
rect 91921 5538 91987 5541
rect 121729 5538 121795 5541
rect 91921 5536 121795 5538
rect 91921 5480 91926 5536
rect 91982 5480 121734 5536
rect 121790 5480 121795 5536
rect 91921 5478 121795 5480
rect 91921 5475 91987 5478
rect 121729 5475 121795 5478
rect 127525 5538 127591 5541
rect 130009 5538 130075 5541
rect 132726 5538 132786 5614
rect 135805 5611 135871 5614
rect 156965 5611 157031 5614
rect 127525 5536 130075 5538
rect 127525 5480 127530 5536
rect 127586 5480 130014 5536
rect 130070 5480 130075 5536
rect 127525 5478 130075 5480
rect 127525 5475 127591 5478
rect 130009 5475 130075 5478
rect 130150 5478 132786 5538
rect 133045 5538 133111 5541
rect 136909 5538 136975 5541
rect 133045 5536 136975 5538
rect 133045 5480 133050 5536
rect 133106 5480 136914 5536
rect 136970 5480 136975 5536
rect 133045 5478 136975 5480
rect 4071 5472 4137 5473
rect 44071 5472 44137 5473
rect 84071 5472 84137 5473
rect 124071 5472 124137 5473
rect 4066 5408 4072 5472
rect 4136 5408 4142 5472
rect 44066 5408 44072 5472
rect 44136 5408 44142 5472
rect 84066 5408 84072 5472
rect 84136 5408 84142 5472
rect 124066 5408 124072 5472
rect 124136 5408 124142 5472
rect 4071 5407 4137 5408
rect 44071 5407 44137 5408
rect 84071 5407 84137 5408
rect 124071 5407 124137 5408
rect 101213 5402 101279 5405
rect 105169 5402 105235 5405
rect 101213 5400 105235 5402
rect 101213 5344 101218 5400
rect 101274 5344 105174 5400
rect 105230 5344 105235 5400
rect 101213 5342 105235 5344
rect 101213 5339 101279 5342
rect 105169 5339 105235 5342
rect 106641 5402 106707 5405
rect 116945 5402 117011 5405
rect 106641 5400 117011 5402
rect 106641 5344 106646 5400
rect 106702 5344 116950 5400
rect 117006 5344 117011 5400
rect 106641 5342 117011 5344
rect 106641 5339 106707 5342
rect 116945 5339 117011 5342
rect 118509 5402 118575 5405
rect 120441 5402 120507 5405
rect 118509 5400 120507 5402
rect 118509 5344 118514 5400
rect 118570 5344 120446 5400
rect 120502 5344 120507 5400
rect 118509 5342 120507 5344
rect 118509 5339 118575 5342
rect 120441 5339 120507 5342
rect 121269 5402 121335 5405
rect 123569 5402 123635 5405
rect 121269 5400 123635 5402
rect 121269 5344 121274 5400
rect 121330 5344 123574 5400
rect 123630 5344 123635 5400
rect 121269 5342 123635 5344
rect 121269 5339 121335 5342
rect 123569 5339 123635 5342
rect 124254 5340 124260 5404
rect 124324 5402 124330 5404
rect 128169 5402 128235 5405
rect 129733 5402 129799 5405
rect 124324 5342 127082 5402
rect 124324 5340 124330 5342
rect 89989 5266 90055 5269
rect 122925 5266 122991 5269
rect 89989 5264 122991 5266
rect 89989 5208 89994 5264
rect 90050 5208 122930 5264
rect 122986 5208 122991 5264
rect 89989 5206 122991 5208
rect 89989 5203 90055 5206
rect 122925 5203 122991 5206
rect 125685 5266 125751 5269
rect 126789 5266 126855 5269
rect 125685 5264 126855 5266
rect 125685 5208 125690 5264
rect 125746 5208 126794 5264
rect 126850 5208 126855 5264
rect 125685 5206 126855 5208
rect 127022 5266 127082 5342
rect 128169 5400 129799 5402
rect 128169 5344 128174 5400
rect 128230 5344 129738 5400
rect 129794 5344 129799 5400
rect 128169 5342 129799 5344
rect 128169 5339 128235 5342
rect 129733 5339 129799 5342
rect 130150 5266 130210 5478
rect 133045 5475 133111 5478
rect 136909 5475 136975 5478
rect 137645 5538 137711 5541
rect 137921 5538 137987 5541
rect 144453 5538 144519 5541
rect 137645 5536 137987 5538
rect 137645 5480 137650 5536
rect 137706 5480 137926 5536
rect 137982 5480 137987 5536
rect 137645 5478 137987 5480
rect 137645 5475 137711 5478
rect 137921 5475 137987 5478
rect 138062 5536 144519 5538
rect 138062 5480 144458 5536
rect 144514 5480 144519 5536
rect 138062 5478 144519 5480
rect 132401 5402 132467 5405
rect 138062 5402 138122 5478
rect 144453 5475 144519 5478
rect 144637 5538 144703 5541
rect 157241 5538 157307 5541
rect 144637 5536 157307 5538
rect 144637 5480 144642 5536
rect 144698 5480 157246 5536
rect 157302 5480 157307 5536
rect 144637 5478 157307 5480
rect 144637 5475 144703 5478
rect 157241 5475 157307 5478
rect 132401 5400 134442 5402
rect 132401 5344 132406 5400
rect 132462 5344 134442 5400
rect 132401 5342 134442 5344
rect 132401 5339 132467 5342
rect 127022 5206 130210 5266
rect 131297 5266 131363 5269
rect 133965 5266 134031 5269
rect 131297 5264 134031 5266
rect 131297 5208 131302 5264
rect 131358 5208 133970 5264
rect 134026 5208 134031 5264
rect 131297 5206 134031 5208
rect 134382 5266 134442 5342
rect 134750 5342 138122 5402
rect 138289 5402 138355 5405
rect 157006 5402 157012 5404
rect 138289 5400 157012 5402
rect 138289 5344 138294 5400
rect 138350 5344 157012 5400
rect 138289 5342 157012 5344
rect 134750 5266 134810 5342
rect 138289 5339 138355 5342
rect 157006 5340 157012 5342
rect 157076 5340 157082 5404
rect 185666 5345 185672 5409
rect 185736 5345 185742 5409
rect 134382 5206 134810 5266
rect 135161 5266 135227 5269
rect 156137 5266 156203 5269
rect 135161 5264 156203 5266
rect 135161 5208 135166 5264
rect 135222 5208 156142 5264
rect 156198 5208 156203 5264
rect 164466 5223 164472 5287
rect 164536 5223 164542 5287
rect 135161 5206 156203 5208
rect 125685 5203 125751 5206
rect 126789 5203 126855 5206
rect 131297 5203 131363 5206
rect 133965 5203 134031 5206
rect 135161 5203 135227 5206
rect 156137 5203 156203 5206
rect 105077 5130 105143 5133
rect 107009 5130 107075 5133
rect 105077 5128 107075 5130
rect 105077 5072 105082 5128
rect 105138 5072 107014 5128
rect 107070 5072 107075 5128
rect 105077 5070 107075 5072
rect 105077 5067 105143 5070
rect 107009 5067 107075 5070
rect 108113 5130 108179 5133
rect 138565 5130 138631 5133
rect 108113 5128 138631 5130
rect 108113 5072 108118 5128
rect 108174 5072 138570 5128
rect 138626 5072 138631 5128
rect 108113 5070 138631 5072
rect 108113 5067 108179 5070
rect 138565 5067 138631 5070
rect 140681 5130 140747 5133
rect 144453 5130 144519 5133
rect 157057 5130 157123 5133
rect 140681 5128 144378 5130
rect 140681 5072 140686 5128
rect 140742 5072 144378 5128
rect 140681 5070 144378 5072
rect 140681 5067 140747 5070
rect 106365 4994 106431 4997
rect 106641 4994 106707 4997
rect 106365 4992 106707 4994
rect 106365 4936 106370 4992
rect 106426 4936 106646 4992
rect 106702 4936 106707 4992
rect 106365 4934 106707 4936
rect 106365 4931 106431 4934
rect 106641 4931 106707 4934
rect 106917 4994 106983 4997
rect 108389 4994 108455 4997
rect 106917 4992 108455 4994
rect 106917 4936 106922 4992
rect 106978 4936 108394 4992
rect 108450 4936 108455 4992
rect 106917 4934 108455 4936
rect 106917 4931 106983 4934
rect 108389 4931 108455 4934
rect 110413 4994 110479 4997
rect 140405 4994 140471 4997
rect 110413 4992 140471 4994
rect 110413 4936 110418 4992
rect 110474 4936 140410 4992
rect 140466 4936 140471 4992
rect 110413 4934 140471 4936
rect 144318 4994 144378 5070
rect 144453 5128 157123 5130
rect 144453 5072 144458 5128
rect 144514 5072 157062 5128
rect 157118 5072 157123 5128
rect 144453 5070 157123 5072
rect 144453 5067 144519 5070
rect 157057 5067 157123 5070
rect 157006 4994 157012 4996
rect 144318 4934 157012 4994
rect 110413 4931 110479 4934
rect 140405 4931 140471 4934
rect 157006 4932 157012 4934
rect 157076 4932 157082 4996
rect 185266 4945 185272 5009
rect 185336 4945 185342 5009
rect 24071 4928 24137 4929
rect 64071 4928 64137 4929
rect 104071 4928 104137 4929
rect 144071 4928 144137 4929
rect 24066 4864 24072 4928
rect 24136 4864 24142 4928
rect 64066 4864 64072 4928
rect 64136 4864 64142 4928
rect 104066 4864 104072 4928
rect 104136 4864 104142 4928
rect 144066 4864 144072 4928
rect 144136 4864 144142 4928
rect 24071 4863 24137 4864
rect 64071 4863 64137 4864
rect 104071 4863 104137 4864
rect 144071 4863 144137 4864
rect 106273 4858 106339 4861
rect 106641 4858 106707 4861
rect 106273 4856 106707 4858
rect 106273 4800 106278 4856
rect 106334 4800 106646 4856
rect 106702 4800 106707 4856
rect 106273 4798 106707 4800
rect 106273 4795 106339 4798
rect 106641 4795 106707 4798
rect 107561 4858 107627 4861
rect 110505 4858 110571 4861
rect 107561 4856 110571 4858
rect 107561 4800 107566 4856
rect 107622 4800 110510 4856
rect 110566 4800 110571 4856
rect 107561 4798 110571 4800
rect 107561 4795 107627 4798
rect 110505 4795 110571 4798
rect 110873 4858 110939 4861
rect 117589 4858 117655 4861
rect 110873 4856 117655 4858
rect 110873 4800 110878 4856
rect 110934 4800 117594 4856
rect 117650 4800 117655 4856
rect 110873 4798 117655 4800
rect 110873 4795 110939 4798
rect 117589 4795 117655 4798
rect 119337 4858 119403 4861
rect 127341 4858 127407 4861
rect 119337 4856 127407 4858
rect 119337 4800 119342 4856
rect 119398 4800 127346 4856
rect 127402 4800 127407 4856
rect 119337 4798 127407 4800
rect 119337 4795 119403 4798
rect 127341 4795 127407 4798
rect 128537 4858 128603 4861
rect 132677 4858 132743 4861
rect 128537 4856 132743 4858
rect 128537 4800 128542 4856
rect 128598 4800 132682 4856
rect 132738 4800 132743 4856
rect 128537 4798 132743 4800
rect 128537 4795 128603 4798
rect 132677 4795 132743 4798
rect 132953 4858 133019 4861
rect 140957 4858 141023 4861
rect 132953 4856 141023 4858
rect 132953 4800 132958 4856
rect 133014 4800 140962 4856
rect 141018 4800 141023 4856
rect 132953 4798 141023 4800
rect 132953 4795 133019 4798
rect 140957 4795 141023 4798
rect 102869 4722 102935 4725
rect 107929 4722 107995 4725
rect 102869 4720 107995 4722
rect 102869 4664 102874 4720
rect 102930 4664 107934 4720
rect 107990 4664 107995 4720
rect 102869 4662 107995 4664
rect 102869 4659 102935 4662
rect 107929 4659 107995 4662
rect 111609 4722 111675 4725
rect 136909 4722 136975 4725
rect 156965 4722 157031 4725
rect 111609 4720 136834 4722
rect 111609 4664 111614 4720
rect 111670 4664 136834 4720
rect 111609 4662 136834 4664
rect 111609 4659 111675 4662
rect 70301 4586 70367 4589
rect 117405 4586 117471 4589
rect 70301 4584 117471 4586
rect 70301 4528 70306 4584
rect 70362 4528 117410 4584
rect 117466 4528 117471 4584
rect 70301 4526 117471 4528
rect 70301 4523 70367 4526
rect 117405 4523 117471 4526
rect 119613 4586 119679 4589
rect 123753 4586 123819 4589
rect 119613 4584 123819 4586
rect 119613 4528 119618 4584
rect 119674 4528 123758 4584
rect 123814 4528 123819 4584
rect 119613 4526 123819 4528
rect 119613 4523 119679 4526
rect 123753 4523 123819 4526
rect 124121 4586 124187 4589
rect 136633 4586 136699 4589
rect 124121 4584 136699 4586
rect 124121 4528 124126 4584
rect 124182 4528 136638 4584
rect 136694 4528 136699 4584
rect 124121 4526 136699 4528
rect 124121 4523 124187 4526
rect 136633 4523 136699 4526
rect 106549 4450 106615 4453
rect 110413 4450 110479 4453
rect 106549 4448 110479 4450
rect 106549 4392 106554 4448
rect 106610 4392 110418 4448
rect 110474 4392 110479 4448
rect 106549 4390 110479 4392
rect 106549 4387 106615 4390
rect 110413 4387 110479 4390
rect 111241 4450 111307 4453
rect 113633 4450 113699 4453
rect 111241 4448 113699 4450
rect 111241 4392 111246 4448
rect 111302 4392 113638 4448
rect 113694 4392 113699 4448
rect 111241 4390 113699 4392
rect 111241 4387 111307 4390
rect 113633 4387 113699 4390
rect 116945 4450 117011 4453
rect 118969 4450 119035 4453
rect 116945 4448 119035 4450
rect 116945 4392 116950 4448
rect 117006 4392 118974 4448
rect 119030 4392 119035 4448
rect 116945 4390 119035 4392
rect 116945 4387 117011 4390
rect 118969 4387 119035 4390
rect 124213 4450 124279 4453
rect 133321 4450 133387 4453
rect 135345 4450 135411 4453
rect 124213 4448 133154 4450
rect 124213 4392 124218 4448
rect 124274 4392 133154 4448
rect 124213 4390 133154 4392
rect 124213 4387 124279 4390
rect 4071 4384 4137 4385
rect 44071 4384 44137 4385
rect 84071 4384 84137 4385
rect 124071 4384 124137 4385
rect 4066 4320 4072 4384
rect 4136 4320 4142 4384
rect 44066 4320 44072 4384
rect 44136 4320 44142 4384
rect 84066 4320 84072 4384
rect 84136 4320 84142 4384
rect 124066 4320 124072 4384
rect 124136 4320 124142 4384
rect 4071 4319 4137 4320
rect 44071 4319 44137 4320
rect 84071 4319 84137 4320
rect 124071 4319 124137 4320
rect 105353 4314 105419 4317
rect 105905 4314 105971 4317
rect 105353 4312 105971 4314
rect 105353 4256 105358 4312
rect 105414 4256 105910 4312
rect 105966 4256 105971 4312
rect 105353 4254 105971 4256
rect 105353 4251 105419 4254
rect 105905 4251 105971 4254
rect 121177 4314 121243 4317
rect 123937 4314 124003 4317
rect 121177 4312 124003 4314
rect 121177 4256 121182 4312
rect 121238 4256 123942 4312
rect 123998 4256 124003 4312
rect 121177 4254 124003 4256
rect 121177 4251 121243 4254
rect 123937 4251 124003 4254
rect 124213 4314 124279 4317
rect 132953 4314 133019 4317
rect 124213 4312 133019 4314
rect 124213 4256 124218 4312
rect 124274 4256 132958 4312
rect 133014 4256 133019 4312
rect 124213 4254 133019 4256
rect 133094 4314 133154 4390
rect 133321 4448 135411 4450
rect 133321 4392 133326 4448
rect 133382 4392 135350 4448
rect 135406 4392 135411 4448
rect 133321 4390 135411 4392
rect 136774 4450 136834 4662
rect 136909 4720 157031 4722
rect 136909 4664 136914 4720
rect 136970 4664 156970 4720
rect 157026 4664 157031 4720
rect 136909 4662 157031 4664
rect 136909 4659 136975 4662
rect 156965 4659 157031 4662
rect 165666 4617 165672 4681
rect 165736 4617 165742 4681
rect 137185 4586 137251 4589
rect 137645 4586 137711 4589
rect 137185 4584 137711 4586
rect 137185 4528 137190 4584
rect 137246 4528 137650 4584
rect 137706 4528 137711 4584
rect 137185 4526 137711 4528
rect 137185 4523 137251 4526
rect 137645 4523 137711 4526
rect 138013 4586 138079 4589
rect 139761 4586 139827 4589
rect 138013 4584 139827 4586
rect 138013 4528 138018 4584
rect 138074 4528 139766 4584
rect 139822 4528 139827 4584
rect 138013 4526 139827 4528
rect 138013 4523 138079 4526
rect 139761 4523 139827 4526
rect 141509 4586 141575 4589
rect 157190 4586 157196 4588
rect 141509 4584 157196 4586
rect 141509 4528 141514 4584
rect 141570 4528 157196 4584
rect 141509 4526 157196 4528
rect 141509 4523 141575 4526
rect 157190 4524 157196 4526
rect 157260 4524 157266 4588
rect 184466 4494 184472 4558
rect 184536 4494 184542 4558
rect 142429 4450 142495 4453
rect 136774 4448 142495 4450
rect 136774 4392 142434 4448
rect 142490 4392 142495 4448
rect 136774 4390 142495 4392
rect 133321 4387 133387 4390
rect 135345 4387 135411 4390
rect 142429 4387 142495 4390
rect 141509 4314 141575 4317
rect 133094 4312 141575 4314
rect 133094 4256 141514 4312
rect 141570 4256 141575 4312
rect 133094 4254 141575 4256
rect 124213 4251 124279 4254
rect 132953 4251 133019 4254
rect 141509 4251 141575 4254
rect 145046 4252 145052 4316
rect 145116 4314 145122 4316
rect 145281 4314 145347 4317
rect 145116 4312 145347 4314
rect 145116 4256 145286 4312
rect 145342 4256 145347 4312
rect 145116 4254 145347 4256
rect 145116 4252 145122 4254
rect 145281 4251 145347 4254
rect 165266 4217 165272 4281
rect 165336 4217 165342 4281
rect 105445 4178 105511 4181
rect 109677 4178 109743 4181
rect 105445 4176 109743 4178
rect 105445 4120 105450 4176
rect 105506 4120 109682 4176
rect 109738 4120 109743 4176
rect 105445 4118 109743 4120
rect 105445 4115 105511 4118
rect 109677 4115 109743 4118
rect 111057 4178 111123 4181
rect 140773 4178 140839 4181
rect 111057 4176 140839 4178
rect 111057 4120 111062 4176
rect 111118 4120 140778 4176
rect 140834 4120 140839 4176
rect 111057 4118 140839 4120
rect 111057 4115 111123 4118
rect 140773 4115 140839 4118
rect 141325 4178 141391 4181
rect 156229 4178 156295 4181
rect 141325 4176 156295 4178
rect 141325 4120 141330 4176
rect 141386 4120 156234 4176
rect 156290 4120 156295 4176
rect 141325 4118 156295 4120
rect 141325 4115 141391 4118
rect 156229 4115 156295 4118
rect 60641 4042 60707 4045
rect 109585 4042 109651 4045
rect 60641 4040 109651 4042
rect 60641 3984 60646 4040
rect 60702 3984 109590 4040
rect 109646 3984 109651 4040
rect 60641 3982 109651 3984
rect 60641 3979 60707 3982
rect 109585 3979 109651 3982
rect 110321 4042 110387 4045
rect 113449 4042 113515 4045
rect 110321 4040 113515 4042
rect 110321 3984 110326 4040
rect 110382 3984 113454 4040
rect 113510 3984 113515 4040
rect 110321 3982 113515 3984
rect 110321 3979 110387 3982
rect 113449 3979 113515 3982
rect 118509 4042 118575 4045
rect 119981 4042 120047 4045
rect 118509 4040 120047 4042
rect 118509 3984 118514 4040
rect 118570 3984 119986 4040
rect 120042 3984 120047 4040
rect 118509 3982 120047 3984
rect 118509 3979 118575 3982
rect 119981 3979 120047 3982
rect 126237 4042 126303 4045
rect 128721 4042 128787 4045
rect 126237 4040 128787 4042
rect 126237 3984 126242 4040
rect 126298 3984 128726 4040
rect 128782 3984 128787 4040
rect 126237 3982 128787 3984
rect 126237 3979 126303 3982
rect 128721 3979 128787 3982
rect 131021 4042 131087 4045
rect 136633 4042 136699 4045
rect 156597 4042 156663 4045
rect 131021 4040 136699 4042
rect 131021 3984 131026 4040
rect 131082 3984 136638 4040
rect 136694 3984 136699 4040
rect 131021 3982 136699 3984
rect 131021 3979 131087 3982
rect 136633 3979 136699 3982
rect 136774 4040 156663 4042
rect 136774 3984 156602 4040
rect 156658 3984 156663 4040
rect 136774 3982 156663 3984
rect 107653 3906 107719 3909
rect 111057 3906 111123 3909
rect 107653 3904 111123 3906
rect 107653 3848 107658 3904
rect 107714 3848 111062 3904
rect 111118 3848 111123 3904
rect 107653 3846 111123 3848
rect 107653 3843 107719 3846
rect 111057 3843 111123 3846
rect 111701 3906 111767 3909
rect 115381 3906 115447 3909
rect 111701 3904 115447 3906
rect 111701 3848 111706 3904
rect 111762 3848 115386 3904
rect 115442 3848 115447 3904
rect 111701 3846 115447 3848
rect 111701 3843 111767 3846
rect 115381 3843 115447 3846
rect 116853 3906 116919 3909
rect 119613 3906 119679 3909
rect 126053 3906 126119 3909
rect 116853 3904 119538 3906
rect 116853 3848 116858 3904
rect 116914 3848 119538 3904
rect 116853 3846 119538 3848
rect 116853 3843 116919 3846
rect 24071 3840 24137 3841
rect 64071 3840 64137 3841
rect 104071 3840 104137 3841
rect 24066 3776 24072 3840
rect 24136 3776 24142 3840
rect 64066 3776 64072 3840
rect 64136 3776 64142 3840
rect 104066 3776 104072 3840
rect 104136 3776 104142 3840
rect 24071 3775 24137 3776
rect 64071 3775 64137 3776
rect 104071 3775 104137 3776
rect 109585 3770 109651 3773
rect 113725 3770 113791 3773
rect 109585 3768 113791 3770
rect 109585 3712 109590 3768
rect 109646 3712 113730 3768
rect 113786 3712 113791 3768
rect 109585 3710 113791 3712
rect 109585 3707 109651 3710
rect 113725 3707 113791 3710
rect 118509 3770 118575 3773
rect 119245 3770 119311 3773
rect 118509 3768 119311 3770
rect 118509 3712 118514 3768
rect 118570 3712 119250 3768
rect 119306 3712 119311 3768
rect 118509 3710 119311 3712
rect 119478 3770 119538 3846
rect 119613 3904 126119 3906
rect 119613 3848 119618 3904
rect 119674 3848 126058 3904
rect 126114 3848 126119 3904
rect 119613 3846 126119 3848
rect 119613 3843 119679 3846
rect 126053 3843 126119 3846
rect 126789 3906 126855 3909
rect 133321 3906 133387 3909
rect 126789 3904 133387 3906
rect 126789 3848 126794 3904
rect 126850 3848 133326 3904
rect 133382 3848 133387 3904
rect 126789 3846 133387 3848
rect 126789 3843 126855 3846
rect 133321 3843 133387 3846
rect 133597 3906 133663 3909
rect 134793 3906 134859 3909
rect 133597 3904 134859 3906
rect 133597 3848 133602 3904
rect 133658 3848 134798 3904
rect 134854 3848 134859 3904
rect 133597 3846 134859 3848
rect 133597 3843 133663 3846
rect 134793 3843 134859 3846
rect 123937 3770 124003 3773
rect 119478 3768 124003 3770
rect 119478 3712 123942 3768
rect 123998 3712 124003 3768
rect 119478 3710 124003 3712
rect 118509 3707 118575 3710
rect 119245 3707 119311 3710
rect 123937 3707 124003 3710
rect 125961 3770 126027 3773
rect 128629 3770 128695 3773
rect 125961 3768 128695 3770
rect 125961 3712 125966 3768
rect 126022 3712 128634 3768
rect 128690 3712 128695 3768
rect 125961 3710 128695 3712
rect 125961 3707 126027 3710
rect 128629 3707 128695 3710
rect 131849 3770 131915 3773
rect 136774 3770 136834 3982
rect 156597 3979 156663 3982
rect 156781 4042 156847 4045
rect 156781 4040 156890 4042
rect 156781 3984 156786 4040
rect 156842 3984 156890 4040
rect 156781 3979 156890 3984
rect 136909 3906 136975 3909
rect 143901 3906 143967 3909
rect 151261 3906 151327 3909
rect 136909 3904 143967 3906
rect 136909 3848 136914 3904
rect 136970 3848 143906 3904
rect 143962 3848 143967 3904
rect 136909 3846 143967 3848
rect 136909 3843 136975 3846
rect 143901 3843 143967 3846
rect 144318 3904 151327 3906
rect 144318 3848 151266 3904
rect 151322 3848 151327 3904
rect 156830 3876 156890 3979
rect 144318 3846 151327 3848
rect 144071 3840 144137 3841
rect 144066 3776 144072 3840
rect 144136 3776 144142 3840
rect 144071 3775 144137 3776
rect 131849 3768 136834 3770
rect 131849 3712 131854 3768
rect 131910 3712 136834 3768
rect 131849 3710 136834 3712
rect 137001 3770 137067 3773
rect 138105 3770 138171 3773
rect 137001 3768 138171 3770
rect 137001 3712 137006 3768
rect 137062 3712 138110 3768
rect 138166 3712 138171 3768
rect 137001 3710 138171 3712
rect 131849 3707 131915 3710
rect 137001 3707 137067 3710
rect 138105 3707 138171 3710
rect 138473 3770 138539 3773
rect 142245 3770 142311 3773
rect 138473 3768 142311 3770
rect 138473 3712 138478 3768
rect 138534 3712 142250 3768
rect 142306 3712 142311 3768
rect 138473 3710 142311 3712
rect 138473 3707 138539 3710
rect 142245 3707 142311 3710
rect 79041 3634 79107 3637
rect 119061 3634 119127 3637
rect 79041 3632 119127 3634
rect 79041 3576 79046 3632
rect 79102 3576 119066 3632
rect 119122 3576 119127 3632
rect 79041 3574 119127 3576
rect 79041 3571 79107 3574
rect 119061 3571 119127 3574
rect 120165 3634 120231 3637
rect 125501 3634 125567 3637
rect 120165 3632 125567 3634
rect 120165 3576 120170 3632
rect 120226 3576 125506 3632
rect 125562 3576 125567 3632
rect 120165 3574 125567 3576
rect 120165 3571 120231 3574
rect 125501 3571 125567 3574
rect 125961 3634 126027 3637
rect 133321 3634 133387 3637
rect 144318 3634 144378 3846
rect 151261 3843 151327 3846
rect 144545 3770 144611 3773
rect 153929 3770 153995 3773
rect 144545 3768 153995 3770
rect 144545 3712 144550 3768
rect 144606 3712 153934 3768
rect 153990 3712 153995 3768
rect 164466 3766 164472 3830
rect 164536 3766 164542 3830
rect 144545 3710 153995 3712
rect 144545 3707 144611 3710
rect 153929 3707 153995 3710
rect 125961 3632 132970 3634
rect 125961 3576 125966 3632
rect 126022 3576 132970 3632
rect 125961 3574 132970 3576
rect 125961 3571 126027 3574
rect 97625 3498 97691 3501
rect 105813 3498 105879 3501
rect 97625 3496 105879 3498
rect 97625 3440 97630 3496
rect 97686 3440 105818 3496
rect 105874 3440 105879 3496
rect 97625 3438 105879 3440
rect 97625 3435 97691 3438
rect 105813 3435 105879 3438
rect 106641 3498 106707 3501
rect 114185 3498 114251 3501
rect 106641 3496 114251 3498
rect 106641 3440 106646 3496
rect 106702 3440 114190 3496
rect 114246 3440 114251 3496
rect 106641 3438 114251 3440
rect 106641 3435 106707 3438
rect 114185 3435 114251 3438
rect 115933 3498 115999 3501
rect 128261 3498 128327 3501
rect 128445 3498 128511 3501
rect 115933 3496 128186 3498
rect 115933 3440 115938 3496
rect 115994 3440 128186 3496
rect 115933 3438 128186 3440
rect 115933 3435 115999 3438
rect 89621 3362 89687 3365
rect 112437 3362 112503 3365
rect 89621 3360 112503 3362
rect 89621 3304 89626 3360
rect 89682 3304 112442 3360
rect 112498 3304 112503 3360
rect 89621 3302 112503 3304
rect 89621 3299 89687 3302
rect 112437 3299 112503 3302
rect 116485 3362 116551 3365
rect 117313 3362 117379 3365
rect 116485 3360 117379 3362
rect 116485 3304 116490 3360
rect 116546 3304 117318 3360
rect 117374 3304 117379 3360
rect 116485 3302 117379 3304
rect 116485 3299 116551 3302
rect 117313 3299 117379 3302
rect 117497 3362 117563 3365
rect 118693 3362 118759 3365
rect 117497 3360 118759 3362
rect 117497 3304 117502 3360
rect 117558 3304 118698 3360
rect 118754 3304 118759 3360
rect 117497 3302 118759 3304
rect 128126 3362 128186 3438
rect 128261 3496 128511 3498
rect 128261 3440 128266 3496
rect 128322 3440 128450 3496
rect 128506 3440 128511 3496
rect 128261 3438 128511 3440
rect 128261 3435 128327 3438
rect 128445 3435 128511 3438
rect 129917 3498 129983 3501
rect 132493 3498 132559 3501
rect 129917 3496 132559 3498
rect 129917 3440 129922 3496
rect 129978 3440 132498 3496
rect 132554 3440 132559 3496
rect 129917 3438 132559 3440
rect 132910 3498 132970 3574
rect 133321 3632 144378 3634
rect 133321 3576 133326 3632
rect 133382 3576 144378 3632
rect 133321 3574 144378 3576
rect 144453 3634 144519 3637
rect 153101 3634 153167 3637
rect 144453 3632 153167 3634
rect 144453 3576 144458 3632
rect 144514 3576 153106 3632
rect 153162 3576 153167 3632
rect 144453 3574 153167 3576
rect 133321 3571 133387 3574
rect 144453 3571 144519 3574
rect 153101 3571 153167 3574
rect 153285 3634 153351 3637
rect 153285 3632 157258 3634
rect 153285 3576 153290 3632
rect 153346 3576 157258 3632
rect 153285 3574 157258 3576
rect 153285 3571 153351 3574
rect 151629 3498 151695 3501
rect 132910 3496 151695 3498
rect 132910 3440 151634 3496
rect 151690 3440 151695 3496
rect 132910 3438 151695 3440
rect 129917 3435 129983 3438
rect 132493 3435 132559 3438
rect 151629 3435 151695 3438
rect 152365 3498 152431 3501
rect 153561 3498 153627 3501
rect 152365 3496 153627 3498
rect 152365 3440 152370 3496
rect 152426 3440 153566 3496
rect 153622 3440 153627 3496
rect 152365 3438 153627 3440
rect 157198 3498 157258 3574
rect 157374 3572 157380 3636
rect 157444 3634 157450 3636
rect 172462 3634 172468 3636
rect 157444 3574 172468 3634
rect 157444 3572 157450 3574
rect 172462 3572 172468 3574
rect 172532 3572 172538 3636
rect 161606 3498 161612 3500
rect 157198 3438 161612 3498
rect 152365 3435 152431 3438
rect 153561 3435 153627 3438
rect 161606 3436 161612 3438
rect 161676 3436 161682 3500
rect 161790 3436 161796 3500
rect 161860 3498 161866 3500
rect 167310 3498 167316 3500
rect 161860 3438 167316 3498
rect 161860 3436 161866 3438
rect 167310 3436 167316 3438
rect 167380 3436 167386 3500
rect 167494 3436 167500 3500
rect 167564 3498 167570 3500
rect 176326 3498 176332 3500
rect 167564 3438 176332 3498
rect 167564 3436 167570 3438
rect 176326 3436 176332 3438
rect 176396 3436 176402 3500
rect 129273 3362 129339 3365
rect 128126 3360 129339 3362
rect 128126 3304 129278 3360
rect 129334 3304 129339 3360
rect 128126 3302 129339 3304
rect 117497 3299 117563 3302
rect 118693 3299 118759 3302
rect 129273 3299 129339 3302
rect 129733 3362 129799 3365
rect 136909 3362 136975 3365
rect 129733 3360 136975 3362
rect 129733 3304 129738 3360
rect 129794 3304 136914 3360
rect 136970 3304 136975 3360
rect 129733 3302 136975 3304
rect 129733 3299 129799 3302
rect 136909 3299 136975 3302
rect 137185 3362 137251 3365
rect 137318 3362 137324 3364
rect 137185 3360 137324 3362
rect 137185 3304 137190 3360
rect 137246 3304 137324 3360
rect 137185 3302 137324 3304
rect 137185 3299 137251 3302
rect 137318 3300 137324 3302
rect 137388 3300 137394 3364
rect 137461 3362 137527 3365
rect 142981 3362 143047 3365
rect 144545 3362 144611 3365
rect 137461 3360 142906 3362
rect 137461 3304 137466 3360
rect 137522 3304 142906 3360
rect 137461 3302 142906 3304
rect 137461 3299 137527 3302
rect 4071 3296 4137 3297
rect 44071 3296 44137 3297
rect 84071 3296 84137 3297
rect 124071 3296 124137 3297
rect 4066 3232 4072 3296
rect 4136 3232 4142 3296
rect 44066 3232 44072 3296
rect 44136 3232 44142 3296
rect 84066 3232 84072 3296
rect 84136 3232 84142 3296
rect 124066 3232 124072 3296
rect 124136 3232 124142 3296
rect 4071 3231 4137 3232
rect 44071 3231 44137 3232
rect 84071 3231 84137 3232
rect 124071 3231 124137 3232
rect 109217 3226 109283 3229
rect 112069 3226 112135 3229
rect 109217 3224 112135 3226
rect 109217 3168 109222 3224
rect 109278 3168 112074 3224
rect 112130 3168 112135 3224
rect 109217 3166 112135 3168
rect 109217 3163 109283 3166
rect 112069 3163 112135 3166
rect 115841 3226 115907 3229
rect 118325 3226 118391 3229
rect 115841 3224 118391 3226
rect 115841 3168 115846 3224
rect 115902 3168 118330 3224
rect 118386 3168 118391 3224
rect 115841 3166 118391 3168
rect 115841 3163 115907 3166
rect 118325 3163 118391 3166
rect 119797 3226 119863 3229
rect 123569 3226 123635 3229
rect 119797 3224 123635 3226
rect 119797 3168 119802 3224
rect 119858 3168 123574 3224
rect 123630 3168 123635 3224
rect 119797 3166 123635 3168
rect 119797 3163 119863 3166
rect 123569 3163 123635 3166
rect 128721 3226 128787 3229
rect 142705 3226 142771 3229
rect 128721 3224 142771 3226
rect 128721 3168 128726 3224
rect 128782 3168 142710 3224
rect 142766 3168 142771 3224
rect 128721 3166 142771 3168
rect 142846 3226 142906 3302
rect 142981 3360 144611 3362
rect 142981 3304 142986 3360
rect 143042 3304 144550 3360
rect 144606 3304 144611 3360
rect 142981 3302 144611 3304
rect 142981 3299 143047 3302
rect 144545 3299 144611 3302
rect 144729 3362 144795 3365
rect 163078 3362 163084 3364
rect 144729 3360 163084 3362
rect 144729 3304 144734 3360
rect 144790 3304 163084 3360
rect 144729 3302 163084 3304
rect 144729 3299 144795 3302
rect 163078 3300 163084 3302
rect 163148 3300 163154 3364
rect 169480 3302 180442 3362
rect 153285 3226 153351 3229
rect 142846 3224 153351 3226
rect 142846 3168 153290 3224
rect 153346 3168 153351 3224
rect 142846 3166 153351 3168
rect 128721 3163 128787 3166
rect 142705 3163 142771 3166
rect 153285 3163 153351 3166
rect 153561 3226 153627 3229
rect 157006 3226 157012 3228
rect 153561 3224 157012 3226
rect 153561 3168 153566 3224
rect 153622 3168 157012 3224
rect 153561 3166 157012 3168
rect 153561 3163 153627 3166
rect 157006 3164 157012 3166
rect 157076 3164 157082 3228
rect 162894 3226 162900 3228
rect 157244 3166 162900 3226
rect 113817 3090 113883 3093
rect 133505 3090 133571 3093
rect 113817 3088 133571 3090
rect 113817 3032 113822 3088
rect 113878 3032 133510 3088
rect 133566 3032 133571 3088
rect 113817 3030 133571 3032
rect 113817 3027 113883 3030
rect 133505 3027 133571 3030
rect 133689 3090 133755 3093
rect 137461 3090 137527 3093
rect 133689 3088 137527 3090
rect 133689 3032 133694 3088
rect 133750 3032 137466 3088
rect 137522 3032 137527 3088
rect 133689 3030 137527 3032
rect 133689 3027 133755 3030
rect 137461 3027 137527 3030
rect 137686 3028 137692 3092
rect 137756 3090 137762 3092
rect 141785 3090 141851 3093
rect 151854 3090 151860 3092
rect 137756 3088 141851 3090
rect 137756 3032 141790 3088
rect 141846 3032 141851 3088
rect 137756 3030 141851 3032
rect 137756 3028 137762 3030
rect 141785 3027 141851 3030
rect 142846 3030 151860 3090
rect 81249 2954 81315 2957
rect 113541 2954 113607 2957
rect 81249 2952 113607 2954
rect 81249 2896 81254 2952
rect 81310 2896 113546 2952
rect 113602 2896 113607 2952
rect 81249 2894 113607 2896
rect 81249 2891 81315 2894
rect 113541 2891 113607 2894
rect 116669 2954 116735 2957
rect 118601 2954 118667 2957
rect 116669 2952 118667 2954
rect 116669 2896 116674 2952
rect 116730 2896 118606 2952
rect 118662 2896 118667 2952
rect 116669 2894 118667 2896
rect 116669 2891 116735 2894
rect 118601 2891 118667 2894
rect 125133 2954 125199 2957
rect 128445 2954 128511 2957
rect 135621 2954 135687 2957
rect 125133 2952 128511 2954
rect 125133 2896 125138 2952
rect 125194 2896 128450 2952
rect 128506 2896 128511 2952
rect 125133 2894 128511 2896
rect 125133 2891 125199 2894
rect 128445 2891 128511 2894
rect 132910 2952 135687 2954
rect 132910 2896 135626 2952
rect 135682 2896 135687 2952
rect 132910 2894 135687 2896
rect 107009 2818 107075 2821
rect 110505 2818 110571 2821
rect 107009 2816 110571 2818
rect 107009 2760 107014 2816
rect 107070 2760 110510 2816
rect 110566 2760 110571 2816
rect 107009 2758 110571 2760
rect 107009 2755 107075 2758
rect 110505 2755 110571 2758
rect 116853 2818 116919 2821
rect 122557 2818 122623 2821
rect 116853 2816 122623 2818
rect 116853 2760 116858 2816
rect 116914 2760 122562 2816
rect 122618 2760 122623 2816
rect 116853 2758 122623 2760
rect 116853 2755 116919 2758
rect 122557 2755 122623 2758
rect 123937 2818 124003 2821
rect 132910 2818 132970 2894
rect 135621 2891 135687 2894
rect 135897 2954 135963 2957
rect 142846 2954 142906 3030
rect 151854 3028 151860 3030
rect 151924 3028 151930 3092
rect 151997 3090 152063 3093
rect 157244 3090 157304 3166
rect 162894 3164 162900 3166
rect 162964 3164 162970 3228
rect 164734 3164 164740 3228
rect 164804 3226 164810 3228
rect 166758 3226 166764 3228
rect 164804 3166 166764 3226
rect 164804 3164 164810 3166
rect 166758 3164 166764 3166
rect 166828 3164 166834 3228
rect 151997 3088 157304 3090
rect 151997 3032 152002 3088
rect 152058 3032 157304 3088
rect 151997 3030 157304 3032
rect 151997 3027 152063 3030
rect 157374 3028 157380 3092
rect 157444 3090 157450 3092
rect 161790 3090 161796 3092
rect 157444 3030 161796 3090
rect 157444 3028 157450 3030
rect 161790 3028 161796 3030
rect 161860 3028 161866 3092
rect 161974 3028 161980 3092
rect 162044 3090 162050 3092
rect 168966 3090 168972 3092
rect 162044 3030 168972 3090
rect 162044 3028 162050 3030
rect 168966 3028 168972 3030
rect 169036 3028 169042 3092
rect 169480 2957 169540 3302
rect 169886 3164 169892 3228
rect 169956 3226 169962 3228
rect 169956 3166 176210 3226
rect 169956 3164 169962 3166
rect 145189 2954 145255 2957
rect 162209 2954 162275 2957
rect 135897 2952 142906 2954
rect 135897 2896 135902 2952
rect 135958 2896 142906 2952
rect 135897 2894 142906 2896
rect 143904 2894 144378 2954
rect 135897 2891 135963 2894
rect 123937 2816 132970 2818
rect 123937 2760 123942 2816
rect 123998 2760 132970 2816
rect 123937 2758 132970 2760
rect 133505 2818 133571 2821
rect 141417 2818 141483 2821
rect 133505 2816 141483 2818
rect 133505 2760 133510 2816
rect 133566 2760 141422 2816
rect 141478 2760 141483 2816
rect 133505 2758 141483 2760
rect 123937 2755 124003 2758
rect 133505 2755 133571 2758
rect 141417 2755 141483 2758
rect 24071 2752 24137 2753
rect 64071 2752 64137 2753
rect 104071 2752 104137 2753
rect 24066 2688 24072 2752
rect 24136 2688 24142 2752
rect 64066 2688 64072 2752
rect 64136 2688 64142 2752
rect 104066 2688 104072 2752
rect 104136 2688 104142 2752
rect 24071 2687 24137 2688
rect 64071 2687 64137 2688
rect 104071 2687 104137 2688
rect 104617 2682 104683 2685
rect 118233 2682 118299 2685
rect 104617 2680 118299 2682
rect 104617 2624 104622 2680
rect 104678 2624 118238 2680
rect 118294 2624 118299 2680
rect 104617 2622 118299 2624
rect 104617 2619 104683 2622
rect 118233 2619 118299 2622
rect 122097 2682 122163 2685
rect 125409 2682 125475 2685
rect 122097 2680 125475 2682
rect 122097 2624 122102 2680
rect 122158 2624 125414 2680
rect 125470 2624 125475 2680
rect 122097 2622 125475 2624
rect 122097 2619 122163 2622
rect 125409 2619 125475 2622
rect 128813 2682 128879 2685
rect 132033 2682 132099 2685
rect 128813 2680 132099 2682
rect 128813 2624 128818 2680
rect 128874 2624 132038 2680
rect 132094 2624 132099 2680
rect 128813 2622 132099 2624
rect 128813 2619 128879 2622
rect 132033 2619 132099 2622
rect 132217 2682 132283 2685
rect 138197 2682 138263 2685
rect 132217 2680 138263 2682
rect 132217 2624 132222 2680
rect 132278 2624 138202 2680
rect 138258 2624 138263 2680
rect 132217 2622 138263 2624
rect 132217 2619 132283 2622
rect 138197 2619 138263 2622
rect 138422 2620 138428 2684
rect 138492 2682 138498 2684
rect 140037 2682 140103 2685
rect 138492 2680 140103 2682
rect 138492 2624 140042 2680
rect 140098 2624 140103 2680
rect 138492 2622 140103 2624
rect 138492 2620 138498 2622
rect 140037 2619 140103 2622
rect 141601 2682 141667 2685
rect 143904 2682 143964 2894
rect 144071 2752 144137 2753
rect 144066 2688 144072 2752
rect 144136 2688 144142 2752
rect 144071 2687 144137 2688
rect 141601 2680 143964 2682
rect 141601 2624 141606 2680
rect 141662 2624 143964 2680
rect 141601 2622 143964 2624
rect 144318 2682 144378 2894
rect 145189 2952 162275 2954
rect 145189 2896 145194 2952
rect 145250 2896 162214 2952
rect 162270 2896 162275 2952
rect 145189 2894 162275 2896
rect 145189 2891 145255 2894
rect 162209 2891 162275 2894
rect 162342 2892 162348 2956
rect 162412 2954 162418 2956
rect 165337 2954 165403 2957
rect 165521 2956 165587 2957
rect 162412 2952 165403 2954
rect 162412 2896 165342 2952
rect 165398 2896 165403 2952
rect 162412 2894 165403 2896
rect 162412 2892 162418 2894
rect 165337 2891 165403 2894
rect 165470 2892 165476 2956
rect 165540 2954 165587 2956
rect 167269 2954 167335 2957
rect 168046 2954 168052 2956
rect 165540 2952 165632 2954
rect 165582 2896 165632 2952
rect 165540 2894 165632 2896
rect 167269 2952 168052 2954
rect 167269 2896 167274 2952
rect 167330 2896 168052 2952
rect 167269 2894 168052 2896
rect 165540 2892 165587 2894
rect 165521 2891 165587 2892
rect 167269 2891 167335 2894
rect 168046 2892 168052 2894
rect 168116 2892 168122 2956
rect 169477 2952 169543 2957
rect 169753 2956 169819 2957
rect 169477 2896 169482 2952
rect 169538 2896 169543 2952
rect 169477 2891 169543 2896
rect 169702 2892 169708 2956
rect 169772 2954 169819 2956
rect 170029 2956 170095 2957
rect 171685 2956 171751 2957
rect 174905 2956 174971 2957
rect 169772 2952 169864 2954
rect 169814 2896 169864 2952
rect 169772 2894 169864 2896
rect 170029 2952 170076 2956
rect 170140 2954 170146 2956
rect 171685 2954 171732 2956
rect 170029 2896 170034 2952
rect 169772 2892 169819 2894
rect 169753 2891 169819 2892
rect 170029 2892 170076 2896
rect 170140 2894 170186 2954
rect 171640 2952 171732 2954
rect 171640 2896 171690 2952
rect 171640 2894 171732 2896
rect 170140 2892 170146 2894
rect 171685 2892 171732 2894
rect 171796 2892 171802 2956
rect 174854 2892 174860 2956
rect 174924 2954 174971 2956
rect 175917 2956 175983 2957
rect 175917 2954 175964 2956
rect 174924 2952 175016 2954
rect 174966 2896 175016 2952
rect 174924 2894 175016 2896
rect 175872 2952 175964 2954
rect 175872 2896 175922 2952
rect 175872 2894 175964 2896
rect 174924 2892 174971 2894
rect 170029 2891 170095 2892
rect 171685 2891 171751 2892
rect 174905 2891 174971 2892
rect 175917 2892 175964 2894
rect 176028 2892 176034 2956
rect 176150 2954 176210 3166
rect 180382 2957 180442 3302
rect 176469 2954 176535 2957
rect 176150 2952 176535 2954
rect 176150 2896 176474 2952
rect 176530 2896 176535 2952
rect 176150 2894 176535 2896
rect 175917 2891 175983 2892
rect 176469 2891 176535 2894
rect 176745 2954 176811 2957
rect 177849 2956 177915 2957
rect 177062 2954 177068 2956
rect 176745 2952 177068 2954
rect 176745 2896 176750 2952
rect 176806 2896 177068 2952
rect 176745 2894 177068 2896
rect 176745 2891 176811 2894
rect 177062 2892 177068 2894
rect 177132 2892 177138 2956
rect 177798 2892 177804 2956
rect 177868 2954 177915 2956
rect 177868 2952 177960 2954
rect 177910 2896 177960 2952
rect 177868 2894 177960 2896
rect 180382 2952 180491 2957
rect 180382 2896 180430 2952
rect 180486 2896 180491 2952
rect 180382 2894 180491 2896
rect 177868 2892 177915 2894
rect 177849 2891 177915 2892
rect 180425 2891 180491 2894
rect 144453 2818 144519 2821
rect 162485 2818 162551 2821
rect 163773 2818 163839 2821
rect 144453 2816 162551 2818
rect 144453 2760 144458 2816
rect 144514 2760 162490 2816
rect 162546 2760 162551 2816
rect 144453 2758 162551 2760
rect 144453 2755 144519 2758
rect 162485 2755 162551 2758
rect 162718 2816 163839 2818
rect 162718 2760 163778 2816
rect 163834 2760 163839 2816
rect 162718 2758 163839 2760
rect 157057 2682 157123 2685
rect 161974 2682 161980 2684
rect 144318 2622 153762 2682
rect 141601 2619 141667 2622
rect 90265 2546 90331 2549
rect 115197 2546 115263 2549
rect 90265 2544 115263 2546
rect 90265 2488 90270 2544
rect 90326 2488 115202 2544
rect 115258 2488 115263 2544
rect 90265 2486 115263 2488
rect 90265 2483 90331 2486
rect 115197 2483 115263 2486
rect 120993 2546 121059 2549
rect 125225 2546 125291 2549
rect 120993 2544 125291 2546
rect 120993 2488 120998 2544
rect 121054 2488 125230 2544
rect 125286 2488 125291 2544
rect 120993 2486 125291 2488
rect 120993 2483 121059 2486
rect 125225 2483 125291 2486
rect 125685 2546 125751 2549
rect 153561 2546 153627 2549
rect 125685 2544 153627 2546
rect 125685 2488 125690 2544
rect 125746 2488 153566 2544
rect 153622 2488 153627 2544
rect 125685 2486 153627 2488
rect 125685 2483 125751 2486
rect 153561 2483 153627 2486
rect 79133 2410 79199 2413
rect 112345 2410 112411 2413
rect 79133 2408 112411 2410
rect 79133 2352 79138 2408
rect 79194 2352 112350 2408
rect 112406 2352 112411 2408
rect 79133 2350 112411 2352
rect 79133 2347 79199 2350
rect 112345 2347 112411 2350
rect 120165 2410 120231 2413
rect 124673 2410 124739 2413
rect 151169 2410 151235 2413
rect 120165 2408 124322 2410
rect 120165 2352 120170 2408
rect 120226 2352 124322 2408
rect 120165 2350 124322 2352
rect 120165 2347 120231 2350
rect 106641 2274 106707 2277
rect 108757 2274 108823 2277
rect 106641 2272 108823 2274
rect 106641 2216 106646 2272
rect 106702 2216 108762 2272
rect 108818 2216 108823 2272
rect 106641 2214 108823 2216
rect 106641 2211 106707 2214
rect 108757 2211 108823 2214
rect 109033 2274 109099 2277
rect 110965 2274 111031 2277
rect 116301 2274 116367 2277
rect 109033 2272 111031 2274
rect 109033 2216 109038 2272
rect 109094 2216 110970 2272
rect 111026 2216 111031 2272
rect 109033 2214 111031 2216
rect 109033 2211 109099 2214
rect 110965 2211 111031 2214
rect 111382 2272 116367 2274
rect 111382 2216 116306 2272
rect 116362 2216 116367 2272
rect 111382 2214 116367 2216
rect 4071 2208 4137 2209
rect 44071 2208 44137 2209
rect 84071 2208 84137 2209
rect 4066 2144 4072 2208
rect 4136 2144 4142 2208
rect 44066 2144 44072 2208
rect 44136 2144 44142 2208
rect 84066 2144 84072 2208
rect 84136 2144 84142 2208
rect 4071 2143 4137 2144
rect 44071 2143 44137 2144
rect 84071 2143 84137 2144
rect 101121 2138 101187 2141
rect 105445 2138 105511 2141
rect 101121 2136 105511 2138
rect 101121 2080 101126 2136
rect 101182 2080 105450 2136
rect 105506 2080 105511 2136
rect 101121 2078 105511 2080
rect 101121 2075 101187 2078
rect 105445 2075 105511 2078
rect 108389 2138 108455 2141
rect 109217 2138 109283 2141
rect 108389 2136 109283 2138
rect 108389 2080 108394 2136
rect 108450 2080 109222 2136
rect 109278 2080 109283 2136
rect 108389 2078 109283 2080
rect 108389 2075 108455 2078
rect 109217 2075 109283 2078
rect 109493 2138 109559 2141
rect 111382 2138 111442 2214
rect 116301 2211 116367 2214
rect 117129 2274 117195 2277
rect 120809 2274 120875 2277
rect 117129 2272 120875 2274
rect 117129 2216 117134 2272
rect 117190 2216 120814 2272
rect 120870 2216 120875 2272
rect 117129 2214 120875 2216
rect 124262 2274 124322 2350
rect 124673 2408 151235 2410
rect 124673 2352 124678 2408
rect 124734 2352 151174 2408
rect 151230 2352 151235 2408
rect 124673 2350 151235 2352
rect 153702 2410 153762 2622
rect 157057 2680 161980 2682
rect 157057 2624 157062 2680
rect 157118 2624 161980 2680
rect 157057 2622 161980 2624
rect 157057 2619 157123 2622
rect 161974 2620 161980 2622
rect 162044 2620 162050 2684
rect 162209 2682 162275 2685
rect 162718 2682 162778 2758
rect 163773 2755 163839 2758
rect 164325 2818 164391 2821
rect 164734 2818 164740 2820
rect 164325 2816 164740 2818
rect 164325 2760 164330 2816
rect 164386 2760 164740 2816
rect 164325 2758 164740 2760
rect 164325 2755 164391 2758
rect 164734 2756 164740 2758
rect 164804 2756 164810 2820
rect 165102 2756 165108 2820
rect 165172 2818 165178 2820
rect 166574 2818 166580 2820
rect 165172 2758 166580 2818
rect 165172 2756 165178 2758
rect 166574 2756 166580 2758
rect 166644 2756 166650 2820
rect 166717 2818 166783 2821
rect 167862 2818 167868 2820
rect 166717 2816 167868 2818
rect 166717 2760 166722 2816
rect 166778 2760 167868 2816
rect 166717 2758 167868 2760
rect 166717 2755 166783 2758
rect 167862 2756 167868 2758
rect 167932 2756 167938 2820
rect 168557 2818 168623 2821
rect 169661 2818 169727 2821
rect 169886 2818 169892 2820
rect 168557 2816 169586 2818
rect 168557 2760 168562 2816
rect 168618 2760 169586 2816
rect 168557 2758 169586 2760
rect 168557 2755 168623 2758
rect 162209 2680 162778 2682
rect 162209 2624 162214 2680
rect 162270 2624 162778 2680
rect 162209 2622 162778 2624
rect 162209 2619 162275 2622
rect 162894 2620 162900 2684
rect 162964 2682 162970 2684
rect 165245 2682 165311 2685
rect 162964 2680 165311 2682
rect 162964 2624 165250 2680
rect 165306 2624 165311 2680
rect 162964 2622 165311 2624
rect 162964 2620 162970 2622
rect 165245 2619 165311 2622
rect 165429 2682 165495 2685
rect 166022 2682 166028 2684
rect 165429 2680 166028 2682
rect 165429 2624 165434 2680
rect 165490 2624 166028 2680
rect 165429 2622 166028 2624
rect 165429 2619 165495 2622
rect 166022 2620 166028 2622
rect 166092 2620 166098 2684
rect 167269 2682 167335 2685
rect 167729 2684 167795 2685
rect 167494 2682 167500 2684
rect 167269 2680 167500 2682
rect 167269 2624 167274 2680
rect 167330 2624 167500 2680
rect 167269 2622 167500 2624
rect 167269 2619 167335 2622
rect 167494 2620 167500 2622
rect 167564 2620 167570 2684
rect 167678 2620 167684 2684
rect 167748 2682 167795 2684
rect 169526 2682 169586 2758
rect 169661 2816 169892 2818
rect 169661 2760 169666 2816
rect 169722 2760 169892 2816
rect 169661 2758 169892 2760
rect 169661 2755 169727 2758
rect 169886 2756 169892 2758
rect 169956 2756 169962 2820
rect 171358 2818 171364 2820
rect 170078 2758 171364 2818
rect 170078 2682 170138 2758
rect 171358 2756 171364 2758
rect 171428 2756 171434 2820
rect 173249 2818 173315 2821
rect 173382 2818 173388 2820
rect 173249 2816 173388 2818
rect 173249 2760 173254 2816
rect 173310 2760 173388 2816
rect 173249 2758 173388 2760
rect 173249 2755 173315 2758
rect 173382 2756 173388 2758
rect 173452 2756 173458 2820
rect 173750 2756 173756 2820
rect 173820 2818 173826 2820
rect 175273 2818 175339 2821
rect 176561 2820 176627 2821
rect 176510 2818 176516 2820
rect 173820 2816 175339 2818
rect 173820 2760 175278 2816
rect 175334 2760 175339 2816
rect 173820 2758 175339 2760
rect 176470 2758 176516 2818
rect 176580 2816 176627 2820
rect 176622 2760 176627 2816
rect 173820 2756 173826 2758
rect 175273 2755 175339 2758
rect 176510 2756 176516 2758
rect 176580 2756 176627 2760
rect 176561 2755 176627 2756
rect 184071 2752 184137 2753
rect 184066 2688 184072 2752
rect 184136 2688 184142 2752
rect 184071 2687 184137 2688
rect 171133 2684 171199 2685
rect 171133 2682 171180 2684
rect 167748 2680 167840 2682
rect 167790 2624 167840 2680
rect 167748 2622 167840 2624
rect 169526 2622 170138 2682
rect 171088 2680 171180 2682
rect 171088 2624 171138 2680
rect 171088 2622 171180 2624
rect 167748 2620 167795 2622
rect 167729 2619 167795 2620
rect 171133 2620 171180 2622
rect 171244 2620 171250 2684
rect 171317 2682 171383 2685
rect 171317 2680 181362 2682
rect 171317 2624 171322 2680
rect 171378 2624 181362 2680
rect 171317 2622 181362 2624
rect 171133 2619 171199 2620
rect 171317 2619 171383 2622
rect 157057 2546 157123 2549
rect 180742 2546 180748 2548
rect 157057 2544 180748 2546
rect 157057 2488 157062 2544
rect 157118 2488 180748 2544
rect 157057 2486 180748 2488
rect 157057 2483 157123 2486
rect 180742 2484 180748 2486
rect 180812 2484 180818 2548
rect 181302 2546 181362 2622
rect 186037 2546 186103 2549
rect 181302 2544 186103 2546
rect 181302 2488 186042 2544
rect 186098 2488 186103 2544
rect 181302 2486 186103 2488
rect 186037 2483 186103 2486
rect 162945 2410 163011 2413
rect 153702 2408 163011 2410
rect 153702 2352 162950 2408
rect 163006 2352 163011 2408
rect 153702 2350 163011 2352
rect 124673 2347 124739 2350
rect 151169 2347 151235 2350
rect 162945 2347 163011 2350
rect 163129 2410 163195 2413
rect 163681 2410 163747 2413
rect 165889 2410 165955 2413
rect 171317 2410 171383 2413
rect 163129 2408 163747 2410
rect 163129 2352 163134 2408
rect 163190 2352 163686 2408
rect 163742 2352 163747 2408
rect 163129 2350 163747 2352
rect 163129 2347 163195 2350
rect 163681 2347 163747 2350
rect 163822 2408 165955 2410
rect 163822 2352 165894 2408
rect 165950 2352 165955 2408
rect 163822 2350 165955 2352
rect 138054 2274 138060 2276
rect 124262 2214 138060 2274
rect 117129 2211 117195 2214
rect 120809 2211 120875 2214
rect 138054 2212 138060 2214
rect 138124 2212 138130 2276
rect 138238 2212 138244 2276
rect 138308 2274 138314 2276
rect 146109 2274 146175 2277
rect 138308 2272 146175 2274
rect 138308 2216 146114 2272
rect 146170 2216 146175 2272
rect 138308 2214 146175 2216
rect 138308 2212 138314 2214
rect 146109 2211 146175 2214
rect 146385 2274 146451 2277
rect 159449 2274 159515 2277
rect 146385 2272 159515 2274
rect 146385 2216 146390 2272
rect 146446 2216 159454 2272
rect 159510 2216 159515 2272
rect 146385 2214 159515 2216
rect 146385 2211 146451 2214
rect 159449 2211 159515 2214
rect 159725 2274 159791 2277
rect 161749 2274 161815 2277
rect 163822 2274 163882 2350
rect 165889 2347 165955 2350
rect 166030 2408 171383 2410
rect 166030 2352 171322 2408
rect 171378 2352 171383 2408
rect 166030 2350 171383 2352
rect 159725 2272 161674 2274
rect 159725 2216 159730 2272
rect 159786 2216 161674 2272
rect 159725 2214 161674 2216
rect 159725 2211 159791 2214
rect 124071 2208 124137 2209
rect 124066 2144 124072 2208
rect 124136 2144 124142 2208
rect 124071 2143 124137 2144
rect 109493 2136 111442 2138
rect 109493 2080 109498 2136
rect 109554 2080 111442 2136
rect 109493 2078 111442 2080
rect 111517 2138 111583 2141
rect 124213 2138 124279 2141
rect 127433 2138 127499 2141
rect 111517 2136 122850 2138
rect 111517 2080 111522 2136
rect 111578 2080 122850 2136
rect 111517 2078 122850 2080
rect 109493 2075 109559 2078
rect 111517 2075 111583 2078
rect 92013 2002 92079 2005
rect 113541 2002 113607 2005
rect 92013 2000 113607 2002
rect 92013 1944 92018 2000
rect 92074 1944 113546 2000
rect 113602 1944 113607 2000
rect 92013 1942 113607 1944
rect 92013 1939 92079 1942
rect 113541 1939 113607 1942
rect -400 1866 800 1896
rect 4061 1866 4127 1869
rect -400 1864 4127 1866
rect -400 1808 4066 1864
rect 4122 1808 4127 1864
rect -400 1806 4127 1808
rect -400 1776 800 1806
rect 4061 1803 4127 1806
rect 86769 1866 86835 1869
rect 112069 1866 112135 1869
rect 86769 1864 112135 1866
rect 86769 1808 86774 1864
rect 86830 1808 112074 1864
rect 112130 1808 112135 1864
rect 86769 1806 112135 1808
rect 86769 1803 86835 1806
rect 112069 1803 112135 1806
rect 112253 1866 112319 1869
rect 119153 1866 119219 1869
rect 112253 1864 119219 1866
rect 112253 1808 112258 1864
rect 112314 1808 119158 1864
rect 119214 1808 119219 1864
rect 112253 1806 119219 1808
rect 122790 1866 122850 2078
rect 124213 2136 127499 2138
rect 124213 2080 124218 2136
rect 124274 2080 127438 2136
rect 127494 2080 127499 2136
rect 124213 2078 127499 2080
rect 124213 2075 124279 2078
rect 127433 2075 127499 2078
rect 127617 2138 127683 2141
rect 131481 2138 131547 2141
rect 127617 2136 131547 2138
rect 127617 2080 127622 2136
rect 127678 2080 131486 2136
rect 131542 2080 131547 2136
rect 127617 2078 131547 2080
rect 127617 2075 127683 2078
rect 131481 2075 131547 2078
rect 131757 2138 131823 2141
rect 137737 2138 137803 2141
rect 131757 2136 137803 2138
rect 131757 2080 131762 2136
rect 131818 2080 137742 2136
rect 137798 2080 137803 2136
rect 131757 2078 137803 2080
rect 131757 2075 131823 2078
rect 137737 2075 137803 2078
rect 137870 2076 137876 2140
rect 137940 2138 137946 2140
rect 139485 2138 139551 2141
rect 137940 2136 139551 2138
rect 137940 2080 139490 2136
rect 139546 2080 139551 2136
rect 137940 2078 139551 2080
rect 137940 2076 137946 2078
rect 139485 2075 139551 2078
rect 140037 2138 140103 2141
rect 145557 2138 145623 2141
rect 140037 2136 145623 2138
rect 140037 2080 140042 2136
rect 140098 2080 145562 2136
rect 145618 2080 145623 2136
rect 140037 2078 145623 2080
rect 140037 2075 140103 2078
rect 145557 2075 145623 2078
rect 145833 2138 145899 2141
rect 160829 2138 160895 2141
rect 161422 2138 161428 2140
rect 145833 2136 159466 2138
rect 145833 2080 145838 2136
rect 145894 2080 159466 2136
rect 145833 2078 159466 2080
rect 145833 2075 145899 2078
rect 123753 2002 123819 2005
rect 125317 2002 125383 2005
rect 123753 2000 125383 2002
rect 123753 1944 123758 2000
rect 123814 1944 125322 2000
rect 125378 1944 125383 2000
rect 123753 1942 125383 1944
rect 123753 1939 123819 1942
rect 125317 1939 125383 1942
rect 125777 2002 125843 2005
rect 152181 2002 152247 2005
rect 125777 2000 152247 2002
rect 125777 1944 125782 2000
rect 125838 1944 152186 2000
rect 152242 1944 152247 2000
rect 125777 1942 152247 1944
rect 125777 1939 125843 1942
rect 152181 1939 152247 1942
rect 155769 2002 155835 2005
rect 158529 2002 158595 2005
rect 155769 2000 158595 2002
rect 155769 1944 155774 2000
rect 155830 1944 158534 2000
rect 158590 1944 158595 2000
rect 155769 1942 158595 1944
rect 155769 1939 155835 1942
rect 158529 1939 158595 1942
rect 158713 2002 158779 2005
rect 158846 2002 158852 2004
rect 158713 2000 158852 2002
rect 158713 1944 158718 2000
rect 158774 1944 158852 2000
rect 158713 1942 158852 1944
rect 158713 1939 158779 1942
rect 158846 1940 158852 1942
rect 158916 1940 158922 2004
rect 159406 2002 159466 2078
rect 160829 2136 161428 2138
rect 160829 2080 160834 2136
rect 160890 2080 161428 2136
rect 160829 2078 161428 2080
rect 160829 2075 160895 2078
rect 161422 2076 161428 2078
rect 161492 2076 161498 2140
rect 161614 2138 161674 2214
rect 161749 2272 163882 2274
rect 161749 2216 161754 2272
rect 161810 2216 163882 2272
rect 161749 2214 163882 2216
rect 164233 2274 164299 2277
rect 166030 2274 166090 2350
rect 171317 2347 171383 2350
rect 171910 2348 171916 2412
rect 171980 2410 171986 2412
rect 175774 2410 175780 2412
rect 171980 2350 175780 2410
rect 171980 2348 171986 2350
rect 175774 2348 175780 2350
rect 175844 2348 175850 2412
rect 176285 2410 176351 2413
rect 179505 2410 179571 2413
rect 176285 2408 179571 2410
rect 176285 2352 176290 2408
rect 176346 2352 179510 2408
rect 179566 2352 179571 2408
rect 176285 2350 179571 2352
rect 176285 2347 176351 2350
rect 179505 2347 179571 2350
rect 182541 2410 182607 2413
rect 185669 2410 185735 2413
rect 187509 2410 187575 2413
rect 182541 2408 185735 2410
rect 182541 2352 182546 2408
rect 182602 2352 185674 2408
rect 185730 2352 185735 2408
rect 182541 2350 185735 2352
rect 182541 2347 182607 2350
rect 185669 2347 185735 2350
rect 185902 2408 187575 2410
rect 185902 2352 187514 2408
rect 187570 2352 187575 2408
rect 185902 2350 187575 2352
rect 164233 2272 166090 2274
rect 164233 2216 164238 2272
rect 164294 2216 166090 2272
rect 164233 2214 166090 2216
rect 166993 2274 167059 2277
rect 168649 2274 168715 2277
rect 166993 2272 168715 2274
rect 166993 2216 166998 2272
rect 167054 2216 168654 2272
rect 168710 2216 168715 2272
rect 166993 2214 168715 2216
rect 161749 2211 161815 2214
rect 164233 2211 164299 2214
rect 166993 2211 167059 2214
rect 168649 2211 168715 2214
rect 169518 2212 169524 2276
rect 169588 2274 169594 2276
rect 169753 2274 169819 2277
rect 169588 2272 169819 2274
rect 169588 2216 169758 2272
rect 169814 2216 169819 2272
rect 169588 2214 169819 2216
rect 169588 2212 169594 2214
rect 169753 2211 169819 2214
rect 170806 2212 170812 2276
rect 170876 2274 170882 2276
rect 176193 2274 176259 2277
rect 170876 2272 176259 2274
rect 170876 2216 176198 2272
rect 176254 2216 176259 2272
rect 170876 2214 176259 2216
rect 170876 2212 170882 2214
rect 176193 2211 176259 2214
rect 176326 2212 176332 2276
rect 176396 2274 176402 2276
rect 177021 2274 177087 2277
rect 176396 2272 177087 2274
rect 176396 2216 177026 2272
rect 177082 2216 177087 2272
rect 176396 2214 177087 2216
rect 176396 2212 176402 2214
rect 177021 2211 177087 2214
rect 184933 2274 184999 2277
rect 185902 2274 185962 2350
rect 187509 2347 187575 2350
rect 184933 2272 185962 2274
rect 184933 2216 184938 2272
rect 184994 2216 185962 2272
rect 184933 2214 185962 2216
rect 186313 2274 186379 2277
rect 189809 2274 189875 2277
rect 186313 2272 189875 2274
rect 186313 2216 186318 2272
rect 186374 2216 189814 2272
rect 189870 2216 189875 2272
rect 186313 2214 189875 2216
rect 184933 2211 184999 2214
rect 186313 2211 186379 2214
rect 189809 2211 189875 2214
rect 164071 2208 164137 2209
rect 164066 2144 164072 2208
rect 164136 2144 164142 2208
rect 164071 2143 164137 2144
rect 163865 2138 163931 2141
rect 161614 2136 163931 2138
rect 161614 2080 163870 2136
rect 163926 2080 163931 2136
rect 161614 2078 163931 2080
rect 163865 2075 163931 2078
rect 164233 2138 164299 2141
rect 165838 2138 165844 2140
rect 164233 2136 165844 2138
rect 164233 2080 164238 2136
rect 164294 2080 165844 2136
rect 164233 2078 165844 2080
rect 164233 2075 164299 2078
rect 165838 2076 165844 2078
rect 165908 2076 165914 2140
rect 166901 2138 166967 2141
rect 171317 2138 171383 2141
rect 178309 2138 178375 2141
rect 181989 2140 182055 2141
rect 181989 2138 182036 2140
rect 166901 2136 171383 2138
rect 166901 2080 166906 2136
rect 166962 2080 171322 2136
rect 171378 2080 171383 2136
rect 166901 2078 171383 2080
rect 166901 2075 166967 2078
rect 171317 2075 171383 2078
rect 171734 2136 178375 2138
rect 171734 2080 178314 2136
rect 178370 2080 178375 2136
rect 171734 2078 178375 2080
rect 181944 2136 182036 2138
rect 181944 2080 181994 2136
rect 181944 2078 182036 2080
rect 171734 2002 171794 2078
rect 178309 2075 178375 2078
rect 181989 2076 182036 2078
rect 182100 2076 182106 2140
rect 186129 2138 186195 2141
rect 186405 2138 186471 2141
rect 186129 2136 186471 2138
rect 186129 2080 186134 2136
rect 186190 2080 186410 2136
rect 186466 2080 186471 2136
rect 186129 2078 186471 2080
rect 181989 2075 182055 2076
rect 186129 2075 186195 2078
rect 186405 2075 186471 2078
rect 187325 2138 187391 2141
rect 192661 2138 192727 2141
rect 187325 2136 192727 2138
rect 187325 2080 187330 2136
rect 187386 2080 192666 2136
rect 192722 2080 192727 2136
rect 187325 2078 192727 2080
rect 187325 2075 187391 2078
rect 192661 2075 192727 2078
rect 159406 1942 171794 2002
rect 171869 2002 171935 2005
rect 193305 2002 193371 2005
rect 171869 2000 193371 2002
rect 171869 1944 171874 2000
rect 171930 1944 193310 2000
rect 193366 1944 193371 2000
rect 171869 1942 193371 1944
rect 171869 1939 171935 1942
rect 193305 1939 193371 1942
rect 126881 1866 126947 1869
rect 122790 1864 126947 1866
rect 122790 1808 126886 1864
rect 126942 1808 126947 1864
rect 122790 1806 126947 1808
rect 112253 1803 112319 1806
rect 119153 1803 119219 1806
rect 126881 1803 126947 1806
rect 127341 1866 127407 1869
rect 132309 1866 132375 1869
rect 127341 1864 132375 1866
rect 127341 1808 127346 1864
rect 127402 1808 132314 1864
rect 132370 1808 132375 1864
rect 127341 1806 132375 1808
rect 127341 1803 127407 1806
rect 132309 1803 132375 1806
rect 134425 1866 134491 1869
rect 137093 1866 137159 1869
rect 134425 1864 137159 1866
rect 134425 1808 134430 1864
rect 134486 1808 137098 1864
rect 137154 1808 137159 1864
rect 134425 1806 137159 1808
rect 134425 1803 134491 1806
rect 137093 1803 137159 1806
rect 137277 1866 137343 1869
rect 137553 1866 137619 1869
rect 137277 1864 137619 1866
rect 137277 1808 137282 1864
rect 137338 1808 137558 1864
rect 137614 1808 137619 1864
rect 137277 1806 137619 1808
rect 137277 1803 137343 1806
rect 137553 1803 137619 1806
rect 137737 1866 137803 1869
rect 139301 1866 139367 1869
rect 137737 1864 139367 1866
rect 137737 1808 137742 1864
rect 137798 1808 139306 1864
rect 139362 1808 139367 1864
rect 137737 1806 139367 1808
rect 137737 1803 137803 1806
rect 139301 1803 139367 1806
rect 139485 1866 139551 1869
rect 161197 1866 161263 1869
rect 139485 1864 161263 1866
rect 139485 1808 139490 1864
rect 139546 1808 161202 1864
rect 161258 1808 161263 1864
rect 139485 1806 161263 1808
rect 139485 1803 139551 1806
rect 161197 1803 161263 1806
rect 161473 1866 161539 1869
rect 163681 1866 163747 1869
rect 161473 1864 163747 1866
rect 161473 1808 161478 1864
rect 161534 1808 163686 1864
rect 163742 1808 163747 1864
rect 161473 1806 163747 1808
rect 161473 1803 161539 1806
rect 163681 1803 163747 1806
rect 163865 1866 163931 1869
rect 165102 1866 165108 1868
rect 163865 1864 165108 1866
rect 163865 1808 163870 1864
rect 163926 1808 165108 1864
rect 163865 1806 165108 1808
rect 163865 1803 163931 1806
rect 165102 1804 165108 1806
rect 165172 1804 165178 1868
rect 165521 1866 165587 1869
rect 169385 1866 169451 1869
rect 173157 1866 173223 1869
rect 165521 1864 169218 1866
rect 165521 1808 165526 1864
rect 165582 1808 169218 1864
rect 165521 1806 169218 1808
rect 165521 1803 165587 1806
rect 107285 1730 107351 1733
rect 109677 1730 109743 1733
rect 107285 1728 109743 1730
rect 107285 1672 107290 1728
rect 107346 1672 109682 1728
rect 109738 1672 109743 1728
rect 107285 1670 109743 1672
rect 107285 1667 107351 1670
rect 109677 1667 109743 1670
rect 120073 1730 120139 1733
rect 138054 1730 138060 1732
rect 120073 1728 138060 1730
rect 120073 1672 120078 1728
rect 120134 1672 138060 1728
rect 120073 1670 138060 1672
rect 120073 1667 120139 1670
rect 138054 1668 138060 1670
rect 138124 1668 138130 1732
rect 138197 1730 138263 1733
rect 142245 1730 142311 1733
rect 138197 1728 142311 1730
rect 138197 1672 138202 1728
rect 138258 1672 142250 1728
rect 142306 1672 142311 1728
rect 138197 1670 142311 1672
rect 138197 1667 138263 1670
rect 142245 1667 142311 1670
rect 144269 1730 144335 1733
rect 165705 1730 165771 1733
rect 144269 1728 165771 1730
rect 144269 1672 144274 1728
rect 144330 1672 165710 1728
rect 165766 1672 165771 1728
rect 144269 1670 165771 1672
rect 144269 1667 144335 1670
rect 165705 1667 165771 1670
rect 165889 1730 165955 1733
rect 169017 1730 169083 1733
rect 165889 1728 169083 1730
rect 165889 1672 165894 1728
rect 165950 1672 169022 1728
rect 169078 1672 169083 1728
rect 165889 1670 169083 1672
rect 169158 1730 169218 1806
rect 169385 1864 173223 1866
rect 169385 1808 169390 1864
rect 169446 1808 173162 1864
rect 173218 1808 173223 1864
rect 169385 1806 173223 1808
rect 169385 1803 169451 1806
rect 173157 1803 173223 1806
rect 177113 1866 177179 1869
rect 183369 1866 183435 1869
rect 177113 1864 183435 1866
rect 177113 1808 177118 1864
rect 177174 1808 183374 1864
rect 183430 1808 183435 1864
rect 177113 1806 183435 1808
rect 177113 1803 177179 1806
rect 183369 1803 183435 1806
rect 186037 1866 186103 1869
rect 189441 1866 189507 1869
rect 186037 1864 189507 1866
rect 186037 1808 186042 1864
rect 186098 1808 189446 1864
rect 189502 1808 189507 1864
rect 186037 1806 189507 1808
rect 186037 1803 186103 1806
rect 189441 1803 189507 1806
rect 175590 1730 175596 1732
rect 169158 1670 175596 1730
rect 165889 1667 165955 1670
rect 169017 1667 169083 1670
rect 175590 1668 175596 1670
rect 175660 1668 175666 1732
rect 176009 1730 176075 1733
rect 181345 1730 181411 1733
rect 176009 1728 181411 1730
rect 176009 1672 176014 1728
rect 176070 1672 181350 1728
rect 181406 1672 181411 1728
rect 176009 1670 181411 1672
rect 176009 1667 176075 1670
rect 181345 1667 181411 1670
rect 24071 1664 24137 1665
rect 64071 1664 64137 1665
rect 104071 1664 104137 1665
rect 144071 1664 144137 1665
rect 184071 1664 184137 1665
rect 24066 1600 24072 1664
rect 24136 1600 24142 1664
rect 64066 1600 64072 1664
rect 64136 1600 64142 1664
rect 104066 1600 104072 1664
rect 104136 1600 104142 1664
rect 144066 1600 144072 1664
rect 144136 1600 144142 1664
rect 184066 1600 184072 1664
rect 184136 1600 184142 1664
rect 24071 1599 24137 1600
rect 64071 1599 64137 1600
rect 104071 1599 104137 1600
rect 144071 1599 144137 1600
rect 184071 1599 184137 1600
rect 109033 1594 109099 1597
rect 109769 1594 109835 1597
rect 109033 1592 109835 1594
rect 109033 1536 109038 1592
rect 109094 1536 109774 1592
rect 109830 1536 109835 1592
rect 109033 1534 109835 1536
rect 109033 1531 109099 1534
rect 109769 1531 109835 1534
rect 110137 1594 110203 1597
rect 124213 1594 124279 1597
rect 110137 1592 124279 1594
rect 110137 1536 110142 1592
rect 110198 1536 124218 1592
rect 124274 1536 124279 1592
rect 110137 1534 124279 1536
rect 110137 1531 110203 1534
rect 124213 1531 124279 1534
rect 125041 1594 125107 1597
rect 143901 1594 143967 1597
rect 149145 1594 149211 1597
rect 125041 1592 143967 1594
rect 125041 1536 125046 1592
rect 125102 1536 143906 1592
rect 143962 1536 143967 1592
rect 125041 1534 143967 1536
rect 125041 1531 125107 1534
rect 143901 1531 143967 1534
rect 144318 1592 149211 1594
rect 144318 1536 149150 1592
rect 149206 1536 149211 1592
rect 144318 1534 149211 1536
rect 80973 1458 81039 1461
rect 110689 1458 110755 1461
rect 80973 1456 110755 1458
rect 80973 1400 80978 1456
rect 81034 1400 110694 1456
rect 110750 1400 110755 1456
rect 80973 1398 110755 1400
rect 80973 1395 81039 1398
rect 110689 1395 110755 1398
rect 111977 1458 112043 1461
rect 120165 1458 120231 1461
rect 111977 1456 120231 1458
rect 111977 1400 111982 1456
rect 112038 1400 120170 1456
rect 120226 1400 120231 1456
rect 111977 1398 120231 1400
rect 111977 1395 112043 1398
rect 120165 1395 120231 1398
rect 124857 1458 124923 1461
rect 144318 1458 144378 1534
rect 149145 1531 149211 1534
rect 151169 1594 151235 1597
rect 154849 1594 154915 1597
rect 151169 1592 154915 1594
rect 151169 1536 151174 1592
rect 151230 1536 154854 1592
rect 154910 1536 154915 1592
rect 151169 1534 154915 1536
rect 151169 1531 151235 1534
rect 154849 1531 154915 1534
rect 156597 1594 156663 1597
rect 159633 1594 159699 1597
rect 156597 1592 159699 1594
rect 156597 1536 156602 1592
rect 156658 1536 159638 1592
rect 159694 1536 159699 1592
rect 156597 1534 159699 1536
rect 156597 1531 156663 1534
rect 159633 1531 159699 1534
rect 159950 1532 159956 1596
rect 160020 1594 160026 1596
rect 161013 1594 161079 1597
rect 164233 1594 164299 1597
rect 160020 1592 161079 1594
rect 160020 1536 161018 1592
rect 161074 1536 161079 1592
rect 160020 1534 161079 1536
rect 160020 1532 160026 1534
rect 161013 1531 161079 1534
rect 161200 1592 164299 1594
rect 161200 1536 164238 1592
rect 164294 1536 164299 1592
rect 161200 1534 164299 1536
rect 150525 1458 150591 1461
rect 124857 1456 144378 1458
rect 124857 1400 124862 1456
rect 124918 1400 144378 1456
rect 124857 1398 144378 1400
rect 144456 1456 150591 1458
rect 144456 1400 150530 1456
rect 150586 1400 150591 1456
rect 144456 1398 150591 1400
rect 124857 1395 124923 1398
rect 93669 1322 93735 1325
rect 142429 1322 142495 1325
rect 93669 1320 142495 1322
rect 93669 1264 93674 1320
rect 93730 1264 142434 1320
rect 142490 1264 142495 1320
rect 93669 1262 142495 1264
rect 93669 1259 93735 1262
rect 142429 1259 142495 1262
rect 143901 1322 143967 1325
rect 144456 1322 144516 1398
rect 150525 1395 150591 1398
rect 156781 1458 156847 1461
rect 161200 1458 161260 1534
rect 164233 1531 164299 1534
rect 164509 1594 164575 1597
rect 183553 1596 183619 1597
rect 177614 1594 177620 1596
rect 164509 1592 177620 1594
rect 164509 1536 164514 1592
rect 164570 1536 177620 1592
rect 164509 1534 177620 1536
rect 164509 1531 164575 1534
rect 177614 1532 177620 1534
rect 177684 1532 177690 1596
rect 183502 1532 183508 1596
rect 183572 1594 183619 1596
rect 183572 1592 183664 1594
rect 183614 1536 183664 1592
rect 183572 1534 183664 1536
rect 183572 1532 183619 1534
rect 183553 1531 183619 1532
rect 164693 1460 164759 1461
rect 156781 1456 161260 1458
rect 156781 1400 156786 1456
rect 156842 1400 161260 1456
rect 156781 1398 161260 1400
rect 161982 1398 164618 1458
rect 156781 1395 156847 1398
rect 143901 1320 144516 1322
rect 143901 1264 143906 1320
rect 143962 1264 144516 1320
rect 143901 1262 144516 1264
rect 144637 1322 144703 1325
rect 145741 1322 145807 1325
rect 144637 1320 145807 1322
rect 144637 1264 144642 1320
rect 144698 1264 145746 1320
rect 145802 1264 145807 1320
rect 144637 1262 145807 1264
rect 143901 1259 143967 1262
rect 144637 1259 144703 1262
rect 145741 1259 145807 1262
rect 156505 1322 156571 1325
rect 161982 1322 162042 1398
rect 164558 1322 164618 1398
rect 164693 1456 164740 1460
rect 164804 1458 164810 1460
rect 164693 1400 164698 1456
rect 164693 1396 164740 1400
rect 164804 1398 164850 1458
rect 164804 1396 164810 1398
rect 165102 1396 165108 1460
rect 165172 1458 165178 1460
rect 166758 1458 166764 1460
rect 165172 1398 166764 1458
rect 165172 1396 165178 1398
rect 166758 1396 166764 1398
rect 166828 1396 166834 1460
rect 167361 1458 167427 1461
rect 170990 1458 170996 1460
rect 167361 1456 170996 1458
rect 167361 1400 167366 1456
rect 167422 1400 170996 1456
rect 167361 1398 170996 1400
rect 164693 1395 164759 1396
rect 167361 1395 167427 1398
rect 170990 1396 170996 1398
rect 171060 1396 171066 1460
rect 171133 1458 171199 1461
rect 198825 1458 198891 1461
rect 171133 1456 198891 1458
rect 171133 1400 171138 1456
rect 171194 1400 198830 1456
rect 198886 1400 198891 1456
rect 171133 1398 198891 1400
rect 171133 1395 171199 1398
rect 198825 1395 198891 1398
rect 182214 1322 182220 1324
rect 156505 1320 162042 1322
rect 156505 1264 156510 1320
rect 156566 1264 162042 1320
rect 156505 1262 162042 1264
rect 162166 1262 164434 1322
rect 164558 1262 182220 1322
rect 156505 1259 156571 1262
rect 116853 1186 116919 1189
rect 121269 1186 121335 1189
rect 116853 1184 121335 1186
rect 116853 1128 116858 1184
rect 116914 1128 121274 1184
rect 121330 1128 121335 1184
rect 116853 1126 121335 1128
rect 116853 1123 116919 1126
rect 121269 1123 121335 1126
rect 132033 1186 132099 1189
rect 137686 1186 137692 1188
rect 132033 1184 137692 1186
rect 132033 1128 132038 1184
rect 132094 1128 137692 1184
rect 132033 1126 137692 1128
rect 132033 1123 132099 1126
rect 137686 1124 137692 1126
rect 137756 1124 137762 1188
rect 137870 1124 137876 1188
rect 137940 1186 137946 1188
rect 162166 1186 162226 1262
rect 137940 1126 162226 1186
rect 137940 1124 137946 1126
rect 162342 1124 162348 1188
rect 162412 1186 162418 1188
rect 163865 1186 163931 1189
rect 162412 1184 163931 1186
rect 162412 1128 163870 1184
rect 163926 1128 163931 1184
rect 162412 1126 163931 1128
rect 164374 1186 164434 1262
rect 182214 1260 182220 1262
rect 182284 1260 182290 1324
rect 175222 1186 175228 1188
rect 164374 1126 175228 1186
rect 162412 1124 162418 1126
rect 163865 1123 163931 1126
rect 175222 1124 175228 1126
rect 175292 1124 175298 1188
rect 4071 1120 4137 1121
rect 44071 1120 44137 1121
rect 84071 1120 84137 1121
rect 124071 1120 124137 1121
rect 164071 1120 164137 1121
rect 4066 1056 4072 1120
rect 4136 1056 4142 1120
rect 44066 1056 44072 1120
rect 44136 1056 44142 1120
rect 84066 1056 84072 1120
rect 84136 1056 84142 1120
rect 124066 1056 124072 1120
rect 124136 1056 124142 1120
rect 164066 1056 164072 1120
rect 164136 1056 164142 1120
rect 4071 1055 4137 1056
rect 44071 1055 44137 1056
rect 84071 1055 84137 1056
rect 124071 1055 124137 1056
rect 164071 1055 164137 1056
rect 128905 1050 128971 1053
rect 137134 1050 137140 1052
rect 128905 1048 137140 1050
rect 128905 992 128910 1048
rect 128966 992 137140 1048
rect 128905 990 137140 992
rect 128905 987 128971 990
rect 137134 988 137140 990
rect 137204 988 137210 1052
rect 137553 1050 137619 1053
rect 141785 1050 141851 1053
rect 137553 1048 141851 1050
rect 137553 992 137558 1048
rect 137614 992 141790 1048
rect 141846 992 141851 1048
rect 137553 990 141851 992
rect 137553 987 137619 990
rect 141785 987 141851 990
rect 142429 1050 142495 1053
rect 146753 1050 146819 1053
rect 142429 1048 146819 1050
rect 142429 992 142434 1048
rect 142490 992 146758 1048
rect 146814 992 146819 1048
rect 142429 990 146819 992
rect 142429 987 142495 990
rect 146753 987 146819 990
rect 151854 988 151860 1052
rect 151924 1050 151930 1052
rect 163865 1050 163931 1053
rect 151924 1048 163931 1050
rect 151924 992 163870 1048
rect 163926 992 163931 1048
rect 151924 990 163931 992
rect 151924 988 151930 990
rect 163865 987 163931 990
rect 164233 1050 164299 1053
rect 168097 1050 168163 1053
rect 164233 1048 168163 1050
rect 164233 992 164238 1048
rect 164294 992 168102 1048
rect 168158 992 168163 1048
rect 164233 990 168163 992
rect 164233 987 164299 990
rect 168097 987 168163 990
rect 168281 1050 168347 1053
rect 181529 1050 181595 1053
rect 168281 1048 181595 1050
rect 168281 992 168286 1048
rect 168342 992 181534 1048
rect 181590 992 181595 1048
rect 168281 990 181595 992
rect 168281 987 168347 990
rect 181529 987 181595 990
rect 123845 914 123911 917
rect 164969 914 165035 917
rect 123845 912 165035 914
rect 123845 856 123850 912
rect 123906 856 164974 912
rect 165030 856 165035 912
rect 123845 854 165035 856
rect 123845 851 123911 854
rect 164969 851 165035 854
rect 165429 914 165495 917
rect 170949 914 171015 917
rect 165429 912 171015 914
rect 165429 856 165434 912
rect 165490 856 170954 912
rect 171010 856 171015 912
rect 165429 854 171015 856
rect 165429 851 165495 854
rect 170949 851 171015 854
rect 110045 778 110111 781
rect 146661 778 146727 781
rect 110045 776 146727 778
rect 110045 720 110050 776
rect 110106 720 146666 776
rect 146722 720 146727 776
rect 110045 718 146727 720
rect 110045 715 110111 718
rect 146661 715 146727 718
rect 156413 778 156479 781
rect 160829 778 160895 781
rect 162301 778 162367 781
rect 156413 776 160895 778
rect 156413 720 156418 776
rect 156474 720 160834 776
rect 160890 720 160895 776
rect 156413 718 160895 720
rect 156413 715 156479 718
rect 160829 715 160895 718
rect 161430 776 162367 778
rect 161430 720 162306 776
rect 162362 720 162367 776
rect 161430 718 162367 720
rect 130561 642 130627 645
rect 161430 642 161490 718
rect 162301 715 162367 718
rect 162485 778 162551 781
rect 169109 778 169175 781
rect 162485 776 169175 778
rect 162485 720 162490 776
rect 162546 720 169114 776
rect 169170 720 169175 776
rect 162485 718 169175 720
rect 162485 715 162551 718
rect 169109 715 169175 718
rect 130561 640 161490 642
rect 130561 584 130566 640
rect 130622 584 161490 640
rect 130561 582 161490 584
rect 130561 579 130627 582
rect 161606 580 161612 644
rect 161676 642 161682 644
rect 166073 642 166139 645
rect 161676 640 166139 642
rect 161676 584 166078 640
rect 166134 584 166139 640
rect 161676 582 166139 584
rect 161676 580 161682 582
rect 166073 579 166139 582
rect 131941 506 132007 509
rect 162117 506 162183 509
rect 131941 504 162183 506
rect 131941 448 131946 504
rect 132002 448 162122 504
rect 162178 448 162183 504
rect 131941 446 162183 448
rect 131941 443 132007 446
rect 162117 443 162183 446
rect 163078 444 163084 508
rect 163148 506 163154 508
rect 163221 506 163287 509
rect 163148 504 163287 506
rect 163148 448 163226 504
rect 163282 448 163287 504
rect 163148 446 163287 448
rect 163148 444 163154 446
rect 163221 443 163287 446
rect 163446 444 163452 508
rect 163516 506 163522 508
rect 166901 506 166967 509
rect 163516 504 166967 506
rect 163516 448 166906 504
rect 166962 448 166967 504
rect 163516 446 166967 448
rect 163516 444 163522 446
rect 166901 443 166967 446
rect 127157 370 127223 373
rect 163313 370 163379 373
rect 127157 368 163379 370
rect 127157 312 127162 368
rect 127218 312 163318 368
rect 163374 312 163379 368
rect 127157 310 163379 312
rect 127157 307 127223 310
rect 163313 307 163379 310
rect 163681 370 163747 373
rect 170397 370 170463 373
rect 163681 368 170463 370
rect 163681 312 163686 368
rect 163742 312 170402 368
rect 170458 312 170463 368
rect 163681 310 170463 312
rect 163681 307 163747 310
rect 170397 307 170463 310
rect 98361 234 98427 237
rect 145046 234 145052 236
rect 98361 232 145052 234
rect 98361 176 98366 232
rect 98422 176 145052 232
rect 98361 174 145052 176
rect 98361 171 98427 174
rect 145046 172 145052 174
rect 145116 172 145122 236
rect 145189 234 145255 237
rect 154297 234 154363 237
rect 145189 232 154363 234
rect 145189 176 145194 232
rect 145250 176 154302 232
rect 154358 176 154363 232
rect 145189 174 154363 176
rect 145189 171 145255 174
rect 154297 171 154363 174
rect 155217 234 155283 237
rect 159265 234 159331 237
rect 155217 232 159331 234
rect 155217 176 155222 232
rect 155278 176 159270 232
rect 159326 176 159331 232
rect 155217 174 159331 176
rect 155217 171 155283 174
rect 159265 171 159331 174
rect 160645 234 160711 237
rect 161974 234 161980 236
rect 160645 232 161980 234
rect 160645 176 160650 232
rect 160706 176 161980 232
rect 160645 174 161980 176
rect 160645 171 160711 174
rect 161974 172 161980 174
rect 162044 172 162050 236
rect 162301 234 162367 237
rect 166574 234 166580 236
rect 162301 232 166580 234
rect 162301 176 162306 232
rect 162362 176 166580 232
rect 162301 174 166580 176
rect 162301 171 162367 174
rect 166574 172 166580 174
rect 166644 172 166650 236
rect 128353 98 128419 101
rect 132718 98 132724 100
rect 128353 96 132724 98
rect 128353 40 128358 96
rect 128414 40 132724 96
rect 128353 38 132724 40
rect 128353 35 128419 38
rect 132718 36 132724 38
rect 132788 36 132794 100
rect 132861 98 132927 101
rect 137645 98 137711 101
rect 132861 96 137711 98
rect 132861 40 132866 96
rect 132922 40 137650 96
rect 137706 40 137711 96
rect 132861 38 137711 40
rect 132861 35 132927 38
rect 137645 35 137711 38
rect 137870 36 137876 100
rect 137940 98 137946 100
rect 161790 98 161796 100
rect 137940 38 161796 98
rect 137940 36 137946 38
rect 161790 36 161796 38
rect 161860 36 161866 100
rect 162117 98 162183 101
rect 167126 98 167132 100
rect 162117 96 167132 98
rect 162117 40 162122 96
rect 162178 40 167132 96
rect 162117 38 167132 40
rect 162117 35 162183 38
rect 167126 36 167132 38
rect 167196 36 167202 100
rect -334 -344 -328 -280
rect -264 -282 -258 -280
rect 4066 -282 4072 -280
rect -264 -342 4072 -282
rect -264 -344 -258 -342
rect 4066 -344 4072 -342
rect 4136 -282 4142 -280
rect 44066 -282 44072 -280
rect 4136 -342 44072 -282
rect 4136 -344 4142 -342
rect 44066 -344 44072 -342
rect 44136 -282 44142 -280
rect 84066 -282 84072 -280
rect 44136 -342 84072 -282
rect 44136 -344 44142 -342
rect 84066 -344 84072 -342
rect 84136 -282 84142 -280
rect 124066 -282 124072 -280
rect 84136 -342 124072 -282
rect 84136 -344 84142 -342
rect 124066 -344 124072 -342
rect 124136 -282 124142 -280
rect 164066 -282 164072 -280
rect 124136 -342 164072 -282
rect 124136 -344 124142 -342
rect 164066 -344 164072 -342
rect 164136 -282 164142 -280
rect 200174 -282 200180 -280
rect 164136 -342 200180 -282
rect 164136 -344 164142 -342
rect 200174 -344 200180 -342
rect 200244 -344 200250 -280
rect -474 -484 -468 -420
rect -404 -422 -398 -420
rect 24066 -422 24072 -420
rect -404 -482 24072 -422
rect -404 -484 -398 -482
rect 24066 -484 24072 -482
rect 24136 -422 24142 -420
rect 64066 -422 64072 -420
rect 24136 -482 64072 -422
rect 24136 -484 24142 -482
rect 64066 -484 64072 -482
rect 64136 -422 64142 -420
rect 104066 -422 104072 -420
rect 64136 -482 104072 -422
rect 64136 -484 64142 -482
rect 104066 -484 104072 -482
rect 104136 -422 104142 -420
rect 144066 -422 144072 -420
rect 104136 -482 144072 -422
rect 104136 -484 104142 -482
rect 144066 -484 144072 -482
rect 144136 -422 144142 -420
rect 184066 -422 184072 -420
rect 144136 -482 184072 -422
rect 144136 -484 144142 -482
rect 184066 -484 184072 -482
rect 184136 -422 184142 -420
rect 200314 -422 200320 -420
rect 184136 -482 200320 -422
rect 184136 -484 184142 -482
rect 200314 -484 200320 -482
rect 200384 -484 200390 -420
rect -614 -624 -608 -560
rect -544 -562 -538 -560
rect 4466 -562 4472 -560
rect -544 -622 4472 -562
rect -544 -624 -538 -622
rect 4466 -624 4472 -622
rect 4536 -562 4542 -560
rect 44466 -562 44472 -560
rect 4536 -622 44472 -562
rect 4536 -624 4542 -622
rect 44466 -624 44472 -622
rect 44536 -562 44542 -560
rect 84466 -562 84472 -560
rect 44536 -622 84472 -562
rect 44536 -624 44542 -622
rect 84466 -624 84472 -622
rect 84536 -562 84542 -560
rect 124466 -562 124472 -560
rect 84536 -622 124472 -562
rect 84536 -624 84542 -622
rect 124466 -624 124472 -622
rect 124536 -562 124542 -560
rect 164466 -562 164472 -560
rect 124536 -622 164472 -562
rect 124536 -624 124542 -622
rect 164466 -624 164472 -622
rect 164536 -562 164542 -560
rect 200454 -562 200460 -560
rect 164536 -622 200460 -562
rect 164536 -624 164542 -622
rect 200454 -624 200460 -622
rect 200524 -624 200530 -560
rect -754 -764 -748 -700
rect -684 -702 -678 -700
rect 24466 -702 24472 -700
rect -684 -762 24472 -702
rect -684 -764 -678 -762
rect 24466 -764 24472 -762
rect 24536 -702 24542 -700
rect 64466 -702 64472 -700
rect 24536 -762 64472 -702
rect 24536 -764 24542 -762
rect 64466 -764 64472 -762
rect 64536 -702 64542 -700
rect 104466 -702 104472 -700
rect 64536 -762 104472 -702
rect 64536 -764 64542 -762
rect 104466 -764 104472 -762
rect 104536 -702 104542 -700
rect 144466 -702 144472 -700
rect 104536 -762 144472 -702
rect 104536 -764 104542 -762
rect 144466 -764 144472 -762
rect 144536 -702 144542 -700
rect 184466 -702 184472 -700
rect 144536 -762 184472 -702
rect 144536 -764 144542 -762
rect 184466 -764 184472 -762
rect 184536 -702 184542 -700
rect 200594 -702 200600 -700
rect 184536 -762 200600 -702
rect 184536 -764 184542 -762
rect 200594 -764 200600 -762
rect 200664 -764 200670 -700
rect -894 -904 -888 -840
rect -824 -842 -818 -840
rect 4866 -842 4872 -840
rect -824 -902 4872 -842
rect -824 -904 -818 -902
rect 4866 -904 4872 -902
rect 4936 -842 4942 -840
rect 44866 -842 44872 -840
rect 4936 -902 44872 -842
rect 4936 -904 4942 -902
rect 44866 -904 44872 -902
rect 44936 -842 44942 -840
rect 84866 -842 84872 -840
rect 44936 -902 84872 -842
rect 44936 -904 44942 -902
rect 84866 -904 84872 -902
rect 84936 -842 84942 -840
rect 124866 -842 124872 -840
rect 84936 -902 124872 -842
rect 84936 -904 84942 -902
rect 124866 -904 124872 -902
rect 124936 -842 124942 -840
rect 164866 -842 164872 -840
rect 124936 -902 164872 -842
rect 124936 -904 124942 -902
rect 164866 -904 164872 -902
rect 164936 -842 164942 -840
rect 200734 -842 200740 -840
rect 164936 -902 200740 -842
rect 164936 -904 164942 -902
rect 200734 -904 200740 -902
rect 200804 -904 200810 -840
rect -1034 -1044 -1028 -980
rect -964 -982 -958 -980
rect 24866 -982 24872 -980
rect -964 -1042 24872 -982
rect -964 -1044 -958 -1042
rect 24866 -1044 24872 -1042
rect 24936 -982 24942 -980
rect 64866 -982 64872 -980
rect 24936 -1042 64872 -982
rect 24936 -1044 24942 -1042
rect 64866 -1044 64872 -1042
rect 64936 -982 64942 -980
rect 104866 -982 104872 -980
rect 64936 -1042 104872 -982
rect 64936 -1044 64942 -1042
rect 104866 -1044 104872 -1042
rect 104936 -982 104942 -980
rect 144866 -982 144872 -980
rect 104936 -1042 144872 -982
rect 104936 -1044 104942 -1042
rect 144866 -1044 144872 -1042
rect 144936 -982 144942 -980
rect 184866 -982 184872 -980
rect 144936 -1042 184872 -982
rect 144936 -1044 144942 -1042
rect 184866 -1044 184872 -1042
rect 184936 -982 184942 -980
rect 200874 -982 200880 -980
rect 184936 -1042 200880 -982
rect 184936 -1044 184942 -1042
rect 200874 -1044 200880 -1042
rect 200944 -1044 200950 -980
rect -1174 -1184 -1168 -1120
rect -1104 -1122 -1098 -1120
rect 5266 -1122 5272 -1120
rect -1104 -1182 5272 -1122
rect -1104 -1184 -1098 -1182
rect 5266 -1184 5272 -1182
rect 5336 -1122 5342 -1120
rect 45266 -1122 45272 -1120
rect 5336 -1182 45272 -1122
rect 5336 -1184 5342 -1182
rect 45266 -1184 45272 -1182
rect 45336 -1122 45342 -1120
rect 85266 -1122 85272 -1120
rect 45336 -1182 85272 -1122
rect 45336 -1184 45342 -1182
rect 85266 -1184 85272 -1182
rect 85336 -1122 85342 -1120
rect 125266 -1122 125272 -1120
rect 85336 -1182 125272 -1122
rect 85336 -1184 85342 -1182
rect 125266 -1184 125272 -1182
rect 125336 -1122 125342 -1120
rect 165266 -1122 165272 -1120
rect 125336 -1182 165272 -1122
rect 125336 -1184 125342 -1182
rect 165266 -1184 165272 -1182
rect 165336 -1122 165342 -1120
rect 201014 -1122 201020 -1120
rect 165336 -1182 201020 -1122
rect 165336 -1184 165342 -1182
rect 201014 -1184 201020 -1182
rect 201084 -1184 201090 -1120
rect -1314 -1324 -1308 -1260
rect -1244 -1262 -1238 -1260
rect 25266 -1262 25272 -1260
rect -1244 -1322 25272 -1262
rect -1244 -1324 -1238 -1322
rect 25266 -1324 25272 -1322
rect 25336 -1262 25342 -1260
rect 65266 -1262 65272 -1260
rect 25336 -1322 65272 -1262
rect 25336 -1324 25342 -1322
rect 65266 -1324 65272 -1322
rect 65336 -1262 65342 -1260
rect 105266 -1262 105272 -1260
rect 65336 -1322 105272 -1262
rect 65336 -1324 65342 -1322
rect 105266 -1324 105272 -1322
rect 105336 -1262 105342 -1260
rect 145266 -1262 145272 -1260
rect 105336 -1322 145272 -1262
rect 105336 -1324 105342 -1322
rect 145266 -1324 145272 -1322
rect 145336 -1262 145342 -1260
rect 185266 -1262 185272 -1260
rect 145336 -1322 185272 -1262
rect 145336 -1324 145342 -1322
rect 185266 -1324 185272 -1322
rect 185336 -1262 185342 -1260
rect 201154 -1262 201160 -1260
rect 185336 -1322 201160 -1262
rect 185336 -1324 185342 -1322
rect 201154 -1324 201160 -1322
rect 201224 -1324 201230 -1260
rect -1454 -1464 -1448 -1400
rect -1384 -1402 -1378 -1400
rect 5666 -1402 5672 -1400
rect -1384 -1462 5672 -1402
rect -1384 -1464 -1378 -1462
rect 5666 -1464 5672 -1462
rect 5736 -1402 5742 -1400
rect 45666 -1402 45672 -1400
rect 5736 -1462 45672 -1402
rect 5736 -1464 5742 -1462
rect 45666 -1464 45672 -1462
rect 45736 -1402 45742 -1400
rect 85666 -1402 85672 -1400
rect 45736 -1462 85672 -1402
rect 45736 -1464 45742 -1462
rect 85666 -1464 85672 -1462
rect 85736 -1402 85742 -1400
rect 125666 -1402 125672 -1400
rect 85736 -1462 125672 -1402
rect 85736 -1464 85742 -1462
rect 125666 -1464 125672 -1462
rect 125736 -1402 125742 -1400
rect 165666 -1402 165672 -1400
rect 125736 -1462 165672 -1402
rect 125736 -1464 125742 -1462
rect 165666 -1464 165672 -1462
rect 165736 -1402 165742 -1400
rect 201294 -1402 201300 -1400
rect 165736 -1462 201300 -1402
rect 165736 -1464 165742 -1462
rect 201294 -1464 201300 -1462
rect 201364 -1464 201370 -1400
rect -1594 -1604 -1588 -1540
rect -1524 -1542 -1518 -1540
rect 25666 -1542 25672 -1540
rect -1524 -1602 25672 -1542
rect -1524 -1604 -1518 -1602
rect 25666 -1604 25672 -1602
rect 25736 -1542 25742 -1540
rect 65666 -1542 65672 -1540
rect 25736 -1602 65672 -1542
rect 25736 -1604 25742 -1602
rect 65666 -1604 65672 -1602
rect 65736 -1542 65742 -1540
rect 105666 -1542 105672 -1540
rect 65736 -1602 105672 -1542
rect 65736 -1604 65742 -1602
rect 105666 -1604 105672 -1602
rect 105736 -1542 105742 -1540
rect 145666 -1542 145672 -1540
rect 105736 -1602 145672 -1542
rect 105736 -1604 105742 -1602
rect 145666 -1604 145672 -1602
rect 145736 -1542 145742 -1540
rect 185666 -1542 185672 -1540
rect 145736 -1602 185672 -1542
rect 145736 -1604 145742 -1602
rect 185666 -1604 185672 -1602
rect 185736 -1542 185742 -1540
rect 201434 -1542 201440 -1540
rect 185736 -1602 201440 -1542
rect 185736 -1604 185742 -1602
rect 201434 -1604 201440 -1602
rect 201504 -1604 201510 -1540
<< via3 >>
rect -1588 12420 -1524 12484
rect 25672 12420 25736 12484
rect 65672 12420 65736 12484
rect 105672 12420 105736 12484
rect 145672 12420 145736 12484
rect 185672 12420 185736 12484
rect 201440 12420 201504 12484
rect -1448 12280 -1384 12344
rect 5672 12280 5736 12344
rect 45672 12280 45736 12344
rect 85672 12280 85736 12344
rect 125672 12280 125736 12344
rect 165672 12280 165736 12344
rect 201300 12280 201364 12344
rect -1308 12140 -1244 12204
rect 25272 12140 25336 12204
rect 65272 12140 65336 12204
rect 105272 12140 105336 12204
rect 145272 12140 145336 12204
rect 185272 12140 185336 12204
rect 201160 12140 201224 12204
rect -1168 12000 -1104 12064
rect 5272 12000 5336 12064
rect 45272 12000 45336 12064
rect 85272 12000 85336 12064
rect 125272 12000 125336 12064
rect 165272 12000 165336 12064
rect 201020 12000 201084 12064
rect -1028 11860 -964 11924
rect 24872 11860 24936 11924
rect 64872 11860 64936 11924
rect 104872 11860 104936 11924
rect 144872 11860 144936 11924
rect 184872 11860 184936 11924
rect 200880 11860 200944 11924
rect -888 11720 -824 11784
rect 4872 11720 4936 11784
rect 44872 11720 44936 11784
rect 84872 11720 84936 11784
rect 124872 11720 124936 11784
rect 164872 11720 164936 11784
rect 200740 11720 200804 11784
rect -748 11580 -684 11644
rect 24472 11580 24536 11644
rect 64472 11580 64536 11644
rect 104472 11580 104536 11644
rect 144472 11580 144536 11644
rect 184472 11580 184536 11644
rect 200600 11580 200664 11644
rect -608 11440 -544 11504
rect 4472 11440 4536 11504
rect 44472 11440 44536 11504
rect 84472 11440 84536 11504
rect 124472 11440 124536 11504
rect 164472 11440 164536 11504
rect 200460 11440 200524 11504
rect -468 11300 -404 11364
rect 24072 11300 24136 11364
rect 64072 11300 64136 11364
rect 104072 11300 104136 11364
rect 144072 11300 144136 11364
rect 184072 11300 184136 11364
rect 200320 11300 200384 11364
rect -328 11160 -264 11224
rect 4072 11160 4136 11224
rect 44072 11160 44136 11224
rect 84072 11160 84136 11224
rect 124072 11160 124136 11224
rect 164072 11160 164136 11224
rect 200180 11160 200244 11224
rect 4072 9820 4136 9824
rect 4072 9764 4076 9820
rect 4076 9764 4132 9820
rect 4132 9764 4136 9820
rect 4072 9760 4136 9764
rect 44072 9820 44136 9824
rect 44072 9764 44076 9820
rect 44076 9764 44132 9820
rect 44132 9764 44136 9820
rect 44072 9760 44136 9764
rect 84072 9820 84136 9824
rect 84072 9764 84076 9820
rect 84076 9764 84132 9820
rect 84132 9764 84136 9820
rect 84072 9760 84136 9764
rect 124072 9820 124136 9824
rect 124072 9764 124076 9820
rect 124076 9764 124132 9820
rect 124132 9764 124136 9820
rect 124072 9760 124136 9764
rect 164072 9820 164136 9824
rect 164072 9764 164076 9820
rect 164076 9764 164132 9820
rect 164132 9764 164136 9820
rect 164072 9760 164136 9764
rect 157380 9692 157444 9756
rect 24072 9276 24136 9280
rect 24072 9220 24076 9276
rect 24076 9220 24132 9276
rect 24132 9220 24136 9276
rect 24072 9216 24136 9220
rect 64072 9276 64136 9280
rect 64072 9220 64076 9276
rect 64076 9220 64132 9276
rect 64132 9220 64136 9276
rect 64072 9216 64136 9220
rect 104072 9276 104136 9280
rect 104072 9220 104076 9276
rect 104076 9220 104132 9276
rect 104132 9220 104136 9276
rect 104072 9216 104136 9220
rect 144072 9276 144136 9280
rect 144072 9220 144076 9276
rect 144076 9220 144132 9276
rect 144132 9220 144136 9276
rect 144072 9216 144136 9220
rect 184072 9276 184136 9280
rect 184072 9220 184076 9276
rect 184076 9220 184132 9276
rect 184132 9220 184136 9276
rect 184072 9216 184136 9220
rect 167868 9012 167932 9076
rect 173756 9072 173820 9076
rect 173756 9016 173770 9072
rect 173770 9016 173820 9072
rect 173756 9012 173820 9016
rect 168972 8876 169036 8940
rect 157748 8740 157812 8804
rect 4072 8732 4136 8736
rect 4072 8676 4076 8732
rect 4076 8676 4132 8732
rect 4132 8676 4136 8732
rect 4072 8672 4136 8676
rect 44072 8732 44136 8736
rect 44072 8676 44076 8732
rect 44076 8676 44132 8732
rect 44132 8676 44136 8732
rect 44072 8672 44136 8676
rect 84072 8732 84136 8736
rect 84072 8676 84076 8732
rect 84076 8676 84132 8732
rect 84132 8676 84136 8732
rect 84072 8672 84136 8676
rect 124072 8732 124136 8736
rect 124072 8676 124076 8732
rect 124076 8676 124132 8732
rect 124132 8676 124136 8732
rect 124072 8672 124136 8676
rect 164072 8732 164136 8736
rect 164072 8676 164076 8732
rect 164076 8676 164132 8732
rect 164132 8676 164136 8732
rect 164072 8672 164136 8676
rect 157564 8332 157628 8396
rect 165476 8332 165540 8396
rect 169524 8332 169588 8396
rect 170812 8392 170876 8396
rect 170812 8336 170826 8392
rect 170826 8336 170876 8392
rect 170812 8332 170876 8336
rect 175964 8332 176028 8396
rect 177620 8332 177684 8396
rect 24072 8188 24136 8192
rect 24072 8132 24076 8188
rect 24076 8132 24132 8188
rect 24132 8132 24136 8188
rect 24072 8128 24136 8132
rect 64072 8188 64136 8192
rect 64072 8132 64076 8188
rect 64076 8132 64132 8188
rect 64132 8132 64136 8188
rect 64072 8128 64136 8132
rect 104072 8188 104136 8192
rect 104072 8132 104076 8188
rect 104076 8132 104132 8188
rect 104132 8132 104136 8188
rect 104072 8128 104136 8132
rect 144072 8188 144136 8192
rect 144072 8132 144076 8188
rect 144076 8132 144132 8188
rect 144132 8132 144136 8188
rect 144072 8128 144136 8132
rect 161980 8060 162044 8124
rect 184072 8188 184136 8192
rect 184072 8132 184076 8188
rect 184076 8132 184132 8188
rect 184132 8132 184136 8188
rect 184072 8128 184136 8132
rect 157196 7652 157260 7716
rect 167132 7788 167196 7852
rect 167316 7788 167380 7852
rect 175596 7788 175660 7852
rect 4072 7644 4136 7648
rect 4072 7588 4076 7644
rect 4076 7588 4132 7644
rect 4132 7588 4136 7644
rect 4072 7584 4136 7588
rect 44072 7644 44136 7648
rect 44072 7588 44076 7644
rect 44076 7588 44132 7644
rect 44132 7588 44136 7644
rect 44072 7584 44136 7588
rect 84072 7644 84136 7648
rect 84072 7588 84076 7644
rect 84076 7588 84132 7644
rect 84132 7588 84136 7644
rect 84072 7584 84136 7588
rect 124072 7644 124136 7648
rect 124072 7588 124076 7644
rect 124076 7588 124132 7644
rect 124132 7588 124136 7644
rect 124072 7584 124136 7588
rect 183508 7712 183572 7716
rect 183508 7656 183558 7712
rect 183558 7656 183572 7712
rect 183508 7652 183572 7656
rect 164072 7644 164136 7648
rect 164072 7588 164076 7644
rect 164076 7588 164132 7644
rect 164132 7588 164136 7644
rect 164072 7584 164136 7588
rect 165108 7516 165172 7580
rect 166028 7516 166092 7580
rect 157012 7380 157076 7444
rect 158668 7380 158732 7444
rect 158852 7440 158916 7444
rect 158852 7384 158902 7440
rect 158902 7384 158916 7440
rect 158852 7380 158916 7384
rect 159956 7440 160020 7444
rect 159956 7384 159970 7440
rect 159970 7384 160020 7440
rect 159956 7380 160020 7384
rect 161428 7380 161492 7444
rect 164740 7440 164804 7444
rect 164740 7384 164754 7440
rect 164754 7384 164804 7440
rect 164740 7380 164804 7384
rect 165844 7380 165908 7444
rect 124260 7244 124324 7308
rect 157380 7244 157444 7308
rect 175044 7516 175108 7580
rect 176516 7576 176580 7580
rect 176516 7520 176530 7576
rect 176530 7520 176580 7576
rect 176516 7516 176580 7520
rect 167684 7440 167748 7444
rect 167684 7384 167734 7440
rect 167734 7384 167748 7440
rect 167684 7380 167748 7384
rect 169708 7440 169772 7444
rect 169708 7384 169758 7440
rect 169758 7384 169772 7440
rect 169708 7380 169772 7384
rect 170076 7440 170140 7444
rect 170076 7384 170090 7440
rect 170090 7384 170140 7440
rect 170076 7380 170140 7384
rect 171180 7440 171244 7444
rect 171180 7384 171230 7440
rect 171230 7384 171244 7440
rect 171180 7380 171244 7384
rect 171364 7440 171428 7444
rect 171364 7384 171414 7440
rect 171414 7384 171428 7440
rect 171364 7380 171428 7384
rect 171732 7440 171796 7444
rect 171732 7384 171782 7440
rect 171782 7384 171796 7440
rect 171732 7380 171796 7384
rect 172468 7380 172532 7444
rect 173388 7380 173452 7444
rect 174860 7440 174924 7444
rect 174860 7384 174910 7440
rect 174910 7384 174924 7440
rect 174860 7380 174924 7384
rect 175780 7380 175844 7444
rect 177068 7380 177132 7444
rect 180748 7380 180812 7444
rect 182036 7440 182100 7444
rect 182036 7384 182050 7440
rect 182050 7384 182100 7440
rect 182036 7380 182100 7384
rect 182220 7440 182284 7444
rect 182220 7384 182270 7440
rect 182270 7384 182284 7440
rect 182220 7380 182284 7384
rect 182404 7380 182468 7444
rect 177804 7304 177868 7308
rect 177804 7248 177854 7304
rect 177854 7248 177868 7304
rect 177804 7244 177868 7248
rect 24072 7100 24136 7104
rect 24072 7044 24076 7100
rect 24076 7044 24132 7100
rect 24132 7044 24136 7100
rect 24072 7040 24136 7044
rect 64072 7100 64136 7104
rect 64072 7044 64076 7100
rect 64076 7044 64132 7100
rect 64132 7044 64136 7100
rect 64072 7040 64136 7044
rect 104072 7100 104136 7104
rect 104072 7044 104076 7100
rect 104076 7044 104132 7100
rect 104132 7044 104136 7100
rect 104072 7040 104136 7044
rect 144072 7100 144136 7104
rect 144072 7044 144076 7100
rect 144076 7044 144132 7100
rect 144132 7044 144136 7100
rect 144072 7040 144136 7044
rect 124214 6700 124278 6764
rect 134748 6700 134812 6764
rect 168052 7108 168116 7172
rect 158668 6972 158732 7036
rect 182404 6972 182468 7036
rect 4072 6556 4136 6560
rect 4072 6500 4076 6556
rect 4076 6500 4132 6556
rect 4132 6500 4136 6556
rect 4072 6496 4136 6500
rect 44072 6556 44136 6560
rect 44072 6500 44076 6556
rect 44076 6500 44132 6556
rect 44132 6500 44136 6556
rect 44072 6496 44136 6500
rect 84072 6556 84136 6560
rect 84072 6500 84076 6556
rect 84076 6500 84132 6556
rect 84132 6500 84136 6556
rect 84072 6496 84136 6500
rect 124072 6556 124136 6560
rect 124072 6500 124076 6556
rect 124076 6500 124132 6556
rect 124132 6500 124136 6556
rect 124072 6496 124136 6500
rect 135116 6428 135180 6492
rect 124260 6156 124324 6220
rect 185672 6803 185736 6867
rect 164472 6680 164536 6744
rect 185272 6403 185336 6467
rect 165672 6074 165736 6138
rect 24072 6012 24136 6016
rect 24072 5956 24076 6012
rect 24076 5956 24132 6012
rect 24132 5956 24136 6012
rect 24072 5952 24136 5956
rect 64072 6012 64136 6016
rect 64072 5956 64076 6012
rect 64076 5956 64132 6012
rect 64132 5956 64136 6012
rect 64072 5952 64136 5956
rect 104072 6012 104136 6016
rect 104072 5956 104076 6012
rect 104076 5956 104132 6012
rect 104132 5956 104136 6012
rect 104072 5952 104136 5956
rect 144072 6012 144136 6016
rect 144072 5956 144076 6012
rect 144076 5956 144132 6012
rect 144132 5956 144136 6012
rect 144072 5952 144136 5956
rect 184472 5952 184536 6016
rect 165272 5674 165336 5738
rect 4072 5468 4136 5472
rect 4072 5412 4076 5468
rect 4076 5412 4132 5468
rect 4132 5412 4136 5468
rect 4072 5408 4136 5412
rect 44072 5468 44136 5472
rect 44072 5412 44076 5468
rect 44076 5412 44132 5468
rect 44132 5412 44136 5468
rect 44072 5408 44136 5412
rect 84072 5468 84136 5472
rect 84072 5412 84076 5468
rect 84076 5412 84132 5468
rect 84132 5412 84136 5468
rect 84072 5408 84136 5412
rect 124072 5468 124136 5472
rect 124072 5412 124076 5468
rect 124076 5412 124132 5468
rect 124132 5412 124136 5468
rect 124072 5408 124136 5412
rect 124260 5340 124324 5404
rect 157012 5340 157076 5404
rect 185672 5345 185736 5409
rect 164472 5223 164536 5287
rect 157012 4932 157076 4996
rect 185272 4945 185336 5009
rect 24072 4924 24136 4928
rect 24072 4868 24076 4924
rect 24076 4868 24132 4924
rect 24132 4868 24136 4924
rect 24072 4864 24136 4868
rect 64072 4924 64136 4928
rect 64072 4868 64076 4924
rect 64076 4868 64132 4924
rect 64132 4868 64136 4924
rect 64072 4864 64136 4868
rect 104072 4924 104136 4928
rect 104072 4868 104076 4924
rect 104076 4868 104132 4924
rect 104132 4868 104136 4924
rect 104072 4864 104136 4868
rect 144072 4924 144136 4928
rect 144072 4868 144076 4924
rect 144076 4868 144132 4924
rect 144132 4868 144136 4924
rect 144072 4864 144136 4868
rect 4072 4380 4136 4384
rect 4072 4324 4076 4380
rect 4076 4324 4132 4380
rect 4132 4324 4136 4380
rect 4072 4320 4136 4324
rect 44072 4380 44136 4384
rect 44072 4324 44076 4380
rect 44076 4324 44132 4380
rect 44132 4324 44136 4380
rect 44072 4320 44136 4324
rect 84072 4380 84136 4384
rect 84072 4324 84076 4380
rect 84076 4324 84132 4380
rect 84132 4324 84136 4380
rect 84072 4320 84136 4324
rect 124072 4380 124136 4384
rect 124072 4324 124076 4380
rect 124076 4324 124132 4380
rect 124132 4324 124136 4380
rect 124072 4320 124136 4324
rect 165672 4617 165736 4681
rect 157196 4524 157260 4588
rect 184472 4494 184536 4558
rect 145052 4252 145116 4316
rect 165272 4217 165336 4281
rect 24072 3836 24136 3840
rect 24072 3780 24076 3836
rect 24076 3780 24132 3836
rect 24132 3780 24136 3836
rect 24072 3776 24136 3780
rect 64072 3836 64136 3840
rect 64072 3780 64076 3836
rect 64076 3780 64132 3836
rect 64132 3780 64136 3836
rect 64072 3776 64136 3780
rect 104072 3836 104136 3840
rect 104072 3780 104076 3836
rect 104076 3780 104132 3836
rect 104132 3780 104136 3836
rect 104072 3776 104136 3780
rect 144072 3836 144136 3840
rect 144072 3780 144076 3836
rect 144076 3780 144132 3836
rect 144132 3780 144136 3836
rect 144072 3776 144136 3780
rect 164472 3766 164536 3830
rect 157380 3572 157444 3636
rect 172468 3572 172532 3636
rect 161612 3436 161676 3500
rect 161796 3436 161860 3500
rect 167316 3436 167380 3500
rect 167500 3436 167564 3500
rect 176332 3436 176396 3500
rect 137324 3300 137388 3364
rect 4072 3292 4136 3296
rect 4072 3236 4076 3292
rect 4076 3236 4132 3292
rect 4132 3236 4136 3292
rect 4072 3232 4136 3236
rect 44072 3292 44136 3296
rect 44072 3236 44076 3292
rect 44076 3236 44132 3292
rect 44132 3236 44136 3292
rect 44072 3232 44136 3236
rect 84072 3292 84136 3296
rect 84072 3236 84076 3292
rect 84076 3236 84132 3292
rect 84132 3236 84136 3292
rect 84072 3232 84136 3236
rect 124072 3292 124136 3296
rect 124072 3236 124076 3292
rect 124076 3236 124132 3292
rect 124132 3236 124136 3292
rect 124072 3232 124136 3236
rect 163084 3300 163148 3364
rect 157012 3164 157076 3228
rect 137692 3028 137756 3092
rect 151860 3028 151924 3092
rect 162900 3164 162964 3228
rect 164740 3164 164804 3228
rect 166764 3164 166828 3228
rect 157380 3028 157444 3092
rect 161796 3028 161860 3092
rect 161980 3028 162044 3092
rect 168972 3028 169036 3092
rect 169892 3164 169956 3228
rect 24072 2748 24136 2752
rect 24072 2692 24076 2748
rect 24076 2692 24132 2748
rect 24132 2692 24136 2748
rect 24072 2688 24136 2692
rect 64072 2748 64136 2752
rect 64072 2692 64076 2748
rect 64076 2692 64132 2748
rect 64132 2692 64136 2748
rect 64072 2688 64136 2692
rect 104072 2748 104136 2752
rect 104072 2692 104076 2748
rect 104076 2692 104132 2748
rect 104132 2692 104136 2748
rect 104072 2688 104136 2692
rect 138428 2620 138492 2684
rect 144072 2748 144136 2752
rect 144072 2692 144076 2748
rect 144076 2692 144132 2748
rect 144132 2692 144136 2748
rect 144072 2688 144136 2692
rect 162348 2892 162412 2956
rect 165476 2952 165540 2956
rect 165476 2896 165526 2952
rect 165526 2896 165540 2952
rect 165476 2892 165540 2896
rect 168052 2892 168116 2956
rect 169708 2952 169772 2956
rect 169708 2896 169758 2952
rect 169758 2896 169772 2952
rect 169708 2892 169772 2896
rect 170076 2952 170140 2956
rect 170076 2896 170090 2952
rect 170090 2896 170140 2952
rect 170076 2892 170140 2896
rect 171732 2952 171796 2956
rect 171732 2896 171746 2952
rect 171746 2896 171796 2952
rect 171732 2892 171796 2896
rect 174860 2952 174924 2956
rect 174860 2896 174910 2952
rect 174910 2896 174924 2952
rect 174860 2892 174924 2896
rect 175964 2952 176028 2956
rect 175964 2896 175978 2952
rect 175978 2896 176028 2952
rect 175964 2892 176028 2896
rect 177068 2892 177132 2956
rect 177804 2952 177868 2956
rect 177804 2896 177854 2952
rect 177854 2896 177868 2952
rect 177804 2892 177868 2896
rect 4072 2204 4136 2208
rect 4072 2148 4076 2204
rect 4076 2148 4132 2204
rect 4132 2148 4136 2204
rect 4072 2144 4136 2148
rect 44072 2204 44136 2208
rect 44072 2148 44076 2204
rect 44076 2148 44132 2204
rect 44132 2148 44136 2204
rect 44072 2144 44136 2148
rect 84072 2204 84136 2208
rect 84072 2148 84076 2204
rect 84076 2148 84132 2204
rect 84132 2148 84136 2204
rect 84072 2144 84136 2148
rect 161980 2620 162044 2684
rect 164740 2756 164804 2820
rect 165108 2756 165172 2820
rect 166580 2756 166644 2820
rect 167868 2756 167932 2820
rect 162900 2620 162964 2684
rect 166028 2620 166092 2684
rect 167500 2620 167564 2684
rect 167684 2680 167748 2684
rect 169892 2756 169956 2820
rect 171364 2756 171428 2820
rect 173388 2756 173452 2820
rect 173756 2756 173820 2820
rect 176516 2816 176580 2820
rect 176516 2760 176566 2816
rect 176566 2760 176580 2816
rect 176516 2756 176580 2760
rect 184072 2748 184136 2752
rect 184072 2692 184076 2748
rect 184076 2692 184132 2748
rect 184132 2692 184136 2748
rect 184072 2688 184136 2692
rect 167684 2624 167734 2680
rect 167734 2624 167748 2680
rect 167684 2620 167748 2624
rect 171180 2680 171244 2684
rect 171180 2624 171194 2680
rect 171194 2624 171244 2680
rect 171180 2620 171244 2624
rect 180748 2484 180812 2548
rect 138060 2212 138124 2276
rect 138244 2212 138308 2276
rect 124072 2204 124136 2208
rect 124072 2148 124076 2204
rect 124076 2148 124132 2204
rect 124132 2148 124136 2204
rect 124072 2144 124136 2148
rect 137876 2076 137940 2140
rect 158852 1940 158916 2004
rect 161428 2076 161492 2140
rect 171916 2348 171980 2412
rect 175780 2348 175844 2412
rect 169524 2212 169588 2276
rect 170812 2212 170876 2276
rect 176332 2212 176396 2276
rect 164072 2204 164136 2208
rect 164072 2148 164076 2204
rect 164076 2148 164132 2204
rect 164132 2148 164136 2204
rect 164072 2144 164136 2148
rect 165844 2076 165908 2140
rect 182036 2136 182100 2140
rect 182036 2080 182050 2136
rect 182050 2080 182100 2136
rect 182036 2076 182100 2080
rect 165108 1804 165172 1868
rect 138060 1668 138124 1732
rect 175596 1668 175660 1732
rect 24072 1660 24136 1664
rect 24072 1604 24076 1660
rect 24076 1604 24132 1660
rect 24132 1604 24136 1660
rect 24072 1600 24136 1604
rect 64072 1660 64136 1664
rect 64072 1604 64076 1660
rect 64076 1604 64132 1660
rect 64132 1604 64136 1660
rect 64072 1600 64136 1604
rect 104072 1660 104136 1664
rect 104072 1604 104076 1660
rect 104076 1604 104132 1660
rect 104132 1604 104136 1660
rect 104072 1600 104136 1604
rect 144072 1660 144136 1664
rect 144072 1604 144076 1660
rect 144076 1604 144132 1660
rect 144132 1604 144136 1660
rect 144072 1600 144136 1604
rect 184072 1660 184136 1664
rect 184072 1604 184076 1660
rect 184076 1604 184132 1660
rect 184132 1604 184136 1660
rect 184072 1600 184136 1604
rect 159956 1532 160020 1596
rect 177620 1532 177684 1596
rect 183508 1592 183572 1596
rect 183508 1536 183558 1592
rect 183558 1536 183572 1592
rect 183508 1532 183572 1536
rect 164740 1456 164804 1460
rect 164740 1400 164754 1456
rect 164754 1400 164804 1456
rect 164740 1396 164804 1400
rect 165108 1396 165172 1460
rect 166764 1396 166828 1460
rect 170996 1396 171060 1460
rect 137692 1124 137756 1188
rect 137876 1124 137940 1188
rect 162348 1124 162412 1188
rect 182220 1260 182284 1324
rect 175228 1124 175292 1188
rect 4072 1116 4136 1120
rect 4072 1060 4076 1116
rect 4076 1060 4132 1116
rect 4132 1060 4136 1116
rect 4072 1056 4136 1060
rect 44072 1116 44136 1120
rect 44072 1060 44076 1116
rect 44076 1060 44132 1116
rect 44132 1060 44136 1116
rect 44072 1056 44136 1060
rect 84072 1116 84136 1120
rect 84072 1060 84076 1116
rect 84076 1060 84132 1116
rect 84132 1060 84136 1116
rect 84072 1056 84136 1060
rect 124072 1116 124136 1120
rect 124072 1060 124076 1116
rect 124076 1060 124132 1116
rect 124132 1060 124136 1116
rect 124072 1056 124136 1060
rect 164072 1116 164136 1120
rect 164072 1060 164076 1116
rect 164076 1060 164132 1116
rect 164132 1060 164136 1116
rect 164072 1056 164136 1060
rect 137140 988 137204 1052
rect 151860 988 151924 1052
rect 161612 580 161676 644
rect 163084 444 163148 508
rect 163452 444 163516 508
rect 145052 172 145116 236
rect 161980 172 162044 236
rect 166580 172 166644 236
rect 132724 36 132788 100
rect 137876 36 137940 100
rect 161796 36 161860 100
rect 167132 36 167196 100
rect -328 -344 -264 -280
rect 4072 -344 4136 -280
rect 44072 -344 44136 -280
rect 84072 -344 84136 -280
rect 124072 -344 124136 -280
rect 164072 -344 164136 -280
rect 200180 -344 200244 -280
rect -468 -484 -404 -420
rect 24072 -484 24136 -420
rect 64072 -484 64136 -420
rect 104072 -484 104136 -420
rect 144072 -484 144136 -420
rect 184072 -484 184136 -420
rect 200320 -484 200384 -420
rect -608 -624 -544 -560
rect 4472 -624 4536 -560
rect 44472 -624 44536 -560
rect 84472 -624 84536 -560
rect 124472 -624 124536 -560
rect 164472 -624 164536 -560
rect 200460 -624 200524 -560
rect -748 -764 -684 -700
rect 24472 -764 24536 -700
rect 64472 -764 64536 -700
rect 104472 -764 104536 -700
rect 144472 -764 144536 -700
rect 184472 -764 184536 -700
rect 200600 -764 200664 -700
rect -888 -904 -824 -840
rect 4872 -904 4936 -840
rect 44872 -904 44936 -840
rect 84872 -904 84936 -840
rect 124872 -904 124936 -840
rect 164872 -904 164936 -840
rect 200740 -904 200804 -840
rect -1028 -1044 -964 -980
rect 24872 -1044 24936 -980
rect 64872 -1044 64936 -980
rect 104872 -1044 104936 -980
rect 144872 -1044 144936 -980
rect 184872 -1044 184936 -980
rect 200880 -1044 200944 -980
rect -1168 -1184 -1104 -1120
rect 5272 -1184 5336 -1120
rect 45272 -1184 45336 -1120
rect 85272 -1184 85336 -1120
rect 125272 -1184 125336 -1120
rect 165272 -1184 165336 -1120
rect 201020 -1184 201084 -1120
rect -1308 -1324 -1244 -1260
rect 25272 -1324 25336 -1260
rect 65272 -1324 65336 -1260
rect 105272 -1324 105336 -1260
rect 145272 -1324 145336 -1260
rect 185272 -1324 185336 -1260
rect 201160 -1324 201224 -1260
rect -1448 -1464 -1384 -1400
rect 5672 -1464 5736 -1400
rect 45672 -1464 45736 -1400
rect 85672 -1464 85736 -1400
rect 125672 -1464 125736 -1400
rect 165672 -1464 165736 -1400
rect 201300 -1464 201364 -1400
rect -1588 -1604 -1524 -1540
rect 25672 -1604 25736 -1540
rect 65672 -1604 65736 -1540
rect 105672 -1604 105736 -1540
rect 145672 -1604 145736 -1540
rect 185672 -1604 185736 -1540
rect 201440 -1604 201504 -1540
<< metal4 >>
rect -1589 12484 -1523 12485
rect -1589 12420 -1588 12484
rect -1524 12420 -1523 12484
rect 25671 12484 25737 12485
rect -1589 12419 -1523 12420
rect -1586 -1539 -1526 12419
rect 5674 12345 5734 12482
rect 25671 12420 25672 12484
rect 25736 12420 25737 12484
rect 65671 12484 65737 12485
rect 25671 12419 25737 12420
rect -1449 12344 -1383 12345
rect -1449 12280 -1448 12344
rect -1384 12280 -1383 12344
rect -1449 12279 -1383 12280
rect 5671 12344 5737 12345
rect 5671 12280 5672 12344
rect 5736 12280 5737 12344
rect 5671 12279 5737 12280
rect -1446 -1399 -1386 12279
rect -1309 12204 -1243 12205
rect -1309 12140 -1308 12204
rect -1244 12140 -1243 12204
rect -1309 12139 -1243 12140
rect -1306 -1259 -1246 12139
rect 5274 12065 5334 12202
rect -1169 12064 -1103 12065
rect -1169 12000 -1168 12064
rect -1104 12000 -1103 12064
rect -1169 11999 -1103 12000
rect 5271 12064 5337 12065
rect 5271 12000 5272 12064
rect 5336 12000 5337 12064
rect 5271 11999 5337 12000
rect -1166 -1119 -1106 11999
rect -1029 11924 -963 11925
rect -1029 11860 -1028 11924
rect -964 11860 -963 11924
rect -1029 11859 -963 11860
rect -1026 -979 -966 11859
rect 4874 11785 4934 11922
rect -889 11784 -823 11785
rect -889 11720 -888 11784
rect -824 11720 -823 11784
rect -889 11719 -823 11720
rect 4871 11784 4937 11785
rect 4871 11720 4872 11784
rect 4936 11720 4937 11784
rect 4871 11719 4937 11720
rect -886 -839 -826 11719
rect -749 11644 -683 11645
rect -749 11580 -748 11644
rect -684 11580 -683 11644
rect -749 11579 -683 11580
rect -746 -699 -686 11579
rect 4474 11505 4534 11642
rect -609 11504 -543 11505
rect -609 11440 -608 11504
rect -544 11440 -543 11504
rect -609 11439 -543 11440
rect 4471 11504 4537 11505
rect 4471 11440 4472 11504
rect 4536 11440 4537 11504
rect 4471 11439 4537 11440
rect -606 -559 -546 11439
rect -469 11364 -403 11365
rect -469 11300 -468 11364
rect -404 11300 -403 11364
rect -469 11299 -403 11300
rect -466 -419 -406 11299
rect 4074 11225 4134 11362
rect -329 11224 -263 11225
rect -329 11160 -328 11224
rect -264 11160 -263 11224
rect -329 11159 -263 11160
rect 4071 11224 4137 11225
rect 4071 11160 4072 11224
rect 4136 11160 4137 11224
rect 4071 11159 4137 11160
rect -326 -279 -266 11159
rect 4074 9840 4134 11159
rect 4071 9824 4137 9840
rect 4071 9760 4072 9824
rect 4136 9760 4137 9824
rect 4071 9744 4137 9760
rect 4074 8752 4134 9744
rect 4071 8736 4137 8752
rect 4071 8672 4072 8736
rect 4136 8672 4137 8736
rect 4071 8656 4137 8672
rect 4074 7664 4134 8656
rect 4071 7648 4137 7664
rect 4071 7584 4072 7648
rect 4136 7584 4137 7648
rect 4071 7568 4137 7584
rect 4074 6576 4134 7568
rect 4071 6560 4137 6576
rect 4071 6496 4072 6560
rect 4136 6496 4137 6560
rect 4071 6480 4137 6496
rect 4074 5488 4134 6480
rect 4071 5472 4137 5488
rect 4071 5408 4072 5472
rect 4136 5408 4137 5472
rect 4071 5392 4137 5408
rect 4074 4400 4134 5392
rect 4071 4384 4137 4400
rect 4071 4320 4072 4384
rect 4136 4320 4137 4384
rect 4071 4304 4137 4320
rect 4074 3312 4134 4304
rect 4071 3296 4137 3312
rect 4071 3232 4072 3296
rect 4136 3232 4137 3296
rect 4071 3216 4137 3232
rect 4074 2224 4134 3216
rect 4071 2208 4137 2224
rect 4071 2144 4072 2208
rect 4136 2144 4137 2208
rect 4071 2128 4137 2144
rect 4074 1136 4134 2128
rect 4071 1120 4137 1136
rect 4071 1056 4072 1120
rect 4136 1056 4137 1120
rect 4071 1040 4137 1056
rect 4074 -279 4134 1040
rect -329 -280 -263 -279
rect -329 -344 -328 -280
rect -264 -344 -263 -280
rect -329 -345 -263 -344
rect 4071 -280 4137 -279
rect 4071 -344 4072 -280
rect 4136 -344 4137 -280
rect 4071 -345 4137 -344
rect -469 -420 -403 -419
rect -469 -484 -468 -420
rect -404 -484 -403 -420
rect 4074 -482 4134 -345
rect -469 -485 -403 -484
rect 4474 -559 4534 11439
rect -609 -560 -543 -559
rect -609 -624 -608 -560
rect -544 -624 -543 -560
rect -609 -625 -543 -624
rect 4471 -560 4537 -559
rect 4471 -624 4472 -560
rect 4536 -624 4537 -560
rect 4471 -625 4537 -624
rect -749 -700 -683 -699
rect -749 -764 -748 -700
rect -684 -764 -683 -700
rect 4474 -762 4534 -625
rect -749 -765 -683 -764
rect 4874 -839 4934 11719
rect -889 -840 -823 -839
rect -889 -904 -888 -840
rect -824 -904 -823 -840
rect -889 -905 -823 -904
rect 4871 -840 4937 -839
rect 4871 -904 4872 -840
rect 4936 -904 4937 -840
rect 4871 -905 4937 -904
rect -1029 -980 -963 -979
rect -1029 -1044 -1028 -980
rect -964 -1044 -963 -980
rect 4874 -1042 4934 -905
rect -1029 -1045 -963 -1044
rect 5274 -1119 5334 11999
rect -1169 -1120 -1103 -1119
rect -1169 -1184 -1168 -1120
rect -1104 -1184 -1103 -1120
rect -1169 -1185 -1103 -1184
rect 5271 -1120 5337 -1119
rect 5271 -1184 5272 -1120
rect 5336 -1184 5337 -1120
rect 5271 -1185 5337 -1184
rect -1309 -1260 -1243 -1259
rect -1309 -1324 -1308 -1260
rect -1244 -1324 -1243 -1260
rect 5274 -1322 5334 -1185
rect -1309 -1325 -1243 -1324
rect 5674 -1399 5734 12279
rect 25271 12204 25337 12205
rect 25271 12140 25272 12204
rect 25336 12140 25337 12204
rect 25271 12139 25337 12140
rect 24871 11924 24937 11925
rect 24871 11860 24872 11924
rect 24936 11860 24937 11924
rect 24871 11859 24937 11860
rect 24471 11644 24537 11645
rect 24471 11580 24472 11644
rect 24536 11580 24537 11644
rect 24471 11579 24537 11580
rect 24071 11364 24137 11365
rect 24071 11300 24072 11364
rect 24136 11300 24137 11364
rect 24071 11299 24137 11300
rect 24074 9296 24134 11299
rect 24071 9280 24137 9296
rect 24071 9216 24072 9280
rect 24136 9216 24137 9280
rect 24071 9200 24137 9216
rect 24074 8208 24134 9200
rect 24071 8192 24137 8208
rect 24071 8128 24072 8192
rect 24136 8128 24137 8192
rect 24071 8112 24137 8128
rect 24074 7120 24134 8112
rect 24071 7104 24137 7120
rect 24071 7040 24072 7104
rect 24136 7040 24137 7104
rect 24071 7024 24137 7040
rect 24074 6032 24134 7024
rect 24071 6016 24137 6032
rect 24071 5952 24072 6016
rect 24136 5952 24137 6016
rect 24071 5936 24137 5952
rect 24074 4944 24134 5936
rect 24071 4928 24137 4944
rect 24071 4864 24072 4928
rect 24136 4864 24137 4928
rect 24071 4848 24137 4864
rect 24074 3856 24134 4848
rect 24071 3840 24137 3856
rect 24071 3776 24072 3840
rect 24136 3776 24137 3840
rect 24071 3760 24137 3776
rect 24074 2768 24134 3760
rect 24071 2752 24137 2768
rect 24071 2688 24072 2752
rect 24136 2688 24137 2752
rect 24071 2672 24137 2688
rect 24074 1680 24134 2672
rect 24071 1664 24137 1680
rect 24071 1600 24072 1664
rect 24136 1600 24137 1664
rect 24071 1584 24137 1600
rect 24074 -419 24134 1584
rect 24071 -420 24137 -419
rect 24071 -484 24072 -420
rect 24136 -484 24137 -420
rect 24071 -485 24137 -484
rect 24474 -699 24534 11579
rect 24471 -700 24537 -699
rect 24471 -764 24472 -700
rect 24536 -764 24537 -700
rect 24471 -765 24537 -764
rect 24874 -979 24934 11859
rect 24871 -980 24937 -979
rect 24871 -1044 24872 -980
rect 24936 -1044 24937 -980
rect 24871 -1045 24937 -1044
rect 25274 -1259 25334 12139
rect 25271 -1260 25337 -1259
rect 25271 -1324 25272 -1260
rect 25336 -1324 25337 -1260
rect 25271 -1325 25337 -1324
rect -1449 -1400 -1383 -1399
rect -1449 -1464 -1448 -1400
rect -1384 -1464 -1383 -1400
rect -1449 -1465 -1383 -1464
rect 5671 -1400 5737 -1399
rect 5671 -1464 5672 -1400
rect 5736 -1464 5737 -1400
rect 5671 -1465 5737 -1464
rect -1589 -1540 -1523 -1539
rect -1589 -1604 -1588 -1540
rect -1524 -1604 -1523 -1540
rect 5674 -1602 5734 -1465
rect 25674 -1539 25734 12419
rect 45674 12345 45734 12482
rect 65671 12420 65672 12484
rect 65736 12420 65737 12484
rect 105671 12484 105737 12485
rect 65671 12419 65737 12420
rect 45671 12344 45737 12345
rect 45671 12280 45672 12344
rect 45736 12280 45737 12344
rect 45671 12279 45737 12280
rect 45274 12065 45334 12202
rect 45271 12064 45337 12065
rect 45271 12000 45272 12064
rect 45336 12000 45337 12064
rect 45271 11999 45337 12000
rect 44874 11785 44934 11922
rect 44871 11784 44937 11785
rect 44871 11720 44872 11784
rect 44936 11720 44937 11784
rect 44871 11719 44937 11720
rect 44474 11505 44534 11642
rect 44471 11504 44537 11505
rect 44471 11440 44472 11504
rect 44536 11440 44537 11504
rect 44471 11439 44537 11440
rect 44074 11225 44134 11362
rect 44071 11224 44137 11225
rect 44071 11160 44072 11224
rect 44136 11160 44137 11224
rect 44071 11159 44137 11160
rect 44074 9840 44134 11159
rect 44071 9824 44137 9840
rect 44071 9760 44072 9824
rect 44136 9760 44137 9824
rect 44071 9744 44137 9760
rect 44074 8752 44134 9744
rect 44071 8736 44137 8752
rect 44071 8672 44072 8736
rect 44136 8672 44137 8736
rect 44071 8656 44137 8672
rect 44074 7664 44134 8656
rect 44071 7648 44137 7664
rect 44071 7584 44072 7648
rect 44136 7584 44137 7648
rect 44071 7568 44137 7584
rect 44074 6576 44134 7568
rect 44071 6560 44137 6576
rect 44071 6496 44072 6560
rect 44136 6496 44137 6560
rect 44071 6480 44137 6496
rect 44074 5488 44134 6480
rect 44071 5472 44137 5488
rect 44071 5408 44072 5472
rect 44136 5408 44137 5472
rect 44071 5392 44137 5408
rect 44074 4400 44134 5392
rect 44071 4384 44137 4400
rect 44071 4320 44072 4384
rect 44136 4320 44137 4384
rect 44071 4304 44137 4320
rect 44074 3312 44134 4304
rect 44071 3296 44137 3312
rect 44071 3232 44072 3296
rect 44136 3232 44137 3296
rect 44071 3216 44137 3232
rect 44074 2224 44134 3216
rect 44071 2208 44137 2224
rect 44071 2144 44072 2208
rect 44136 2144 44137 2208
rect 44071 2128 44137 2144
rect 44074 1136 44134 2128
rect 44071 1120 44137 1136
rect 44071 1056 44072 1120
rect 44136 1056 44137 1120
rect 44071 1040 44137 1056
rect 44074 -279 44134 1040
rect 44071 -280 44137 -279
rect 44071 -344 44072 -280
rect 44136 -344 44137 -280
rect 44071 -345 44137 -344
rect 44074 -482 44134 -345
rect 44474 -559 44534 11439
rect 44471 -560 44537 -559
rect 44471 -624 44472 -560
rect 44536 -624 44537 -560
rect 44471 -625 44537 -624
rect 44474 -762 44534 -625
rect 44874 -839 44934 11719
rect 44871 -840 44937 -839
rect 44871 -904 44872 -840
rect 44936 -904 44937 -840
rect 44871 -905 44937 -904
rect 44874 -1042 44934 -905
rect 45274 -1119 45334 11999
rect 45271 -1120 45337 -1119
rect 45271 -1184 45272 -1120
rect 45336 -1184 45337 -1120
rect 45271 -1185 45337 -1184
rect 45274 -1322 45334 -1185
rect 45674 -1399 45734 12279
rect 65271 12204 65337 12205
rect 65271 12140 65272 12204
rect 65336 12140 65337 12204
rect 65271 12139 65337 12140
rect 64871 11924 64937 11925
rect 64871 11860 64872 11924
rect 64936 11860 64937 11924
rect 64871 11859 64937 11860
rect 64471 11644 64537 11645
rect 64471 11580 64472 11644
rect 64536 11580 64537 11644
rect 64471 11579 64537 11580
rect 64071 11364 64137 11365
rect 64071 11300 64072 11364
rect 64136 11300 64137 11364
rect 64071 11299 64137 11300
rect 64074 9296 64134 11299
rect 64071 9280 64137 9296
rect 64071 9216 64072 9280
rect 64136 9216 64137 9280
rect 64071 9200 64137 9216
rect 64074 8208 64134 9200
rect 64071 8192 64137 8208
rect 64071 8128 64072 8192
rect 64136 8128 64137 8192
rect 64071 8112 64137 8128
rect 64074 7120 64134 8112
rect 64071 7104 64137 7120
rect 64071 7040 64072 7104
rect 64136 7040 64137 7104
rect 64071 7024 64137 7040
rect 64074 6032 64134 7024
rect 64071 6016 64137 6032
rect 64071 5952 64072 6016
rect 64136 5952 64137 6016
rect 64071 5936 64137 5952
rect 64074 4944 64134 5936
rect 64071 4928 64137 4944
rect 64071 4864 64072 4928
rect 64136 4864 64137 4928
rect 64071 4848 64137 4864
rect 64074 3856 64134 4848
rect 64071 3840 64137 3856
rect 64071 3776 64072 3840
rect 64136 3776 64137 3840
rect 64071 3760 64137 3776
rect 64074 2768 64134 3760
rect 64071 2752 64137 2768
rect 64071 2688 64072 2752
rect 64136 2688 64137 2752
rect 64071 2672 64137 2688
rect 64074 1680 64134 2672
rect 64071 1664 64137 1680
rect 64071 1600 64072 1664
rect 64136 1600 64137 1664
rect 64071 1584 64137 1600
rect 64074 -419 64134 1584
rect 64071 -420 64137 -419
rect 64071 -484 64072 -420
rect 64136 -484 64137 -420
rect 64071 -485 64137 -484
rect 64474 -699 64534 11579
rect 64471 -700 64537 -699
rect 64471 -764 64472 -700
rect 64536 -764 64537 -700
rect 64471 -765 64537 -764
rect 64874 -979 64934 11859
rect 64871 -980 64937 -979
rect 64871 -1044 64872 -980
rect 64936 -1044 64937 -980
rect 64871 -1045 64937 -1044
rect 65274 -1259 65334 12139
rect 65271 -1260 65337 -1259
rect 65271 -1324 65272 -1260
rect 65336 -1324 65337 -1260
rect 65271 -1325 65337 -1324
rect 45671 -1400 45737 -1399
rect 45671 -1464 45672 -1400
rect 45736 -1464 45737 -1400
rect 45671 -1465 45737 -1464
rect 25671 -1540 25737 -1539
rect -1589 -1605 -1523 -1604
rect 25671 -1604 25672 -1540
rect 25736 -1604 25737 -1540
rect 45674 -1602 45734 -1465
rect 65674 -1539 65734 12419
rect 85674 12345 85734 12482
rect 105671 12420 105672 12484
rect 105736 12420 105737 12484
rect 145671 12484 145737 12485
rect 105671 12419 105737 12420
rect 85671 12344 85737 12345
rect 85671 12280 85672 12344
rect 85736 12280 85737 12344
rect 85671 12279 85737 12280
rect 85274 12065 85334 12202
rect 85271 12064 85337 12065
rect 85271 12000 85272 12064
rect 85336 12000 85337 12064
rect 85271 11999 85337 12000
rect 84874 11785 84934 11922
rect 84871 11784 84937 11785
rect 84871 11720 84872 11784
rect 84936 11720 84937 11784
rect 84871 11719 84937 11720
rect 84474 11505 84534 11642
rect 84471 11504 84537 11505
rect 84471 11440 84472 11504
rect 84536 11440 84537 11504
rect 84471 11439 84537 11440
rect 84074 11225 84134 11362
rect 84071 11224 84137 11225
rect 84071 11160 84072 11224
rect 84136 11160 84137 11224
rect 84071 11159 84137 11160
rect 84074 9840 84134 11159
rect 84071 9824 84137 9840
rect 84071 9760 84072 9824
rect 84136 9760 84137 9824
rect 84071 9744 84137 9760
rect 84074 8752 84134 9744
rect 84071 8736 84137 8752
rect 84071 8672 84072 8736
rect 84136 8672 84137 8736
rect 84071 8656 84137 8672
rect 84074 7664 84134 8656
rect 84071 7648 84137 7664
rect 84071 7584 84072 7648
rect 84136 7584 84137 7648
rect 84071 7568 84137 7584
rect 84074 6576 84134 7568
rect 84071 6560 84137 6576
rect 84071 6496 84072 6560
rect 84136 6496 84137 6560
rect 84071 6480 84137 6496
rect 84074 5488 84134 6480
rect 84071 5472 84137 5488
rect 84071 5408 84072 5472
rect 84136 5408 84137 5472
rect 84071 5392 84137 5408
rect 84074 4400 84134 5392
rect 84071 4384 84137 4400
rect 84071 4320 84072 4384
rect 84136 4320 84137 4384
rect 84071 4304 84137 4320
rect 84074 3312 84134 4304
rect 84071 3296 84137 3312
rect 84071 3232 84072 3296
rect 84136 3232 84137 3296
rect 84071 3216 84137 3232
rect 84074 2224 84134 3216
rect 84071 2208 84137 2224
rect 84071 2144 84072 2208
rect 84136 2144 84137 2208
rect 84071 2128 84137 2144
rect 84074 1136 84134 2128
rect 84071 1120 84137 1136
rect 84071 1056 84072 1120
rect 84136 1056 84137 1120
rect 84071 1040 84137 1056
rect 84074 -279 84134 1040
rect 84071 -280 84137 -279
rect 84071 -344 84072 -280
rect 84136 -344 84137 -280
rect 84071 -345 84137 -344
rect 84074 -482 84134 -345
rect 84474 -559 84534 11439
rect 84471 -560 84537 -559
rect 84471 -624 84472 -560
rect 84536 -624 84537 -560
rect 84471 -625 84537 -624
rect 84474 -762 84534 -625
rect 84874 -839 84934 11719
rect 84871 -840 84937 -839
rect 84871 -904 84872 -840
rect 84936 -904 84937 -840
rect 84871 -905 84937 -904
rect 84874 -1042 84934 -905
rect 85274 -1119 85334 11999
rect 85271 -1120 85337 -1119
rect 85271 -1184 85272 -1120
rect 85336 -1184 85337 -1120
rect 85271 -1185 85337 -1184
rect 85274 -1322 85334 -1185
rect 85674 -1399 85734 12279
rect 105271 12204 105337 12205
rect 105271 12140 105272 12204
rect 105336 12140 105337 12204
rect 105271 12139 105337 12140
rect 104871 11924 104937 11925
rect 104871 11860 104872 11924
rect 104936 11860 104937 11924
rect 104871 11859 104937 11860
rect 104471 11644 104537 11645
rect 104471 11580 104472 11644
rect 104536 11580 104537 11644
rect 104471 11579 104537 11580
rect 104071 11364 104137 11365
rect 104071 11300 104072 11364
rect 104136 11300 104137 11364
rect 104071 11299 104137 11300
rect 104074 9296 104134 11299
rect 104071 9280 104137 9296
rect 104071 9216 104072 9280
rect 104136 9216 104137 9280
rect 104071 9200 104137 9216
rect 104074 8208 104134 9200
rect 104071 8192 104137 8208
rect 104071 8128 104072 8192
rect 104136 8128 104137 8192
rect 104071 8112 104137 8128
rect 104074 7120 104134 8112
rect 104071 7104 104137 7120
rect 104071 7040 104072 7104
rect 104136 7040 104137 7104
rect 104071 7024 104137 7040
rect 104074 6032 104134 7024
rect 104071 6016 104137 6032
rect 104071 5952 104072 6016
rect 104136 5952 104137 6016
rect 104071 5936 104137 5952
rect 104074 4944 104134 5936
rect 104071 4928 104137 4944
rect 104071 4864 104072 4928
rect 104136 4864 104137 4928
rect 104071 4848 104137 4864
rect 104074 3856 104134 4848
rect 104071 3840 104137 3856
rect 104071 3776 104072 3840
rect 104136 3776 104137 3840
rect 104071 3760 104137 3776
rect 104074 2768 104134 3760
rect 104071 2752 104137 2768
rect 104071 2688 104072 2752
rect 104136 2688 104137 2752
rect 104071 2672 104137 2688
rect 104074 1680 104134 2672
rect 104071 1664 104137 1680
rect 104071 1600 104072 1664
rect 104136 1600 104137 1664
rect 104071 1584 104137 1600
rect 104074 -419 104134 1584
rect 104071 -420 104137 -419
rect 104071 -484 104072 -420
rect 104136 -484 104137 -420
rect 104071 -485 104137 -484
rect 104474 -699 104534 11579
rect 104471 -700 104537 -699
rect 104471 -764 104472 -700
rect 104536 -764 104537 -700
rect 104471 -765 104537 -764
rect 104874 -979 104934 11859
rect 104871 -980 104937 -979
rect 104871 -1044 104872 -980
rect 104936 -1044 104937 -980
rect 104871 -1045 104937 -1044
rect 105274 -1259 105334 12139
rect 105271 -1260 105337 -1259
rect 105271 -1324 105272 -1260
rect 105336 -1324 105337 -1260
rect 105271 -1325 105337 -1324
rect 85671 -1400 85737 -1399
rect 85671 -1464 85672 -1400
rect 85736 -1464 85737 -1400
rect 85671 -1465 85737 -1464
rect 65671 -1540 65737 -1539
rect 25671 -1605 25737 -1604
rect 65671 -1604 65672 -1540
rect 65736 -1604 65737 -1540
rect 85674 -1602 85734 -1465
rect 105674 -1539 105734 12419
rect 125674 12345 125734 12482
rect 145671 12420 145672 12484
rect 145736 12420 145737 12484
rect 185671 12484 185737 12485
rect 145671 12419 145737 12420
rect 125671 12344 125737 12345
rect 125671 12280 125672 12344
rect 125736 12280 125737 12344
rect 125671 12279 125737 12280
rect 125274 12065 125334 12202
rect 125271 12064 125337 12065
rect 125271 12000 125272 12064
rect 125336 12000 125337 12064
rect 125271 11999 125337 12000
rect 124874 11785 124934 11922
rect 124871 11784 124937 11785
rect 124871 11720 124872 11784
rect 124936 11720 124937 11784
rect 124871 11719 124937 11720
rect 124474 11505 124534 11642
rect 124471 11504 124537 11505
rect 124471 11440 124472 11504
rect 124536 11440 124537 11504
rect 124471 11439 124537 11440
rect 124074 11225 124134 11362
rect 124071 11224 124137 11225
rect 124071 11160 124072 11224
rect 124136 11160 124137 11224
rect 124071 11159 124137 11160
rect 124074 9840 124134 11159
rect 124071 9824 124137 9840
rect 124071 9760 124072 9824
rect 124136 9760 124137 9824
rect 124071 9744 124137 9760
rect 124074 8752 124134 9744
rect 124071 8736 124137 8752
rect 124071 8672 124072 8736
rect 124136 8672 124137 8736
rect 124071 8656 124137 8672
rect 124074 7664 124134 8656
rect 124071 7648 124137 7664
rect 124071 7584 124072 7648
rect 124136 7584 124137 7648
rect 124071 7568 124137 7584
rect 124074 6576 124134 7568
rect 124259 7308 124325 7309
rect 124259 7244 124260 7308
rect 124324 7244 124325 7308
rect 124259 7243 124325 7244
rect 124262 6765 124322 7243
rect 124213 6764 124322 6765
rect 124213 6700 124214 6764
rect 124278 6702 124322 6764
rect 124278 6700 124279 6702
rect 124213 6699 124279 6700
rect 124071 6560 124137 6576
rect 124071 6496 124072 6560
rect 124136 6496 124137 6560
rect 124071 6480 124137 6496
rect 124074 5488 124134 6480
rect 124259 6220 124325 6221
rect 124259 6156 124260 6220
rect 124324 6156 124325 6220
rect 124259 6155 124325 6156
rect 124071 5472 124137 5488
rect 124071 5408 124072 5472
rect 124136 5408 124137 5472
rect 124071 5392 124137 5408
rect 124262 5405 124322 6155
rect 124259 5404 124325 5405
rect 124074 4400 124134 5392
rect 124259 5340 124260 5404
rect 124324 5340 124325 5404
rect 124259 5339 124325 5340
rect 124071 4384 124137 4400
rect 124071 4320 124072 4384
rect 124136 4320 124137 4384
rect 124071 4304 124137 4320
rect 124074 3312 124134 4304
rect 124071 3296 124137 3312
rect 124071 3232 124072 3296
rect 124136 3232 124137 3296
rect 124071 3216 124137 3232
rect 124074 2224 124134 3216
rect 124071 2208 124137 2224
rect 124071 2144 124072 2208
rect 124136 2144 124137 2208
rect 124071 2128 124137 2144
rect 124074 1136 124134 2128
rect 124071 1120 124137 1136
rect 124071 1056 124072 1120
rect 124136 1056 124137 1120
rect 124071 1040 124137 1056
rect 124074 -279 124134 1040
rect 124071 -280 124137 -279
rect 124071 -344 124072 -280
rect 124136 -344 124137 -280
rect 124071 -345 124137 -344
rect 124074 -482 124134 -345
rect 124474 -559 124534 11439
rect 124471 -560 124537 -559
rect 124471 -624 124472 -560
rect 124536 -624 124537 -560
rect 124471 -625 124537 -624
rect 124474 -762 124534 -625
rect 124874 -839 124934 11719
rect 124871 -840 124937 -839
rect 124871 -904 124872 -840
rect 124936 -904 124937 -840
rect 124871 -905 124937 -904
rect 124874 -1042 124934 -905
rect 125274 -1119 125334 11999
rect 125271 -1120 125337 -1119
rect 125271 -1184 125272 -1120
rect 125336 -1184 125337 -1120
rect 125271 -1185 125337 -1184
rect 125274 -1322 125334 -1185
rect 125674 -1399 125734 12279
rect 145271 12204 145337 12205
rect 145271 12140 145272 12204
rect 145336 12140 145337 12204
rect 145271 12139 145337 12140
rect 144871 11924 144937 11925
rect 144871 11860 144872 11924
rect 144936 11860 144937 11924
rect 144871 11859 144937 11860
rect 144471 11644 144537 11645
rect 144471 11580 144472 11644
rect 144536 11580 144537 11644
rect 144471 11579 144537 11580
rect 144071 11364 144137 11365
rect 144071 11300 144072 11364
rect 144136 11300 144137 11364
rect 144071 11299 144137 11300
rect 144074 9296 144134 11299
rect 144071 9280 144137 9296
rect 144071 9216 144072 9280
rect 144136 9216 144137 9280
rect 144071 9200 144137 9216
rect 144074 8208 144134 9200
rect 144071 8192 144137 8208
rect 144071 8128 144072 8192
rect 144136 8128 144137 8192
rect 144071 8112 144137 8128
rect 144074 7120 144134 8112
rect 144071 7104 144137 7120
rect 144071 7040 144072 7104
rect 144136 7040 144137 7104
rect 144071 7024 144137 7040
rect 134747 6764 134813 6765
rect 134747 6700 134748 6764
rect 134812 6700 134813 6764
rect 134747 6699 134813 6700
rect 134750 6490 134810 6699
rect 135115 6492 135181 6493
rect 135115 6490 135116 6492
rect 134750 6430 135116 6490
rect 135115 6428 135116 6430
rect 135180 6428 135181 6492
rect 135115 6427 135181 6428
rect 144074 6032 144134 7024
rect 144071 6016 144137 6032
rect 144071 5952 144072 6016
rect 144136 5952 144137 6016
rect 144071 5936 144137 5952
rect 144074 4944 144134 5936
rect 144071 4928 144137 4944
rect 144071 4864 144072 4928
rect 144136 4864 144137 4928
rect 144071 4848 144137 4864
rect 144074 3856 144134 4848
rect 144071 3840 144137 3856
rect 144071 3776 144072 3840
rect 144136 3776 144137 3840
rect 144071 3760 144137 3776
rect 137323 3364 137389 3365
rect 137323 3300 137324 3364
rect 137388 3300 137389 3364
rect 137323 3299 137389 3300
rect 137326 3090 137386 3299
rect 137691 3092 137757 3093
rect 137691 3090 137692 3092
rect 137326 3030 137692 3090
rect 137691 3028 137692 3030
rect 137756 3028 137757 3092
rect 137691 3027 137757 3028
rect 144074 2768 144134 3760
rect 144071 2752 144137 2768
rect 144071 2688 144072 2752
rect 144136 2688 144137 2752
rect 138427 2684 138493 2685
rect 138427 2682 138428 2684
rect 138062 2622 138428 2682
rect 138062 2277 138122 2622
rect 138427 2620 138428 2622
rect 138492 2620 138493 2684
rect 144071 2672 144137 2688
rect 138427 2619 138493 2620
rect 138059 2276 138125 2277
rect 138059 2212 138060 2276
rect 138124 2212 138125 2276
rect 138059 2211 138125 2212
rect 138243 2276 138309 2277
rect 138243 2212 138244 2276
rect 138308 2212 138309 2276
rect 138243 2211 138309 2212
rect 137875 2140 137941 2141
rect 137875 2076 137876 2140
rect 137940 2076 137941 2140
rect 137875 2075 137941 2076
rect 137878 1730 137938 2075
rect 137694 1670 137938 1730
rect 138059 1732 138125 1733
rect 137694 1189 137754 1670
rect 138059 1668 138060 1732
rect 138124 1730 138125 1732
rect 138246 1730 138306 2211
rect 138124 1670 138306 1730
rect 144074 1680 144134 2672
rect 138124 1668 138125 1670
rect 138059 1667 138125 1668
rect 144071 1664 144137 1680
rect 144071 1600 144072 1664
rect 144136 1600 144137 1664
rect 144071 1584 144137 1600
rect 137691 1188 137757 1189
rect 137691 1124 137692 1188
rect 137756 1124 137757 1188
rect 137691 1123 137757 1124
rect 137875 1188 137941 1189
rect 137875 1124 137876 1188
rect 137940 1124 137941 1188
rect 137875 1123 137941 1124
rect 137139 1052 137205 1053
rect 137139 988 137140 1052
rect 137204 1050 137205 1052
rect 137878 1050 137938 1123
rect 137204 990 137938 1050
rect 137204 988 137205 990
rect 137139 987 137205 988
rect 132726 310 137938 370
rect 132726 101 132786 310
rect 137878 101 137938 310
rect 132723 100 132789 101
rect 132723 36 132724 100
rect 132788 36 132789 100
rect 132723 35 132789 36
rect 137875 100 137941 101
rect 137875 36 137876 100
rect 137940 36 137941 100
rect 137875 35 137941 36
rect 144074 -419 144134 1584
rect 144071 -420 144137 -419
rect 144071 -484 144072 -420
rect 144136 -484 144137 -420
rect 144071 -485 144137 -484
rect 144474 -699 144534 11579
rect 144471 -700 144537 -699
rect 144471 -764 144472 -700
rect 144536 -764 144537 -700
rect 144471 -765 144537 -764
rect 144874 -979 144934 11859
rect 145051 4316 145117 4317
rect 145051 4252 145052 4316
rect 145116 4252 145117 4316
rect 145051 4251 145117 4252
rect 145054 237 145114 4251
rect 145051 236 145117 237
rect 145051 172 145052 236
rect 145116 172 145117 236
rect 145051 171 145117 172
rect 144871 -980 144937 -979
rect 144871 -1044 144872 -980
rect 144936 -1044 144937 -980
rect 144871 -1045 144937 -1044
rect 145274 -1259 145334 12139
rect 145271 -1260 145337 -1259
rect 145271 -1324 145272 -1260
rect 145336 -1324 145337 -1260
rect 145271 -1325 145337 -1324
rect 125671 -1400 125737 -1399
rect 125671 -1464 125672 -1400
rect 125736 -1464 125737 -1400
rect 125671 -1465 125737 -1464
rect 105671 -1540 105737 -1539
rect 65671 -1605 65737 -1604
rect 105671 -1604 105672 -1540
rect 105736 -1604 105737 -1540
rect 125674 -1602 125734 -1465
rect 145674 -1539 145734 12419
rect 165674 12345 165734 12482
rect 185671 12420 185672 12484
rect 185736 12420 185737 12484
rect 185671 12419 185737 12420
rect 201439 12484 201505 12485
rect 201439 12420 201440 12484
rect 201504 12420 201505 12484
rect 201439 12419 201505 12420
rect 165671 12344 165737 12345
rect 165671 12280 165672 12344
rect 165736 12280 165737 12344
rect 165671 12279 165737 12280
rect 165274 12065 165334 12202
rect 165271 12064 165337 12065
rect 165271 12000 165272 12064
rect 165336 12000 165337 12064
rect 165271 11999 165337 12000
rect 164874 11785 164934 11922
rect 164871 11784 164937 11785
rect 164871 11720 164872 11784
rect 164936 11720 164937 11784
rect 164871 11719 164937 11720
rect 164474 11505 164534 11642
rect 164471 11504 164537 11505
rect 164471 11440 164472 11504
rect 164536 11440 164537 11504
rect 164471 11439 164537 11440
rect 164074 11225 164134 11362
rect 164071 11224 164137 11225
rect 164071 11160 164072 11224
rect 164136 11160 164137 11224
rect 164071 11159 164137 11160
rect 164074 9840 164134 11159
rect 164071 9824 164137 9840
rect 164071 9760 164072 9824
rect 164136 9760 164137 9824
rect 157379 9756 157445 9757
rect 157379 9692 157380 9756
rect 157444 9692 157445 9756
rect 164071 9744 164137 9760
rect 157379 9691 157445 9692
rect 157195 7716 157261 7717
rect 157195 7652 157196 7716
rect 157260 7652 157261 7716
rect 157195 7651 157261 7652
rect 157011 7444 157077 7445
rect 157011 7380 157012 7444
rect 157076 7380 157077 7444
rect 157011 7379 157077 7380
rect 157014 5405 157074 7379
rect 157011 5404 157077 5405
rect 157011 5340 157012 5404
rect 157076 5340 157077 5404
rect 157011 5339 157077 5340
rect 157011 4996 157077 4997
rect 157011 4932 157012 4996
rect 157076 4932 157077 4996
rect 157011 4931 157077 4932
rect 157014 4450 157074 4931
rect 157198 4589 157258 7651
rect 157382 7309 157442 9691
rect 157747 8804 157813 8805
rect 157747 8740 157748 8804
rect 157812 8740 157813 8804
rect 164074 8752 164134 9744
rect 157747 8739 157813 8740
rect 157750 8530 157810 8739
rect 164071 8736 164137 8752
rect 164071 8672 164072 8736
rect 164136 8672 164137 8736
rect 164071 8656 164137 8672
rect 157566 8470 157810 8530
rect 157566 8397 157626 8470
rect 157563 8396 157629 8397
rect 157563 8332 157564 8396
rect 157628 8332 157629 8396
rect 157563 8331 157629 8332
rect 161979 8124 162045 8125
rect 161979 8060 161980 8124
rect 162044 8122 162045 8124
rect 162044 8062 162226 8122
rect 162044 8060 162045 8062
rect 161979 8059 162045 8060
rect 158667 7444 158733 7445
rect 158667 7380 158668 7444
rect 158732 7380 158733 7444
rect 158667 7379 158733 7380
rect 158851 7444 158917 7445
rect 158851 7380 158852 7444
rect 158916 7380 158917 7444
rect 158851 7379 158917 7380
rect 159955 7444 160021 7445
rect 159955 7380 159956 7444
rect 160020 7380 160021 7444
rect 159955 7379 160021 7380
rect 161427 7444 161493 7445
rect 161427 7380 161428 7444
rect 161492 7380 161493 7444
rect 161427 7379 161493 7380
rect 157379 7308 157445 7309
rect 157379 7244 157380 7308
rect 157444 7244 157445 7308
rect 157379 7243 157445 7244
rect 158670 7037 158730 7379
rect 158667 7036 158733 7037
rect 158667 6972 158668 7036
rect 158732 6972 158733 7036
rect 158667 6971 158733 6972
rect 157195 4588 157261 4589
rect 157195 4524 157196 4588
rect 157260 4524 157261 4588
rect 157195 4523 157261 4524
rect 157014 4390 157442 4450
rect 157382 3637 157442 4390
rect 157379 3636 157445 3637
rect 157379 3572 157380 3636
rect 157444 3572 157445 3636
rect 157379 3571 157445 3572
rect 157011 3228 157077 3229
rect 157011 3164 157012 3228
rect 157076 3226 157077 3228
rect 157076 3166 157442 3226
rect 157076 3164 157077 3166
rect 157011 3163 157077 3164
rect 157382 3093 157442 3166
rect 151859 3092 151925 3093
rect 151859 3028 151860 3092
rect 151924 3028 151925 3092
rect 151859 3027 151925 3028
rect 157379 3092 157445 3093
rect 157379 3028 157380 3092
rect 157444 3028 157445 3092
rect 157379 3027 157445 3028
rect 151862 1053 151922 3027
rect 158854 2005 158914 7379
rect 158851 2004 158917 2005
rect 158851 1940 158852 2004
rect 158916 1940 158917 2004
rect 158851 1939 158917 1940
rect 159958 1597 160018 7379
rect 161430 2141 161490 7379
rect 161611 3500 161677 3501
rect 161611 3436 161612 3500
rect 161676 3436 161677 3500
rect 161611 3435 161677 3436
rect 161795 3500 161861 3501
rect 161795 3436 161796 3500
rect 161860 3436 161861 3500
rect 161795 3435 161861 3436
rect 161427 2140 161493 2141
rect 161427 2076 161428 2140
rect 161492 2076 161493 2140
rect 161427 2075 161493 2076
rect 159955 1596 160021 1597
rect 159955 1532 159956 1596
rect 160020 1532 160021 1596
rect 159955 1531 160021 1532
rect 151859 1052 151925 1053
rect 151859 988 151860 1052
rect 151924 988 151925 1052
rect 151859 987 151925 988
rect 161614 645 161674 3435
rect 161798 3093 161858 3435
rect 161795 3092 161861 3093
rect 161795 3028 161796 3092
rect 161860 3028 161861 3092
rect 161795 3027 161861 3028
rect 161979 3092 162045 3093
rect 161979 3028 161980 3092
rect 162044 3028 162045 3092
rect 161979 3027 162045 3028
rect 161982 2685 162042 3027
rect 162166 2954 162226 8062
rect 164074 7664 164134 8656
rect 164071 7648 164137 7664
rect 164071 7584 164072 7648
rect 164136 7584 164137 7648
rect 164071 7568 164137 7584
rect 163083 3364 163149 3365
rect 163083 3300 163084 3364
rect 163148 3300 163149 3364
rect 163083 3299 163149 3300
rect 162899 3228 162965 3229
rect 162899 3164 162900 3228
rect 162964 3164 162965 3228
rect 162899 3163 162965 3164
rect 162347 2956 162413 2957
rect 162347 2954 162348 2956
rect 162166 2894 162348 2954
rect 162347 2892 162348 2894
rect 162412 2892 162413 2956
rect 162347 2891 162413 2892
rect 162902 2685 162962 3163
rect 161979 2684 162045 2685
rect 161979 2620 161980 2684
rect 162044 2620 162045 2684
rect 161979 2619 162045 2620
rect 162899 2684 162965 2685
rect 162899 2620 162900 2684
rect 162964 2620 162965 2684
rect 162899 2619 162965 2620
rect 162347 1188 162413 1189
rect 162347 1124 162348 1188
rect 162412 1124 162413 1188
rect 162347 1123 162413 1124
rect 162350 1050 162410 1123
rect 161798 990 162410 1050
rect 161611 644 161677 645
rect 161611 580 161612 644
rect 161676 580 161677 644
rect 161611 579 161677 580
rect 161798 101 161858 990
rect 163086 509 163146 3299
rect 164074 2224 164134 7568
rect 164474 6745 164534 11439
rect 164739 7444 164805 7445
rect 164739 7380 164740 7444
rect 164804 7380 164805 7444
rect 164739 7379 164805 7380
rect 164471 6744 164537 6745
rect 164471 6680 164472 6744
rect 164536 6680 164537 6744
rect 164471 6679 164537 6680
rect 164474 5288 164534 6679
rect 164471 5287 164537 5288
rect 164471 5223 164472 5287
rect 164536 5223 164537 5287
rect 164471 5222 164537 5223
rect 164474 3831 164534 5222
rect 164471 3830 164537 3831
rect 164471 3766 164472 3830
rect 164536 3766 164537 3830
rect 164471 3765 164537 3766
rect 164071 2208 164137 2224
rect 164071 2144 164072 2208
rect 164136 2144 164137 2208
rect 164071 2128 164137 2144
rect 164074 1136 164134 2128
rect 164071 1120 164137 1136
rect 164071 1056 164072 1120
rect 164136 1056 164137 1120
rect 164071 1040 164137 1056
rect 163083 508 163149 509
rect 163083 444 163084 508
rect 163148 444 163149 508
rect 163083 443 163149 444
rect 163451 508 163517 509
rect 163451 444 163452 508
rect 163516 444 163517 508
rect 163451 443 163517 444
rect 163454 370 163514 443
rect 161982 310 163514 370
rect 161982 237 162042 310
rect 161979 236 162045 237
rect 161979 172 161980 236
rect 162044 172 162045 236
rect 161979 171 162045 172
rect 161795 100 161861 101
rect 161795 36 161796 100
rect 161860 36 161861 100
rect 161795 35 161861 36
rect 164074 -279 164134 1040
rect 164071 -280 164137 -279
rect 164071 -344 164072 -280
rect 164136 -344 164137 -280
rect 164071 -345 164137 -344
rect 164074 -482 164134 -345
rect 164474 -559 164534 3765
rect 164742 3229 164802 7379
rect 164739 3228 164805 3229
rect 164739 3164 164740 3228
rect 164804 3164 164805 3228
rect 164739 3163 164805 3164
rect 164739 2820 164805 2821
rect 164739 2756 164740 2820
rect 164804 2756 164805 2820
rect 164739 2755 164805 2756
rect 164742 1461 164802 2755
rect 164739 1460 164805 1461
rect 164739 1396 164740 1460
rect 164804 1396 164805 1460
rect 164739 1395 164805 1396
rect 164471 -560 164537 -559
rect 164471 -624 164472 -560
rect 164536 -624 164537 -560
rect 164471 -625 164537 -624
rect 164474 -762 164534 -625
rect 164874 -839 164934 11719
rect 165107 7580 165173 7581
rect 165107 7516 165108 7580
rect 165172 7516 165173 7580
rect 165107 7515 165173 7516
rect 165110 2821 165170 7515
rect 165274 5739 165334 11999
rect 165475 8396 165541 8397
rect 165475 8332 165476 8396
rect 165540 8332 165541 8396
rect 165475 8331 165541 8332
rect 165271 5738 165337 5739
rect 165271 5674 165272 5738
rect 165336 5674 165337 5738
rect 165271 5673 165337 5674
rect 165274 4282 165334 5673
rect 165271 4281 165337 4282
rect 165271 4217 165272 4281
rect 165336 4217 165337 4281
rect 165271 4216 165337 4217
rect 165107 2820 165173 2821
rect 165107 2756 165108 2820
rect 165172 2756 165173 2820
rect 165107 2755 165173 2756
rect 165107 1868 165173 1869
rect 165107 1804 165108 1868
rect 165172 1804 165173 1868
rect 165107 1803 165173 1804
rect 165110 1461 165170 1803
rect 165107 1460 165173 1461
rect 165107 1396 165108 1460
rect 165172 1396 165173 1460
rect 165107 1395 165173 1396
rect 164871 -840 164937 -839
rect 164871 -904 164872 -840
rect 164936 -904 164937 -840
rect 164871 -905 164937 -904
rect 164874 -1042 164934 -905
rect 165274 -1119 165334 4216
rect 165478 2957 165538 8331
rect 165674 6139 165734 12279
rect 185271 12204 185337 12205
rect 185271 12140 185272 12204
rect 185336 12140 185337 12204
rect 185271 12139 185337 12140
rect 184871 11924 184937 11925
rect 184871 11860 184872 11924
rect 184936 11860 184937 11924
rect 184871 11859 184937 11860
rect 184471 11644 184537 11645
rect 184471 11580 184472 11644
rect 184536 11580 184537 11644
rect 184471 11579 184537 11580
rect 184071 11364 184137 11365
rect 184071 11300 184072 11364
rect 184136 11300 184137 11364
rect 184071 11299 184137 11300
rect 184074 9296 184134 11299
rect 184071 9280 184137 9296
rect 184071 9216 184072 9280
rect 184136 9216 184137 9280
rect 184071 9200 184137 9216
rect 167867 9076 167933 9077
rect 167867 9012 167868 9076
rect 167932 9012 167933 9076
rect 167867 9011 167933 9012
rect 173755 9076 173821 9077
rect 173755 9012 173756 9076
rect 173820 9012 173821 9076
rect 173755 9011 173821 9012
rect 167131 7852 167197 7853
rect 167131 7788 167132 7852
rect 167196 7788 167197 7852
rect 167131 7787 167197 7788
rect 167315 7852 167381 7853
rect 167315 7788 167316 7852
rect 167380 7788 167381 7852
rect 167315 7787 167381 7788
rect 166027 7580 166093 7581
rect 166027 7516 166028 7580
rect 166092 7516 166093 7580
rect 166027 7515 166093 7516
rect 165843 7444 165909 7445
rect 165843 7380 165844 7444
rect 165908 7380 165909 7444
rect 165843 7379 165909 7380
rect 165671 6138 165737 6139
rect 165671 6074 165672 6138
rect 165736 6074 165737 6138
rect 165671 6073 165737 6074
rect 165674 4682 165734 6073
rect 165671 4681 165737 4682
rect 165671 4617 165672 4681
rect 165736 4617 165737 4681
rect 165671 4616 165737 4617
rect 165475 2956 165541 2957
rect 165475 2892 165476 2956
rect 165540 2892 165541 2956
rect 165475 2891 165541 2892
rect 165271 -1120 165337 -1119
rect 165271 -1184 165272 -1120
rect 165336 -1184 165337 -1120
rect 165271 -1185 165337 -1184
rect 165274 -1322 165334 -1185
rect 165674 -1399 165734 4616
rect 165846 2141 165906 7379
rect 166030 2685 166090 7515
rect 166763 3228 166829 3229
rect 166763 3164 166764 3228
rect 166828 3164 166829 3228
rect 166763 3163 166829 3164
rect 166579 2820 166645 2821
rect 166579 2756 166580 2820
rect 166644 2756 166645 2820
rect 166579 2755 166645 2756
rect 166027 2684 166093 2685
rect 166027 2620 166028 2684
rect 166092 2620 166093 2684
rect 166027 2619 166093 2620
rect 165843 2140 165909 2141
rect 165843 2076 165844 2140
rect 165908 2076 165909 2140
rect 165843 2075 165909 2076
rect 166582 237 166642 2755
rect 166766 1461 166826 3163
rect 166763 1460 166829 1461
rect 166763 1396 166764 1460
rect 166828 1396 166829 1460
rect 166763 1395 166829 1396
rect 166579 236 166645 237
rect 166579 172 166580 236
rect 166644 172 166645 236
rect 166579 171 166645 172
rect 167134 101 167194 7787
rect 167318 3501 167378 7787
rect 167683 7444 167749 7445
rect 167683 7380 167684 7444
rect 167748 7380 167749 7444
rect 167683 7379 167749 7380
rect 167315 3500 167381 3501
rect 167315 3436 167316 3500
rect 167380 3436 167381 3500
rect 167315 3435 167381 3436
rect 167499 3500 167565 3501
rect 167499 3436 167500 3500
rect 167564 3436 167565 3500
rect 167499 3435 167565 3436
rect 167502 2685 167562 3435
rect 167686 2685 167746 7379
rect 167870 2821 167930 9011
rect 168971 8940 169037 8941
rect 168971 8876 168972 8940
rect 169036 8876 169037 8940
rect 168971 8875 169037 8876
rect 168051 7172 168117 7173
rect 168051 7108 168052 7172
rect 168116 7108 168117 7172
rect 168051 7107 168117 7108
rect 168054 2957 168114 7107
rect 168974 3093 169034 8875
rect 169523 8396 169589 8397
rect 169523 8332 169524 8396
rect 169588 8332 169589 8396
rect 169523 8331 169589 8332
rect 170811 8396 170877 8397
rect 170811 8332 170812 8396
rect 170876 8332 170877 8396
rect 170811 8331 170877 8332
rect 168971 3092 169037 3093
rect 168971 3028 168972 3092
rect 169036 3028 169037 3092
rect 168971 3027 169037 3028
rect 168051 2956 168117 2957
rect 168051 2892 168052 2956
rect 168116 2892 168117 2956
rect 168051 2891 168117 2892
rect 167867 2820 167933 2821
rect 167867 2756 167868 2820
rect 167932 2756 167933 2820
rect 167867 2755 167933 2756
rect 167499 2684 167565 2685
rect 167499 2620 167500 2684
rect 167564 2620 167565 2684
rect 167499 2619 167565 2620
rect 167683 2684 167749 2685
rect 167683 2620 167684 2684
rect 167748 2620 167749 2684
rect 167683 2619 167749 2620
rect 169526 2277 169586 8331
rect 169707 7444 169773 7445
rect 169707 7380 169708 7444
rect 169772 7380 169773 7444
rect 169707 7379 169773 7380
rect 170075 7444 170141 7445
rect 170075 7380 170076 7444
rect 170140 7380 170141 7444
rect 170075 7379 170141 7380
rect 169710 2957 169770 7379
rect 169891 3228 169957 3229
rect 169891 3164 169892 3228
rect 169956 3164 169957 3228
rect 169891 3163 169957 3164
rect 169707 2956 169773 2957
rect 169707 2892 169708 2956
rect 169772 2892 169773 2956
rect 169707 2891 169773 2892
rect 169894 2821 169954 3163
rect 170078 2957 170138 7379
rect 170075 2956 170141 2957
rect 170075 2892 170076 2956
rect 170140 2892 170141 2956
rect 170075 2891 170141 2892
rect 169891 2820 169957 2821
rect 169891 2756 169892 2820
rect 169956 2756 169957 2820
rect 169891 2755 169957 2756
rect 170814 2277 170874 8331
rect 171179 7444 171245 7445
rect 171179 7380 171180 7444
rect 171244 7380 171245 7444
rect 171179 7379 171245 7380
rect 171363 7444 171429 7445
rect 171363 7380 171364 7444
rect 171428 7380 171429 7444
rect 171363 7379 171429 7380
rect 171731 7444 171797 7445
rect 171731 7380 171732 7444
rect 171796 7380 171797 7444
rect 171731 7379 171797 7380
rect 172467 7444 172533 7445
rect 172467 7380 172468 7444
rect 172532 7380 172533 7444
rect 172467 7379 172533 7380
rect 173387 7444 173453 7445
rect 173387 7380 173388 7444
rect 173452 7380 173453 7444
rect 173387 7379 173453 7380
rect 171182 2685 171242 7379
rect 171366 2821 171426 7379
rect 171734 2957 171794 7379
rect 172470 3637 172530 7379
rect 172467 3636 172533 3637
rect 172467 3572 172468 3636
rect 172532 3572 172533 3636
rect 172467 3571 172533 3572
rect 171731 2956 171797 2957
rect 171731 2892 171732 2956
rect 171796 2892 171797 2956
rect 171731 2891 171797 2892
rect 173390 2821 173450 7379
rect 173758 2821 173818 9011
rect 175963 8396 176029 8397
rect 175963 8332 175964 8396
rect 176028 8332 176029 8396
rect 175963 8331 176029 8332
rect 177619 8396 177685 8397
rect 177619 8332 177620 8396
rect 177684 8332 177685 8396
rect 177619 8331 177685 8332
rect 175595 7852 175661 7853
rect 175595 7788 175596 7852
rect 175660 7788 175661 7852
rect 175595 7787 175661 7788
rect 175043 7580 175109 7581
rect 175043 7516 175044 7580
rect 175108 7516 175109 7580
rect 175043 7515 175109 7516
rect 174859 7444 174925 7445
rect 174859 7380 174860 7444
rect 174924 7380 174925 7444
rect 174859 7379 174925 7380
rect 174862 2957 174922 7379
rect 175046 3090 175106 7515
rect 175046 3030 175290 3090
rect 174859 2956 174925 2957
rect 174859 2892 174860 2956
rect 174924 2892 174925 2956
rect 174859 2891 174925 2892
rect 171363 2820 171429 2821
rect 171363 2756 171364 2820
rect 171428 2756 171429 2820
rect 171363 2755 171429 2756
rect 173387 2820 173453 2821
rect 173387 2756 173388 2820
rect 173452 2756 173453 2820
rect 173387 2755 173453 2756
rect 173755 2820 173821 2821
rect 173755 2756 173756 2820
rect 173820 2756 173821 2820
rect 173755 2755 173821 2756
rect 171179 2684 171245 2685
rect 171179 2620 171180 2684
rect 171244 2620 171245 2684
rect 171179 2619 171245 2620
rect 171915 2412 171981 2413
rect 171915 2410 171916 2412
rect 170998 2350 171916 2410
rect 169523 2276 169589 2277
rect 169523 2212 169524 2276
rect 169588 2212 169589 2276
rect 169523 2211 169589 2212
rect 170811 2276 170877 2277
rect 170811 2212 170812 2276
rect 170876 2212 170877 2276
rect 170811 2211 170877 2212
rect 170998 1461 171058 2350
rect 171915 2348 171916 2350
rect 171980 2348 171981 2412
rect 171915 2347 171981 2348
rect 170995 1460 171061 1461
rect 170995 1396 170996 1460
rect 171060 1396 171061 1460
rect 170995 1395 171061 1396
rect 175230 1189 175290 3030
rect 175598 1733 175658 7787
rect 175779 7444 175845 7445
rect 175779 7380 175780 7444
rect 175844 7380 175845 7444
rect 175779 7379 175845 7380
rect 175782 2413 175842 7379
rect 175966 2957 176026 8331
rect 176515 7580 176581 7581
rect 176515 7516 176516 7580
rect 176580 7516 176581 7580
rect 176515 7515 176581 7516
rect 176331 3500 176397 3501
rect 176331 3436 176332 3500
rect 176396 3436 176397 3500
rect 176331 3435 176397 3436
rect 175963 2956 176029 2957
rect 175963 2892 175964 2956
rect 176028 2892 176029 2956
rect 175963 2891 176029 2892
rect 175779 2412 175845 2413
rect 175779 2348 175780 2412
rect 175844 2348 175845 2412
rect 175779 2347 175845 2348
rect 176334 2277 176394 3435
rect 176518 2821 176578 7515
rect 177067 7444 177133 7445
rect 177067 7380 177068 7444
rect 177132 7380 177133 7444
rect 177067 7379 177133 7380
rect 177070 2957 177130 7379
rect 177067 2956 177133 2957
rect 177067 2892 177068 2956
rect 177132 2892 177133 2956
rect 177067 2891 177133 2892
rect 176515 2820 176581 2821
rect 176515 2756 176516 2820
rect 176580 2756 176581 2820
rect 176515 2755 176581 2756
rect 176331 2276 176397 2277
rect 176331 2212 176332 2276
rect 176396 2212 176397 2276
rect 176331 2211 176397 2212
rect 175595 1732 175661 1733
rect 175595 1668 175596 1732
rect 175660 1668 175661 1732
rect 175595 1667 175661 1668
rect 177622 1597 177682 8331
rect 184074 8208 184134 9200
rect 184071 8192 184137 8208
rect 184071 8128 184072 8192
rect 184136 8128 184137 8192
rect 184071 8112 184137 8128
rect 183507 7716 183573 7717
rect 183507 7652 183508 7716
rect 183572 7652 183573 7716
rect 183507 7651 183573 7652
rect 180747 7444 180813 7445
rect 180747 7380 180748 7444
rect 180812 7380 180813 7444
rect 180747 7379 180813 7380
rect 182035 7444 182101 7445
rect 182035 7380 182036 7444
rect 182100 7380 182101 7444
rect 182035 7379 182101 7380
rect 182219 7444 182285 7445
rect 182219 7380 182220 7444
rect 182284 7380 182285 7444
rect 182219 7379 182285 7380
rect 182403 7444 182469 7445
rect 182403 7380 182404 7444
rect 182468 7380 182469 7444
rect 182403 7379 182469 7380
rect 177803 7308 177869 7309
rect 177803 7244 177804 7308
rect 177868 7244 177869 7308
rect 177803 7243 177869 7244
rect 177806 2957 177866 7243
rect 177803 2956 177869 2957
rect 177803 2892 177804 2956
rect 177868 2892 177869 2956
rect 177803 2891 177869 2892
rect 180750 2549 180810 7379
rect 180747 2548 180813 2549
rect 180747 2484 180748 2548
rect 180812 2484 180813 2548
rect 180747 2483 180813 2484
rect 182038 2141 182098 7379
rect 182035 2140 182101 2141
rect 182035 2076 182036 2140
rect 182100 2076 182101 2140
rect 182035 2075 182101 2076
rect 177619 1596 177685 1597
rect 177619 1532 177620 1596
rect 177684 1532 177685 1596
rect 177619 1531 177685 1532
rect 182222 1325 182282 7379
rect 182406 7037 182466 7379
rect 182403 7036 182469 7037
rect 182403 6972 182404 7036
rect 182468 6972 182469 7036
rect 182403 6971 182469 6972
rect 183510 1597 183570 7651
rect 184074 2768 184134 8112
rect 184474 6017 184534 11579
rect 184471 6016 184537 6017
rect 184471 5952 184472 6016
rect 184536 5952 184537 6016
rect 184471 5951 184537 5952
rect 184474 4559 184534 5951
rect 184471 4558 184537 4559
rect 184471 4494 184472 4558
rect 184536 4494 184537 4558
rect 184471 4493 184537 4494
rect 184071 2752 184137 2768
rect 184071 2688 184072 2752
rect 184136 2688 184137 2752
rect 184071 2672 184137 2688
rect 184074 1680 184134 2672
rect 184071 1664 184137 1680
rect 184071 1600 184072 1664
rect 184136 1600 184137 1664
rect 183507 1596 183573 1597
rect 183507 1532 183508 1596
rect 183572 1532 183573 1596
rect 184071 1584 184137 1600
rect 183507 1531 183573 1532
rect 182219 1324 182285 1325
rect 182219 1260 182220 1324
rect 182284 1260 182285 1324
rect 182219 1259 182285 1260
rect 175227 1188 175293 1189
rect 175227 1124 175228 1188
rect 175292 1124 175293 1188
rect 175227 1123 175293 1124
rect 167131 100 167197 101
rect 167131 36 167132 100
rect 167196 36 167197 100
rect 167131 35 167197 36
rect 184074 -419 184134 1584
rect 184071 -420 184137 -419
rect 184071 -484 184072 -420
rect 184136 -484 184137 -420
rect 184071 -485 184137 -484
rect 184474 -699 184534 4493
rect 184471 -700 184537 -699
rect 184471 -764 184472 -700
rect 184536 -764 184537 -700
rect 184471 -765 184537 -764
rect 184874 -979 184934 11859
rect 185274 6468 185334 12139
rect 185674 6868 185734 12419
rect 201299 12344 201365 12345
rect 201299 12280 201300 12344
rect 201364 12280 201365 12344
rect 201299 12279 201365 12280
rect 201159 12204 201225 12205
rect 201159 12140 201160 12204
rect 201224 12140 201225 12204
rect 201159 12139 201225 12140
rect 201019 12064 201085 12065
rect 201019 12000 201020 12064
rect 201084 12000 201085 12064
rect 201019 11999 201085 12000
rect 200879 11924 200945 11925
rect 200879 11860 200880 11924
rect 200944 11860 200945 11924
rect 200879 11859 200945 11860
rect 200739 11784 200805 11785
rect 200739 11720 200740 11784
rect 200804 11720 200805 11784
rect 200739 11719 200805 11720
rect 200599 11644 200665 11645
rect 200599 11580 200600 11644
rect 200664 11580 200665 11644
rect 200599 11579 200665 11580
rect 200459 11504 200525 11505
rect 200459 11440 200460 11504
rect 200524 11440 200525 11504
rect 200459 11439 200525 11440
rect 200319 11364 200385 11365
rect 200319 11300 200320 11364
rect 200384 11300 200385 11364
rect 200319 11299 200385 11300
rect 200179 11224 200245 11225
rect 200179 11160 200180 11224
rect 200244 11160 200245 11224
rect 200179 11159 200245 11160
rect 185671 6867 185737 6868
rect 185671 6803 185672 6867
rect 185736 6803 185737 6867
rect 185671 6802 185737 6803
rect 185271 6467 185337 6468
rect 185271 6403 185272 6467
rect 185336 6403 185337 6467
rect 185271 6402 185337 6403
rect 185274 5010 185334 6402
rect 185674 5410 185734 6802
rect 185671 5409 185737 5410
rect 185671 5345 185672 5409
rect 185736 5345 185737 5409
rect 185671 5344 185737 5345
rect 185271 5009 185337 5010
rect 185271 4945 185272 5009
rect 185336 4945 185337 5009
rect 185271 4944 185337 4945
rect 184871 -980 184937 -979
rect 184871 -1044 184872 -980
rect 184936 -1044 184937 -980
rect 184871 -1045 184937 -1044
rect 185274 -1259 185334 4944
rect 185271 -1260 185337 -1259
rect 185271 -1324 185272 -1260
rect 185336 -1324 185337 -1260
rect 185271 -1325 185337 -1324
rect 165671 -1400 165737 -1399
rect 165671 -1464 165672 -1400
rect 165736 -1464 165737 -1400
rect 165671 -1465 165737 -1464
rect 145671 -1540 145737 -1539
rect 105671 -1605 105737 -1604
rect 145671 -1604 145672 -1540
rect 145736 -1604 145737 -1540
rect 165674 -1602 165734 -1465
rect 185674 -1539 185734 5344
rect 200182 -279 200242 11159
rect 200179 -280 200245 -279
rect 200179 -344 200180 -280
rect 200244 -344 200245 -280
rect 200179 -345 200245 -344
rect 200322 -419 200382 11299
rect 200319 -420 200385 -419
rect 200319 -484 200320 -420
rect 200384 -484 200385 -420
rect 200319 -485 200385 -484
rect 200462 -559 200522 11439
rect 200459 -560 200525 -559
rect 200459 -624 200460 -560
rect 200524 -624 200525 -560
rect 200459 -625 200525 -624
rect 200602 -699 200662 11579
rect 200599 -700 200665 -699
rect 200599 -764 200600 -700
rect 200664 -764 200665 -700
rect 200599 -765 200665 -764
rect 200742 -839 200802 11719
rect 200739 -840 200805 -839
rect 200739 -904 200740 -840
rect 200804 -904 200805 -840
rect 200739 -905 200805 -904
rect 200882 -979 200942 11859
rect 200879 -980 200945 -979
rect 200879 -1044 200880 -980
rect 200944 -1044 200945 -980
rect 200879 -1045 200945 -1044
rect 201022 -1119 201082 11999
rect 201019 -1120 201085 -1119
rect 201019 -1184 201020 -1120
rect 201084 -1184 201085 -1120
rect 201019 -1185 201085 -1184
rect 201162 -1259 201222 12139
rect 201159 -1260 201225 -1259
rect 201159 -1324 201160 -1260
rect 201224 -1324 201225 -1260
rect 201159 -1325 201225 -1324
rect 201302 -1399 201362 12279
rect 201299 -1400 201365 -1399
rect 201299 -1464 201300 -1400
rect 201364 -1464 201365 -1400
rect 201299 -1465 201365 -1464
rect 201442 -1539 201502 12419
rect 185671 -1540 185737 -1539
rect 145671 -1605 145737 -1604
rect 185671 -1604 185672 -1540
rect 185736 -1604 185737 -1540
rect 185671 -1605 185737 -1604
rect 201439 -1540 201505 -1539
rect 201439 -1604 201440 -1540
rect 201504 -1604 201505 -1540
rect 201439 -1605 201505 -1604
use mgmt_protect_hv  powergood_check
timestamp 1607567185
transform 1 0 156610 0 1 3035
box 0 1 40002 4205
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607567185
transform -1 0 198812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1607567185
transform 1 0 197892 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_2140
timestamp 1607567185
transform 1 0 197984 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_2127
timestamp 1607567185
transform 1 0 196788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[31\]
timestamp 1607567185
transform 1 0 195132 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1607567185
transform 1 0 195040 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2100
timestamp 1607567185
transform 1 0 194304 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[27\]
timestamp 1607567185
transform 1 0 192648 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1607567185
transform 1 0 192188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_2078
timestamp 1607567185
transform 1 0 192280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_2065
timestamp 1607567185
transform 1 0 191084 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[25\]
timestamp 1607567185
transform 1 0 189428 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1607567185
transform 1 0 189336 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_2045
timestamp 1607567185
transform 1 0 189244 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[20\]
timestamp 1607567185
transform 1 0 186852 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2037
timestamp 1607567185
transform 1 0 188508 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1607567185
transform 1 0 186484 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_2007
timestamp 1607567185
transform 1 0 185748 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_2016
timestamp 1607567185
transform 1 0 186576 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[29\]
timestamp 1607567185
transform 1 0 184092 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1607567185
transform 1 0 183632 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1985
timestamp 1607567185
transform 1 0 183724 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1976
timestamp 1607567185
transform 1 0 182896 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[30\]
timestamp 1607567185
transform 1 0 181240 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1607567185
transform 1 0 180780 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1945
timestamp 1607567185
transform 1 0 180044 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1954
timestamp 1607567185
transform 1 0 180872 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[33\]
timestamp 1607567185
transform 1 0 179768 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[35\]
timestamp 1607567185
transform 1 0 178756 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1934
timestamp 1607567185
transform 1 0 179032 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1607567185
transform 1 0 177928 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1913
timestamp 1607567185
transform 1 0 177100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1921
timestamp 1607567185
transform 1 0 177836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1923
timestamp 1607567185
transform 1 0 178020 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[13\]
timestamp 1607567185
transform 1 0 175444 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1607567185
transform 1 0 175076 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1892
timestamp 1607567185
transform 1 0 175168 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1879
timestamp 1607567185
transform 1 0 173972 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[8\]
timestamp 1607567185
transform 1 0 172316 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1607567185
transform 1 0 172224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1852
timestamp 1607567185
transform 1 0 171488 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[15\]
timestamp 1607567185
transform 1 0 169832 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1607567185
transform 1 0 169372 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1817
timestamp 1607567185
transform 1 0 168268 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1830
timestamp 1607567185
transform 1 0 169464 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[7\]
timestamp 1607567185
transform 1 0 166612 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1607567185
transform 1 0 166520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1786
timestamp 1607567185
transform 1 0 165416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[5\]
timestamp 1607567185
transform 1 0 163760 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[40\]
timestamp 1607567185
transform 1 0 162656 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1607567185
transform 1 0 163668 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1759
timestamp 1607567185
transform 1 0 162932 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[46\]
timestamp 1607567185
transform 1 0 161644 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1737
timestamp 1607567185
transform 1 0 160908 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1748
timestamp 1607567185
transform 1 0 161920 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1607567185
transform 1 0 197248 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607567185
transform -1 0 198812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_2135
timestamp 1607567185
transform 1 0 197524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_2143
timestamp 1607567185
transform 1 0 198260 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_2124
timestamp 1607567185
transform 1 0 196512 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[26\]
timestamp 1607567185
transform 1 0 194856 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607567185
transform 1 0 194764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_2104
timestamp 1607567185
transform 1 0 194672 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_2092
timestamp 1607567185
transform 1 0 193568 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[23\]
timestamp 1607567185
transform 1 0 191912 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_2066
timestamp 1607567185
transform 1 0 191176 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[22\]
timestamp 1607567185
transform 1 0 189520 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607567185
transform 1 0 189152 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_2045
timestamp 1607567185
transform 1 0 189244 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[32\]
timestamp 1607567185
transform 1 0 188140 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_2027
timestamp 1607567185
transform 1 0 187588 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_2036
timestamp 1607567185
transform 1 0 188416 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_2015
timestamp 1607567185
transform 1 0 186484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[20\]
timestamp 1607567185
transform 1 0 184828 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[27\]
timestamp 1607567185
transform 1 0 183632 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607567185
transform 1 0 183540 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1987
timestamp 1607567185
transform 1 0 183908 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1995
timestamp 1607567185
transform 1 0 184644 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1969
timestamp 1607567185
transform 1 0 182252 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1981
timestamp 1607567185
transform 1 0 183356 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[17\]
timestamp 1607567185
transform 1 0 180596 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[34\]
timestamp 1607567185
transform 1 0 179584 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1926
timestamp 1607567185
transform 1 0 178296 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1938
timestamp 1607567185
transform 1 0 179400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1943
timestamp 1607567185
transform 1 0 179860 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[22\]
timestamp 1607567185
transform 1 0 176824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[31\]
timestamp 1607567185
transform 1 0 178020 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607567185
transform 1 0 177928 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1907
timestamp 1607567185
transform 1 0 176548 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1913
timestamp 1607567185
transform 1 0 177100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1921
timestamp 1607567185
transform 1 0 177836 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1895
timestamp 1607567185
transform 1 0 175444 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[12\]
timestamp 1607567185
transform 1 0 173788 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1869
timestamp 1607567185
transform 1 0 173052 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[26\]
timestamp 1607567185
transform 1 0 172776 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607567185
transform 1 0 172316 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1853
timestamp 1607567185
transform 1 0 171580 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1862
timestamp 1607567185
transform 1 0 172408 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[12\]
timestamp 1607567185
transform 1 0 169924 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1834
timestamp 1607567185
transform 1 0 169832 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1826
timestamp 1607567185
transform 1 0 169096 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[4\]
timestamp 1607567185
transform 1 0 167440 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607567185
transform 1 0 166704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1801
timestamp 1607567185
transform 1 0 166796 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1807
timestamp 1607567185
transform 1 0 167348 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[14\]
timestamp 1607567185
transform 1 0 165324 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1777
timestamp 1607567185
transform 1 0 164588 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1788
timestamp 1607567185
transform 1 0 165600 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[4\]
timestamp 1607567185
transform 1 0 162932 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[41\]
timestamp 1607567185
transform 1 0 161920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607567185
transform 1 0 161092 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1740
timestamp 1607567185
transform 1 0 161184 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1751
timestamp 1607567185
transform 1 0 162196 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607567185
transform -1 0 198812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607567185
transform 1 0 197524 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2133
timestamp 1607567185
transform 1 0 197340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2136
timestamp 1607567185
transform 1 0 197616 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2144
timestamp 1607567185
transform 1 0 198352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1607567185
transform 1 0 195960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_2121
timestamp 1607567185
transform 1 0 196236 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2110
timestamp 1607567185
transform 1 0 195224 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[26\]
timestamp 1607567185
transform 1 0 193568 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_13_2078
timestamp 1607567185
transform 1 0 192280 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2090
timestamp 1607567185
transform 1 0 193384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1607567185
transform 1 0 192004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607567185
transform 1 0 191912 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_2058
timestamp 1607567185
transform 1 0 190440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2070
timestamp 1607567185
transform 1 0 191544 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[21\]
timestamp 1607567185
transform 1 0 188784 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2032
timestamp 1607567185
transform 1 0 188048 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[30\]
timestamp 1607567185
transform 1 0 186392 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607567185
transform 1 0 186300 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2005
timestamp 1607567185
transform 1 0 185564 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[29\]
timestamp 1607567185
transform 1 0 183908 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1986
timestamp 1607567185
transform 1 0 183816 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1978
timestamp 1607567185
transform 1 0 183080 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[18\]
timestamp 1607567185
transform 1 0 181424 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607567185
transform 1 0 180688 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1949
timestamp 1607567185
transform 1 0 180412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1953
timestamp 1607567185
transform 1 0 180780 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1959
timestamp 1607567185
transform 1 0 181332 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1937
timestamp 1607567185
transform 1 0 179308 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[17\]
timestamp 1607567185
transform 1 0 177652 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1911
timestamp 1607567185
transform 1 0 176916 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[13\]
timestamp 1607567185
transform 1 0 175260 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607567185
transform 1 0 175076 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1892
timestamp 1607567185
transform 1 0 175168 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[20\]
timestamp 1607567185
transform 1 0 174064 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[23\]
timestamp 1607567185
transform 1 0 173052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1872
timestamp 1607567185
transform 1 0 173328 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1883
timestamp 1607567185
transform 1 0 174340 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1861
timestamp 1607567185
transform 1 0 172316 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[10\]
timestamp 1607567185
transform 1 0 170660 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[36\]
timestamp 1607567185
transform 1 0 169648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1831
timestamp 1607567185
transform 1 0 169556 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1835
timestamp 1607567185
transform 1 0 169924 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[37\]
timestamp 1607567185
transform 1 0 168452 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607567185
transform 1 0 169464 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1816
timestamp 1607567185
transform 1 0 168176 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1822
timestamp 1607567185
transform 1 0 168728 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1808
timestamp 1607567185
transform 1 0 167440 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[19\]
timestamp 1607567185
transform 1 0 165784 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[15\]
timestamp 1607567185
transform 1 0 164496 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1779
timestamp 1607567185
transform 1 0 164772 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1787
timestamp 1607567185
transform 1 0 165508 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607567185
transform 1 0 163852 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1761
timestamp 1607567185
transform 1 0 163116 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1770
timestamp 1607567185
transform 1 0 163944 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[10\]
timestamp 1607567185
transform 1 0 161460 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1739
timestamp 1607567185
transform 1 0 161092 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1607567185
transform 1 0 197248 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607567185
transform -1 0 198812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_2135
timestamp 1607567185
transform 1 0 197524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_2143
timestamp 1607567185
transform 1 0 198260 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_2124
timestamp 1607567185
transform 1 0 196512 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[27\]
timestamp 1607567185
transform 1 0 194856 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607567185
transform 1 0 194764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_2101
timestamp 1607567185
transform 1 0 194396 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_2089
timestamp 1607567185
transform 1 0 193292 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[23\]
timestamp 1607567185
transform 1 0 191636 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_2063
timestamp 1607567185
transform 1 0 190900 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[31\]
timestamp 1607567185
transform 1 0 189244 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607567185
transform 1 0 189152 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2043
timestamp 1607567185
transform 1 0 189060 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _467_
timestamp 1607567185
transform 1 0 188048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_2024
timestamp 1607567185
transform 1 0 187312 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_2035
timestamp 1607567185
transform 1 0 188324 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[28\]
timestamp 1607567185
transform 1 0 185656 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_12_2003
timestamp 1607567185
transform 1 0 185380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[30\]
timestamp 1607567185
transform 1 0 184368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607567185
transform 1 0 183540 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1984
timestamp 1607567185
transform 1 0 183632 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1995
timestamp 1607567185
transform 1 0 184644 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1975
timestamp 1607567185
transform 1 0 182804 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[28\]
timestamp 1607567185
transform 1 0 181148 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1953
timestamp 1607567185
transform 1 0 180780 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1941
timestamp 1607567185
transform 1 0 179676 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[21\]
timestamp 1607567185
transform 1 0 178020 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607567185
transform 1 0 177928 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1907
timestamp 1607567185
transform 1 0 176548 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1919
timestamp 1607567185
transform 1 0 177652 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[16\]
timestamp 1607567185
transform 1 0 174892 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1888
timestamp 1607567185
transform 1 0 174800 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1880
timestamp 1607567185
transform 1 0 174064 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[6\]
timestamp 1607567185
transform 1 0 172408 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[18\]
timestamp 1607567185
transform 1 0 171304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607567185
transform 1 0 172316 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1853
timestamp 1607567185
transform 1 0 171580 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[16\]
timestamp 1607567185
transform 1 0 170108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1840
timestamp 1607567185
transform 1 0 170384 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1848
timestamp 1607567185
transform 1 0 171120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1829
timestamp 1607567185
transform 1 0 169372 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[18\]
timestamp 1607567185
transform 1 0 167716 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607567185
transform 1 0 166704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1801
timestamp 1607567185
transform 1 0 166796 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1809
timestamp 1607567185
transform 1 0 167532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1792
timestamp 1607567185
transform 1 0 165968 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[5\]
timestamp 1607567185
transform 1 0 164312 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[29\]
timestamp 1607567185
transform 1 0 163300 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1766
timestamp 1607567185
transform 1 0 163576 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[38\]
timestamp 1607567185
transform 1 0 162288 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[39\]
timestamp 1607567185
transform 1 0 161276 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607567185
transform 1 0 161092 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1738
timestamp 1607567185
transform 1 0 161000 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1740
timestamp 1607567185
transform 1 0 161184 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1744
timestamp 1607567185
transform 1 0 161552 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1755
timestamp 1607567185
transform 1 0 162564 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1607567185
transform 1 0 160816 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[49\]
timestamp 1607567185
transform 1 0 159804 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1717
timestamp 1607567185
transform 1 0 159068 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1728
timestamp 1607567185
transform 1 0 160080 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[54\]
timestamp 1607567185
transform 1 0 158792 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1607567185
transform 1 0 157964 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1706
timestamp 1607567185
transform 1 0 158056 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1693
timestamp 1607567185
transform 1 0 156860 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[8\]
timestamp 1607567185
transform 1 0 155204 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1607567185
transform 1 0 155112 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1662
timestamp 1607567185
transform 1 0 154008 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_sel_buf\[3\]
timestamp 1607567185
transform 1 0 152352 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1607567185
transform 1 0 152260 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[72\]
timestamp 1607567185
transform 1 0 151248 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1628
timestamp 1607567185
transform 1 0 150880 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1635
timestamp 1607567185
transform 1 0 151524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[8\]
timestamp 1607567185
transform 1 0 149500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1607567185
transform 1 0 149408 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1608
timestamp 1607567185
transform 1 0 149040 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1616
timestamp 1607567185
transform 1 0 149776 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[4\]
timestamp 1607567185
transform 1 0 147660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1585
timestamp 1607567185
transform 1 0 146924 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1596
timestamp 1607567185
transform 1 0 147936 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[326\]
timestamp 1607567185
transform 1 0 146648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1607567185
transform 1 0 146556 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1577
timestamp 1607567185
transform 1 0 146188 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[446\]
timestamp 1607567185
transform 1 0 143796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[448\]
timestamp 1607567185
transform 1 0 144808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1607567185
transform 1 0 143704 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1554
timestamp 1607567185
transform 1 0 144072 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1565
timestamp 1607567185
transform 1 0 145084 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[325\]
timestamp 1607567185
transform 1 0 141956 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1534
timestamp 1607567185
transform 1 0 142232 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1546
timestamp 1607567185
transform 1 0 143336 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[320\]
timestamp 1607567185
transform 1 0 140944 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1607567185
transform 1 0 140852 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1515
timestamp 1607567185
transform 1 0 140484 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1523
timestamp 1607567185
transform 1 0 141220 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[312\]
timestamp 1607567185
transform 1 0 139104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1492
timestamp 1607567185
transform 1 0 138368 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1503
timestamp 1607567185
transform 1 0 139380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[309\]
timestamp 1607567185
transform 1 0 138092 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1607567185
transform 1 0 138000 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1472
timestamp 1607567185
transform 1 0 136528 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1484
timestamp 1607567185
transform 1 0 137632 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[305\]
timestamp 1607567185
transform 1 0 135240 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[307\]
timestamp 1607567185
transform 1 0 136252 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1607567185
transform 1 0 135148 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1453
timestamp 1607567185
transform 1 0 134780 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1461
timestamp 1607567185
transform 1 0 135516 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[301\]
timestamp 1607567185
transform 1 0 133400 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1441
timestamp 1607567185
transform 1 0 133676 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[300\]
timestamp 1607567185
transform 1 0 132388 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1607567185
transform 1 0 132296 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1430
timestamp 1607567185
transform 1 0 132664 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1414
timestamp 1607567185
transform 1 0 131192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[118\]
timestamp 1607567185
transform 1 0 129536 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1607567185
transform 1 0 129444 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1387
timestamp 1607567185
transform 1 0 128708 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[98\]
timestamp 1607567185
transform 1 0 127052 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1607567185
transform 1 0 126592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1363
timestamp 1607567185
transform 1 0 126500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1365
timestamp 1607567185
transform 1 0 126684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1355
timestamp 1607567185
transform 1 0 125764 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[296\]
timestamp 1607567185
transform 1 0 122728 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[94\]
timestamp 1607567185
transform 1 0 124108 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1607567185
transform 1 0 123740 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1325
timestamp 1607567185
transform 1 0 123004 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_1334
timestamp 1607567185
transform 1 0 123832 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[298\]
timestamp 1607567185
transform 1 0 120980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1306
timestamp 1607567185
transform 1 0 121256 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1318
timestamp 1607567185
transform 1 0 122360 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[47\]
timestamp 1607567185
transform 1 0 160080 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[52\]
timestamp 1607567185
transform 1 0 159068 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1720
timestamp 1607567185
transform 1 0 159344 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1731
timestamp 1607567185
transform 1 0 160356 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[43\]
timestamp 1607567185
transform 1 0 157964 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1708
timestamp 1607567185
transform 1 0 158240 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1716
timestamp 1607567185
transform 1 0 158976 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1697
timestamp 1607567185
transform 1 0 157228 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[2\]
timestamp 1607567185
transform 1 0 155572 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607567185
transform 1 0 155480 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1670
timestamp 1607567185
transform 1 0 154744 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[1\]
timestamp 1607567185
transform 1 0 153088 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1644
timestamp 1607567185
transform 1 0 152352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[62\]
timestamp 1607567185
transform 1 0 152076 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[65\]
timestamp 1607567185
transform 1 0 151064 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1629
timestamp 1607567185
transform 1 0 150972 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1633
timestamp 1607567185
transform 1 0 151340 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[5\]
timestamp 1607567185
transform 1 0 149960 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607567185
transform 1 0 149868 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1613
timestamp 1607567185
transform 1 0 149500 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1621
timestamp 1607567185
transform 1 0 150236 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1601
timestamp 1607567185
transform 1 0 148396 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_we_buf
timestamp 1607567185
transform 1 0 146740 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1575
timestamp 1607567185
transform 1 0 146004 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_stb_buf
timestamp 1607567185
transform 1 0 144348 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607567185
transform 1 0 144256 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1555
timestamp 1607567185
transform 1 0 144164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[323\]
timestamp 1607567185
transform 1 0 142140 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[327\]
timestamp 1607567185
transform 1 0 143152 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1536
timestamp 1607567185
transform 1 0 142416 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1547
timestamp 1607567185
transform 1 0 143428 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[319\]
timestamp 1607567185
transform 1 0 141128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1514
timestamp 1607567185
transform 1 0 140392 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1525
timestamp 1607567185
transform 1 0 141404 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[125\]
timestamp 1607567185
transform 1 0 138736 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607567185
transform 1 0 138644 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1491
timestamp 1607567185
transform 1 0 138276 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[308\]
timestamp 1607567185
transform 1 0 136896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1479
timestamp 1607567185
transform 1 0 137172 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1468
timestamp 1607567185
transform 1 0 136160 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[292\]
timestamp 1607567185
transform 1 0 133124 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[123\]
timestamp 1607567185
transform 1 0 134504 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1438
timestamp 1607567185
transform 1 0 133400 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[277\]
timestamp 1607567185
transform 1 0 131836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607567185
transform 1 0 133032 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1424
timestamp 1607567185
transform 1 0 132112 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1432
timestamp 1607567185
transform 1 0 132848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[274\]
timestamp 1607567185
transform 1 0 130824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1402
timestamp 1607567185
transform 1 0 130088 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1413
timestamp 1607567185
transform 1 0 131100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[105\]
timestamp 1607567185
transform 1 0 128432 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1382
timestamp 1607567185
transform 1 0 128248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607567185
transform 1 0 127420 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1370
timestamp 1607567185
transform 1 0 127144 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1374
timestamp 1607567185
transform 1 0 127512 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[103\]
timestamp 1607567185
transform 1 0 124384 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1358
timestamp 1607567185
transform 1 0 126040 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1331
timestamp 1607567185
transform 1 0 123556 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1339
timestamp 1607567185
transform 1 0 124292 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[39\]
timestamp 1607567185
transform 1 0 121900 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607567185
transform 1 0 121808 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1309
timestamp 1607567185
transform 1 0 121532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1727
timestamp 1607567185
transform 1 0 159988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[126\]
timestamp 1607567185
transform 1 0 158332 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607567185
transform 1 0 158240 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1700
timestamp 1607567185
transform 1 0 157504 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[12\]
timestamp 1607567185
transform 1 0 156216 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[328\]
timestamp 1607567185
transform 1 0 157228 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1689
timestamp 1607567185
transform 1 0 156492 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1678
timestamp 1607567185
transform 1 0 155480 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[9\]
timestamp 1607567185
transform 1 0 153824 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[11\]
timestamp 1607567185
transform 1 0 152812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607567185
transform 1 0 152628 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1648
timestamp 1607567185
transform 1 0 152720 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1652
timestamp 1607567185
transform 1 0 153088 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[50\]
timestamp 1607567185
transform 1 0 151616 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[68\]
timestamp 1607567185
transform 1 0 150604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1628
timestamp 1607567185
transform 1 0 150880 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1639
timestamp 1607567185
transform 1 0 151892 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[73\]
timestamp 1607567185
transform 1 0 149592 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1606
timestamp 1607567185
transform 1 0 148856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1617
timestamp 1607567185
transform 1 0 149868 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_sel_buf\[2\]
timestamp 1607567185
transform 1 0 147200 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607567185
transform 1 0 147016 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1587
timestamp 1607567185
transform 1 0 147108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1578
timestamp 1607567185
transform 1 0 146280 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[443\]
timestamp 1607567185
transform 1 0 143520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[124\]
timestamp 1607567185
transform 1 0 144624 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1551
timestamp 1607567185
transform 1 0 143796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1559
timestamp 1607567185
transform 1 0 144532 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[322\]
timestamp 1607567185
transform 1 0 142508 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1529
timestamp 1607567185
transform 1 0 141772 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1540
timestamp 1607567185
transform 1 0 142784 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[317\]
timestamp 1607567185
transform 1 0 141496 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607567185
transform 1 0 141404 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1516
timestamp 1607567185
transform 1 0 140576 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1524
timestamp 1607567185
transform 1 0 141312 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[121\]
timestamp 1607567185
transform 1 0 138920 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[120\]
timestamp 1607567185
transform 1 0 136528 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1490
timestamp 1607567185
transform 1 0 138184 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607567185
transform 1 0 135792 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1456
timestamp 1607567185
transform 1 0 135056 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1465
timestamp 1607567185
transform 1 0 135884 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1471
timestamp 1607567185
transform 1 0 136436 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[107\]
timestamp 1607567185
transform 1 0 133400 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1430
timestamp 1607567185
transform 1 0 132664 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[110\]
timestamp 1607567185
transform 1 0 131008 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607567185
transform 1 0 130180 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1404
timestamp 1607567185
transform 1 0 130272 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1395
timestamp 1607567185
transform 1 0 129444 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[75\]
timestamp 1607567185
transform 1 0 127788 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1366
timestamp 1607567185
transform 1 0 126776 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1374
timestamp 1607567185
transform 1 0 127512 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[106\]
timestamp 1607567185
transform 1 0 125120 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607567185
transform 1 0 124568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1343
timestamp 1607567185
transform 1 0 124660 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1347
timestamp 1607567185
transform 1 0 125028 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[266\]
timestamp 1607567185
transform 1 0 123556 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1328
timestamp 1607567185
transform 1 0 123280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1334
timestamp 1607567185
transform 1 0 123832 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[291\]
timestamp 1607567185
transform 1 0 122268 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[297\]
timestamp 1607567185
transform 1 0 121256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1309
timestamp 1607567185
transform 1 0 121532 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1320
timestamp 1607567185
transform 1 0 122544 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1730
timestamp 1607567185
transform 1 0 160264 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[1\]
timestamp 1607567185
transform 1 0 158608 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1709
timestamp 1607567185
transform 1 0 158332 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1697
timestamp 1607567185
transform 1 0 157228 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_cyc_buf
timestamp 1607567185
transform 1 0 155572 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607567185
transform 1 0 155480 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1670
timestamp 1607567185
transform 1 0 154744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[0\]
timestamp 1607567185
transform 1 0 153088 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1644
timestamp 1607567185
transform 1 0 152352 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[3\]
timestamp 1607567185
transform 1 0 152076 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[51\]
timestamp 1607567185
transform 1 0 151064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1633
timestamp 1607567185
transform 1 0 151340 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[71\]
timestamp 1607567185
transform 1 0 150052 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607567185
transform 1 0 149868 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1614
timestamp 1607567185
transform 1 0 149592 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1618
timestamp 1607567185
transform 1 0 149960 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1622
timestamp 1607567185
transform 1 0 150328 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[324\]
timestamp 1607567185
transform 1 0 148212 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1591
timestamp 1607567185
transform 1 0 147476 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1602
timestamp 1607567185
transform 1 0 148488 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[116\]
timestamp 1607567185
transform 1 0 145820 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1572
timestamp 1607567185
transform 1 0 145728 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[444\]
timestamp 1607567185
transform 1 0 144348 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607567185
transform 1 0 144256 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1553
timestamp 1607567185
transform 1 0 143980 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1560
timestamp 1607567185
transform 1 0 144624 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[314\]
timestamp 1607567185
transform 1 0 142600 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1537
timestamp 1607567185
transform 1 0 142508 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1541
timestamp 1607567185
transform 1 0 142876 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[315\]
timestamp 1607567185
transform 1 0 141128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1514
timestamp 1607567185
transform 1 0 140392 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1525
timestamp 1607567185
transform 1 0 141404 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[115\]
timestamp 1607567185
transform 1 0 138736 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1607567185
transform 1 0 138644 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1494
timestamp 1607567185
transform 1 0 138552 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[303\]
timestamp 1607567185
transform 1 0 136528 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[306\]
timestamp 1607567185
transform 1 0 137540 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1475
timestamp 1607567185
transform 1 0 136804 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1486
timestamp 1607567185
transform 1 0 137816 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[302\]
timestamp 1607567185
transform 1 0 135516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1453
timestamp 1607567185
transform 1 0 134780 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1464
timestamp 1607567185
transform 1 0 135792 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[101\]
timestamp 1607567185
transform 1 0 133124 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607567185
transform 1 0 133032 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1423
timestamp 1607567185
transform 1 0 132020 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1431
timestamp 1607567185
transform 1 0 132756 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[100\]
timestamp 1607567185
transform 1 0 130364 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1404
timestamp 1607567185
transform 1 0 130272 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1392
timestamp 1607567185
transform 1 0 129168 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[117\]
timestamp 1607567185
transform 1 0 127512 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607567185
transform 1 0 127420 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1369
timestamp 1607567185
transform 1 0 127052 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[13\]
timestamp 1607567185
transform 1 0 125672 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1346
timestamp 1607567185
transform 1 0 124936 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1357
timestamp 1607567185
transform 1 0 125948 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[89\]
timestamp 1607567185
transform 1 0 123280 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1325
timestamp 1607567185
transform 1 0 123004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[261\]
timestamp 1607567185
transform 1 0 121992 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607567185
transform 1 0 121808 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1308
timestamp 1607567185
transform 1 0 121440 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1313
timestamp 1607567185
transform 1 0 121900 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1317
timestamp 1607567185
transform 1 0 122268 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607567185
transform -1 0 154560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[19\]
timestamp 1607567185
transform 1 0 152904 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607567185
transform 1 0 152628 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1648
timestamp 1607567185
transform 1 0 152720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1653
timestamp 1607567185
transform 1 0 153180 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1639
timestamp 1607567185
transform 1 0 151892 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_sel_buf\[0\]
timestamp 1607567185
transform 1 0 150236 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1611
timestamp 1607567185
transform 1 0 149316 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1619
timestamp 1607567185
transform 1 0 150052 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[7\]
timestamp 1607567185
transform 1 0 147660 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607567185
transform 1 0 147016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1585
timestamp 1607567185
transform 1 0 146924 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1587
timestamp 1607567185
transform 1 0 147108 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[318\]
timestamp 1607567185
transform 1 0 145912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1571
timestamp 1607567185
transform 1 0 145636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1577
timestamp 1607567185
transform 1 0 146188 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[447\]
timestamp 1607567185
transform 1 0 144624 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1552
timestamp 1607567185
transform 1 0 143888 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1563
timestamp 1607567185
transform 1 0 144900 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[112\]
timestamp 1607567185
transform 1 0 142232 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1607567185
transform 1 0 141404 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1517
timestamp 1607567185
transform 1 0 140668 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1526
timestamp 1607567185
transform 1 0 141496 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[127\]
timestamp 1607567185
transform 1 0 139012 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1495
timestamp 1607567185
transform 1 0 138644 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1483
timestamp 1607567185
transform 1 0 137540 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[109\]
timestamp 1607567185
transform 1 0 135884 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607567185
transform 1 0 135792 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1455
timestamp 1607567185
transform 1 0 134964 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1463
timestamp 1607567185
transform 1 0 135700 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[267\]
timestamp 1607567185
transform 1 0 133676 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[283\]
timestamp 1607567185
transform 1 0 134688 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1444
timestamp 1607567185
transform 1 0 133952 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1433
timestamp 1607567185
transform 1 0 132940 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[3\]
timestamp 1607567185
transform 1 0 131284 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[256\]
timestamp 1607567185
transform 1 0 130272 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607567185
transform 1 0 130180 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1401
timestamp 1607567185
transform 1 0 129996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1407
timestamp 1607567185
transform 1 0 130548 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[252\]
timestamp 1607567185
transform 1 0 128616 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1378
timestamp 1607567185
transform 1 0 127880 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1389
timestamp 1607567185
transform 1 0 128892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[64\]
timestamp 1607567185
transform 1 0 126224 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[10\]
timestamp 1607567185
transform 1 0 125212 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607567185
transform 1 0 124568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1343
timestamp 1607567185
transform 1 0 124660 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1352
timestamp 1607567185
transform 1 0 125488 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[253\]
timestamp 1607567185
transform 1 0 123556 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1329
timestamp 1607567185
transform 1 0 123372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1334
timestamp 1607567185
transform 1 0 123832 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1317
timestamp 1607567185
transform 1 0 122268 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607567185
transform -1 0 154560 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607567185
transform -1 0 154560 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1663
timestamp 1607567185
transform 1 0 154100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[42\]
timestamp 1607567185
transform 1 0 153272 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607567185
transform 1 0 152628 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1648
timestamp 1607567185
transform 1 0 152720 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1657
timestamp 1607567185
transform 1 0 153548 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1655
timestamp 1607567185
transform 1 0 153364 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[9\]
timestamp 1607567185
transform 1 0 151708 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[69\]
timestamp 1607567185
transform 1 0 151616 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[6\]
timestamp 1607567185
transform 1 0 150696 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[9\]
timestamp 1607567185
transform 1 0 150604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1628
timestamp 1607567185
transform 1 0 150880 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1639
timestamp 1607567185
transform 1 0 151892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1629
timestamp 1607567185
transform 1 0 150972 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607567185
transform 1 0 149868 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1614
timestamp 1607567185
transform 1 0 149592 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1622
timestamp 1607567185
transform 1 0 150328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1614
timestamp 1607567185
transform 1 0 149592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1618
timestamp 1607567185
transform 1 0 149960 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[17\]
timestamp 1607567185
transform 1 0 147108 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607567185
transform 1 0 147016 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1590
timestamp 1607567185
transform 1 0 147384 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1602
timestamp 1607567185
transform 1 0 148488 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1602
timestamp 1607567185
transform 1 0 148488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[454\]
timestamp 1607567185
transform 1 0 145360 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[122\]
timestamp 1607567185
transform 1 0 146832 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1570
timestamp 1607567185
transform 1 0 145544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1582
timestamp 1607567185
transform 1 0 146648 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1571
timestamp 1607567185
transform 1 0 145636 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1583
timestamp 1607567185
transform 1 0 146740 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[14\]
timestamp 1607567185
transform 1 0 143888 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[450\]
timestamp 1607567185
transform 1 0 144348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607567185
transform 1 0 144256 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1554
timestamp 1607567185
transform 1 0 144072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1560
timestamp 1607567185
transform 1 0 144624 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[329\]
timestamp 1607567185
transform 1 0 142508 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1529
timestamp 1607567185
transform 1 0 141772 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1540
timestamp 1607567185
transform 1 0 142784 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1542
timestamp 1607567185
transform 1 0 142968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[313\]
timestamp 1607567185
transform 1 0 141496 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[113\]
timestamp 1607567185
transform 1 0 141312 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607567185
transform 1 0 141404 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1511
timestamp 1607567185
transform 1 0 140116 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1523
timestamp 1607567185
transform 1 0 141220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1510
timestamp 1607567185
transform 1 0 140024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1522
timestamp 1607567185
transform 1 0 141128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[310\]
timestamp 1607567185
transform 1 0 138736 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[311\]
timestamp 1607567185
transform 1 0 139748 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[84\]
timestamp 1607567185
transform 1 0 138460 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607567185
transform 1 0 138644 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1494
timestamp 1607567185
transform 1 0 138552 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1499
timestamp 1607567185
transform 1 0 139012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[286\]
timestamp 1607567185
transform 1 0 136528 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[304\]
timestamp 1607567185
transform 1 0 137540 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1485
timestamp 1607567185
transform 1 0 137724 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1475
timestamp 1607567185
transform 1 0 136804 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1486
timestamp 1607567185
transform 1 0 137816 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[269\]
timestamp 1607567185
transform 1 0 134780 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[111\]
timestamp 1607567185
transform 1 0 136068 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607567185
transform 1 0 135792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1456
timestamp 1607567185
transform 1 0 135056 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1465
timestamp 1607567185
transform 1 0 135884 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1464
timestamp 1607567185
transform 1 0 135792 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[262\]
timestamp 1607567185
transform 1 0 133768 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[263\]
timestamp 1607567185
transform 1 0 133124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[104\]
timestamp 1607567185
transform 1 0 134136 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1445
timestamp 1607567185
transform 1 0 134044 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1438
timestamp 1607567185
transform 1 0 133400 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[108\]
timestamp 1607567185
transform 1 0 131376 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607567185
transform 1 0 133032 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1434
timestamp 1607567185
transform 1 0 133032 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1422
timestamp 1607567185
transform 1 0 131928 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[21\]
timestamp 1607567185
transform 1 0 130272 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[114\]
timestamp 1607567185
transform 1 0 130272 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607567185
transform 1 0 130180 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1400
timestamp 1607567185
transform 1 0 129904 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1407
timestamp 1607567185
transform 1 0 130548 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1415
timestamp 1607567185
transform 1 0 131284 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[72\]
timestamp 1607567185
transform 1 0 127880 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1388
timestamp 1607567185
transform 1 0 128800 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1396
timestamp 1607567185
transform 1 0 129536 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[57\]
timestamp 1607567185
transform 1 0 127144 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607567185
transform 1 0 127420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1361
timestamp 1607567185
transform 1 0 126316 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1369
timestamp 1607567185
transform 1 0 127052 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1360
timestamp 1607567185
transform 1 0 126224 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1372
timestamp 1607567185
transform 1 0 127328 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1374
timestamp 1607567185
transform 1 0 127512 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[95\]
timestamp 1607567185
transform 1 0 124568 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[96\]
timestamp 1607567185
transform 1 0 124660 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607567185
transform 1 0 124568 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1340
timestamp 1607567185
transform 1 0 124384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1326
timestamp 1607567185
transform 1 0 123096 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1338
timestamp 1607567185
transform 1 0 124200 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1332
timestamp 1607567185
transform 1 0 123648 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[62\]
timestamp 1607567185
transform 1 0 121992 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[93\]
timestamp 1607567185
transform 1 0 121440 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607567185
transform 1 0 121808 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1308
timestamp 1607567185
transform 1 0 121440 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1313
timestamp 1607567185
transform 1 0 121900 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607567185
transform -1 0 154560 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1657
timestamp 1607567185
transform 1 0 153548 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[16\]
timestamp 1607567185
transform 1 0 151892 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1630
timestamp 1607567185
transform 1 0 151064 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1638
timestamp 1607567185
transform 1 0 151800 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607567185
transform 1 0 149868 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1607
timestamp 1607567185
transform 1 0 148948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1615
timestamp 1607567185
transform 1 0 149684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1618
timestamp 1607567185
transform 1 0 149960 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1595
timestamp 1607567185
transform 1 0 147844 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[56\]
timestamp 1607567185
transform 1 0 145360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1571
timestamp 1607567185
transform 1 0 145636 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1583
timestamp 1607567185
transform 1 0 146740 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[45\]
timestamp 1607567185
transform 1 0 144348 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607567185
transform 1 0 144256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1548
timestamp 1607567185
transform 1 0 143520 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1560
timestamp 1607567185
transform 1 0 144624 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[24\]
timestamp 1607567185
transform 1 0 143244 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[445\]
timestamp 1607567185
transform 1 0 142140 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1536
timestamp 1607567185
transform 1 0 142416 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1544
timestamp 1607567185
transform 1 0 143152 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[316\]
timestamp 1607567185
transform 1 0 141128 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1514
timestamp 1607567185
transform 1 0 140392 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1525
timestamp 1607567185
transform 1 0 141404 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[87\]
timestamp 1607567185
transform 1 0 138736 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607567185
transform 1 0 138644 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1491
timestamp 1607567185
transform 1 0 138276 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1479
timestamp 1607567185
transform 1 0 137172 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[102\]
timestamp 1607567185
transform 1 0 135516 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1453
timestamp 1607567185
transform 1 0 134780 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[11\]
timestamp 1607567185
transform 1 0 133124 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607567185
transform 1 0 133032 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1426
timestamp 1607567185
transform 1 0 132296 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[119\]
timestamp 1607567185
transform 1 0 130640 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1405
timestamp 1607567185
transform 1 0 130364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1393
timestamp 1607567185
transform 1 0 129260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _655_
timestamp 1607567185
transform 1 0 126408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[3\]
timestamp 1607567185
transform 1 0 127604 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607567185
transform 1 0 127420 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1365
timestamp 1607567185
transform 1 0 126684 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1374
timestamp 1607567185
transform 1 0 127512 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1344
timestamp 1607567185
transform 1 0 124752 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1356
timestamp 1607567185
transform 1 0 125856 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[59\]
timestamp 1607567185
transform 1 0 123096 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[237\]
timestamp 1607567185
transform 1 0 122084 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607567185
transform 1 0 121808 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1304
timestamp 1607567185
transform 1 0 121072 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1313
timestamp 1607567185
transform 1 0 121900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1318
timestamp 1607567185
transform 1 0 122360 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1607567185
transform 1 0 120888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1290
timestamp 1607567185
transform 1 0 119784 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[97\]
timestamp 1607567185
transform 1 0 118128 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1607567185
transform 1 0 118036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1267
timestamp 1607567185
transform 1 0 117668 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[290\]
timestamp 1607567185
transform 1 0 116288 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1255
timestamp 1607567185
transform 1 0 116564 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[273\]
timestamp 1607567185
transform 1 0 115276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1607567185
transform 1 0 115184 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1228
timestamp 1607567185
transform 1 0 114080 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1244
timestamp 1607567185
transform 1 0 115552 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[92\]
timestamp 1607567185
transform 1 0 112424 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1607567185
transform 1 0 112332 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1201
timestamp 1607567185
transform 1 0 111596 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[91\]
timestamp 1607567185
transform 1 0 109940 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1607567185
transform 1 0 109480 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1170
timestamp 1607567185
transform 1 0 108744 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1179
timestamp 1607567185
transform 1 0 109572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[287\]
timestamp 1607567185
transform 1 0 108468 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[293\]
timestamp 1607567185
transform 1 0 107456 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1159
timestamp 1607567185
transform 1 0 107732 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1607567185
transform 1 0 106628 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1143
timestamp 1607567185
transform 1 0 106260 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1148
timestamp 1607567185
transform 1 0 106720 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[433\]
timestamp 1607567185
transform 1 0 103868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[435\]
timestamp 1607567185
transform 1 0 104880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1607567185
transform 1 0 103776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1120
timestamp 1607567185
transform 1 0 104144 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1131
timestamp 1607567185
transform 1 0 105156 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[429\]
timestamp 1607567185
transform 1 0 102028 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1100
timestamp 1607567185
transform 1 0 102304 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1112
timestamp 1607567185
transform 1 0 103408 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[427\]
timestamp 1607567185
transform 1 0 101016 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1607567185
transform 1 0 100924 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1081
timestamp 1607567185
transform 1 0 100556 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1089
timestamp 1607567185
transform 1 0 101292 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[416\]
timestamp 1607567185
transform 1 0 99176 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1058
timestamp 1607567185
transform 1 0 98440 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1069
timestamp 1607567185
transform 1 0 99452 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[268\]
timestamp 1607567185
transform 1 0 96876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[275\]
timestamp 1607567185
transform 1 0 98164 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1607567185
transform 1 0 98072 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1044
timestamp 1607567185
transform 1 0 97152 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1052
timestamp 1607567185
transform 1 0 97888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[97\]
timestamp 1607567185
transform 1 0 95312 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1607567185
transform 1 0 95220 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1033
timestamp 1607567185
transform 1 0 96140 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1015
timestamp 1607567185
transform 1 0 94484 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[78\]
timestamp 1607567185
transform 1 0 92828 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1607567185
transform 1 0 92368 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_983
timestamp 1607567185
transform 1 0 91540 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_991
timestamp 1607567185
transform 1 0 92276 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_993
timestamp 1607567185
transform 1 0 92460 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[280\]
timestamp 1607567185
transform 1 0 91264 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_965
timestamp 1607567185
transform 1 0 89884 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_977
timestamp 1607567185
transform 1 0 90988 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[410\]
timestamp 1607567185
transform 1 0 89608 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1607567185
transform 1 0 89516 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_945
timestamp 1607567185
transform 1 0 88044 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_957
timestamp 1607567185
transform 1 0 89148 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[403\]
timestamp 1607567185
transform 1 0 86756 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[406\]
timestamp 1607567185
transform 1 0 87768 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1607567185
transform 1 0 86664 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_926
timestamp 1607567185
transform 1 0 86296 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_934
timestamp 1607567185
transform 1 0 87032 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[398\]
timestamp 1607567185
transform 1 0 84916 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_914
timestamp 1607567185
transform 1 0 85192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[392\]
timestamp 1607567185
transform 1 0 83904 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1607567185
transform 1 0 83812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_889
timestamp 1607567185
transform 1 0 82892 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_897
timestamp 1607567185
transform 1 0 83628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_903
timestamp 1607567185
transform 1 0 84180 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[389\]
timestamp 1607567185
transform 1 0 82616 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[73\]
timestamp 1607567185
transform 1 0 81052 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_878
timestamp 1607567185
transform 1 0 81880 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[241\]
timestamp 1607567185
transform 1 0 120520 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1290
timestamp 1607567185
transform 1 0 119784 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1301
timestamp 1607567185
transform 1 0 120796 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[69\]
timestamp 1607567185
transform 1 0 118128 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1264
timestamp 1607567185
transform 1 0 117392 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[271\]
timestamp 1607567185
transform 1 0 117116 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607567185
transform 1 0 116196 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1246
timestamp 1607567185
transform 1 0 115736 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1250
timestamp 1607567185
transform 1 0 116104 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1252
timestamp 1607567185
transform 1 0 116288 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1260
timestamp 1607567185
transform 1 0 117024 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1234
timestamp 1607567185
transform 1 0 114632 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[80\]
timestamp 1607567185
transform 1 0 112976 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1212
timestamp 1607567185
transform 1 0 112608 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[116\]
timestamp 1607567185
transform 1 0 110676 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607567185
transform 1 0 110584 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1200
timestamp 1607567185
transform 1 0 111504 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[282\]
timestamp 1607567185
transform 1 0 109572 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1182
timestamp 1607567185
transform 1 0 109848 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[113\]
timestamp 1607567185
transform 1 0 107640 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1167
timestamp 1607567185
transform 1 0 108468 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[278\]
timestamp 1607567185
transform 1 0 106628 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[294\]
timestamp 1607567185
transform 1 0 105616 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1139
timestamp 1607567185
transform 1 0 105892 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1150
timestamp 1607567185
transform 1 0 106904 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607567185
transform 1 0 104972 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1123
timestamp 1607567185
transform 1 0 104420 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1130
timestamp 1607567185
transform 1 0 105064 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[284\]
timestamp 1607567185
transform 1 0 102028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[430\]
timestamp 1607567185
transform 1 0 103040 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_1095
timestamp 1607567185
transform 1 0 101844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1100
timestamp 1607567185
transform 1 0 102304 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1111
timestamp 1607567185
transform 1 0 103316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[417\]
timestamp 1607567185
transform 1 0 100464 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1083
timestamp 1607567185
transform 1 0 100740 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[206\]
timestamp 1607567185
transform 1 0 99452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607567185
transform 1 0 99360 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1059
timestamp 1607567185
transform 1 0 98532 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1067
timestamp 1607567185
transform 1 0 99268 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1072
timestamp 1607567185
transform 1 0 99728 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[99\]
timestamp 1607567185
transform 1 0 97704 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1042
timestamp 1607567185
transform 1 0 96968 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[74\]
timestamp 1607567185
transform 1 0 95312 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1023
timestamp 1607567185
transform 1 0 95220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[276\]
timestamp 1607567185
transform 1 0 93840 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607567185
transform 1 0 93748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1003
timestamp 1607567185
transform 1 0 93380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1011
timestamp 1607567185
transform 1 0 94116 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[86\]
timestamp 1607567185
transform 1 0 91448 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_991
timestamp 1607567185
transform 1 0 92276 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[409\]
timestamp 1607567185
transform 1 0 90344 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_969
timestamp 1607567185
transform 1 0 90252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_973
timestamp 1607567185
transform 1 0 90620 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_981
timestamp 1607567185
transform 1 0 91356 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[404\]
timestamp 1607567185
transform 1 0 88228 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[407\]
timestamp 1607567185
transform 1 0 89240 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607567185
transform 1 0 88136 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_950
timestamp 1607567185
transform 1 0 88504 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_961
timestamp 1607567185
transform 1 0 89516 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[401\]
timestamp 1607567185
transform 1 0 86756 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_934
timestamp 1607567185
transform 1 0 87032 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_923
timestamp 1607567185
transform 1 0 86020 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[49\]
timestamp 1607567185
transform 1 0 84364 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_14_889
timestamp 1607567185
transform 1 0 82892 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_901
timestamp 1607567185
transform 1 0 83996 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[384\]
timestamp 1607567185
transform 1 0 82616 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[388\]
timestamp 1607567185
transform 1 0 81052 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607567185
transform 1 0 82524 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_872
timestamp 1607567185
transform 1 0 81328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_884
timestamp 1607567185
transform 1 0 82432 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[264\]
timestamp 1607567185
transform 1 0 120244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1285
timestamp 1607567185
transform 1 0 119324 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1293
timestamp 1607567185
transform 1 0 120060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1298
timestamp 1607567185
transform 1 0 120520 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[272\]
timestamp 1607567185
transform 1 0 117392 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[295\]
timestamp 1607567185
transform 1 0 119048 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607567185
transform 1 0 118956 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1267
timestamp 1607567185
transform 1 0 117668 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1279
timestamp 1607567185
transform 1 0 118772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1252
timestamp 1607567185
transform 1 0 116288 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[71\]
timestamp 1607567185
transform 1 0 114632 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1232
timestamp 1607567185
transform 1 0 114448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[248\]
timestamp 1607567185
transform 1 0 113436 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607567185
transform 1 0 113344 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1208
timestamp 1607567185
transform 1 0 112240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1224
timestamp 1607567185
transform 1 0 113712 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[118\]
timestamp 1607567185
transform 1 0 111412 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1191
timestamp 1607567185
transform 1 0 110676 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[76\]
timestamp 1607567185
transform 1 0 109020 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1171
timestamp 1607567185
transform 1 0 108836 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[246\]
timestamp 1607567185
transform 1 0 107824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607567185
transform 1 0 107732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1163
timestamp 1607567185
transform 1 0 108100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[125\]
timestamp 1607567185
transform 1 0 105800 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1137
timestamp 1607567185
transform 1 0 105708 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1147
timestamp 1607567185
transform 1 0 106628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1129
timestamp 1607567185
transform 1 0 104972 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[281\]
timestamp 1607567185
transform 1 0 102212 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[82\]
timestamp 1607567185
transform 1 0 103316 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607567185
transform 1 0 102120 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1095
timestamp 1607567185
transform 1 0 101844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1102
timestamp 1607567185
transform 1 0 102488 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1110
timestamp 1607567185
transform 1 0 103224 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1083
timestamp 1607567185
transform 1 0 100740 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[4\]
timestamp 1607567185
transform 1 0 99084 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1059
timestamp 1607567185
transform 1 0 98532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[110\]
timestamp 1607567185
transform 1 0 96600 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1047
timestamp 1607567185
transform 1 0 97428 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607567185
transform 1 0 96508 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1026
timestamp 1607567185
transform 1 0 95496 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1034
timestamp 1607567185
transform 1 0 96232 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[91\]
timestamp 1607567185
transform 1 0 94668 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1009
timestamp 1607567185
transform 1 0 93932 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[77\]
timestamp 1607567185
transform 1 0 92276 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_13_989
timestamp 1607567185
transform 1 0 92092 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[279\]
timestamp 1607567185
transform 1 0 91080 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607567185
transform 1 0 90896 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_971
timestamp 1607567185
transform 1 0 90436 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_975
timestamp 1607567185
transform 1 0 90804 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_977
timestamp 1607567185
transform 1 0 90988 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_981
timestamp 1607567185
transform 1 0 91356 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[82\]
timestamp 1607567185
transform 1 0 88504 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_959
timestamp 1607567185
transform 1 0 89332 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[80\]
timestamp 1607567185
transform 1 0 86940 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_925
timestamp 1607567185
transform 1 0 86204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_942
timestamp 1607567185
transform 1 0 87768 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[76\]
timestamp 1607567185
transform 1 0 85376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607567185
transform 1 0 85284 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_911
timestamp 1607567185
transform 1 0 84916 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[251\]
timestamp 1607567185
transform 1 0 83536 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1607567185
transform 1 0 83444 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_899
timestamp 1607567185
transform 1 0 83812 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_883
timestamp 1607567185
transform 1 0 82340 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1296
timestamp 1607567185
transform 1 0 120336 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[258\]
timestamp 1607567185
transform 1 0 117668 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[70\]
timestamp 1607567185
transform 1 0 118680 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1270
timestamp 1607567185
transform 1 0 117944 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[288\]
timestamp 1607567185
transform 1 0 116288 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607567185
transform 1 0 116196 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1249
timestamp 1607567185
transform 1 0 116012 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1255
timestamp 1607567185
transform 1 0 116564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1241
timestamp 1607567185
transform 1 0 115276 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[47\]
timestamp 1607567185
transform 1 0 113620 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1215
timestamp 1607567185
transform 1 0 112884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[85\]
timestamp 1607567185
transform 1 0 111228 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607567185
transform 1 0 110584 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1189
timestamp 1607567185
transform 1 0 110492 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1191
timestamp 1607567185
transform 1 0 110676 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[115\]
timestamp 1607567185
transform 1 0 108928 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1181
timestamp 1607567185
transform 1 0 109756 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[114\]
timestamp 1607567185
transform 1 0 107364 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1151
timestamp 1607567185
transform 1 0 106996 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1164
timestamp 1607567185
transform 1 0 108192 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1139
timestamp 1607567185
transform 1 0 105892 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[123\]
timestamp 1607567185
transform 1 0 105064 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607567185
transform 1 0 104972 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1119
timestamp 1607567185
transform 1 0 104052 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1127
timestamp 1607567185
transform 1 0 104788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[79\]
timestamp 1607567185
transform 1 0 102396 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1095
timestamp 1607567185
transform 1 0 101844 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[421\]
timestamp 1607567185
transform 1 0 100464 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1083
timestamp 1607567185
transform 1 0 100740 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[414\]
timestamp 1607567185
transform 1 0 99452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607567185
transform 1 0 99360 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1060
timestamp 1607567185
transform 1 0 98624 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1072
timestamp 1607567185
transform 1 0 99728 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[73\]
timestamp 1607567185
transform 1 0 96968 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[95\]
timestamp 1607567185
transform 1 0 95404 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1034
timestamp 1607567185
transform 1 0 96232 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[94\]
timestamp 1607567185
transform 1 0 93840 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607567185
transform 1 0 93748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1017
timestamp 1607567185
transform 1 0 94668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[87\]
timestamp 1607567185
transform 1 0 92184 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_982
timestamp 1607567185
transform 1 0 91448 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_999
timestamp 1607567185
transform 1 0 93012 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[96\]
timestamp 1607567185
transform 1 0 90620 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_968
timestamp 1607567185
transform 1 0 90160 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_972
timestamp 1607567185
transform 1 0 90528 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[81\]
timestamp 1607567185
transform 1 0 88228 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607567185
transform 1 0 88136 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_945
timestamp 1607567185
transform 1 0 88044 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_956
timestamp 1607567185
transform 1 0 89056 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[78\]
timestamp 1607567185
transform 1 0 86480 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_937
timestamp 1607567185
transform 1 0 87308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[75\]
timestamp 1607567185
transform 1 0 84916 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_907
timestamp 1607567185
transform 1 0 84548 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_920
timestamp 1607567185
transform 1 0 85744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_895
timestamp 1607567185
transform 1 0 83444 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[74\]
timestamp 1607567185
transform 1 0 82616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607567185
transform 1 0 82524 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_869
timestamp 1607567185
transform 1 0 81052 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_881
timestamp 1607567185
transform 1 0 82156 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[257\]
timestamp 1607567185
transform 1 0 119508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[55\]
timestamp 1607567185
transform 1 0 120612 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1286
timestamp 1607567185
transform 1 0 119416 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1290
timestamp 1607567185
transform 1 0 119784 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1298
timestamp 1607567185
transform 1 0 120520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607567185
transform 1 0 118956 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1273
timestamp 1607567185
transform 1 0 118220 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1282
timestamp 1607567185
transform 1 0 119048 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[88\]
timestamp 1607567185
transform 1 0 116564 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1254
timestamp 1607567185
transform 1 0 116472 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1242
timestamp 1607567185
transform 1 0 115368 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[46\]
timestamp 1607567185
transform 1 0 113712 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607567185
transform 1 0 113344 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1209
timestamp 1607567185
transform 1 0 112332 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1217
timestamp 1607567185
transform 1 0 113068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1221
timestamp 1607567185
transform 1 0 113436 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[249\]
timestamp 1607567185
transform 1 0 112056 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1198
timestamp 1607567185
transform 1 0 111320 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[44\]
timestamp 1607567185
transform 1 0 109664 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1177
timestamp 1607567185
transform 1 0 109388 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[120\]
timestamp 1607567185
transform 1 0 107824 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607567185
transform 1 0 107732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1156
timestamp 1607567185
transform 1 0 107456 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1169
timestamp 1607567185
transform 1 0 108652 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[121\]
timestamp 1607567185
transform 1 0 105892 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1148
timestamp 1607567185
transform 1 0 106720 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[112\]
timestamp 1607567185
transform 1 0 104328 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1114
timestamp 1607567185
transform 1 0 103592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1131
timestamp 1607567185
transform 1 0 105156 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[111\]
timestamp 1607567185
transform 1 0 102764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607567185
transform 1 0 102120 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1096
timestamp 1607567185
transform 1 0 101936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1099
timestamp 1607567185
transform 1 0 102212 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[424\]
timestamp 1607567185
transform 1 0 100924 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1077
timestamp 1607567185
transform 1 0 100188 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1088
timestamp 1607567185
transform 1 0 101200 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[98\]
timestamp 1607567185
transform 1 0 99360 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1060
timestamp 1607567185
transform 1 0 98624 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[66\]
timestamp 1607567185
transform 1 0 96968 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1038
timestamp 1607567185
transform 1 0 96600 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607567185
transform 1 0 96508 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1024
timestamp 1607567185
transform 1 0 95312 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1036
timestamp 1607567185
transform 1 0 96416 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[102\]
timestamp 1607567185
transform 1 0 94484 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1003
timestamp 1607567185
transform 1 0 93380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[93\]
timestamp 1607567185
transform 1 0 92552 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_986
timestamp 1607567185
transform 1 0 91816 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[88\]
timestamp 1607567185
transform 1 0 90988 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607567185
transform 1 0 90896 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_968
timestamp 1607567185
transform 1 0 90160 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[84\]
timestamp 1607567185
transform 1 0 89332 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_954
timestamp 1607567185
transform 1 0 88872 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_958
timestamp 1607567185
transform 1 0 89240 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[77\]
timestamp 1607567185
transform 1 0 86940 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_925
timestamp 1607567185
transform 1 0 86204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_942
timestamp 1607567185
transform 1 0 87768 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[68\]
timestamp 1607567185
transform 1 0 85376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607567185
transform 1 0 85284 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_909
timestamp 1607567185
transform 1 0 84732 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[69\]
timestamp 1607567185
transform 1 0 82800 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_897
timestamp 1607567185
transform 1 0 83628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[54\]
timestamp 1607567185
transform 1 0 81236 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_870
timestamp 1607567185
transform 1 0 81144 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_880
timestamp 1607567185
transform 1 0 82064 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1300
timestamp 1607567185
transform 1 0 120704 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1296
timestamp 1607567185
transform 1 0 120336 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[250\]
timestamp 1607567185
transform 1 0 117760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[48\]
timestamp 1607567185
transform 1 0 118680 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[56\]
timestamp 1607567185
transform 1 0 119048 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607567185
transform 1 0 118956 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1266
timestamp 1607567185
transform 1 0 117576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1271
timestamp 1607567185
transform 1 0 118036 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1279
timestamp 1607567185
transform 1 0 118772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1270
timestamp 1607567185
transform 1 0 117944 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[86\]
timestamp 1607567185
transform 1 0 116288 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607567185
transform 1 0 116196 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1254
timestamp 1607567185
transform 1 0 116472 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1248
timestamp 1607567185
transform 1 0 115920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[36\]
timestamp 1607567185
transform 1 0 114816 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1228
timestamp 1607567185
transform 1 0 114080 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1240
timestamp 1607567185
transform 1 0 115184 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[40\]
timestamp 1607567185
transform 1 0 113528 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1221
timestamp 1607567185
transform 1 0 113436 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1221
timestamp 1607567185
transform 1 0 113436 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1219
timestamp 1607567185
transform 1 0 113252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607567185
transform 1 0 113344 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[238\]
timestamp 1607567185
transform 1 0 113804 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1213
timestamp 1607567185
transform 1 0 112700 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1208
timestamp 1607567185
transform 1 0 112240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1215
timestamp 1607567185
transform 1 0 112884 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[242\]
timestamp 1607567185
transform 1 0 112424 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[119\]
timestamp 1607567185
transform 1 0 110676 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[126\]
timestamp 1607567185
transform 1 0 110952 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607567185
transform 1 0 110584 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1203
timestamp 1607567185
transform 1 0 111780 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1200
timestamp 1607567185
transform 1 0 111504 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[117\]
timestamp 1607567185
transform 1 0 109388 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1186
timestamp 1607567185
transform 1 0 110216 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1176
timestamp 1607567185
transform 1 0 109296 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1188
timestamp 1607567185
transform 1 0 110400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[109\]
timestamp 1607567185
transform 1 0 107824 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[41\]
timestamp 1607567185
transform 1 0 107640 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607567185
transform 1 0 107732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1158
timestamp 1607567185
transform 1 0 107640 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1169
timestamp 1607567185
transform 1 0 108652 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[243\]
timestamp 1607567185
transform 1 0 106260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[28\]
timestamp 1607567185
transform 1 0 105248 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1135
timestamp 1607567185
transform 1 0 105524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1146
timestamp 1607567185
transform 1 0 106536 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1150
timestamp 1607567185
transform 1 0 106904 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[17\]
timestamp 1607567185
transform 1 0 103868 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607567185
transform 1 0 104972 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1116
timestamp 1607567185
transform 1 0 103776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1119
timestamp 1607567185
transform 1 0 104052 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1127
timestamp 1607567185
transform 1 0 104788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1130
timestamp 1607567185
transform 1 0 105064 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[108\]
timestamp 1607567185
transform 1 0 102212 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[42\]
timestamp 1607567185
transform 1 0 102396 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607567185
transform 1 0 102120 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1097
timestamp 1607567185
transform 1 0 102028 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1108
timestamp 1607567185
transform 1 0 103040 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1098
timestamp 1607567185
transform 1 0 102120 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[244\]
timestamp 1607567185
transform 1 0 100740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[422\]
timestamp 1607567185
transform 1 0 101016 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1078
timestamp 1607567185
transform 1 0 100280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1089
timestamp 1607567185
transform 1 0 101292 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1080
timestamp 1607567185
transform 1 0 100464 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1086
timestamp 1607567185
transform 1 0 101016 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[418\]
timestamp 1607567185
transform 1 0 99452 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[419\]
timestamp 1607567185
transform 1 0 100004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[104\]
timestamp 1607567185
transform 1 0 98440 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607567185
transform 1 0 99360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1067
timestamp 1607567185
transform 1 0 99268 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1059
timestamp 1607567185
transform 1 0 98532 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1067
timestamp 1607567185
transform 1 0 99268 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1072
timestamp 1607567185
transform 1 0 99728 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[101\]
timestamp 1607567185
transform 1 0 96876 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[105\]
timestamp 1607567185
transform 1 0 97704 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1038
timestamp 1607567185
transform 1 0 96600 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1050
timestamp 1607567185
transform 1 0 97704 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1042
timestamp 1607567185
transform 1 0 96968 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[103\]
timestamp 1607567185
transform 1 0 96140 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607567185
transform 1 0 96508 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1027
timestamp 1607567185
transform 1 0 95588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1035
timestamp 1607567185
transform 1 0 96324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1024
timestamp 1607567185
transform 1 0 95312 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1032
timestamp 1607567185
transform 1 0 96048 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[100\]
timestamp 1607567185
transform 1 0 94484 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[90\]
timestamp 1607567185
transform 1 0 94760 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607567185
transform 1 0 93748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1007
timestamp 1607567185
transform 1 0 93748 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1015
timestamp 1607567185
transform 1 0 94484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1005
timestamp 1607567185
transform 1 0 93564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1008
timestamp 1607567185
transform 1 0 93840 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1014
timestamp 1607567185
transform 1 0 94392 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[83\]
timestamp 1607567185
transform 1 0 92920 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[89\]
timestamp 1607567185
transform 1 0 91632 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_987
timestamp 1607567185
transform 1 0 91908 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_995
timestamp 1607567185
transform 1 0 92644 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_993
timestamp 1607567185
transform 1 0 92460 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[79\]
timestamp 1607567185
transform 1 0 90068 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[92\]
timestamp 1607567185
transform 1 0 91080 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607567185
transform 1 0 90896 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_973
timestamp 1607567185
transform 1 0 90620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_977
timestamp 1607567185
transform 1 0 90988 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_966
timestamp 1607567185
transform 1 0 89976 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_976
timestamp 1607567185
transform 1 0 90896 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[393\]
timestamp 1607567185
transform 1 0 88228 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[72\]
timestamp 1607567185
transform 1 0 88688 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607567185
transform 1 0 88136 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_944
timestamp 1607567185
transform 1 0 87952 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_961
timestamp 1607567185
transform 1 0 89516 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_945
timestamp 1607567185
transform 1 0 88044 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_950
timestamp 1607567185
transform 1 0 88504 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_962
timestamp 1607567185
transform 1 0 89608 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[391\]
timestamp 1607567185
transform 1 0 86664 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[70\]
timestamp 1607567185
transform 1 0 87124 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_925
timestamp 1607567185
transform 1 0 86204 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_933
timestamp 1607567185
transform 1 0 86940 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_933
timestamp 1607567185
transform 1 0 86940 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[63\]
timestamp 1607567185
transform 1 0 85100 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[67\]
timestamp 1607567185
transform 1 0 85376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607567185
transform 1 0 85284 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_910
timestamp 1607567185
transform 1 0 84824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_914
timestamp 1607567185
transform 1 0 85192 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_907
timestamp 1607567185
transform 1 0 84548 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_922
timestamp 1607567185
transform 1 0 85928 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[53\]
timestamp 1607567185
transform 1 0 82892 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_898
timestamp 1607567185
transform 1 0 83720 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_895
timestamp 1607567185
transform 1 0 83444 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[50\]
timestamp 1607567185
transform 1 0 81328 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[59\]
timestamp 1607567185
transform 1 0 82616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607567185
transform 1 0 82524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_881
timestamp 1607567185
transform 1 0 82156 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_876
timestamp 1607567185
transform 1 0 81696 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_884
timestamp 1607567185
transform 1 0 82432 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[254\]
timestamp 1607567185
transform 1 0 120796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1292
timestamp 1607567185
transform 1 0 119968 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1300
timestamp 1607567185
transform 1 0 120704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[53\]
timestamp 1607567185
transform 1 0 118312 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1266
timestamp 1607567185
transform 1 0 117576 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[240\]
timestamp 1607567185
transform 1 0 116288 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[255\]
timestamp 1607567185
transform 1 0 117300 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607567185
transform 1 0 116196 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1247
timestamp 1607567185
transform 1 0 115828 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1255
timestamp 1607567185
transform 1 0 116564 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1235
timestamp 1607567185
transform 1 0 114724 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[24\]
timestamp 1607567185
transform 1 0 113068 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1209
timestamp 1607567185
transform 1 0 112332 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[34\]
timestamp 1607567185
transform 1 0 110676 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607567185
transform 1 0 110584 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1189
timestamp 1607567185
transform 1 0 110492 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1177
timestamp 1607567185
transform 1 0 109388 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[124\]
timestamp 1607567185
transform 1 0 108560 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1160
timestamp 1607567185
transform 1 0 107824 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[20\]
timestamp 1607567185
transform 1 0 106168 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1133
timestamp 1607567185
transform 1 0 105340 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1141
timestamp 1607567185
transform 1 0 106076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[230\]
timestamp 1607567185
transform 1 0 105064 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607567185
transform 1 0 104972 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1121
timestamp 1607567185
transform 1 0 104236 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[219\]
timestamp 1607567185
transform 1 0 101844 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[106\]
timestamp 1607567185
transform 1 0 103408 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1098
timestamp 1607567185
transform 1 0 102120 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1110
timestamp 1607567185
transform 1 0 103224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[423\]
timestamp 1607567185
transform 1 0 100464 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1083
timestamp 1607567185
transform 1 0 100740 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[218\]
timestamp 1607567185
transform 1 0 99452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607567185
transform 1 0 99360 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1059
timestamp 1607567185
transform 1 0 98532 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1067
timestamp 1607567185
transform 1 0 99268 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1072
timestamp 1607567185
transform 1 0 99728 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[2\]
timestamp 1607567185
transform 1 0 96876 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1038
timestamp 1607567185
transform 1 0 96600 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1030
timestamp 1607567185
transform 1 0 95864 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[18\]
timestamp 1607567185
transform 1 0 94208 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607567185
transform 1 0 93748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1001
timestamp 1607567185
transform 1 0 93196 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1008
timestamp 1607567185
transform 1 0 93840 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_989
timestamp 1607567185
transform 1 0 92092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[85\]
timestamp 1607567185
transform 1 0 91264 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_965
timestamp 1607567185
transform 1 0 89884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_977
timestamp 1607567185
transform 1 0 90988 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[11\]
timestamp 1607567185
transform 1 0 88228 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607567185
transform 1 0 88136 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[213\]
timestamp 1607567185
transform 1 0 86756 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_929
timestamp 1607567185
transform 1 0 86572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_934
timestamp 1607567185
transform 1 0 87032 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[397\]
timestamp 1607567185
transform 1 0 85192 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_906
timestamp 1607567185
transform 1 0 84456 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_917
timestamp 1607567185
transform 1 0 85468 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[387\]
timestamp 1607567185
transform 1 0 84180 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_895
timestamp 1607567185
transform 1 0 83444 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[57\]
timestamp 1607567185
transform 1 0 82616 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607567185
transform 1 0 82524 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_875
timestamp 1607567185
transform 1 0 81604 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_883
timestamp 1607567185
transform 1 0 82340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1607567185
transform 1 0 80960 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[247\]
timestamp 1607567185
transform 1 0 79672 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_853
timestamp 1607567185
transform 1 0 79580 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_857
timestamp 1607567185
transform 1 0 79948 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_865
timestamp 1607567185
transform 1 0 80684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[382\]
timestamp 1607567185
transform 1 0 78200 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1607567185
transform 1 0 78108 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_833
timestamp 1607567185
transform 1 0 77740 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_841
timestamp 1607567185
transform 1 0 78476 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[374\]
timestamp 1607567185
transform 1 0 76360 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_821
timestamp 1607567185
transform 1 0 76636 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[362\]
timestamp 1607567185
transform 1 0 74152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[369\]
timestamp 1607567185
transform 1 0 75348 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1607567185
transform 1 0 75256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_793
timestamp 1607567185
transform 1 0 74060 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_797
timestamp 1607567185
transform 1 0 74428 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_805
timestamp 1607567185
transform 1 0 75164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_810
timestamp 1607567185
transform 1 0 75624 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[270\]
timestamp 1607567185
transform 1 0 73048 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1607567185
transform 1 0 72404 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_774
timestamp 1607567185
transform 1 0 72312 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_776
timestamp 1607567185
transform 1 0 72496 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_785
timestamp 1607567185
transform 1 0 73324 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[355\]
timestamp 1607567185
transform 1 0 70932 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_758
timestamp 1607567185
transform 1 0 70840 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_762
timestamp 1607567185
transform 1 0 71208 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[365\]
timestamp 1607567185
transform 1 0 69828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1607567185
transform 1 0 69552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_736
timestamp 1607567185
transform 1 0 68816 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_745
timestamp 1607567185
transform 1 0 69644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_750
timestamp 1607567185
transform 1 0 70104 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[370\]
timestamp 1607567185
transform 1 0 68540 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[371\]
timestamp 1607567185
transform 1 0 67528 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_725
timestamp 1607567185
transform 1 0 67804 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[375\]
timestamp 1607567185
transform 1 0 65688 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1607567185
transform 1 0 66700 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_705
timestamp 1607567185
transform 1 0 65964 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_714
timestamp 1607567185
transform 1 0 66792 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[390\]
timestamp 1607567185
transform 1 0 64676 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1607567185
transform 1 0 63848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_680
timestamp 1607567185
transform 1 0 63664 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_683
timestamp 1607567185
transform 1 0 63940 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_694
timestamp 1607567185
transform 1 0 64952 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[341\]
timestamp 1607567185
transform 1 0 62652 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_661
timestamp 1607567185
transform 1 0 61916 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_672
timestamp 1607567185
transform 1 0 62928 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[9\]
timestamp 1607567185
transform 1 0 61088 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1607567185
transform 1 0 60996 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_649
timestamp 1607567185
transform 1 0 60812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[336\]
timestamp 1607567185
transform 1 0 59800 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_633
timestamp 1607567185
transform 1 0 59340 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_637
timestamp 1607567185
transform 1 0 59708 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_641
timestamp 1607567185
transform 1 0 60076 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1607567185
transform 1 0 58144 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_614
timestamp 1607567185
transform 1 0 57592 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_621
timestamp 1607567185
transform 1 0 58236 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1607567185
transform 1 0 55292 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_590
timestamp 1607567185
transform 1 0 55384 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_602
timestamp 1607567185
transform 1 0 56488 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_571
timestamp 1607567185
transform 1 0 53636 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_583
timestamp 1607567185
transform 1 0 54740 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1607567185
transform 1 0 52440 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_552
timestamp 1607567185
transform 1 0 51888 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_559
timestamp 1607567185
transform 1 0 52532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_540
timestamp 1607567185
transform 1 0 50784 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1607567185
transform 1 0 49588 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_511
timestamp 1607567185
transform 1 0 48116 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_523
timestamp 1607567185
transform 1 0 49220 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_528
timestamp 1607567185
transform 1 0 49680 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[164\]
timestamp 1607567185
transform 1 0 46828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[171\]
timestamp 1607567185
transform 1 0 47840 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1607567185
transform 1 0 46736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_500
timestamp 1607567185
transform 1 0 47104 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_484
timestamp 1607567185
transform 1 0 45632 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[96\]
timestamp 1607567185
transform 1 0 43976 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1607567185
transform 1 0 43884 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_455
timestamp 1607567185
transform 1 0 42964 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_463
timestamp 1607567185
transform 1 0 43700 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[168\]
timestamp 1607567185
transform 1 0 42688 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_435
timestamp 1607567185
transform 1 0 41124 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_447
timestamp 1607567185
transform 1 0 42228 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_451
timestamp 1607567185
transform 1 0 42596 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[71\]
timestamp 1607567185
transform 1 0 79488 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_861
timestamp 1607567185
transform 1 0 80316 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_834
timestamp 1607567185
transform 1 0 77832 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_846
timestamp 1607567185
transform 1 0 78936 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[65\]
timestamp 1607567185
transform 1 0 77004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607567185
transform 1 0 76912 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_819
timestamp 1607567185
transform 1 0 76452 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_823
timestamp 1607567185
transform 1 0 76820 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_807
timestamp 1607567185
transform 1 0 75348 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[68\]
timestamp 1607567185
transform 1 0 73692 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_14_785
timestamp 1607567185
transform 1 0 73324 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[45\]
timestamp 1607567185
transform 1 0 71392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607567185
transform 1 0 71300 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_755
timestamp 1607567185
transform 1 0 70564 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_773
timestamp 1607567185
transform 1 0 72220 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[358\]
timestamp 1607567185
transform 1 0 70288 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[360\]
timestamp 1607567185
transform 1 0 69276 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_738
timestamp 1607567185
transform 1 0 69000 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_744
timestamp 1607567185
transform 1 0 69552 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[352\]
timestamp 1607567185
transform 1 0 67988 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_719
timestamp 1607567185
transform 1 0 67252 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_730
timestamp 1607567185
transform 1 0 68264 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[193\]
timestamp 1607567185
transform 1 0 66976 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[372\]
timestamp 1607567185
transform 1 0 65964 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607567185
transform 1 0 65688 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_703
timestamp 1607567185
transform 1 0 65780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_708
timestamp 1607567185
transform 1 0 66240 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[344\]
timestamp 1607567185
transform 1 0 63756 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_684
timestamp 1607567185
transform 1 0 64032 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_696
timestamp 1607567185
transform 1 0 65136 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[339\]
timestamp 1607567185
transform 1 0 62744 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_662
timestamp 1607567185
transform 1 0 62008 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_673
timestamp 1607567185
transform 1 0 63020 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[187\]
timestamp 1607567185
transform 1 0 61732 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[8\]
timestamp 1607567185
transform 1 0 60168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_651
timestamp 1607567185
transform 1 0 60996 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[186\]
timestamp 1607567185
transform 1 0 59064 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607567185
transform 1 0 60076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_629
timestamp 1607567185
transform 1 0 58972 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_633
timestamp 1607567185
transform 1 0 59340 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_605
timestamp 1607567185
transform 1 0 56764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_617
timestamp 1607567185
transform 1 0 57868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[108\]
timestamp 1607567185
transform 1 0 55108 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607567185
transform 1 0 54464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_571
timestamp 1607567185
transform 1 0 53636 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_579
timestamp 1607567185
transform 1 0 54372 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1607567185
transform 1 0 54556 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_559
timestamp 1607567185
transform 1 0 52532 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_535
timestamp 1607567185
transform 1 0 50324 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_547
timestamp 1607567185
transform 1 0 51428 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[176\]
timestamp 1607567185
transform 1 0 48944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607567185
transform 1 0 48852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_523
timestamp 1607567185
transform 1 0 49220 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_507
timestamp 1607567185
transform 1 0 47748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[97\]
timestamp 1607567185
transform 1 0 46092 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_481
timestamp 1607567185
transform 1 0 45356 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[88\]
timestamp 1607567185
transform 1 0 43700 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607567185
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_459
timestamp 1607567185
transform 1 0 43332 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_450
timestamp 1607567185
transform 1 0 42504 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[45\]
timestamp 1607567185
transform 1 0 80684 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607567185
transform 1 0 79672 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_853
timestamp 1607567185
transform 1 0 79580 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_855
timestamp 1607567185
transform 1 0 79764 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_863
timestamp 1607567185
transform 1 0 80500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[381\]
timestamp 1607567185
transform 1 0 78568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_841
timestamp 1607567185
transform 1 0 78476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_845
timestamp 1607567185
transform 1 0 78844 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[58\]
timestamp 1607567185
transform 1 0 76544 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_818
timestamp 1607567185
transform 1 0 76360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_829
timestamp 1607567185
transform 1 0 77372 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[60\]
timestamp 1607567185
transform 1 0 74428 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607567185
transform 1 0 74060 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_794
timestamp 1607567185
transform 1 0 74152 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_806
timestamp 1607567185
transform 1 0 75256 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[40\]
timestamp 1607567185
transform 1 0 72496 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_785
timestamp 1607567185
transform 1 0 73324 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[42\]
timestamp 1607567185
transform 1 0 70932 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_768
timestamp 1607567185
transform 1 0 71760 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[351\]
timestamp 1607567185
transform 1 0 69000 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_737
timestamp 1607567185
transform 1 0 68908 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_741
timestamp 1607567185
transform 1 0 69276 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_753
timestamp 1607567185
transform 1 0 70380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607567185
transform 1 0 68448 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_724
timestamp 1607567185
transform 1 0 67712 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_733
timestamp 1607567185
transform 1 0 68540 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[119\]
timestamp 1607567185
transform 1 0 66056 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_13_705
timestamp 1607567185
transform 1 0 65964 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[340\]
timestamp 1607567185
transform 1 0 63940 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[343\]
timestamp 1607567185
transform 1 0 64952 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_686
timestamp 1607567185
transform 1 0 64216 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_697
timestamp 1607567185
transform 1 0 65228 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[338\]
timestamp 1607567185
transform 1 0 62928 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607567185
transform 1 0 62836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1607567185
transform 1 0 62284 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_675
timestamp 1607567185
transform 1 0 63204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_653
timestamp 1607567185
transform 1 0 61180 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[112\]
timestamp 1607567185
transform 1 0 59524 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[337\]
timestamp 1607567185
transform 1 0 58512 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_623
timestamp 1607567185
transform 1 0 58420 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_627
timestamp 1607567185
transform 1 0 58788 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607567185
transform 1 0 57224 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_608
timestamp 1607567185
transform 1 0 57040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_611
timestamp 1607567185
transform 1 0 57316 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_600
timestamp 1607567185
transform 1 0 56304 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[107\]
timestamp 1607567185
transform 1 0 54648 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[196\]
timestamp 1607567185
transform 1 0 53636 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_570
timestamp 1607567185
transform 1 0 53544 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_574
timestamp 1607567185
transform 1 0 53912 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607567185
transform 1 0 51612 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_550
timestamp 1607567185
transform 1 0 51704 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_562
timestamp 1607567185
transform 1 0 52808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[179\]
timestamp 1607567185
transform 1 0 49956 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_534
timestamp 1607567185
transform 1 0 50232 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_546
timestamp 1607567185
transform 1 0 51336 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_523
timestamp 1607567185
transform 1 0 49220 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[102\]
timestamp 1607567185
transform 1 0 47564 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_13_492
timestamp 1607567185
transform 1 0 46368 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_504
timestamp 1607567185
transform 1 0 47472 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[162\]
timestamp 1607567185
transform 1 0 46092 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607567185
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1607567185
transform 1 0 44620 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_485
timestamp 1607567185
transform 1 0 45724 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[159\]
timestamp 1607567185
transform 1 0 44344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_462
timestamp 1607567185
transform 1 0 43608 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[81\]
timestamp 1607567185
transform 1 0 41952 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_13_436
timestamp 1607567185
transform 1 0 41216 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[62\]
timestamp 1607567185
transform 1 0 80224 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_857
timestamp 1607567185
transform 1 0 79948 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[52\]
timestamp 1607567185
transform 1 0 78016 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_845
timestamp 1607567185
transform 1 0 78844 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[366\]
timestamp 1607567185
transform 1 0 77004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607567185
transform 1 0 76912 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_812
timestamp 1607567185
transform 1 0 75808 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_828
timestamp 1607567185
transform 1 0 77280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[64\]
timestamp 1607567185
transform 1 0 74980 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_792
timestamp 1607567185
transform 1 0 73968 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_800
timestamp 1607567185
transform 1 0 74704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[32\]
timestamp 1607567185
transform 1 0 73140 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_781
timestamp 1607567185
transform 1 0 72956 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[41\]
timestamp 1607567185
transform 1 0 71392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607567185
transform 1 0 71300 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_761
timestamp 1607567185
transform 1 0 71116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_773
timestamp 1607567185
transform 1 0 72220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[349\]
timestamp 1607567185
transform 1 0 69092 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[353\]
timestamp 1607567185
transform 1 0 70104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_742
timestamp 1607567185
transform 1 0 69368 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_753
timestamp 1607567185
transform 1 0 70380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[22\]
timestamp 1607567185
transform 1 0 67528 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_718
timestamp 1607567185
transform 1 0 67160 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_731
timestamp 1607567185
transform 1 0 68356 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[347\]
timestamp 1607567185
transform 1 0 65780 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607567185
transform 1 0 65688 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_706
timestamp 1607567185
transform 1 0 66056 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[13\]
timestamp 1607567185
transform 1 0 64124 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_694
timestamp 1607567185
transform 1 0 64952 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[10\]
timestamp 1607567185
transform 1 0 62560 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_677
timestamp 1607567185
transform 1 0 63388 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[113\]
timestamp 1607567185
transform 1 0 60168 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_660
timestamp 1607567185
transform 1 0 61824 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[7\]
timestamp 1607567185
transform 1 0 58512 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607567185
transform 1 0 60076 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_633
timestamp 1607567185
transform 1 0 59340 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_610
timestamp 1607567185
transform 1 0 57224 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_622
timestamp 1607567185
transform 1 0 58328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[182\]
timestamp 1607567185
transform 1 0 55844 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_587
timestamp 1607567185
transform 1 0 55108 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_598
timestamp 1607567185
transform 1 0 56120 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[181\]
timestamp 1607567185
transform 1 0 54832 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607567185
transform 1 0 54464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_576
timestamp 1607567185
transform 1 0 54096 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_581
timestamp 1607567185
transform 1 0 54556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[174\]
timestamp 1607567185
transform 1 0 52716 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[188\]
timestamp 1607567185
transform 1 0 51704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_553
timestamp 1607567185
transform 1 0 51980 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_564
timestamp 1607567185
transform 1 0 52992 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[167\]
timestamp 1607567185
transform 1 0 49956 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_534
timestamp 1607567185
transform 1 0 50232 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_546
timestamp 1607567185
transform 1 0 51336 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[163\]
timestamp 1607567185
transform 1 0 48944 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607567185
transform 1 0 48852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_517
timestamp 1607567185
transform 1 0 48668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_523
timestamp 1607567185
transform 1 0 49220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[91\]
timestamp 1607567185
transform 1 0 46276 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_509
timestamp 1607567185
transform 1 0 47932 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_483
timestamp 1607567185
transform 1 0 45540 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[85\]
timestamp 1607567185
transform 1 0 43884 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607567185
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_459
timestamp 1607567185
transform 1 0 43332 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[155\]
timestamp 1607567185
transform 1 0 42228 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_437
timestamp 1607567185
transform 1 0 41308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_445
timestamp 1607567185
transform 1 0 42044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_450
timestamp 1607567185
transform 1 0 42504 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[378\]
timestamp 1607567185
transform 1 0 79764 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607567185
transform 1 0 79672 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_852
timestamp 1607567185
transform 1 0 79488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_858
timestamp 1607567185
transform 1 0 80040 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[48\]
timestamp 1607567185
transform 1 0 77556 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_830
timestamp 1607567185
transform 1 0 77464 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_840
timestamp 1607567185
transform 1 0 78384 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[359\]
timestamp 1607567185
transform 1 0 76084 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_818
timestamp 1607567185
transform 1 0 76360 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[44\]
timestamp 1607567185
transform 1 0 74520 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607567185
transform 1 0 74060 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_794
timestamp 1607567185
transform 1 0 74152 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_807
timestamp 1607567185
transform 1 0 75348 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[39\]
timestamp 1607567185
transform 1 0 72496 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_775
timestamp 1607567185
transform 1 0 72404 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_785
timestamp 1607567185
transform 1 0 73324 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_759
timestamp 1607567185
transform 1 0 70932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_771
timestamp 1607567185
transform 1 0 72036 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[25\]
timestamp 1607567185
transform 1 0 70104 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_742
timestamp 1607567185
transform 1 0 69368 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[348\]
timestamp 1607567185
transform 1 0 67068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[19\]
timestamp 1607567185
transform 1 0 68540 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607567185
transform 1 0 68448 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_720
timestamp 1607567185
transform 1 0 67344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[342\]
timestamp 1607567185
transform 1 0 66056 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_698
timestamp 1607567185
transform 1 0 65320 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_709
timestamp 1607567185
transform 1 0 66332 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[17\]
timestamp 1607567185
transform 1 0 64492 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_681
timestamp 1607567185
transform 1 0 63756 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[12\]
timestamp 1607567185
transform 1 0 62928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607567185
transform 1 0 62836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_662
timestamp 1607567185
transform 1 0 62008 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_670
timestamp 1607567185
transform 1 0 62744 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[11\]
timestamp 1607567185
transform 1 0 61180 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_645
timestamp 1607567185
transform 1 0 60444 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[4\]
timestamp 1607567185
transform 1 0 59616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_628
timestamp 1607567185
transform 1 0 58880 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[6\]
timestamp 1607567185
transform 1 0 58052 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607567185
transform 1 0 57224 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_606
timestamp 1607567185
transform 1 0 56856 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_611
timestamp 1607567185
transform 1 0 57316 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_594
timestamp 1607567185
transform 1 0 55752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[122\]
timestamp 1607567185
transform 1 0 54096 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_11_568
timestamp 1607567185
transform 1 0 53360 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[114\]
timestamp 1607567185
transform 1 0 51704 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607567185
transform 1 0 51612 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_541
timestamp 1607567185
transform 1 0 50876 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[93\]
timestamp 1607567185
transform 1 0 49220 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_11_519
timestamp 1607567185
transform 1 0 48852 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_507
timestamp 1607567185
transform 1 0 47748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[90\]
timestamp 1607567185
transform 1 0 46092 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607567185
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_472
timestamp 1607567185
transform 1 0 44528 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_484
timestamp 1607567185
transform 1 0 45632 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[83\]
timestamp 1607567185
transform 1 0 42872 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[165\]
timestamp 1607567185
transform 1 0 41860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_440
timestamp 1607567185
transform 1 0 41584 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_446
timestamp 1607567185
transform 1 0 42136 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[373\]
timestamp 1607567185
transform 1 0 79856 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[49\]
timestamp 1607567185
transform 1 0 79764 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[61\]
timestamp 1607567185
transform 1 0 80868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607567185
transform 1 0 79672 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_864
timestamp 1607567185
transform 1 0 80592 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_859
timestamp 1607567185
transform 1 0 80132 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[368\]
timestamp 1607567185
transform 1 0 78844 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[51\]
timestamp 1607567185
transform 1 0 78108 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_835
timestamp 1607567185
transform 1 0 77924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_846
timestamp 1607567185
transform 1 0 78936 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_837
timestamp 1607567185
transform 1 0 78108 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_848
timestamp 1607567185
transform 1 0 79120 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[43\]
timestamp 1607567185
transform 1 0 77280 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[46\]
timestamp 1607567185
transform 1 0 76360 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607567185
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_827
timestamp 1607567185
transform 1 0 77188 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_815
timestamp 1607567185
transform 1 0 76084 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_823
timestamp 1607567185
transform 1 0 76820 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_825
timestamp 1607567185
transform 1 0 77004 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[36\]
timestamp 1607567185
transform 1 0 74796 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[38\]
timestamp 1607567185
transform 1 0 75256 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607567185
transform 1 0 74060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_792
timestamp 1607567185
transform 1 0 73968 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_794
timestamp 1607567185
transform 1 0 74152 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_800
timestamp 1607567185
transform 1 0 74704 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_810
timestamp 1607567185
transform 1 0 75624 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_802
timestamp 1607567185
transform 1 0 74888 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[29\]
timestamp 1607567185
transform 1 0 72956 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_776
timestamp 1607567185
transform 1 0 72496 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_788
timestamp 1607567185
transform 1 0 73600 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_790
timestamp 1607567185
transform 1 0 73784 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[27\]
timestamp 1607567185
transform 1 0 71668 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[28\]
timestamp 1607567185
transform 1 0 71392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607567185
transform 1 0 71300 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_759
timestamp 1607567185
transform 1 0 70932 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_760
timestamp 1607567185
transform 1 0 71024 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_773
timestamp 1607567185
transform 1 0 72220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[21\]
timestamp 1607567185
transform 1 0 69092 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[24\]
timestamp 1607567185
transform 1 0 70104 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_742
timestamp 1607567185
transform 1 0 69368 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_748
timestamp 1607567185
transform 1 0 69920 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[350\]
timestamp 1607567185
transform 1 0 67160 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[20\]
timestamp 1607567185
transform 1 0 67528 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[23\]
timestamp 1607567185
transform 1 0 68540 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607567185
transform 1 0 68448 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_721
timestamp 1607567185
transform 1 0 67436 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_729
timestamp 1607567185
transform 1 0 68172 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_731
timestamp 1607567185
transform 1 0 68356 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[345\]
timestamp 1607567185
transform 1 0 66148 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[18\]
timestamp 1607567185
transform 1 0 65964 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607567185
transform 1 0 65688 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_699
timestamp 1607567185
transform 1 0 65412 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_710
timestamp 1607567185
transform 1 0 66424 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_703
timestamp 1607567185
transform 1 0 65780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_714
timestamp 1607567185
transform 1 0 66792 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[334\]
timestamp 1607567185
transform 1 0 65136 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[15\]
timestamp 1607567185
transform 1 0 63756 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[16\]
timestamp 1607567185
transform 1 0 63572 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_688
timestamp 1607567185
transform 1 0 64400 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_690
timestamp 1607567185
transform 1 0 64584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[14\]
timestamp 1607567185
transform 1 0 62192 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607567185
transform 1 0 62836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_668
timestamp 1607567185
transform 1 0 62560 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_672
timestamp 1607567185
transform 1 0 62928 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_678
timestamp 1607567185
transform 1 0 63480 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_663
timestamp 1607567185
transform 1 0 62100 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_673
timestamp 1607567185
transform 1 0 63020 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[201\]
timestamp 1607567185
transform 1 0 61548 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[2\]
timestamp 1607567185
transform 1 0 60168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_649
timestamp 1607567185
transform 1 0 60812 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_660
timestamp 1607567185
transform 1 0 61824 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_651
timestamp 1607567185
transform 1 0 60996 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[127\]
timestamp 1607567185
transform 1 0 59156 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[0\]
timestamp 1607567185
transform 1 0 58512 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607567185
transform 1 0 60076 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_626
timestamp 1607567185
transform 1 0 58696 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_630
timestamp 1607567185
transform 1 0 59064 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_633
timestamp 1607567185
transform 1 0 59340 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[190\]
timestamp 1607567185
transform 1 0 57316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607567185
transform 1 0 57224 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_605
timestamp 1607567185
transform 1 0 56764 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_609
timestamp 1607567185
transform 1 0 57132 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_614
timestamp 1607567185
transform 1 0 57592 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_616
timestamp 1607567185
transform 1 0 57776 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[116\]
timestamp 1607567185
transform 1 0 56120 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[195\]
timestamp 1607567185
transform 1 0 55384 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_593
timestamp 1607567185
transform 1 0 55660 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_596
timestamp 1607567185
transform 1 0 55936 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[191\]
timestamp 1607567185
transform 1 0 54556 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607567185
transform 1 0 54464 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_582
timestamp 1607567185
transform 1 0 54648 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_569
timestamp 1607567185
transform 1 0 53452 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_577
timestamp 1607567185
transform 1 0 54188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_584
timestamp 1607567185
transform 1 0 54832 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[100\]
timestamp 1607567185
transform 1 0 51796 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[117\]
timestamp 1607567185
transform 1 0 52992 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[185\]
timestamp 1607567185
transform 1 0 51704 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607567185
transform 1 0 51612 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_553
timestamp 1607567185
transform 1 0 51980 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_561
timestamp 1607567185
transform 1 0 52716 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_550
timestamp 1607567185
transform 1 0 51704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_533
timestamp 1607567185
transform 1 0 50140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_545
timestamp 1607567185
transform 1 0 51244 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_538
timestamp 1607567185
transform 1 0 50600 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[105\]
timestamp 1607567185
transform 1 0 48944 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[109\]
timestamp 1607567185
transform 1 0 48484 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607567185
transform 1 0 48852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_510
timestamp 1607567185
transform 1 0 48024 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_518
timestamp 1607567185
transform 1 0 48760 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  la_buf\[89\]
timestamp 1607567185
transform 1 0 46368 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_9_507
timestamp 1607567185
transform 1 0 47748 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[87\]
timestamp 1607567185
transform 1 0 46092 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607567185
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_480
timestamp 1607567185
transform 1 0 45264 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_484
timestamp 1607567185
transform 1 0 45632 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[101\]
timestamp 1607567185
transform 1 0 43976 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[79\]
timestamp 1607567185
transform 1 0 43608 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607567185
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_454
timestamp 1607567185
transform 1 0 42872 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_459
timestamp 1607567185
transform 1 0 43332 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_465
timestamp 1607567185
transform 1 0 43884 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[157\]
timestamp 1607567185
transform 1 0 42228 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[175\]
timestamp 1607567185
transform 1 0 42596 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_440
timestamp 1607567185
transform 1 0 41584 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_448
timestamp 1607567185
transform 1 0 42320 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_441
timestamp 1607567185
transform 1 0 41676 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_450
timestamp 1607567185
transform 1 0 42504 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[6\]
timestamp 1607567185
transform 1 0 79948 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_849
timestamp 1607567185
transform 1 0 79212 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[13\]
timestamp 1607567185
transform 1 0 77556 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607567185
transform 1 0 76912 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_816
timestamp 1607567185
transform 1 0 76176 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_825
timestamp 1607567185
transform 1 0 77004 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[47\]
timestamp 1607567185
transform 1 0 75348 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_799
timestamp 1607567185
transform 1 0 74612 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[35\]
timestamp 1607567185
transform 1 0 73784 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_782
timestamp 1607567185
transform 1 0 73048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[5\]
timestamp 1607567185
transform 1 0 71392 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607567185
transform 1 0 71300 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_762
timestamp 1607567185
transform 1 0 71208 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[207\]
timestamp 1607567185
transform 1 0 70196 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_739
timestamp 1607567185
transform 1 0 69092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_754
timestamp 1607567185
transform 1 0 70472 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[12\]
timestamp 1607567185
transform 1 0 67436 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[356\]
timestamp 1607567185
transform 1 0 66424 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607567185
transform 1 0 65688 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_703
timestamp 1607567185
transform 1 0 65780 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_709
timestamp 1607567185
transform 1 0 66332 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_713
timestamp 1607567185
transform 1 0 66700 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[333\]
timestamp 1607567185
transform 1 0 64308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_679
timestamp 1607567185
transform 1 0 63572 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_690
timestamp 1607567185
transform 1 0 64584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[3\]
timestamp 1607567185
transform 1 0 62744 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_662
timestamp 1607567185
transform 1 0 62008 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[3\]
timestamp 1607567185
transform 1 0 60352 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_8_642
timestamp 1607567185
transform 1 0 60168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607567185
transform 1 0 60076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_633
timestamp 1607567185
transform 1 0 59340 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[7\]
timestamp 1607567185
transform 1 0 57684 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_8_611
timestamp 1607567185
transform 1 0 57316 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_599
timestamp 1607567185
transform 1 0 56212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[121\]
timestamp 1607567185
transform 1 0 54556 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607567185
transform 1 0 54464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_566
timestamp 1607567185
transform 1 0 53176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_578
timestamp 1607567185
transform 1 0 54280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[192\]
timestamp 1607567185
transform 1 0 52900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_555
timestamp 1607567185
transform 1 0 52164 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[111\]
timestamp 1607567185
transform 1 0 50508 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_8_535
timestamp 1607567185
transform 1 0 50324 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[178\]
timestamp 1607567185
transform 1 0 48944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607567185
transform 1 0 48852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_518
timestamp 1607567185
transform 1 0 48760 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_523
timestamp 1607567185
transform 1 0 49220 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[161\]
timestamp 1607567185
transform 1 0 47380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_495
timestamp 1607567185
transform 1 0 46644 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_506
timestamp 1607567185
transform 1 0 47656 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[104\]
timestamp 1607567185
transform 1 0 44988 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[153\]
timestamp 1607567185
transform 1 0 43976 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607567185
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_455
timestamp 1607567185
transform 1 0 42964 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_459
timestamp 1607567185
transform 1 0 43332 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_465
timestamp 1607567185
transform 1 0 43884 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_469
timestamp 1607567185
transform 1 0 44252 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[173\]
timestamp 1607567185
transform 1 0 41952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_439
timestamp 1607567185
transform 1 0 41492 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_443
timestamp 1607567185
transform 1 0 41860 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_447
timestamp 1607567185
transform 1 0 42228 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1607567185
transform 1 0 41032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_416
timestamp 1607567185
transform 1 0 39376 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_428
timestamp 1607567185
transform 1 0 40480 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1607567185
transform 1 0 38180 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_397
timestamp 1607567185
transform 1 0 37628 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_404
timestamp 1607567185
transform 1 0 38272 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_385
timestamp 1607567185
transform 1 0 36524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1607567185
transform 1 0 35328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_366
timestamp 1607567185
transform 1 0 34776 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1607567185
transform 1 0 35420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1607567185
transform 1 0 32476 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_342
timestamp 1607567185
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_354
timestamp 1607567185
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_323
timestamp 1607567185
transform 1 0 30820 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_335
timestamp 1607567185
transform 1 0 31924 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1607567185
transform 1 0 29624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_302
timestamp 1607567185
transform 1 0 28888 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_311
timestamp 1607567185
transform 1 0 29716 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[141\]
timestamp 1607567185
transform 1 0 27508 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_286
timestamp 1607567185
transform 1 0 27416 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_290
timestamp 1607567185
transform 1 0 27784 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1607567185
transform 1 0 26772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1607567185
transform 1 0 26220 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_280
timestamp 1607567185
transform 1 0 26864 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607567185
transform 1 0 23920 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1607567185
transform 1 0 24012 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1607567185
transform 1 0 25116 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_230
timestamp 1607567185
transform 1 0 22264 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_242
timestamp 1607567185
transform 1 0 23368 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607567185
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_211
timestamp 1607567185
transform 1 0 20516 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_218
timestamp 1607567185
transform 1 0 21160 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_199
timestamp 1607567185
transform 1 0 19412 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607567185
transform 1 0 18216 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_174
timestamp 1607567185
transform 1 0 17112 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_187
timestamp 1607567185
transform 1 0 18308 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[5\]
timestamp 1607567185
transform 1 0 15456 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607567185
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_152
timestamp 1607567185
transform 1 0 15088 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_140
timestamp 1607567185
transform 1 0 13984 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[80\]
timestamp 1607567185
transform 1 0 12604 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607567185
transform 1 0 12512 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_118
timestamp 1607567185
transform 1 0 11960 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_128
timestamp 1607567185
transform 1 0 12880 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_106
timestamp 1607567185
transform 1 0 10856 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607567185
transform 1 0 9660 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1607567185
transform 1 0 8556 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1607567185
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_rstn_buf
timestamp 1607567185
transform 1 0 6900 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607567185
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_54
timestamp 1607567185
transform 1 0 6072 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1607567185
transform 1 0 2944 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  mprj_clk_buf
timestamp 1607567185
transform 1 0 4416 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607567185
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_19
timestamp 1607567185
transform 1 0 2852 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_23
timestamp 1607567185
transform 1 0 3220 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1607567185
transform 1 0 4048 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607567185
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607567185
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1607567185
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[94\]
timestamp 1607567185
transform 1 0 40848 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_14_416
timestamp 1607567185
transform 1 0 39376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_428
timestamp 1607567185
transform 1 0 40480 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[86\]
timestamp 1607567185
transform 1 0 37720 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607567185
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_387
timestamp 1607567185
transform 1 0 36708 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_395
timestamp 1607567185
transform 1 0 37444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_363
timestamp 1607567185
transform 1 0 34500 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_375
timestamp 1607567185
transform 1 0 35604 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[136\]
timestamp 1607567185
transform 1 0 33120 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_340
timestamp 1607567185
transform 1 0 32384 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_351
timestamp 1607567185
transform 1 0 33396 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[135\]
timestamp 1607567185
transform 1 0 32108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607567185
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1607567185
transform 1 0 30636 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_333
timestamp 1607567185
transform 1 0 31740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1607567185
transform 1 0 29532 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[67\]
timestamp 1607567185
transform 1 0 27876 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_283
timestamp 1607567185
transform 1 0 27140 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[142\]
timestamp 1607567185
transform 1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607567185
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1607567185
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_276
timestamp 1607567185
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_247
timestamp 1607567185
transform 1 0 23828 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_259
timestamp 1607567185
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_235
timestamp 1607567185
transform 1 0 22724 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[115\]
timestamp 1607567185
transform 1 0 21344 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607567185
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1607567185
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1607567185
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1607567185
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_223
timestamp 1607567185
transform 1 0 21620 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_195
timestamp 1607567185
transform 1 0 19044 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_207
timestamp 1607567185
transform 1 0 20148 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_183
timestamp 1607567185
transform 1 0 17940 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[4\]
timestamp 1607567185
transform 1 0 16284 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[79\]
timestamp 1607567185
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607567185
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_157
timestamp 1607567185
transform 1 0 15548 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[96\]
timestamp 1607567185
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1607567185
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1607567185
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_128
timestamp 1607567185
transform 1 0 12880 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[6\]
timestamp 1607567185
transform 1 0 11224 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_14_105
timestamp 1607567185
transform 1 0 10764 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_109
timestamp 1607567185
transform 1 0 11132 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607567185
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_78
timestamp 1607567185
transform 1 0 8280 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1607567185
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1607567185
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1607567185
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[2\]
timestamp 1607567185
transform 1 0 8004 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_67
timestamp 1607567185
transform 1 0 7268 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[9\]
timestamp 1607567185
transform 1 0 4600 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_14_56
timestamp 1607567185
transform 1 0 6256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[0\]
timestamp 1607567185
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607567185
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1607567185
transform 1 0 2852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1607567185
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1607567185
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607567185
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607567185
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1607567185
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[170\]
timestamp 1607567185
transform 1 0 40940 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607567185
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_416
timestamp 1607567185
transform 1 0 39376 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_424
timestamp 1607567185
transform 1 0 40112 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_428
timestamp 1607567185
transform 1 0 40480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_432
timestamp 1607567185
transform 1 0 40848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[160\]
timestamp 1607567185
transform 1 0 39100 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_405
timestamp 1607567185
transform 1 0 38364 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[74\]
timestamp 1607567185
transform 1 0 36708 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_13_382
timestamp 1607567185
transform 1 0 36248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_386
timestamp 1607567185
transform 1 0 36616 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[150\]
timestamp 1607567185
transform 1 0 34868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607567185
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_365
timestamp 1607567185
transform 1 0 34684 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_370
timestamp 1607567185
transform 1 0 35144 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_353
timestamp 1607567185
transform 1 0 33580 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[62\]
timestamp 1607567185
transform 1 0 31924 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_13_324
timestamp 1607567185
transform 1 0 30912 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_332
timestamp 1607567185
transform 1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[68\]
timestamp 1607567185
transform 1 0 29256 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607567185
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_304
timestamp 1607567185
transform 1 0 29072 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[129\]
timestamp 1607567185
transform 1 0 27324 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_288
timestamp 1607567185
transform 1 0 27600 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_300
timestamp 1607567185
transform 1 0 28704 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_277
timestamp 1607567185
transform 1 0 26588 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[60\]
timestamp 1607567185
transform 1 0 24932 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1607567185
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_257
timestamp 1607567185
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607567185
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_228
timestamp 1607567185
transform 1 0 22080 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1607567185
transform 1 0 23184 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[41\]
timestamp 1607567185
transform 1 0 20424 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_13_208
timestamp 1607567185
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1607567185
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[78\]
timestamp 1607567185
transform 1 0 16744 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607567185
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_173
timestamp 1607567185
transform 1 0 17020 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1607567185
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1607567185
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_162
timestamp 1607567185
transform 1 0 16008 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[22\]
timestamp 1607567185
transform 1 0 14352 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_13_138
timestamp 1607567185
transform 1 0 13800 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[75\]
timestamp 1607567185
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607567185
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1607567185
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_126
timestamp 1607567185
transform 1 0 12696 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[74\]
timestamp 1607567185
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_104
timestamp 1607567185
transform 1 0 10672 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_110
timestamp 1607567185
transform 1 0 11224 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_80
timestamp 1607567185
transform 1 0 8464 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_92
timestamp 1607567185
transform 1 0 9568 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_clk2_buf
timestamp 1607567185
transform 1 0 6808 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607567185
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1607567185
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[7\]
timestamp 1607567185
transform 1 0 4324 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[1\]
timestamp 1607567185
transform 1 0 3312 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_23
timestamp 1607567185
transform 1 0 3220 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1607567185
transform 1 0 3588 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607567185
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607567185
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1607567185
transform 1 0 2484 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_425
timestamp 1607567185
transform 1 0 40204 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[148\]
timestamp 1607567185
transform 1 0 37720 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607567185
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1607567185
transform 1 0 37996 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_413
timestamp 1607567185
transform 1 0 39100 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_381
timestamp 1607567185
transform 1 0 36156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_393
timestamp 1607567185
transform 1 0 37260 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[76\]
timestamp 1607567185
transform 1 0 34500 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_355
timestamp 1607567185
transform 1 0 33764 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[61\]
timestamp 1607567185
transform 1 0 32108 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607567185
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_323
timestamp 1607567185
transform 1 0 30820 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_335
timestamp 1607567185
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[125\]
timestamp 1607567185
transform 1 0 29532 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[128\]
timestamp 1607567185
transform 1 0 30544 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_306
timestamp 1607567185
transform 1 0 29256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_312
timestamp 1607567185
transform 1 0 29808 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_298
timestamp 1607567185
transform 1 0 28520 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[55\]
timestamp 1607567185
transform 1 0 26864 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607567185
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_273
timestamp 1607567185
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1607567185
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[110\]
timestamp 1607567185
transform 1 0 24840 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[134\]
timestamp 1607567185
transform 1 0 23828 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_246
timestamp 1607567185
transform 1 0 23736 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_250
timestamp 1607567185
transform 1 0 24104 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_261
timestamp 1607567185
transform 1 0 25116 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[124\]
timestamp 1607567185
transform 1 0 22724 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_227
timestamp 1607567185
transform 1 0 21988 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_238
timestamp 1607567185
transform 1 0 23000 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[120\]
timestamp 1607567185
transform 1 0 21712 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607567185
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1607567185
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_223
timestamp 1607567185
transform 1 0 21620 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[121\]
timestamp 1607567185
transform 1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_190
timestamp 1607567185
transform 1 0 18584 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_198
timestamp 1607567185
transform 1 0 19320 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1607567185
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[32\]
timestamp 1607567185
transform 1 0 16928 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[109\]
timestamp 1607567185
transform 1 0 15548 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607567185
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1607567185
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_160
timestamp 1607567185
transform 1 0 15824 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[77\]
timestamp 1607567185
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_133
timestamp 1607567185
transform 1 0 13340 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1607567185
transform 1 0 14076 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1607567185
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[76\]
timestamp 1607567185
transform 1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_122
timestamp 1607567185
transform 1 0 12328 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[1\]
timestamp 1607567185
transform 1 0 10672 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_12_96
timestamp 1607567185
transform 1 0 9936 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[95\]
timestamp 1607567185
transform 1 0 8372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[98\]
timestamp 1607567185
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607567185
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_82
timestamp 1607567185
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1607567185
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[81\]
timestamp 1607567185
transform 1 0 7360 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_60
timestamp 1607567185
transform 1 0 6624 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_71
timestamp 1607567185
transform 1 0 7636 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[8\]
timestamp 1607567185
transform 1 0 4968 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_12_40
timestamp 1607567185
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[86\]
timestamp 1607567185
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607567185
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp 1607567185
transform 1 0 2852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1607567185
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1607567185
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607567185
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607567185
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1607567185
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607567185
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_418
timestamp 1607567185
transform 1 0 39560 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_426
timestamp 1607567185
transform 1 0 40296 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_428
timestamp 1607567185
transform 1 0 40480 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_406
timestamp 1607567185
transform 1 0 38456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[72\]
timestamp 1607567185
transform 1 0 36800 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_11_379
timestamp 1607567185
transform 1 0 35972 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_387
timestamp 1607567185
transform 1 0 36708 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607567185
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_364
timestamp 1607567185
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1607567185
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_352
timestamp 1607567185
transform 1 0 33488 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[54\]
timestamp 1607567185
transform 1 0 31832 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_11_326
timestamp 1607567185
transform 1 0 31096 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[51\]
timestamp 1607567185
transform 1 0 29440 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607567185
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_306
timestamp 1607567185
transform 1 0 29256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[131\]
timestamp 1607567185
transform 1 0 27232 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_287
timestamp 1607567185
transform 1 0 27508 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_299
timestamp 1607567185
transform 1 0 28612 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_276
timestamp 1607567185
transform 1 0 26496 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[36\]
timestamp 1607567185
transform 1 0 24840 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[127\]
timestamp 1607567185
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_248
timestamp 1607567185
transform 1 0 23920 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_256
timestamp 1607567185
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607567185
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_228
timestamp 1607567185
transform 1 0 22080 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_240
timestamp 1607567185
transform 1 0 23184 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[47\]
timestamp 1607567185
transform 1 0 20424 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_11_202
timestamp 1607567185
transform 1 0 19688 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[34\]
timestamp 1607567185
transform 1 0 18032 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607567185
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1607567185
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_167
timestamp 1607567185
transform 1 0 16468 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[3\]
timestamp 1607567185
transform 1 0 14812 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_11_141
timestamp 1607567185
transform 1 0 14076 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[2\]
timestamp 1607567185
transform 1 0 12420 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607567185
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_114
timestamp 1607567185
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[0\]
timestamp 1607567185
transform 1 0 9936 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_11_85
timestamp 1607567185
transform 1 0 8924 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_93
timestamp 1607567185
transform 1 0 9660 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[21\]
timestamp 1607567185
transform 1 0 7268 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607567185
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1607567185
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_66
timestamp 1607567185
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_53
timestamp 1607567185
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[12\]
timestamp 1607567185
transform 1 0 4324 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[82\]
timestamp 1607567185
transform 1 0 3312 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 1607567185
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_27
timestamp 1607567185
transform 1 0 3588 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607567185
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607567185
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 1607567185
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607567185
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_417
timestamp 1607567185
transform 1 0 39468 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_425
timestamp 1607567185
transform 1 0 40204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_428
timestamp 1607567185
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_417
timestamp 1607567185
transform 1 0 39468 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_429
timestamp 1607567185
transform 1 0 40572 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[82\]
timestamp 1607567185
transform 1 0 37812 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[146\]
timestamp 1607567185
transform 1 0 38088 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607567185
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_398
timestamp 1607567185
transform 1 0 37720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_405
timestamp 1607567185
transform 1 0 38364 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[156\]
timestamp 1607567185
transform 1 0 36616 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_391
timestamp 1607567185
transform 1 0 37076 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_378
timestamp 1607567185
transform 1 0 35880 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_389
timestamp 1607567185
transform 1 0 36892 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[77\]
timestamp 1607567185
transform 1 0 35420 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[139\]
timestamp 1607567185
transform 1 0 34500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607567185
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_367
timestamp 1607567185
transform 1 0 34868 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_366
timestamp 1607567185
transform 1 0 34776 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_354
timestamp 1607567185
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1607567185
transform 1 0 33764 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[58\]
timestamp 1607567185
transform 1 0 32016 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[65\]
timestamp 1607567185
transform 1 0 32108 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[137\]
timestamp 1607567185
transform 1 0 31004 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607567185
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp 1607567185
transform 1 0 31280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_328
timestamp 1607567185
transform 1 0 31280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[63\]
timestamp 1607567185
transform 1 0 29624 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[126\]
timestamp 1607567185
transform 1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607567185
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_306
timestamp 1607567185
transform 1 0 29256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_305
timestamp 1607567185
transform 1 0 29164 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_317
timestamp 1607567185
transform 1 0 30268 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_297
timestamp 1607567185
transform 1 0 28428 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_294
timestamp 1607567185
transform 1 0 28152 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[56\]
timestamp 1607567185
transform 1 0 26772 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[57\]
timestamp 1607567185
transform 1 0 26496 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607567185
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1607567185
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[50\]
timestamp 1607567185
transform 1 0 23644 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[53\]
timestamp 1607567185
transform 1 0 23644 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_9_263
timestamp 1607567185
transform 1 0 25300 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1607567185
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607567185
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1607567185
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_237
timestamp 1607567185
transform 1 0 22908 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[43\]
timestamp 1607567185
transform 1 0 20792 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[46\]
timestamp 1607567185
transform 1 0 21252 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607567185
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1607567185
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[108\]
timestamp 1607567185
transform 1 0 18676 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_202
timestamp 1607567185
transform 1 0 19688 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_194
timestamp 1607567185
transform 1 0 18952 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_206
timestamp 1607567185
transform 1 0 20056 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[38\]
timestamp 1607567185
transform 1 0 18032 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[106\]
timestamp 1607567185
transform 1 0 17664 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607567185
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1607567185
transform 1 0 17204 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_172
timestamp 1607567185
transform 1 0 16928 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_183
timestamp 1607567185
transform 1 0 17940 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[35\]
timestamp 1607567185
transform 1 0 15548 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[37\]
timestamp 1607567185
transform 1 0 15272 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607567185
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1607567185
transform 1 0 15180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1607567185
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[107\]
timestamp 1607567185
transform 1 0 13984 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_141
timestamp 1607567185
transform 1 0 14076 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 1607567185
transform 1 0 13248 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_143
timestamp 1607567185
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[30\]
timestamp 1607567185
transform 1 0 12420 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[111\]
timestamp 1607567185
transform 1 0 12972 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607567185
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1607567185
transform 1 0 11592 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_121
timestamp 1607567185
transform 1 0 12236 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[24\]
timestamp 1607567185
transform 1 0 10580 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[104\]
timestamp 1607567185
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[94\]
timestamp 1607567185
transform 1 0 10212 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1607567185
transform 1 0 10488 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_110
timestamp 1607567185
transform 1 0 11224 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1607567185
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[91\]
timestamp 1607567185
transform 1 0 9200 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607567185
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_80
timestamp 1607567185
transform 1 0 8464 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_91
timestamp 1607567185
transform 1 0 9476 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_83
timestamp 1607567185
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1607567185
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1607567185
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[15\]
timestamp 1607567185
transform 1 0 6808 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[18\]
timestamp 1607567185
transform 1 0 7084 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607567185
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_57
timestamp 1607567185
transform 1 0 6348 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[11\]
timestamp 1607567185
transform 1 0 4692 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1607567185
transform 1 0 5980 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1607567185
transform 1 0 4600 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1607567185
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[16\]
timestamp 1607567185
transform 1 0 4324 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[83\]
timestamp 1607567185
transform 1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607567185
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_23
timestamp 1607567185
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1607567185
transform 1 0 3588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_19
timestamp 1607567185
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1607567185
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1607567185
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607567185
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607567185
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607567185
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1607567185
transform 1 0 2484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1607567185
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1607567185
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[172\]
timestamp 1607567185
transform 1 0 40112 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_416
timestamp 1607567185
transform 1 0 39376 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_427
timestamp 1607567185
transform 1 0 40388 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[80\]
timestamp 1607567185
transform 1 0 37720 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607567185
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[151\]
timestamp 1607567185
transform 1 0 36064 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_377
timestamp 1607567185
transform 1 0 35788 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_383
timestamp 1607567185
transform 1 0 36340 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_395
timestamp 1607567185
transform 1 0 37444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_369
timestamp 1607567185
transform 1 0 35052 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[71\]
timestamp 1607567185
transform 1 0 33396 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[132\]
timestamp 1607567185
transform 1 0 32384 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_343
timestamp 1607567185
transform 1 0 32660 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[144\]
timestamp 1607567185
transform 1 0 31004 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607567185
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_328
timestamp 1607567185
transform 1 0 31280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_337
timestamp 1607567185
transform 1 0 32108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_317
timestamp 1607567185
transform 1 0 30268 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[52\]
timestamp 1607567185
transform 1 0 28612 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[130\]
timestamp 1607567185
transform 1 0 27600 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_287
timestamp 1607567185
transform 1 0 27508 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_291
timestamp 1607567185
transform 1 0 27876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[123\]
timestamp 1607567185
transform 1 0 26496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607567185
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_279
timestamp 1607567185
transform 1 0 26772 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[49\]
timestamp 1607567185
transform 1 0 23644 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1607567185
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_237
timestamp 1607567185
transform 1 0 22908 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[44\]
timestamp 1607567185
transform 1 0 21252 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607567185
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1607567185
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_206
timestamp 1607567185
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[42\]
timestamp 1607567185
transform 1 0 18400 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_8_172
timestamp 1607567185
transform 1 0 16928 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1607567185
transform 1 0 18032 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[33\]
timestamp 1607567185
transform 1 0 15272 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607567185
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_137
timestamp 1607567185
transform 1 0 13708 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1607567185
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_8  la_buf\[28\]
timestamp 1607567185
transform 1 0 12052 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_111
timestamp 1607567185
transform 1 0 11316 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[20\]
timestamp 1607567185
transform 1 0 9660 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[89\]
timestamp 1607567185
transform 1 0 8280 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607567185
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_81
timestamp 1607567185
transform 1 0 8556 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1607567185
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[85\]
timestamp 1607567185
transform 1 0 7268 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_59
timestamp 1607567185
transform 1 0 6532 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_70
timestamp 1607567185
transform 1 0 7544 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[13\]
timestamp 1607567185
transform 1 0 4876 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_8_40
timestamp 1607567185
transform 1 0 4784 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[87\]
timestamp 1607567185
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607567185
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1607567185
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1607567185
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[90\]
timestamp 1607567185
transform 1 0 1932 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607567185
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1607567185
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_12
timestamp 1607567185
transform 1 0 2208 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607567185
transform -1 0 198812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_2143
timestamp 1607567185
transform 1 0 198260 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 1607567185
transform 1 0 195868 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp 1607567185
transform 1 0 196880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2120
timestamp 1607567185
transform 1 0 196144 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_2131
timestamp 1607567185
transform 1 0 197156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1607567185
transform 1 0 194856 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1607567185
transform 1 0 194764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2097
timestamp 1607567185
transform 1 0 194028 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2109
timestamp 1607567185
transform 1 0 195132 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1607567185
transform 1 0 193752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1607567185
transform 1 0 192556 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2084
timestamp 1607567185
transform 1 0 192832 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_2092
timestamp 1607567185
transform 1 0 193568 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1607567185
transform 1 0 190532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1607567185
transform 1 0 191544 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2062
timestamp 1607567185
transform 1 0 190808 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2073
timestamp 1607567185
transform 1 0 191820 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1607567185
transform 1 0 189244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1607567185
transform 1 0 189152 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2040
timestamp 1607567185
transform 1 0 188784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2048
timestamp 1607567185
transform 1 0 189520 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_2056
timestamp 1607567185
transform 1 0 190256 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_2028
timestamp 1607567185
transform 1 0 187680 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[22\]
timestamp 1607567185
transform 1 0 186024 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2002
timestamp 1607567185
transform 1 0 185288 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[25\]
timestamp 1607567185
transform 1 0 183632 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1607567185
transform 1 0 183540 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1975
timestamp 1607567185
transform 1 0 182804 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[24\]
timestamp 1607567185
transform 1 0 181148 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1949
timestamp 1607567185
transform 1 0 180412 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[24\]
timestamp 1607567185
transform 1 0 178756 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1607567185
transform 1 0 176916 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1607567185
transform 1 0 177928 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1910
timestamp 1607567185
transform 1 0 176824 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1914
timestamp 1607567185
transform 1 0 177192 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1923
timestamp 1607567185
transform 1 0 178020 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1607567185
transform 1 0 174800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1607567185
transform 1 0 175812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1891
timestamp 1607567185
transform 1 0 175076 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1902
timestamp 1607567185
transform 1 0 176088 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1880
timestamp 1607567185
transform 1 0 174064 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[6\]
timestamp 1607567185
transform 1 0 172408 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1607567185
transform 1 0 172316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1851
timestamp 1607567185
transform 1 0 171396 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1859
timestamp 1607567185
transform 1 0 172132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1607567185
transform 1 0 171120 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1842
timestamp 1607567185
transform 1 0 170568 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1607567185
transform 1 0 169188 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1813
timestamp 1607567185
transform 1 0 167900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1825
timestamp 1607567185
transform 1 0 169004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1830
timestamp 1607567185
transform 1 0 169464 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[28\]
timestamp 1607567185
transform 1 0 167624 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1607567185
transform 1 0 166704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1801
timestamp 1607567185
transform 1 0 166796 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1809
timestamp 1607567185
transform 1 0 167532 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1607567185
transform 1 0 164680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[57\]
timestamp 1607567185
transform 1 0 165692 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1776
timestamp 1607567185
transform 1 0 164496 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1781
timestamp 1607567185
transform 1 0 164956 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1792
timestamp 1607567185
transform 1 0 165968 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1607567185
transform 1 0 163116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1764
timestamp 1607567185
transform 1 0 163392 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1607567185
transform 1 0 161184 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1607567185
transform 1 0 161092 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1743
timestamp 1607567185
transform 1 0 161460 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1755
timestamp 1607567185
transform 1 0 162564 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607567185
transform -1 0 198812 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607567185
transform -1 0 198812 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1607567185
transform 1 0 197892 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1607567185
transform 1 0 197524 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2133
timestamp 1607567185
transform 1 0 197340 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2140
timestamp 1607567185
transform 1 0 197984 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2134
timestamp 1607567185
transform 1 0 197432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2136
timestamp 1607567185
transform 1 0 197616 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2144
timestamp 1607567185
transform 1 0 198352 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1607567185
transform 1 0 195684 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_2121
timestamp 1607567185
transform 1 0 196236 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_2118
timestamp 1607567185
transform 1 0 195960 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2130
timestamp 1607567185
transform 1 0 197064 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  mprj2_pwrgood
timestamp 1607567185
transform 1 0 193844 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  mprj_pwrgood
timestamp 1607567185
transform 1 0 195132 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1607567185
transform 1 0 195040 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2100
timestamp 1607567185
transform 1 0 194304 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2107
timestamp 1607567185
transform 1 0 194948 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1607567185
transform 1 0 192832 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  mprj2_vdd_pwrgood
timestamp 1607567185
transform 1 0 193200 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1607567185
transform 1 0 192188 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2078
timestamp 1607567185
transform 1 0 192280 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2086
timestamp 1607567185
transform 1 0 193016 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2083
timestamp 1607567185
transform 1 0 192740 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2087
timestamp 1607567185
transform 1 0 193108 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1607567185
transform 1 0 191176 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1607567185
transform 1 0 190532 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1607567185
transform 1 0 191912 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2062
timestamp 1607567185
transform 1 0 190808 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2069
timestamp 1607567185
transform 1 0 191452 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_2062
timestamp 1607567185
transform 1 0 190808 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2075
timestamp 1607567185
transform 1 0 192004 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1607567185
transform 1 0 189520 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1607567185
transform 1 0 189428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1607567185
transform 1 0 189336 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2045
timestamp 1607567185
transform 1 0 189244 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_2050
timestamp 1607567185
transform 1 0 189704 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_2045
timestamp 1607567185
transform 1 0 189244 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2051
timestamp 1607567185
transform 1 0 189796 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1607567185
transform 1 0 187864 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1607567185
transform 1 0 188232 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1607567185
transform 1 0 187220 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2022
timestamp 1607567185
transform 1 0 187128 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2026
timestamp 1607567185
transform 1 0 187496 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2037
timestamp 1607567185
transform 1 0 188508 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2029
timestamp 1607567185
transform 1 0 187772 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_2033
timestamp 1607567185
transform 1 0 188140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1607567185
transform 1 0 186392 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1607567185
transform 1 0 185288 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1607567185
transform 1 0 186484 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1607567185
transform 1 0 186300 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2009
timestamp 1607567185
transform 1 0 185932 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2016
timestamp 1607567185
transform 1 0 186576 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2005
timestamp 1607567185
transform 1 0 185564 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_2017
timestamp 1607567185
transform 1 0 186668 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1607567185
transform 1 0 183632 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1607567185
transform 1 0 184552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1607567185
transform 1 0 183632 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1985
timestamp 1607567185
transform 1 0 183724 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1993
timestamp 1607567185
transform 1 0 184460 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1997
timestamp 1607567185
transform 1 0 184828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1987
timestamp 1607567185
transform 1 0 183908 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1999
timestamp 1607567185
transform 1 0 185012 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1607567185
transform 1 0 181884 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1607567185
transform 1 0 182252 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1972
timestamp 1607567185
transform 1 0 182528 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1968
timestamp 1607567185
transform 1 0 182160 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1980
timestamp 1607567185
transform 1 0 183264 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1957
timestamp 1607567185
transform 1 0 181148 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1953
timestamp 1607567185
transform 1 0 180780 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1961
timestamp 1607567185
transform 1 0 181516 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1954
timestamp 1607567185
transform 1 0 180872 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1607567185
transform 1 0 180780 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1607567185
transform 1 0 181240 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1607567185
transform 1 0 180872 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1949
timestamp 1607567185
transform 1 0 180412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1950
timestamp 1607567185
transform 1 0 180504 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1607567185
transform 1 0 180688 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1607567185
transform 1 0 178388 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1607567185
transform 1 0 179400 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1607567185
transform 1 0 179124 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1927
timestamp 1607567185
transform 1 0 178388 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1938
timestamp 1607567185
transform 1 0 179400 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1930
timestamp 1607567185
transform 1 0 178664 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1941
timestamp 1607567185
transform 1 0 179676 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1607567185
transform 1 0 178112 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1607567185
transform 1 0 177100 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1607567185
transform 1 0 177928 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1906
timestamp 1607567185
transform 1 0 176456 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1918
timestamp 1607567185
transform 1 0 177560 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1923
timestamp 1607567185
transform 1 0 178020 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1907
timestamp 1607567185
transform 1 0 176548 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1916
timestamp 1607567185
transform 1 0 177376 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1924
timestamp 1607567185
transform 1 0 178112 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1607567185
transform 1 0 175168 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1607567185
transform 1 0 175168 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1607567185
transform 1 0 176180 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1607567185
transform 1 0 175076 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1607567185
transform 1 0 175076 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1895
timestamp 1607567185
transform 1 0 175444 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1888
timestamp 1607567185
transform 1 0 174800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1895
timestamp 1607567185
transform 1 0 175444 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1607567185
transform 1 0 173328 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1607567185
transform 1 0 173788 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1875
timestamp 1607567185
transform 1 0 173604 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1887
timestamp 1607567185
transform 1 0 174708 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1869
timestamp 1607567185
transform 1 0 173052 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1880
timestamp 1607567185
transform 1 0 174064 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1607567185
transform 1 0 172316 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[19\]
timestamp 1607567185
transform 1 0 171396 0 1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1607567185
transform 1 0 172224 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1852
timestamp 1607567185
transform 1 0 171488 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1864
timestamp 1607567185
transform 1 0 172592 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1850
timestamp 1607567185
transform 1 0 171304 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1607567185
transform 1 0 169740 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1607567185
transform 1 0 169556 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1607567185
transform 1 0 171212 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1836
timestamp 1607567185
transform 1 0 170016 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1848
timestamp 1607567185
transform 1 0 171120 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1834
timestamp 1607567185
transform 1 0 169832 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1846
timestamp 1607567185
transform 1 0 170936 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1607567185
transform 1 0 168452 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[458\]
timestamp 1607567185
transform 1 0 168360 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1607567185
transform 1 0 169372 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1607567185
transform 1 0 169464 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1821
timestamp 1607567185
transform 1 0 168636 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1830
timestamp 1607567185
transform 1 0 169464 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1822
timestamp 1607567185
transform 1 0 168728 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[48\]
timestamp 1607567185
transform 1 0 167440 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[55\]
timestamp 1607567185
transform 1 0 167348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1607567185
transform 1 0 166520 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1799
timestamp 1607567185
transform 1 0 166612 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1810
timestamp 1607567185
transform 1 0 167624 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1803
timestamp 1607567185
transform 1 0 166980 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1807
timestamp 1607567185
transform 1 0 167348 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1811
timestamp 1607567185
transform 1 0 167716 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1607567185
transform 1 0 164588 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1607567185
transform 1 0 165600 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[59\]
timestamp 1607567185
transform 1 0 165508 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[60\]
timestamp 1607567185
transform 1 0 164496 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1779
timestamp 1607567185
transform 1 0 164772 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1790
timestamp 1607567185
transform 1 0 165784 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1776
timestamp 1607567185
transform 1 0 164496 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1780
timestamp 1607567185
transform 1 0 164864 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1791
timestamp 1607567185
transform 1 0 165876 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1607567185
transform 1 0 162656 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1607567185
transform 1 0 162748 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1607567185
transform 1 0 163668 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1607567185
transform 1 0 163852 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1759
timestamp 1607567185
transform 1 0 162932 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1768
timestamp 1607567185
transform 1 0 163760 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1760
timestamp 1607567185
transform 1 0 163024 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1768
timestamp 1607567185
transform 1 0 163760 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1770
timestamp 1607567185
transform 1 0 163944 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1607567185
transform 1 0 160908 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1607567185
transform 1 0 161736 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1740
timestamp 1607567185
transform 1 0 161184 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1752
timestamp 1607567185
transform 1 0 162288 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1738
timestamp 1607567185
transform 1 0 161000 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1749
timestamp 1607567185
transform 1 0 162012 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607567185
transform -1 0 154560 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1657
timestamp 1607567185
transform 1 0 153548 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1648
timestamp 1607567185
transform 1 0 152720 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607567185
transform 1 0 152628 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[58\]
timestamp 1607567185
transform 1 0 153272 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1635
timestamp 1607567185
transform 1 0 151524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1623
timestamp 1607567185
transform 1 0 150420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1611
timestamp 1607567185
transform 1 0 149316 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1599
timestamp 1607567185
transform 1 0 148212 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1587
timestamp 1607567185
transform 1 0 147108 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607567185
transform 1 0 147016 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1574
timestamp 1607567185
transform 1 0 145912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1562
timestamp 1607567185
transform 1 0 144808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1541
timestamp 1607567185
transform 1 0 142876 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1529
timestamp 1607567185
transform 1 0 141772 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[14\]
timestamp 1607567185
transform 1 0 143152 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1521
timestamp 1607567185
transform 1 0 141036 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607567185
transform 1 0 141404 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[449\]
timestamp 1607567185
transform 1 0 141496 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1509
timestamp 1607567185
transform 1 0 139932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[83\]
timestamp 1607567185
transform 1 0 138276 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1483
timestamp 1607567185
transform 1 0 137540 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1461
timestamp 1607567185
transform 1 0 135516 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1453
timestamp 1607567185
transform 1 0 134780 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607567185
transform 1 0 135792 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[81\]
timestamp 1607567185
transform 1 0 135884 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1442
timestamp 1607567185
transform 1 0 133768 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[260\]
timestamp 1607567185
transform 1 0 134504 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[259\]
timestamp 1607567185
transform 1 0 133492 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1431
timestamp 1607567185
transform 1 0 132756 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1412
timestamp 1607567185
transform 1 0 131008 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1404
timestamp 1607567185
transform 1 0 130272 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1401
timestamp 1607567185
transform 1 0 129996 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607567185
transform 1 0 130180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[11\]
timestamp 1607567185
transform 1 0 131100 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1389
timestamp 1607567185
transform 1 0 128892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1369
timestamp 1607567185
transform 1 0 127052 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1361
timestamp 1607567185
transform 1 0 126316 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[50\]
timestamp 1607567185
transform 1 0 127236 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607567185
transform 1 0 124568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[52\]
timestamp 1607567185
transform 1 0 124660 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1334
timestamp 1607567185
transform 1 0 123832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1325
timestamp 1607567185
transform 1 0 123004 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1607567185
transform 1 0 123556 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1313
timestamp 1607567185
transform 1 0 121900 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1662
timestamp 1607567185
transform 1 0 154008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607567185
transform -1 0 154560 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1654
timestamp 1607567185
transform 1 0 153272 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1642
timestamp 1607567185
transform 1 0 152168 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1630
timestamp 1607567185
transform 1 0 151064 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1618
timestamp 1607567185
transform 1 0 149960 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1605
timestamp 1607567185
transform 1 0 148764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607567185
transform 1 0 149868 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1593
timestamp 1607567185
transform 1 0 147660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1581
timestamp 1607567185
transform 1 0 146556 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1569
timestamp 1607567185
transform 1 0 145452 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1557
timestamp 1607567185
transform 1 0 144348 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1555
timestamp 1607567185
transform 1 0 144164 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1551
timestamp 1607567185
transform 1 0 143796 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607567185
transform 1 0 144256 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1539
timestamp 1607567185
transform 1 0 142692 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[456\]
timestamp 1607567185
transform 1 0 142416 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1528
timestamp 1607567185
transform 1 0 141680 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[15\]
timestamp 1607567185
transform 1 0 140024 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1507
timestamp 1607567185
transform 1 0 139748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1499
timestamp 1607567185
transform 1 0 139012 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1492
timestamp 1607567185
transform 1 0 138368 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607567185
transform 1 0 138644 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[289\]
timestamp 1607567185
transform 1 0 138736 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1484
timestamp 1607567185
transform 1 0 137632 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1473
timestamp 1607567185
transform 1 0 136620 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[285\]
timestamp 1607567185
transform 1 0 137356 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1454
timestamp 1607567185
transform 1 0 134872 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[60\]
timestamp 1607567185
transform 1 0 134964 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1446
timestamp 1607567185
transform 1 0 134136 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1435
timestamp 1607567185
transform 1 0 133124 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _660_
timestamp 1607567185
transform 1 0 133860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1431
timestamp 1607567185
transform 1 0 132756 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1423
timestamp 1607567185
transform 1 0 132020 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607567185
transform 1 0 133032 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _656_
timestamp 1607567185
transform 1 0 131744 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1412
timestamp 1607567185
transform 1 0 131008 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1401
timestamp 1607567185
transform 1 0 129996 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _651_
timestamp 1607567185
transform 1 0 130732 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1382
timestamp 1607567185
transform 1 0 128248 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_adr_buf\[0\]
timestamp 1607567185
transform 1 0 128340 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1374
timestamp 1607567185
transform 1 0 127512 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1365
timestamp 1607567185
transform 1 0 126684 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607567185
transform 1 0 127420 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[51\]
timestamp 1607567185
transform 1 0 125028 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1339
timestamp 1607567185
transform 1 0 124292 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1313
timestamp 1607567185
transform 1 0 121900 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1311
timestamp 1607567185
transform 1 0 121716 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1307
timestamp 1607567185
transform 1 0 121348 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607567185
transform 1 0 121808 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_sel_buf\[1\]
timestamp 1607567185
transform 1 0 122636 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1664
timestamp 1607567185
transform 1 0 154192 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1662
timestamp 1607567185
transform 1 0 154008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607567185
transform -1 0 154560 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607567185
transform -1 0 154560 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1660
timestamp 1607567185
transform 1 0 153824 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1648
timestamp 1607567185
transform 1 0 152720 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1654
timestamp 1607567185
transform 1 0 153272 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1642
timestamp 1607567185
transform 1 0 152168 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607567185
transform 1 0 152628 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1635
timestamp 1607567185
transform 1 0 151524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1623
timestamp 1607567185
transform 1 0 150420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1630
timestamp 1607567185
transform 1 0 151064 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1611
timestamp 1607567185
transform 1 0 149316 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1618
timestamp 1607567185
transform 1 0 149960 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1609
timestamp 1607567185
transform 1 0 149132 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1607567185
transform 1 0 149868 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1607567185
transform 1 0 148856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1599
timestamp 1607567185
transform 1 0 148212 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1587
timestamp 1607567185
transform 1 0 147108 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1598
timestamp 1607567185
transform 1 0 148120 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1586
timestamp 1607567185
transform 1 0 147016 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607567185
transform 1 0 147016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1584
timestamp 1607567185
transform 1 0 146832 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1576
timestamp 1607567185
transform 1 0 146096 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1574
timestamp 1607567185
transform 1 0 145912 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1564
timestamp 1607567185
transform 1 0 144992 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1552
timestamp 1607567185
transform 1 0 143888 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1562
timestamp 1607567185
transform 1 0 144808 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1548
timestamp 1607567185
transform 1 0 143520 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1607567185
transform 1 0 144624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1607567185
transform 1 0 144256 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1607567185
transform 1 0 144348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1540
timestamp 1607567185
transform 1 0 142784 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1529
timestamp 1607567185
transform 1 0 141772 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1536
timestamp 1607567185
transform 1 0 142416 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[53\]
timestamp 1607567185
transform 1 0 142508 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1607567185
transform 1 0 142140 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1517
timestamp 1607567185
transform 1 0 140668 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1521
timestamp 1607567185
transform 1 0 141036 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1510
timestamp 1607567185
transform 1 0 140024 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607567185
transform 1 0 141404 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[455\]
timestamp 1607567185
transform 1 0 140760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[453\]
timestamp 1607567185
transform 1 0 141496 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[25\]
timestamp 1607567185
transform 1 0 140392 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1506
timestamp 1607567185
transform 1 0 139656 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1499
timestamp 1607567185
transform 1 0 139012 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1494
timestamp 1607567185
transform 1 0 138552 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1607567185
transform 1 0 138644 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[44\]
timestamp 1607567185
transform 1 0 139748 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[321\]
timestamp 1607567185
transform 1 0 138736 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1487
timestamp 1607567185
transform 1 0 137908 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1479
timestamp 1607567185
transform 1 0 137172 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1486
timestamp 1607567185
transform 1 0 137816 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1475
timestamp 1607567185
transform 1 0 136804 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1607567185
transform 1 0 137356 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[63\]
timestamp 1607567185
transform 1 0 138000 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[265\]
timestamp 1607567185
transform 1 0 136896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1607567185
transform 1 0 137540 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1468
timestamp 1607567185
transform 1 0 136160 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1462
timestamp 1607567185
transform 1 0 135608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607567185
transform 1 0 135792 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[58\]
timestamp 1607567185
transform 1 0 135148 0 -1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _659_
timestamp 1607567185
transform 1 0 135884 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1450
timestamp 1607567185
transform 1 0 134504 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1449
timestamp 1607567185
transform 1 0 134412 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1438
timestamp 1607567185
transform 1 0 133400 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _658_
timestamp 1607567185
transform 1 0 134136 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1607567185
transform 1 0 133124 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1424
timestamp 1607567185
transform 1 0 132112 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1433
timestamp 1607567185
transform 1 0 132940 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1429
timestamp 1607567185
transform 1 0 132572 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1417
timestamp 1607567185
transform 1 0 131468 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1607567185
transform 1 0 133032 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[65\]
timestamp 1607567185
transform 1 0 132848 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1404
timestamp 1607567185
transform 1 0 130272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1402
timestamp 1607567185
transform 1 0 130088 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1398
timestamp 1607567185
transform 1 0 129720 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607567185
transform 1 0 130180 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[61\]
timestamp 1607567185
transform 1 0 130456 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[54\]
timestamp 1607567185
transform 1 0 129812 0 -1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1386
timestamp 1607567185
transform 1 0 128616 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1387
timestamp 1607567185
transform 1 0 128708 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1382
timestamp 1607567185
transform 1 0 128248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1607567185
transform 1 0 128432 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1607567185
transform 1 0 128340 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1375
timestamp 1607567185
transform 1 0 127604 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1374
timestamp 1607567185
transform 1 0 127512 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1372
timestamp 1607567185
transform 1 0 127328 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1360
timestamp 1607567185
transform 1 0 126224 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1607567185
transform 1 0 127420 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  mprj_dat_buf\[2\]
timestamp 1607567185
transform 1 0 125948 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1607567185
transform 1 0 125948 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1607567185
transform 1 0 125764 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1354
timestamp 1607567185
transform 1 0 125672 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1607567185
transform 1 0 124936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607567185
transform 1 0 124568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1348
timestamp 1607567185
transform 1 0 125120 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1341
timestamp 1607567185
transform 1 0 124476 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1343
timestamp 1607567185
transform 1 0 124660 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1349
timestamp 1607567185
transform 1 0 125212 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1333
timestamp 1607567185
transform 1 0 123740 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1327
timestamp 1607567185
transform 1 0 123188 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[35\]
timestamp 1607567185
transform 1 0 123464 0 -1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1607567185
transform 1 0 123464 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1315
timestamp 1607567185
transform 1 0 122084 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1318
timestamp 1607567185
transform 1 0 122360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1313
timestamp 1607567185
transform 1 0 121900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1310
timestamp 1607567185
transform 1 0 121624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1607567185
transform 1 0 121808 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _638_
timestamp 1607567185
transform 1 0 122084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1664
timestamp 1607567185
transform 1 0 154192 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607567185
transform -1 0 154560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1660
timestamp 1607567185
transform 1 0 153824 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1648
timestamp 1607567185
transform 1 0 152720 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1644
timestamp 1607567185
transform 1 0 152352 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1607567185
transform 1 0 152628 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1636
timestamp 1607567185
transform 1 0 151616 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1631
timestamp 1607567185
transform 1 0 151156 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1623
timestamp 1607567185
transform 1 0 150420 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1607567185
transform 1 0 151340 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1611
timestamp 1607567185
transform 1 0 149316 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1599
timestamp 1607567185
transform 1 0 148212 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1587
timestamp 1607567185
transform 1 0 147108 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1607567185
transform 1 0 147016 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1580
timestamp 1607567185
transform 1 0 146464 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1568
timestamp 1607567185
transform 1 0 145360 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1561
timestamp 1607567185
transform 1 0 144716 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1553
timestamp 1607567185
transform 1 0 143980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1607567185
transform 1 0 144900 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1607567185
transform 1 0 145084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1541
timestamp 1607567185
transform 1 0 142876 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1529
timestamp 1607567185
transform 1 0 141772 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1517
timestamp 1607567185
transform 1 0 140668 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1607567185
transform 1 0 141404 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[7\]
timestamp 1607567185
transform 1 0 141496 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[457\]
timestamp 1607567185
transform 1 0 140392 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1506
timestamp 1607567185
transform 1 0 139656 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1495
timestamp 1607567185
transform 1 0 138644 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[452\]
timestamp 1607567185
transform 1 0 139380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1607567185
transform 1 0 138368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1484
timestamp 1607567185
transform 1 0 137632 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1476
timestamp 1607567185
transform 1 0 136896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1607567185
transform 1 0 137172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1607567185
transform 1 0 137356 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1468
timestamp 1607567185
transform 1 0 136160 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1456
timestamp 1607567185
transform 1 0 135056 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1607567185
transform 1 0 135792 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp 1607567185
transform 1 0 134780 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1607567185
transform 1 0 135884 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1445
timestamp 1607567185
transform 1 0 134044 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1425
timestamp 1607567185
transform 1 0 132204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1417
timestamp 1607567185
transform 1 0 131468 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[67\]
timestamp 1607567185
transform 1 0 132388 0 1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1412
timestamp 1607567185
transform 1 0 131008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1404
timestamp 1607567185
transform 1 0 130272 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1607567185
transform 1 0 130180 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1607567185
transform 1 0 131192 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1391
timestamp 1607567185
transform 1 0 129076 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1380
timestamp 1607567185
transform 1 0 128064 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1607567185
transform 1 0 128616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1607567185
transform 1 0 128800 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[99\]
timestamp 1607567185
transform 1 0 126408 0 1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1354
timestamp 1607567185
transform 1 0 125672 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1343
timestamp 1607567185
transform 1 0 124660 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1341
timestamp 1607567185
transform 1 0 124476 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1607567185
transform 1 0 124568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _634_
timestamp 1607567185
transform 1 0 125396 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1333
timestamp 1607567185
transform 1 0 123740 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1324
timestamp 1607567185
transform 1 0 122912 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1607567185
transform 1 0 123464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1312
timestamp 1607567185
transform 1 0 121808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _633_
timestamp 1607567185
transform 1 0 121532 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1731
timestamp 1607567185
transform 1 0 160356 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1720
timestamp 1607567185
transform 1 0 159344 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[63\]
timestamp 1607567185
transform 1 0 159068 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[61\]
timestamp 1607567185
transform 1 0 160080 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1709
timestamp 1607567185
transform 1 0 158332 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1698
timestamp 1607567185
transform 1 0 157320 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[66\]
timestamp 1607567185
transform 1 0 158056 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1691
timestamp 1607567185
transform 1 0 156676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[70\]
timestamp 1607567185
transform 1 0 157044 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1679
timestamp 1607567185
transform 1 0 155572 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1666
timestamp 1607567185
transform 1 0 154376 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1607567185
transform 1 0 155480 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1654
timestamp 1607567185
transform 1 0 153272 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1642
timestamp 1607567185
transform 1 0 152168 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1630
timestamp 1607567185
transform 1 0 151064 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1618
timestamp 1607567185
transform 1 0 149960 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1616
timestamp 1607567185
transform 1 0 149776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1610
timestamp 1607567185
transform 1 0 149224 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1607567185
transform 1 0 149868 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1598
timestamp 1607567185
transform 1 0 148120 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1586
timestamp 1607567185
transform 1 0 147016 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1574
timestamp 1607567185
transform 1 0 145912 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1562
timestamp 1607567185
transform 1 0 144808 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1557
timestamp 1607567185
transform 1 0 144348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1554
timestamp 1607567185
transform 1 0 144072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1607567185
transform 1 0 144256 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1607567185
transform 1 0 144532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1546
timestamp 1607567185
transform 1 0 143336 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1534
timestamp 1607567185
transform 1 0 142232 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1522
timestamp 1607567185
transform 1 0 141128 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1510
timestamp 1607567185
transform 1 0 140024 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1499
timestamp 1607567185
transform 1 0 139012 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1607567185
transform 1 0 138644 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1607567185
transform 1 0 139748 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1607567185
transform 1 0 138736 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1487
timestamp 1607567185
transform 1 0 137908 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1480
timestamp 1607567185
transform 1 0 137264 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1607567185
transform 1 0 137632 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1468
timestamp 1607567185
transform 1 0 136160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1438
timestamp 1607567185
transform 1 0 133400 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[90\]
timestamp 1607567185
transform 1 0 134504 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _649_
timestamp 1607567185
transform 1 0 133124 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1432
timestamp 1607567185
transform 1 0 132848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1424
timestamp 1607567185
transform 1 0 132112 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1607567185
transform 1 0 133032 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1607567185
transform 1 0 131836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1413
timestamp 1607567185
transform 1 0 131100 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1407
timestamp 1607567185
transform 1 0 130548 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1399
timestamp 1607567185
transform 1 0 129812 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1607567185
transform 1 0 130824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1388
timestamp 1607567185
transform 1 0 128800 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1607567185
transform 1 0 129352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1607567185
transform 1 0 129536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1607567185
transform 1 0 128524 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1377
timestamp 1607567185
transform 1 0 127788 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1369
timestamp 1607567185
transform 1 0 127052 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1607567185
transform 1 0 127420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1607567185
transform 1 0 127512 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1357
timestamp 1607567185
transform 1 0 125948 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1346
timestamp 1607567185
transform 1 0 124936 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1607567185
transform 1 0 124476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1607567185
transform 1 0 125488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1607567185
transform 1 0 124660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1607567185
transform 1 0 125672 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1335
timestamp 1607567185
transform 1 0 123924 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1328
timestamp 1607567185
transform 1 0 123280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1607567185
transform 1 0 123648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1316
timestamp 1607567185
transform 1 0 122176 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1310
timestamp 1607567185
transform 1 0 121624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1607567185
transform 1 0 121808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _628_
timestamp 1607567185
transform 1 0 121900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1607567185
transform 1 0 160816 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1727
timestamp 1607567185
transform 1 0 159988 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1728
timestamp 1607567185
transform 1 0 160080 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[64\]
timestamp 1607567185
transform 1 0 159712 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1607567185
transform 1 0 160724 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  mprj_vdd_pwrgood
timestamp 1607567185
transform 1 0 158976 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[67\]
timestamp 1607567185
transform 1 0 158700 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1607567185
transform 1 0 158240 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1714
timestamp 1607567185
transform 1 0 158792 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1709
timestamp 1607567185
transform 1 0 158332 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1716
timestamp 1607567185
transform 1 0 158976 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1607567185
transform 1 0 157964 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1702
timestamp 1607567185
transform 1 0 157688 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1706
timestamp 1607567185
transform 1 0 158056 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1700
timestamp 1607567185
transform 1 0 157504 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1696
timestamp 1607567185
transform 1 0 157136 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1684
timestamp 1607567185
transform 1 0 156032 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1690
timestamp 1607567185
transform 1 0 156584 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1607567185
transform 1 0 157228 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1607567185
transform 1 0 155756 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1679
timestamp 1607567185
transform 1 0 155572 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1667
timestamp 1607567185
transform 1 0 154468 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1678
timestamp 1607567185
transform 1 0 155480 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1666
timestamp 1607567185
transform 1 0 154376 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1607567185
transform 1 0 155112 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _447_
timestamp 1607567185
transform 1 0 155204 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1607567185
transform 1 0 154100 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1647
timestamp 1607567185
transform 1 0 152628 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1655
timestamp 1607567185
transform 1 0 153364 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1607567185
transform 1 0 153088 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1659
timestamp 1607567185
transform 1 0 153732 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1607567185
transform 1 0 152352 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1607567185
transform 1 0 152260 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1607567185
transform 1 0 152628 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1642
timestamp 1607567185
transform 1 0 152168 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1645
timestamp 1607567185
transform 1 0 152444 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1648
timestamp 1607567185
transform 1 0 152720 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1637
timestamp 1607567185
transform 1 0 151708 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1625
timestamp 1607567185
transform 1 0 150604 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1636
timestamp 1607567185
transform 1 0 151616 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1624
timestamp 1607567185
transform 1 0 150512 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1613
timestamp 1607567185
transform 1 0 149500 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1613
timestamp 1607567185
transform 1 0 149500 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1609
timestamp 1607567185
transform 1 0 149132 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1607567185
transform 1 0 149408 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1607567185
transform 1 0 150236 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1601
timestamp 1607567185
transform 1 0 148396 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1590
timestamp 1607567185
transform 1 0 147384 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1597
timestamp 1607567185
transform 1 0 148028 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1585
timestamp 1607567185
transform 1 0 146924 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1607567185
transform 1 0 147016 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1607567185
transform 1 0 148120 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1607567185
transform 1 0 147108 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1578
timestamp 1607567185
transform 1 0 146280 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1574
timestamp 1607567185
transform 1 0 145912 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1579
timestamp 1607567185
transform 1 0 146372 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1567
timestamp 1607567185
transform 1 0 145268 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1607567185
transform 1 0 146556 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1607567185
transform 1 0 146648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1607567185
transform 1 0 146004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1566
timestamp 1607567185
transform 1 0 145176 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1607567185
transform 1 0 144900 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1607567185
transform 1 0 144992 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1607567185
transform 1 0 143980 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1607567185
transform 1 0 143888 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1607567185
transform 1 0 143704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1549
timestamp 1607567185
transform 1 0 143612 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1551
timestamp 1607567185
transform 1 0 143796 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1556
timestamp 1607567185
transform 1 0 144256 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1550
timestamp 1607567185
transform 1 0 143704 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1555
timestamp 1607567185
transform 1 0 144164 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1538
timestamp 1607567185
transform 1 0 142600 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1537
timestamp 1607567185
transform 1 0 142508 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1526
timestamp 1607567185
transform 1 0 141496 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1517
timestamp 1607567185
transform 1 0 140668 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1525
timestamp 1607567185
transform 1 0 141404 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1520
timestamp 1607567185
transform 1 0 140944 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1513
timestamp 1607567185
transform 1 0 140300 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1607567185
transform 1 0 141404 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1607567185
transform 1 0 140852 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1607567185
transform 1 0 141128 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1607567185
transform 1 0 140392 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1506
timestamp 1607567185
transform 1 0 139656 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1495
timestamp 1607567185
transform 1 0 138644 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1501
timestamp 1607567185
transform 1 0 139196 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1497
timestamp 1607567185
transform 1 0 138828 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1607567185
transform 1 0 138920 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1607567185
transform 1 0 139380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1607567185
transform 1 0 138368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1484
timestamp 1607567185
transform 1 0 137632 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1480
timestamp 1607567185
transform 1 0 137264 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1489
timestamp 1607567185
transform 1 0 138092 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1484
timestamp 1607567185
transform 1 0 137632 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1472
timestamp 1607567185
transform 1 0 136528 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1607567185
transform 1 0 138000 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1607567185
transform 1 0 137356 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1468
timestamp 1607567185
transform 1 0 136160 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1607567185
transform 1 0 135884 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _657_
timestamp 1607567185
transform 1 0 136252 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1607567185
transform 1 0 135792 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1607567185
transform 1 0 134780 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _653_
timestamp 1607567185
transform 1 0 135240 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1607567185
transform 1 0 135148 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1453
timestamp 1607567185
transform 1 0 134780 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1461
timestamp 1607567185
transform 1 0 135516 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1456
timestamp 1607567185
transform 1 0 135056 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1445
timestamp 1607567185
transform 1 0 134044 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1441
timestamp 1607567185
transform 1 0 133676 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1607567185
transform 1 0 133216 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _650_
timestamp 1607567185
transform 1 0 133768 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1607567185
transform 1 0 133400 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1434
timestamp 1607567185
transform 1 0 133032 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1430
timestamp 1607567185
transform 1 0 132664 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1418
timestamp 1607567185
transform 1 0 131560 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1430
timestamp 1607567185
transform 1 0 132664 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1422
timestamp 1607567185
transform 1 0 131928 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1607567185
transform 1 0 132296 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1607567185
transform 1 0 132756 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1607567185
transform 1 0 132388 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1407
timestamp 1607567185
transform 1 0 130548 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1401
timestamp 1607567185
transform 1 0 129996 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1410
timestamp 1607567185
transform 1 0 130824 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1399
timestamp 1607567185
transform 1 0 129812 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1607567185
transform 1 0 130180 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1607567185
transform 1 0 130272 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1607567185
transform 1 0 130548 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1607567185
transform 1 0 131284 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1393
timestamp 1607567185
transform 1 0 129260 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1382
timestamp 1607567185
transform 1 0 128248 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1387
timestamp 1607567185
transform 1 0 128708 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1607567185
transform 1 0 129444 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1607567185
transform 1 0 128432 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1607567185
transform 1 0 129536 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1607567185
transform 1 0 128984 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1607567185
transform 1 0 127972 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1377
timestamp 1607567185
transform 1 0 127788 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1369
timestamp 1607567185
transform 1 0 127052 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1376
timestamp 1607567185
transform 1 0 127696 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1365
timestamp 1607567185
transform 1 0 126684 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1360
timestamp 1607567185
transform 1 0 126224 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1607567185
transform 1 0 126592 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1607567185
transform 1 0 126592 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1607567185
transform 1 0 126776 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1607567185
transform 1 0 127420 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1348
timestamp 1607567185
transform 1 0 125120 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1607567185
transform 1 0 125764 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1607567185
transform 1 0 125580 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1352
timestamp 1607567185
transform 1 0 125488 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1358
timestamp 1607567185
transform 1 0 126040 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1607567185
transform 1 0 124844 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1607567185
transform 1 0 124660 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1607567185
transform 1 0 124568 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1607567185
transform 1 0 124936 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1341
timestamp 1607567185
transform 1 0 124476 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1348
timestamp 1607567185
transform 1 0 125120 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1333
timestamp 1607567185
transform 1 0 123740 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1322
timestamp 1607567185
transform 1 0 122728 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1337
timestamp 1607567185
transform 1 0 124108 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1325
timestamp 1607567185
transform 1 0 123004 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1607567185
transform 1 0 123740 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1607567185
transform 1 0 122728 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1607567185
transform 1 0 123464 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1607567185
transform 1 0 123832 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1316
timestamp 1607567185
transform 1 0 122176 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1308
timestamp 1607567185
transform 1 0 121440 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1310
timestamp 1607567185
transform 1 0 121624 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1303
timestamp 1607567185
transform 1 0 120980 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _636_
timestamp 1607567185
transform 1 0 122452 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _625_
timestamp 1607567185
transform 1 0 121164 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1607567185
transform 1 0 121348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _647_
timestamp 1607567185
transform 1 0 119968 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[245\]
timestamp 1607567185
transform 1 0 119232 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[43\]
timestamp 1607567185
transform 1 0 120244 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1291
timestamp 1607567185
transform 1 0 119876 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1295
timestamp 1607567185
transform 1 0 120244 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1287
timestamp 1607567185
transform 1 0 119508 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607567185
transform 1 0 118956 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1279
timestamp 1607567185
transform 1 0 118772 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1266
timestamp 1607567185
transform 1 0 117576 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1278
timestamp 1607567185
transform 1 0 118680 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1282
timestamp 1607567185
transform 1 0 119048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[33\]
timestamp 1607567185
transform 1 0 117116 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[38\]
timestamp 1607567185
transform 1 0 115920 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607567185
transform 1 0 116196 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1252
timestamp 1607567185
transform 1 0 116288 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1260
timestamp 1607567185
transform 1 0 117024 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1247
timestamp 1607567185
transform 1 0 115828 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[239\]
timestamp 1607567185
transform 1 0 114816 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1228
timestamp 1607567185
transform 1 0 114080 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1239
timestamp 1607567185
transform 1 0 115092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1239
timestamp 1607567185
transform 1 0 115092 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[226\]
timestamp 1607567185
transform 1 0 112332 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[29\]
timestamp 1607567185
transform 1 0 112424 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[31\]
timestamp 1607567185
transform 1 0 113436 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607567185
transform 1 0 113344 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1212
timestamp 1607567185
transform 1 0 112608 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[233\]
timestamp 1607567185
transform 1 0 111412 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607567185
transform 1 0 110584 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1189
timestamp 1607567185
transform 1 0 110492 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1191
timestamp 1607567185
transform 1 0 110676 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1202
timestamp 1607567185
transform 1 0 111688 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1195
timestamp 1607567185
transform 1 0 111044 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1207
timestamp 1607567185
transform 1 0 112148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[127\]
timestamp 1607567185
transform 1 0 110216 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1177
timestamp 1607567185
transform 1 0 109388 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1181
timestamp 1607567185
transform 1 0 109756 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1185
timestamp 1607567185
transform 1 0 110124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[122\]
timestamp 1607567185
transform 1 0 107824 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[30\]
timestamp 1607567185
transform 1 0 107732 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607567185
transform 1 0 107732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1151
timestamp 1607567185
transform 1 0 106996 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1169
timestamp 1607567185
transform 1 0 108652 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[222\]
timestamp 1607567185
transform 1 0 106352 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[232\]
timestamp 1607567185
transform 1 0 106720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1139
timestamp 1607567185
transform 1 0 105892 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1607567185
transform 1 0 106628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1136
timestamp 1607567185
transform 1 0 105616 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1147
timestamp 1607567185
transform 1 0 106628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[107\]
timestamp 1607567185
transform 1 0 105064 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[21\]
timestamp 1607567185
transform 1 0 103960 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607567185
transform 1 0 104972 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1120
timestamp 1607567185
transform 1 0 104144 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1128
timestamp 1607567185
transform 1 0 104880 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[223\]
timestamp 1607567185
transform 1 0 102948 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[23\]
timestamp 1607567185
transform 1 0 102488 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607567185
transform 1 0 102120 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1099
timestamp 1607567185
transform 1 0 102212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1097
timestamp 1607567185
transform 1 0 102028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1099
timestamp 1607567185
transform 1 0 102212 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1110
timestamp 1607567185
transform 1 0 103224 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1087
timestamp 1607567185
transform 1 0 101108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1089
timestamp 1607567185
transform 1 0 101292 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[229\]
timestamp 1607567185
transform 1 0 98348 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[16\]
timestamp 1607567185
transform 1 0 99636 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[27\]
timestamp 1607567185
transform 1 0 99452 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607567185
transform 1 0 99360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1060
timestamp 1607567185
transform 1 0 98624 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1058
timestamp 1607567185
transform 1 0 98440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1070
timestamp 1607567185
transform 1 0 99544 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[204\]
timestamp 1607567185
transform 1 0 98164 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[86\]
timestamp 1607567185
transform 1 0 96600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1047
timestamp 1607567185
transform 1 0 97428 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1055
timestamp 1607567185
transform 1 0 98164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1047
timestamp 1607567185
transform 1 0 97428 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[25\]
timestamp 1607567185
transform 1 0 95772 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607567185
transform 1 0 96508 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1020
timestamp 1607567185
transform 1 0 94944 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1032
timestamp 1607567185
transform 1 0 96048 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1036
timestamp 1607567185
transform 1 0 96416 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[82\]
timestamp 1607567185
transform 1 0 93840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[14\]
timestamp 1607567185
transform 1 0 93288 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607567185
transform 1 0 93748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1001
timestamp 1607567185
transform 1 0 93196 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1017
timestamp 1607567185
transform 1 0 94668 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_989
timestamp 1607567185
transform 1 0 92092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_986
timestamp 1607567185
transform 1 0 91816 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_998
timestamp 1607567185
transform 1 0 92920 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[89\]
timestamp 1607567185
transform 1 0 90988 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[19\]
timestamp 1607567185
transform 1 0 90436 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607567185
transform 1 0 90896 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_968
timestamp 1607567185
transform 1 0 90160 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_968
timestamp 1607567185
transform 1 0 90160 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[92\]
timestamp 1607567185
transform 1 0 88228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[22\]
timestamp 1607567185
transform 1 0 88504 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607567185
transform 1 0 88136 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_956
timestamp 1607567185
transform 1 0 89056 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_946
timestamp 1607567185
transform 1 0 88136 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[224\]
timestamp 1607567185
transform 1 0 87124 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_926
timestamp 1607567185
transform 1 0 86296 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_934
timestamp 1607567185
transform 1 0 87032 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_938
timestamp 1607567185
transform 1 0 87400 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_934
timestamp 1607567185
transform 1 0 87032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[66\]
timestamp 1607567185
transform 1 0 85468 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[8\]
timestamp 1607567185
transform 1 0 85376 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607567185
transform 1 0 85284 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_909
timestamp 1607567185
transform 1 0 84732 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_907
timestamp 1607567185
transform 1 0 84548 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[210\]
timestamp 1607567185
transform 1 0 84272 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[380\]
timestamp 1607567185
transform 1 0 82892 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[60\]
timestamp 1607567185
transform 1 0 83904 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_889
timestamp 1607567185
transform 1 0 82892 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_897
timestamp 1607567185
transform 1 0 83628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_892
timestamp 1607567185
transform 1 0 83168 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[383\]
timestamp 1607567185
transform 1 0 82616 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[56\]
timestamp 1607567185
transform 1 0 81328 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607567185
transform 1 0 82524 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_870
timestamp 1607567185
transform 1 0 81144 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_882
timestamp 1607567185
transform 1 0 82248 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_881
timestamp 1607567185
transform 1 0 82156 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[234\]
timestamp 1607567185
transform 1 0 119416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[32\]
timestamp 1607567185
transform 1 0 120428 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1289
timestamp 1607567185
transform 1 0 119692 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[235\]
timestamp 1607567185
transform 1 0 117944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607567185
transform 1 0 118956 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1273
timestamp 1607567185
transform 1 0 118220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1282
timestamp 1607567185
transform 1 0 119048 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _645_
timestamp 1607567185
transform 1 0 116932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1251
timestamp 1607567185
transform 1 0 116196 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1262
timestamp 1607567185
transform 1 0 117208 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[37\]
timestamp 1607567185
transform 1 0 114540 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1232
timestamp 1607567185
transform 1 0 114448 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _648_
timestamp 1607567185
transform 1 0 113436 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607567185
transform 1 0 113344 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1208
timestamp 1607567185
transform 1 0 112240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1224
timestamp 1607567185
transform 1 0 113712 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[231\]
timestamp 1607567185
transform 1 0 111964 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1191
timestamp 1607567185
transform 1 0 110676 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1203
timestamp 1607567185
transform 1 0 111780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[236\]
timestamp 1607567185
transform 1 0 109388 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[437\]
timestamp 1607567185
transform 1 0 110400 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1180
timestamp 1607567185
transform 1 0 109664 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[114\]
timestamp 1607567185
transform 1 0 107824 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607567185
transform 1 0 107732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1151
timestamp 1607567185
transform 1 0 106996 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1169
timestamp 1607567185
transform 1 0 108652 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[436\]
timestamp 1607567185
transform 1 0 106720 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1140
timestamp 1607567185
transform 1 0 105984 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[26\]
timestamp 1607567185
transform 1 0 104328 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1114
timestamp 1607567185
transform 1 0 103592 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[225\]
timestamp 1607567185
transform 1 0 102212 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[228\]
timestamp 1607567185
transform 1 0 103316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607567185
transform 1 0 102120 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1102
timestamp 1607567185
transform 1 0 102488 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1110
timestamp 1607567185
transform 1 0 103224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[98\]
timestamp 1607567185
transform 1 0 100556 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1090
timestamp 1607567185
transform 1 0 101384 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[91\]
timestamp 1607567185
transform 1 0 98992 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1062
timestamp 1607567185
transform 1 0 98808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1073
timestamp 1607567185
transform 1 0 99820 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[87\]
timestamp 1607567185
transform 1 0 96876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1038
timestamp 1607567185
transform 1 0 96600 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1050
timestamp 1607567185
transform 1 0 97704 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[220\]
timestamp 1607567185
transform 1 0 94944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607567185
transform 1 0 96508 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1023
timestamp 1607567185
transform 1 0 95220 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1035
timestamp 1607567185
transform 1 0 96324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[216\]
timestamp 1607567185
transform 1 0 93932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1001
timestamp 1607567185
transform 1 0 93196 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1012
timestamp 1607567185
transform 1 0 94208 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[80\]
timestamp 1607567185
transform 1 0 92368 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[221\]
timestamp 1607567185
transform 1 0 90988 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607567185
transform 1 0 90896 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_963
timestamp 1607567185
transform 1 0 89700 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_975
timestamp 1607567185
transform 1 0 90804 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_980
timestamp 1607567185
transform 1 0 91264 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[73\]
timestamp 1607567185
transform 1 0 88872 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_946
timestamp 1607567185
transform 1 0 88136 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[71\]
timestamp 1607567185
transform 1 0 87308 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_931
timestamp 1607567185
transform 1 0 86756 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[396\]
timestamp 1607567185
transform 1 0 85376 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607567185
transform 1 0 85284 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_912
timestamp 1607567185
transform 1 0 85008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_919
timestamp 1607567185
transform 1 0 85652 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[64\]
timestamp 1607567185
transform 1 0 83444 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_894
timestamp 1607567185
transform 1 0 83352 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_904
timestamp 1607567185
transform 1 0 84272 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[386\]
timestamp 1607567185
transform 1 0 81972 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_871
timestamp 1607567185
transform 1 0 81236 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_882
timestamp 1607567185
transform 1 0 82248 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _629_
timestamp 1607567185
transform 1 0 119232 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _646_
timestamp 1607567185
transform 1 0 120244 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1287
timestamp 1607567185
transform 1 0 119508 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1298
timestamp 1607567185
transform 1 0 120520 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _654_
timestamp 1607567185
transform 1 0 118036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1274
timestamp 1607567185
transform 1 0 118312 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1282
timestamp 1607567185
transform 1 0 119048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _643_
timestamp 1607567185
transform 1 0 117024 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1607567185
transform 1 0 116196 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1252
timestamp 1607567185
transform 1 0 116288 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1263
timestamp 1607567185
transform 1 0 117300 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[299\]
timestamp 1607567185
transform 1 0 115184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1227
timestamp 1607567185
transform 1 0 113988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1239
timestamp 1607567185
transform 1 0 115092 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1243
timestamp 1607567185
transform 1 0 115460 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _641_
timestamp 1607567185
transform 1 0 113712 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _644_
timestamp 1607567185
transform 1 0 112700 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1216
timestamp 1607567185
transform 1 0 112976 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _616_
timestamp 1607567185
transform 1 0 110676 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[438\]
timestamp 1607567185
transform 1 0 111688 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1607567185
transform 1 0 110584 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1194
timestamp 1607567185
transform 1 0 110952 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1205
timestamp 1607567185
transform 1 0 111964 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1174
timestamp 1607567185
transform 1 0 109112 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1186
timestamp 1607567185
transform 1 0 110216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[115\]
timestamp 1607567185
transform 1 0 108284 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1157
timestamp 1607567185
transform 1 0 107548 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[113\]
timestamp 1607567185
transform 1 0 106720 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1140
timestamp 1607567185
transform 1 0 105984 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[109\]
timestamp 1607567185
transform 1 0 105156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1607567185
transform 1 0 104972 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1123
timestamp 1607567185
transform 1 0 104420 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1130
timestamp 1607567185
transform 1 0 105064 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[432\]
timestamp 1607567185
transform 1 0 102028 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[434\]
timestamp 1607567185
transform 1 0 103040 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1100
timestamp 1607567185
transform 1 0 102304 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1111
timestamp 1607567185
transform 1 0 103316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[431\]
timestamp 1607567185
transform 1 0 101016 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1078
timestamp 1607567185
transform 1 0 100280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1089
timestamp 1607567185
transform 1 0 101292 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[95\]
timestamp 1607567185
transform 1 0 99452 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1607567185
transform 1 0 99360 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1057
timestamp 1607567185
transform 1 0 98348 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1065
timestamp 1607567185
transform 1 0 99084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[105\]
timestamp 1607567185
transform 1 0 97520 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1039
timestamp 1607567185
transform 1 0 96692 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1047
timestamp 1607567185
transform 1 0 97428 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[227\]
timestamp 1607567185
transform 1 0 95404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[420\]
timestamp 1607567185
transform 1 0 96416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1028
timestamp 1607567185
transform 1 0 95680 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[96\]
timestamp 1607567185
transform 1 0 93840 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1607567185
transform 1 0 93748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1003
timestamp 1607567185
transform 1 0 93380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1017
timestamp 1607567185
transform 1 0 94668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[81\]
timestamp 1607567185
transform 1 0 91448 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_991
timestamp 1607567185
transform 1 0 92276 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_964
timestamp 1607567185
transform 1 0 89792 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_976
timestamp 1607567185
transform 1 0 90896 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[74\]
timestamp 1607567185
transform 1 0 88964 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1607567185
transform 1 0 88136 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_945
timestamp 1607567185
transform 1 0 88044 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_947
timestamp 1607567185
transform 1 0 88228 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_929
timestamp 1607567185
transform 1 0 86572 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_941
timestamp 1607567185
transform 1 0 87676 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[69\]
timestamp 1607567185
transform 1 0 85744 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_912
timestamp 1607567185
transform 1 0 85008 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[405\]
timestamp 1607567185
transform 1 0 83168 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[65\]
timestamp 1607567185
transform 1 0 84180 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_895
timestamp 1607567185
transform 1 0 83444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1607567185
transform 1 0 82524 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_869
timestamp 1607567185
transform 1 0 81052 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_881
timestamp 1607567185
transform 1 0 82156 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_886
timestamp 1607567185
transform 1 0 82616 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _622_
timestamp 1607567185
transform 1 0 119508 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1607567185
transform 1 0 120520 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1286
timestamp 1607567185
transform 1 0 119416 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1290
timestamp 1607567185
transform 1 0 119784 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1301
timestamp 1607567185
transform 1 0 120796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1607567185
transform 1 0 117668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1607567185
transform 1 0 118956 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1264
timestamp 1607567185
transform 1 0 117392 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1270
timestamp 1607567185
transform 1 0 117944 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1278
timestamp 1607567185
transform 1 0 118680 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1282
timestamp 1607567185
transform 1 0 119048 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _635_
timestamp 1607567185
transform 1 0 116380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1250
timestamp 1607567185
transform 1 0 116104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1256
timestamp 1607567185
transform 1 0 116656 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _624_
timestamp 1607567185
transform 1 0 115092 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1238
timestamp 1607567185
transform 1 0 115000 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1242
timestamp 1607567185
transform 1 0 115368 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1607567185
transform 1 0 113436 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1607567185
transform 1 0 113344 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1607567185
transform 1 0 113712 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1208
timestamp 1607567185
transform 1 0 112240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1226
timestamp 1607567185
transform 1 0 113896 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _611_
timestamp 1607567185
transform 1 0 110952 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _617_
timestamp 1607567185
transform 1 0 111964 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1197
timestamp 1607567185
transform 1 0 111228 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[117\]
timestamp 1607567185
transform 1 0 109388 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1186
timestamp 1607567185
transform 1 0 110216 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[116\]
timestamp 1607567185
transform 1 0 107824 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1607567185
transform 1 0 107732 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1158
timestamp 1607567185
transform 1 0 107640 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1169
timestamp 1607567185
transform 1 0 108652 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[122\]
timestamp 1607567185
transform 1 0 105708 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1136
timestamp 1607567185
transform 1 0 105616 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1146
timestamp 1607567185
transform 1 0 106536 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _603_
timestamp 1607567185
transform 1 0 104604 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1123
timestamp 1607567185
transform 1 0 104420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1128
timestamp 1607567185
transform 1 0 104880 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[106\]
timestamp 1607567185
transform 1 0 102488 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1607567185
transform 1 0 102120 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1095
timestamp 1607567185
transform 1 0 101844 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1099
timestamp 1607567185
transform 1 0 102212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1111
timestamp 1607567185
transform 1 0 103316 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1083
timestamp 1607567185
transform 1 0 100740 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[108\]
timestamp 1607567185
transform 1 0 99912 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1064
timestamp 1607567185
transform 1 0 98992 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1072
timestamp 1607567185
transform 1 0 99728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[426\]
timestamp 1607567185
transform 1 0 96600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[104\]
timestamp 1607567185
transform 1 0 98164 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1041
timestamp 1607567185
transform 1 0 96876 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1053
timestamp 1607567185
transform 1 0 97980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1607567185
transform 1 0 96508 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1024
timestamp 1607567185
transform 1 0 95312 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1036
timestamp 1607567185
transform 1 0 96416 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[94\]
timestamp 1607567185
transform 1 0 94484 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1007
timestamp 1607567185
transform 1 0 93748 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[100\]
timestamp 1607567185
transform 1 0 92920 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_986
timestamp 1607567185
transform 1 0 91816 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[402\]
timestamp 1607567185
transform 1 0 89700 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[88\]
timestamp 1607567185
transform 1 0 90988 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1607567185
transform 1 0 90896 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_966
timestamp 1607567185
transform 1 0 89976 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_974
timestamp 1607567185
transform 1 0 90712 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[77\]
timestamp 1607567185
transform 1 0 88136 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_955
timestamp 1607567185
transform 1 0 88964 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[400\]
timestamp 1607567185
transform 1 0 87124 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_925
timestamp 1607567185
transform 1 0 86204 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_933
timestamp 1607567185
transform 1 0 86940 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_938
timestamp 1607567185
transform 1 0 87400 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[67\]
timestamp 1607567185
transform 1 0 85376 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1607567185
transform 1 0 85284 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_914
timestamp 1607567185
transform 1 0 85192 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[62\]
timestamp 1607567185
transform 1 0 83260 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_902
timestamp 1607567185
transform 1 0 84088 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[399\]
timestamp 1607567185
transform 1 0 81328 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_875
timestamp 1607567185
transform 1 0 81604 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_887
timestamp 1607567185
transform 1 0 82708 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1607567185
transform 1 0 119140 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1607567185
transform 1 0 120244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1607567185
transform 1 0 120060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1286
timestamp 1607567185
transform 1 0 119416 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1292
timestamp 1607567185
transform 1 0 119968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1298
timestamp 1607567185
transform 1 0 120520 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1607567185
transform 1 0 118128 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1264
timestamp 1607567185
transform 1 0 117392 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1275
timestamp 1607567185
transform 1 0 118404 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _620_
timestamp 1607567185
transform 1 0 117116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1607567185
transform 1 0 116196 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1250
timestamp 1607567185
transform 1 0 116104 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1252
timestamp 1607567185
transform 1 0 116288 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1260
timestamp 1607567185
transform 1 0 117024 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _613_
timestamp 1607567185
transform 1 0 114080 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _621_
timestamp 1607567185
transform 1 0 115092 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1227
timestamp 1607567185
transform 1 0 113988 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1231
timestamp 1607567185
transform 1 0 114356 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1242
timestamp 1607567185
transform 1 0 115368 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _612_
timestamp 1607567185
transform 1 0 112240 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1211
timestamp 1607567185
transform 1 0 112516 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1223
timestamp 1607567185
transform 1 0 113620 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[127\]
timestamp 1607567185
transform 1 0 110676 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1607567185
transform 1 0 110584 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1189
timestamp 1607567185
transform 1 0 110492 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1200
timestamp 1607567185
transform 1 0 111504 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[118\]
timestamp 1607567185
transform 1 0 108928 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1181
timestamp 1607567185
transform 1 0 109756 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1154
timestamp 1607567185
transform 1 0 107272 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1166
timestamp 1607567185
transform 1 0 108376 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[121\]
timestamp 1607567185
transform 1 0 106444 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1134
timestamp 1607567185
transform 1 0 105432 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1142
timestamp 1607567185
transform 1 0 106168 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _606_
timestamp 1607567185
transform 1 0 105156 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1607567185
transform 1 0 104972 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1124
timestamp 1607567185
transform 1 0 104512 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1128
timestamp 1607567185
transform 1 0 104880 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1130
timestamp 1607567185
transform 1 0 105064 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[125\]
timestamp 1607567185
transform 1 0 102580 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1095
timestamp 1607567185
transform 1 0 101844 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1112
timestamp 1607567185
transform 1 0 103408 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[107\]
timestamp 1607567185
transform 1 0 101016 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1078
timestamp 1607567185
transform 1 0 100280 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[99\]
timestamp 1607567185
transform 1 0 99452 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1607567185
transform 1 0 99360 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1064
timestamp 1607567185
transform 1 0 98992 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[101\]
timestamp 1607567185
transform 1 0 97060 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1052
timestamp 1607567185
transform 1 0 97888 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[428\]
timestamp 1607567185
transform 1 0 96048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1024
timestamp 1607567185
transform 1 0 95312 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1035
timestamp 1607567185
transform 1 0 96324 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[102\]
timestamp 1607567185
transform 1 0 94484 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1607567185
transform 1 0 93748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1005
timestamp 1607567185
transform 1 0 93564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1008
timestamp 1607567185
transform 1 0 93840 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1014
timestamp 1607567185
transform 1 0 94392 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[413\]
timestamp 1607567185
transform 1 0 92552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_986
timestamp 1607567185
transform 1 0 91816 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_997
timestamp 1607567185
transform 1 0 92828 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[84\]
timestamp 1607567185
transform 1 0 90988 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_969
timestamp 1607567185
transform 1 0 90252 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[412\]
timestamp 1607567185
transform 1 0 88228 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[76\]
timestamp 1607567185
transform 1 0 89424 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1607567185
transform 1 0 88136 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_945
timestamp 1607567185
transform 1 0 88044 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_950
timestamp 1607567185
transform 1 0 88504 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_958
timestamp 1607567185
transform 1 0 89240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_933
timestamp 1607567185
transform 1 0 86940 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[75\]
timestamp 1607567185
transform 1 0 86112 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_910
timestamp 1607567185
transform 1 0 84824 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_922
timestamp 1607567185
transform 1 0 85928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[408\]
timestamp 1607567185
transform 1 0 82984 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[61\]
timestamp 1607567185
transform 1 0 83996 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_893
timestamp 1607567185
transform 1 0 83260 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1607567185
transform 1 0 82524 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_869
timestamp 1607567185
transform 1 0 81052 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_881
timestamp 1607567185
transform 1 0 82156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_886
timestamp 1607567185
transform 1 0 82616 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1607567185
transform 1 0 120888 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1607567185
transform 1 0 120152 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _623_
timestamp 1607567185
transform 1 0 119140 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1607567185
transform 1 0 119968 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1286
timestamp 1607567185
transform 1 0 119416 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1298
timestamp 1607567185
transform 1 0 120520 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1285
timestamp 1607567185
transform 1 0 119324 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1291
timestamp 1607567185
transform 1 0 119876 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1297
timestamp 1607567185
transform 1 0 120428 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1607567185
transform 1 0 119048 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _619_
timestamp 1607567185
transform 1 0 118128 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1607567185
transform 1 0 118036 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1607567185
transform 1 0 118956 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1267
timestamp 1607567185
transform 1 0 117668 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1275
timestamp 1607567185
transform 1 0 118404 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1266
timestamp 1607567185
transform 1 0 117576 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1278
timestamp 1607567185
transform 1 0 118680 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1607567185
transform 1 0 117300 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _615_
timestamp 1607567185
transform 1 0 116104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1607567185
transform 1 0 116288 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1607567185
transform 1 0 117116 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1255
timestamp 1607567185
transform 1 0 116564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1253
timestamp 1607567185
transform 1 0 116380 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1607567185
transform 1 0 115276 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1607567185
transform 1 0 115092 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _627_
timestamp 1607567185
transform 1 0 114172 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1607567185
transform 1 0 115184 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1232
timestamp 1607567185
transform 1 0 114448 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1244
timestamp 1607567185
transform 1 0 115552 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1236
timestamp 1607567185
transform 1 0 114816 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1242
timestamp 1607567185
transform 1 0 115368 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _610_
timestamp 1607567185
transform 1 0 112424 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _618_
timestamp 1607567185
transform 1 0 113436 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1607567185
transform 1 0 112332 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1607567185
transform 1 0 113344 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1213
timestamp 1607567185
transform 1 0 112700 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1225
timestamp 1607567185
transform 1 0 113804 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1208
timestamp 1607567185
transform 1 0 112240 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1224
timestamp 1607567185
transform 1 0 113712 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _605_
timestamp 1607567185
transform 1 0 110584 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _607_
timestamp 1607567185
transform 1 0 111964 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1193
timestamp 1607567185
transform 1 0 110860 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1205
timestamp 1607567185
transform 1 0 111964 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1190
timestamp 1607567185
transform 1 0 110584 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1202
timestamp 1607567185
transform 1 0 111688 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _601_
timestamp 1607567185
transform 1 0 109572 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[119\]
timestamp 1607567185
transform 1 0 109756 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1607567185
transform 1 0 109480 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1170
timestamp 1607567185
transform 1 0 108744 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1182
timestamp 1607567185
transform 1 0 109848 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _604_
timestamp 1607567185
transform 1 0 108468 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[124\]
timestamp 1607567185
transform 1 0 107824 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1607567185
transform 1 0 107732 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1157
timestamp 1607567185
transform 1 0 107548 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1165
timestamp 1607567185
transform 1 0 108284 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1151
timestamp 1607567185
transform 1 0 106996 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1169
timestamp 1607567185
transform 1 0 108652 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _609_
timestamp 1607567185
transform 1 0 105616 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[120\]
timestamp 1607567185
transform 1 0 106168 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[123\]
timestamp 1607567185
transform 1 0 106720 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1607567185
transform 1 0 106628 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1139
timestamp 1607567185
transform 1 0 105892 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1134
timestamp 1607567185
transform 1 0 105432 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _614_
timestamp 1607567185
transform 1 0 104604 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[126\]
timestamp 1607567185
transform 1 0 104604 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1607567185
transform 1 0 103776 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1115
timestamp 1607567185
transform 1 0 103684 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1117
timestamp 1607567185
transform 1 0 103868 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1128
timestamp 1607567185
transform 1 0 104880 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1120
timestamp 1607567185
transform 1 0 104144 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1124
timestamp 1607567185
transform 1 0 104512 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[111\]
timestamp 1607567185
transform 1 0 102212 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1607567185
transform 1 0 102120 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1099
timestamp 1607567185
transform 1 0 102212 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1111
timestamp 1607567185
transform 1 0 103316 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1108
timestamp 1607567185
transform 1 0 103040 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _600_
timestamp 1607567185
transform 1 0 101108 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _608_
timestamp 1607567185
transform 1 0 100096 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[112\]
timestamp 1607567185
transform 1 0 101384 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1607567185
transform 1 0 100924 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1080
timestamp 1607567185
transform 1 0 100464 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1084
timestamp 1607567185
transform 1 0 100832 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1086
timestamp 1607567185
transform 1 0 101016 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1079
timestamp 1607567185
transform 1 0 100372 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1090
timestamp 1607567185
transform 1 0 101384 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _599_
timestamp 1607567185
transform 1 0 99084 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[110\]
timestamp 1607567185
transform 1 0 98440 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1063
timestamp 1607567185
transform 1 0 98900 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_1068
timestamp 1607567185
transform 1 0 99360 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1067
timestamp 1607567185
transform 1 0 99268 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1075
timestamp 1607567185
transform 1 0 100004 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _602_
timestamp 1607567185
transform 1 0 96876 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[97\]
timestamp 1607567185
transform 1 0 96600 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1607567185
transform 1 0 98072 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1044
timestamp 1607567185
transform 1 0 97152 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1052
timestamp 1607567185
transform 1 0 97888 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1055
timestamp 1607567185
transform 1 0 98164 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1047
timestamp 1607567185
transform 1 0 97428 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1055
timestamp 1607567185
transform 1 0 98164 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[90\]
timestamp 1607567185
transform 1 0 95312 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1607567185
transform 1 0 95220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1607567185
transform 1 0 96508 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1021
timestamp 1607567185
transform 1 0 95036 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1033
timestamp 1607567185
transform 1 0 96140 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1027
timestamp 1607567185
transform 1 0 95588 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1035
timestamp 1607567185
transform 1 0 96324 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[425\]
timestamp 1607567185
transform 1 0 94024 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[103\]
timestamp 1607567185
transform 1 0 94760 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1002
timestamp 1607567185
transform 1 0 93288 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1013
timestamp 1607567185
transform 1 0 94300 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1003
timestamp 1607567185
transform 1 0 93380 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1015
timestamp 1607567185
transform 1 0 94484 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[83\]
timestamp 1607567185
transform 1 0 92460 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[93\]
timestamp 1607567185
transform 1 0 92552 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1607567185
transform 1 0 92368 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_982
timestamp 1607567185
transform 1 0 91448 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_990
timestamp 1607567185
transform 1 0 92184 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_986
timestamp 1607567185
transform 1 0 91816 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[415\]
timestamp 1607567185
transform 1 0 91172 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[85\]
timestamp 1607567185
transform 1 0 90988 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1607567185
transform 1 0 90896 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_971
timestamp 1607567185
transform 1 0 90436 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_973
timestamp 1607567185
transform 1 0 90620 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[439\]
timestamp 1607567185
transform 1 0 88504 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[78\]
timestamp 1607567185
transform 1 0 88688 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[79\]
timestamp 1607567185
transform 1 0 89608 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1607567185
transform 1 0 89516 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_948
timestamp 1607567185
transform 1 0 88320 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_953
timestamp 1607567185
transform 1 0 88780 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_944
timestamp 1607567185
transform 1 0 87952 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_961
timestamp 1607567185
transform 1 0 89516 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[70\]
timestamp 1607567185
transform 1 0 86756 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[72\]
timestamp 1607567185
transform 1 0 87124 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1607567185
transform 1 0 86664 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_929
timestamp 1607567185
transform 1 0 86572 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_940
timestamp 1607567185
transform 1 0 87584 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_925
timestamp 1607567185
transform 1 0 86204 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_933
timestamp 1607567185
transform 1 0 86940 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[411\]
timestamp 1607567185
transform 1 0 85560 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[68\]
timestamp 1607567185
transform 1 0 85376 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1607567185
transform 1 0 85284 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_909
timestamp 1607567185
transform 1 0 84732 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_917
timestamp 1607567185
transform 1 0 85468 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_921
timestamp 1607567185
transform 1 0 85836 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_910
timestamp 1607567185
transform 1 0 84824 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_914
timestamp 1607567185
transform 1 0 85192 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[440\]
timestamp 1607567185
transform 1 0 82800 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[63\]
timestamp 1607567185
transform 1 0 82892 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[66\]
timestamp 1607567185
transform 1 0 83904 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1607567185
transform 1 0 83812 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_891
timestamp 1607567185
transform 1 0 83076 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_898
timestamp 1607567185
transform 1 0 83720 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[441\]
timestamp 1607567185
transform 1 0 81788 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[59\]
timestamp 1607567185
transform 1 0 81328 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_869
timestamp 1607567185
transform 1 0 81052 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_880
timestamp 1607567185
transform 1 0 82064 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_881
timestamp 1607567185
transform 1 0 82156 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[55\]
timestamp 1607567185
transform 1 0 79764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[15\]
timestamp 1607567185
transform 1 0 79488 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607567185
transform 1 0 79672 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_864
timestamp 1607567185
transform 1 0 80592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[45\]
timestamp 1607567185
transform 1 0 78108 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_834
timestamp 1607567185
transform 1 0 77832 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_846
timestamp 1607567185
transform 1 0 78936 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_846
timestamp 1607567185
transform 1 0 78936 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[208\]
timestamp 1607567185
transform 1 0 77096 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[215\]
timestamp 1607567185
transform 1 0 76084 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[42\]
timestamp 1607567185
transform 1 0 77004 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607567185
transform 1 0 76912 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_818
timestamp 1607567185
transform 1 0 76360 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_818
timestamp 1607567185
transform 1 0 76360 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_829
timestamp 1607567185
transform 1 0 77372 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[40\]
timestamp 1607567185
transform 1 0 74428 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[37\]
timestamp 1607567185
transform 1 0 74152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607567185
transform 1 0 74060 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_794
timestamp 1607567185
transform 1 0 74152 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_806
timestamp 1607567185
transform 1 0 75256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_792
timestamp 1607567185
transform 1 0 73968 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_803
timestamp 1607567185
transform 1 0 74980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_782
timestamp 1607567185
transform 1 0 73048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_780
timestamp 1607567185
transform 1 0 72864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[34\]
timestamp 1607567185
transform 1 0 72036 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[10\]
timestamp 1607567185
transform 1 0 71392 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607567185
transform 1 0 71300 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_755
timestamp 1607567185
transform 1 0 70564 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_763
timestamp 1607567185
transform 1 0 71300 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[30\]
timestamp 1607567185
transform 1 0 70472 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[31\]
timestamp 1607567185
transform 1 0 68908 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[9\]
timestamp 1607567185
transform 1 0 68908 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_7_746
timestamp 1607567185
transform 1 0 69736 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[211\]
timestamp 1607567185
transform 1 0 67896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607567185
transform 1 0 68448 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_718
timestamp 1607567185
transform 1 0 67160 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_729
timestamp 1607567185
transform 1 0 68172 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_724
timestamp 1607567185
transform 1 0 67712 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_733
timestamp 1607567185
transform 1 0 68540 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[214\]
timestamp 1607567185
transform 1 0 66884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[363\]
timestamp 1607567185
transform 1 0 65872 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[26\]
timestamp 1607567185
transform 1 0 66884 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607567185
transform 1 0 65688 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_703
timestamp 1607567185
transform 1 0 65780 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_707
timestamp 1607567185
transform 1 0 66148 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[335\]
timestamp 1607567185
transform 1 0 63572 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[346\]
timestamp 1607567185
transform 1 0 64492 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_682
timestamp 1607567185
transform 1 0 63848 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_694
timestamp 1607567185
transform 1 0 64952 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_681
timestamp 1607567185
transform 1 0 63756 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_692
timestamp 1607567185
transform 1 0 64768 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[332\]
timestamp 1607567185
transform 1 0 62560 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[5\]
timestamp 1607567185
transform 1 0 62928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607567185
transform 1 0 62836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_671
timestamp 1607567185
transform 1 0 62836 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_663
timestamp 1607567185
transform 1 0 62100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[125\]
timestamp 1607567185
transform 1 0 60168 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[200\]
timestamp 1607567185
transform 1 0 61824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_660
timestamp 1607567185
transform 1 0 61824 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_652
timestamp 1607567185
transform 1 0 61088 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[126\]
timestamp 1607567185
transform 1 0 59432 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[199\]
timestamp 1607567185
transform 1 0 59064 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607567185
transform 1 0 60076 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_633
timestamp 1607567185
transform 1 0 59340 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_626
timestamp 1607567185
transform 1 0 58696 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[198\]
timestamp 1607567185
transform 1 0 57040 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[203\]
timestamp 1607567185
transform 1 0 58052 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[1\]
timestamp 1607567185
transform 1 0 57868 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607567185
transform 1 0 57224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_611
timestamp 1607567185
transform 1 0 57316 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_622
timestamp 1607567185
transform 1 0 58328 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_611
timestamp 1607567185
transform 1 0 57316 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_600
timestamp 1607567185
transform 1 0 56304 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_602
timestamp 1607567185
transform 1 0 56488 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[124\]
timestamp 1607567185
transform 1 0 54832 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[0\]
timestamp 1607567185
transform 1 0 54648 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607567185
transform 1 0 54464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_568
timestamp 1607567185
transform 1 0 53360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_581
timestamp 1607567185
transform 1 0 54556 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_574
timestamp 1607567185
transform 1 0 53912 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_582
timestamp 1607567185
transform 1 0 54648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_8  la_buf\[118\]
timestamp 1607567185
transform 1 0 52256 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[120\]
timestamp 1607567185
transform 1 0 51704 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607567185
transform 1 0 51612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_550
timestamp 1607567185
transform 1 0 51704 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[194\]
timestamp 1607567185
transform 1 0 50600 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_538
timestamp 1607567185
transform 1 0 50600 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_541
timestamp 1607567185
transform 1 0 50876 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[115\]
timestamp 1607567185
transform 1 0 48944 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[183\]
timestamp 1607567185
transform 1 0 49220 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607567185
transform 1 0 48852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_519
timestamp 1607567185
transform 1 0 48852 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_526
timestamp 1607567185
transform 1 0 49496 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[177\]
timestamp 1607567185
transform 1 0 47472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_496
timestamp 1607567185
transform 1 0 46736 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_507
timestamp 1607567185
transform 1 0 47748 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_507
timestamp 1607567185
transform 1 0 47748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[103\]
timestamp 1607567185
transform 1 0 46092 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[106\]
timestamp 1607567185
transform 1 0 45080 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607567185
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_474
timestamp 1607567185
transform 1 0 44712 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_480
timestamp 1607567185
transform 1 0 45264 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _567_
timestamp 1607567185
transform 1 0 43332 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  la_buf\[110\]
timestamp 1607567185
transform 1 0 43608 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607567185
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_457
timestamp 1607567185
transform 1 0 43148 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_462
timestamp 1607567185
transform 1 0 43608 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_458
timestamp 1607567185
transform 1 0 43240 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_449
timestamp 1607567185
transform 1 0 42412 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_446
timestamp 1607567185
transform 1 0 42136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[379\]
timestamp 1607567185
transform 1 0 80960 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[217\]
timestamp 1607567185
transform 1 0 79764 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607567185
transform 1 0 79672 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_858
timestamp 1607567185
transform 1 0 80040 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_866
timestamp 1607567185
transform 1 0 80776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[56\]
timestamp 1607567185
transform 1 0 78108 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_834
timestamp 1607567185
transform 1 0 77832 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_846
timestamp 1607567185
transform 1 0 78936 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[41\]
timestamp 1607567185
transform 1 0 75900 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_811
timestamp 1607567185
transform 1 0 75716 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_822
timestamp 1607567185
transform 1 0 76728 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[39\]
timestamp 1607567185
transform 1 0 74152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607567185
transform 1 0 74060 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_803
timestamp 1607567185
transform 1 0 74980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[357\]
timestamp 1607567185
transform 1 0 72680 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_781
timestamp 1607567185
transform 1 0 72956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[354\]
timestamp 1607567185
transform 1 0 71668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_759
timestamp 1607567185
transform 1 0 70932 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_770
timestamp 1607567185
transform 1 0 71944 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  user_to_mprj_in_gates\[33\]
timestamp 1607567185
transform 1 0 70104 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_742
timestamp 1607567185
transform 1 0 69368 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[364\]
timestamp 1607567185
transform 1 0 67436 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[22\]
timestamp 1607567185
transform 1 0 68540 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607567185
transform 1 0 68448 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_724
timestamp 1607567185
transform 1 0 67712 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_709
timestamp 1607567185
transform 1 0 66332 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_685
timestamp 1607567185
transform 1 0 64124 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_697
timestamp 1607567185
transform 1 0 65228 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[12\]
timestamp 1607567185
transform 1 0 63296 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607567185
transform 1 0 62836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_661
timestamp 1607567185
transform 1 0 61916 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_669
timestamp 1607567185
transform 1 0 62652 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_672
timestamp 1607567185
transform 1 0 62928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[331\]
timestamp 1607567185
transform 1 0 61640 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_650
timestamp 1607567185
transform 1 0 60904 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  user_to_mprj_oen_buffers\[1\]
timestamp 1607567185
transform 1 0 59248 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_5_624
timestamp 1607567185
transform 1 0 58512 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[7\]
timestamp 1607567185
transform 1 0 57684 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607567185
transform 1 0 57224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_609
timestamp 1607567185
transform 1 0 57132 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_611
timestamp 1607567185
transform 1 0 57316 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1607567185
transform 1 0 55108 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _590_
timestamp 1607567185
transform 1 0 56120 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_590
timestamp 1607567185
transform 1 0 55384 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_601
timestamp 1607567185
transform 1 0 56396 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1607567185
transform 1 0 54096 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_568
timestamp 1607567185
transform 1 0 53360 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_579
timestamp 1607567185
transform 1 0 54372 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[123\]
timestamp 1607567185
transform 1 0 51704 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607567185
transform 1 0 51612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[197\]
timestamp 1607567185
transform 1 0 50600 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_531
timestamp 1607567185
transform 1 0 49956 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_537
timestamp 1607567185
transform 1 0 50508 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_541
timestamp 1607567185
transform 1 0 50876 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[189\]
timestamp 1607567185
transform 1 0 48576 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_514
timestamp 1607567185
transform 1 0 48392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_519
timestamp 1607567185
transform 1 0 48852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _573_
timestamp 1607567185
transform 1 0 46368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[184\]
timestamp 1607567185
transform 1 0 47380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_495
timestamp 1607567185
transform 1 0 46644 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_506
timestamp 1607567185
transform 1 0 47656 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[169\]
timestamp 1607567185
transform 1 0 44712 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607567185
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_473
timestamp 1607567185
transform 1 0 44620 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_477
timestamp 1607567185
transform 1 0 44988 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_485
timestamp 1607567185
transform 1 0 45724 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_489
timestamp 1607567185
transform 1 0 46092 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_465
timestamp 1607567185
transform 1 0 43884 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[99\]
timestamp 1607567185
transform 1 0 42228 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1607567185
transform 1 0 41860 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[58\]
timestamp 1607567185
transform 1 0 80224 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_852
timestamp 1607567185
transform 1 0 79488 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[49\]
timestamp 1607567185
transform 1 0 78660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_840
timestamp 1607567185
transform 1 0 78384 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[376\]
timestamp 1607567185
transform 1 0 77004 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1607567185
transform 1 0 76912 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_816
timestamp 1607567185
transform 1 0 76176 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_828
timestamp 1607567185
transform 1 0 77280 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[44\]
timestamp 1607567185
transform 1 0 75348 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_803
timestamp 1607567185
transform 1 0 74980 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[367\]
timestamp 1607567185
transform 1 0 73600 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_780
timestamp 1607567185
transform 1 0 72864 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_791
timestamp 1607567185
transform 1 0 73876 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[38\]
timestamp 1607567185
transform 1 0 72036 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1607567185
transform 1 0 71300 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_762
timestamp 1607567185
transform 1 0 71208 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_764
timestamp 1607567185
transform 1 0 71392 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_770
timestamp 1607567185
transform 1 0 71944 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[212\]
timestamp 1607567185
transform 1 0 69828 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[361\]
timestamp 1607567185
transform 1 0 68816 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_739
timestamp 1607567185
transform 1 0 69092 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_750
timestamp 1607567185
transform 1 0 70104 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_725
timestamp 1607567185
transform 1 0 67804 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_733
timestamp 1607567185
transform 1 0 68540 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[26\]
timestamp 1607567185
transform 1 0 65872 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1607567185
transform 1 0 65688 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_701
timestamp 1607567185
transform 1 0 65596 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_703
timestamp 1607567185
transform 1 0 65780 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_713
timestamp 1607567185
transform 1 0 66700 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_689
timestamp 1607567185
transform 1 0 64492 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_665
timestamp 1607567185
transform 1 0 62284 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_677
timestamp 1607567185
transform 1 0 63388 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[205\]
timestamp 1607567185
transform 1 0 60168 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[11\]
timestamp 1607567185
transform 1 0 61456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_645
timestamp 1607567185
transform 1 0 60444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_653
timestamp 1607567185
transform 1 0 61180 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[330\]
timestamp 1607567185
transform 1 0 59064 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1607567185
transform 1 0 60076 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_624
timestamp 1607567185
transform 1 0 58512 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_633
timestamp 1607567185
transform 1 0 59340 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[209\]
timestamp 1607567185
transform 1 0 57132 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_606
timestamp 1607567185
transform 1 0 56856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_612
timestamp 1607567185
transform 1 0 57408 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _593_
timestamp 1607567185
transform 1 0 55476 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_589
timestamp 1607567185
transform 1 0 55292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_594
timestamp 1607567185
transform 1 0 55752 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1607567185
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_566
timestamp 1607567185
transform 1 0 53176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_578
timestamp 1607567185
transform 1 0 54280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_581
timestamp 1607567185
transform 1 0 54556 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _578_
timestamp 1607567185
transform 1 0 51888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _579_
timestamp 1607567185
transform 1 0 52900 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_555
timestamp 1607567185
transform 1 0 52164 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[202\]
timestamp 1607567185
transform 1 0 50876 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_532
timestamp 1607567185
transform 1 0 50048 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_540
timestamp 1607567185
transform 1 0 50784 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_544
timestamp 1607567185
transform 1 0 51152 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1607567185
transform 1 0 48852 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_515
timestamp 1607567185
transform 1 0 48484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_520
timestamp 1607567185
transform 1 0 48944 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_491
timestamp 1607567185
transform 1 0 46276 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_503
timestamp 1607567185
transform 1 0 47380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[95\]
timestamp 1607567185
transform 1 0 44620 0 -1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _565_
timestamp 1607567185
transform 1 0 43332 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1607567185
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_462
timestamp 1607567185
transform 1 0 43608 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_470
timestamp 1607567185
transform 1 0 44344 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _562_
timestamp 1607567185
transform 1 0 41308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_440
timestamp 1607567185
transform 1 0 41584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_452
timestamp 1607567185
transform 1 0 42688 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[57\]
timestamp 1607567185
transform 1 0 79764 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1607567185
transform 1 0 79672 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_864
timestamp 1607567185
transform 1 0 80592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[385\]
timestamp 1607567185
transform 1 0 78660 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_835
timestamp 1607567185
transform 1 0 77924 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_846
timestamp 1607567185
transform 1 0 78936 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[48\]
timestamp 1607567185
transform 1 0 77096 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_818
timestamp 1607567185
transform 1 0 76360 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[377\]
timestamp 1607567185
transform 1 0 74152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[43\]
timestamp 1607567185
transform 1 0 75532 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1607567185
transform 1 0 74060 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_792
timestamp 1607567185
transform 1 0 73968 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_797
timestamp 1607567185
transform 1 0 74428 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_780
timestamp 1607567185
transform 1 0 72864 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[36\]
timestamp 1607567185
transform 1 0 72036 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_763
timestamp 1607567185
transform 1 0 71300 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[30\]
timestamp 1607567185
transform 1 0 70472 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_742
timestamp 1607567185
transform 1 0 69368 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[29\]
timestamp 1607567185
transform 1 0 68540 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1607567185
transform 1 0 68448 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_718
timestamp 1607567185
transform 1 0 67160 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_730
timestamp 1607567185
transform 1 0 68264 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[24\]
timestamp 1607567185
transform 1 0 66332 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_701
timestamp 1607567185
transform 1 0 65596 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[13\]
timestamp 1607567185
transform 1 0 64768 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_681
timestamp 1607567185
transform 1 0 63756 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_689
timestamp 1607567185
transform 1 0 64492 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[10\]
timestamp 1607567185
transform 1 0 62928 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1607567185
transform 1 0 62836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_664
timestamp 1607567185
transform 1 0 62192 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_670
timestamp 1607567185
transform 1 0 62744 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[6\]
timestamp 1607567185
transform 1 0 60260 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_652
timestamp 1607567185
transform 1 0 61088 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_631
timestamp 1607567185
transform 1 0 59156 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _597_
timestamp 1607567185
transform 1 0 57776 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1607567185
transform 1 0 57224 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_607
timestamp 1607567185
transform 1 0 56948 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_611
timestamp 1607567185
transform 1 0 57316 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1607567185
transform 1 0 57684 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_619
timestamp 1607567185
transform 1 0 58052 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_595
timestamp 1607567185
transform 1 0 55844 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _589_
timestamp 1607567185
transform 1 0 53452 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _595_
timestamp 1607567185
transform 1 0 54464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_572
timestamp 1607567185
transform 1 0 53728 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_583
timestamp 1607567185
transform 1 0 54740 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[3\]
timestamp 1607567185
transform 1 0 51888 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1607567185
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_550
timestamp 1607567185
transform 1 0 51704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_561
timestamp 1607567185
transform 1 0 52716 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _594_
timestamp 1607567185
transform 1 0 50600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_530
timestamp 1607567185
transform 1 0 49864 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_541
timestamp 1607567185
transform 1 0 50876 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _576_
timestamp 1607567185
transform 1 0 48484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_512
timestamp 1607567185
transform 1 0 48208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_518
timestamp 1607567185
transform 1 0 48760 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_492
timestamp 1607567185
transform 1 0 46368 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_504
timestamp 1607567185
transform 1 0 47472 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _574_
timestamp 1607567185
transform 1 0 46092 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[180\]
timestamp 1607567185
transform 1 0 44712 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1607567185
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_477
timestamp 1607567185
transform 1 0 44988 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_485
timestamp 1607567185
transform 1 0 45724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _568_
timestamp 1607567185
transform 1 0 43700 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_455
timestamp 1607567185
transform 1 0 42964 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_466
timestamp 1607567185
transform 1 0 43976 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _559_
timestamp 1607567185
transform 1 0 41124 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _561_
timestamp 1607567185
transform 1 0 42688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_438
timestamp 1607567185
transform 1 0 41400 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_450
timestamp 1607567185
transform 1 0 42504 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[54\]
timestamp 1607567185
transform 1 0 80224 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_852
timestamp 1607567185
transform 1 0 79488 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[52\]
timestamp 1607567185
transform 1 0 78660 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_835
timestamp 1607567185
transform 1 0 77924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[46\]
timestamp 1607567185
transform 1 0 77096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1607567185
transform 1 0 76912 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_811
timestamp 1607567185
transform 1 0 75716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_823
timestamp 1607567185
transform 1 0 76820 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_825
timestamp 1607567185
transform 1 0 77004 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[394\]
timestamp 1607567185
transform 1 0 75440 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_800
timestamp 1607567185
transform 1 0 74704 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[37\]
timestamp 1607567185
transform 1 0 73876 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_780
timestamp 1607567185
transform 1 0 72864 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_788
timestamp 1607567185
transform 1 0 73600 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[35\]
timestamp 1607567185
transform 1 0 72036 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1607567185
transform 1 0 71300 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_755
timestamp 1607567185
transform 1 0 70564 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_764
timestamp 1607567185
transform 1 0 71392 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_770
timestamp 1607567185
transform 1 0 71944 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[28\]
timestamp 1607567185
transform 1 0 69736 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_736
timestamp 1607567185
transform 1 0 68816 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_744
timestamp 1607567185
transform 1 0 69552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[25\]
timestamp 1607567185
transform 1 0 67988 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_719
timestamp 1607567185
transform 1 0 67252 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[20\]
timestamp 1607567185
transform 1 0 66424 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1607567185
transform 1 0 65688 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_699
timestamp 1607567185
transform 1 0 65412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_703
timestamp 1607567185
transform 1 0 65780 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_709
timestamp 1607567185
transform 1 0 66332 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_679
timestamp 1607567185
transform 1 0 63572 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_691
timestamp 1607567185
transform 1 0 64676 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[17\]
timestamp 1607567185
transform 1 0 62744 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_667
timestamp 1607567185
transform 1 0 62468 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[8\]
timestamp 1607567185
transform 1 0 60536 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_642
timestamp 1607567185
transform 1 0 60168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_655
timestamp 1607567185
transform 1 0 61364 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1607567185
transform 1 0 60076 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_630
timestamp 1607567185
transform 1 0 59064 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_638
timestamp 1607567185
transform 1 0 59800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[1\]
timestamp 1607567185
transform 1 0 57132 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_608
timestamp 1607567185
transform 1 0 57040 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_618
timestamp 1607567185
transform 1 0 57960 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _598_
timestamp 1607567185
transform 1 0 55660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_585
timestamp 1607567185
transform 1 0 54924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_596
timestamp 1607567185
transform 1 0 55936 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _591_
timestamp 1607567185
transform 1 0 54648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1607567185
transform 1 0 54464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_576
timestamp 1607567185
transform 1 0 54096 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_581
timestamp 1607567185
transform 1 0 54556 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _585_
timestamp 1607567185
transform 1 0 51704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1607567185
transform 1 0 52716 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_553
timestamp 1607567185
transform 1 0 51980 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_564
timestamp 1607567185
transform 1 0 52992 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1607567185
transform 1 0 50324 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_532
timestamp 1607567185
transform 1 0 50048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_538
timestamp 1607567185
transform 1 0 50600 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1607567185
transform 1 0 48852 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_517
timestamp 1607567185
transform 1 0 48668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_520
timestamp 1607567185
transform 1 0 48944 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1607567185
transform 1 0 46644 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1607567185
transform 1 0 47656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_498
timestamp 1607567185
transform 1 0 46920 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_509
timestamp 1607567185
transform 1 0 47932 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _563_
timestamp 1607567185
transform 1 0 44620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _572_
timestamp 1607567185
transform 1 0 45632 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_476
timestamp 1607567185
transform 1 0 44896 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_487
timestamp 1607567185
transform 1 0 45908 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _560_
timestamp 1607567185
transform 1 0 43332 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1607567185
transform 1 0 43240 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_462
timestamp 1607567185
transform 1 0 43608 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_470
timestamp 1607567185
transform 1 0 44344 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _570_
timestamp 1607567185
transform 1 0 42228 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_438
timestamp 1607567185
transform 1 0 41400 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_446
timestamp 1607567185
transform 1 0 42136 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_450
timestamp 1607567185
transform 1 0 42504 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1607567185
transform 1 0 80960 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[442\]
timestamp 1607567185
transform 1 0 79948 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[55\]
timestamp 1607567185
transform 1 0 79764 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1607567185
transform 1 0 79672 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_855
timestamp 1607567185
transform 1 0 79764 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_860
timestamp 1607567185
transform 1 0 80224 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_852
timestamp 1607567185
transform 1 0 79488 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_864
timestamp 1607567185
transform 1 0 80592 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[51\]
timestamp 1607567185
transform 1 0 77556 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[53\]
timestamp 1607567185
transform 1 0 78200 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1607567185
transform 1 0 78108 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_847
timestamp 1607567185
transform 1 0 79028 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_840
timestamp 1607567185
transform 1 0 78384 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[451\]
timestamp 1607567185
transform 1 0 77096 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[50\]
timestamp 1607567185
transform 1 0 75992 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_816
timestamp 1607567185
transform 1 0 76176 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_824
timestamp 1607567185
transform 1 0 76912 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_829
timestamp 1607567185
transform 1 0 77372 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_811
timestamp 1607567185
transform 1 0 75716 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_823
timestamp 1607567185
transform 1 0 76820 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[395\]
timestamp 1607567185
transform 1 0 74060 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[32\]
timestamp 1607567185
transform 1 0 74152 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[47\]
timestamp 1607567185
transform 1 0 75348 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1607567185
transform 1 0 75256 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1607567185
transform 1 0 74060 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_796
timestamp 1607567185
transform 1 0 74336 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_804
timestamp 1607567185
transform 1 0 75072 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_792
timestamp 1607567185
transform 1 0 73968 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_803
timestamp 1607567185
transform 1 0 74980 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[33\]
timestamp 1607567185
transform 1 0 72496 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1607567185
transform 1 0 72404 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_774
timestamp 1607567185
transform 1 0 72312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_785
timestamp 1607567185
transform 1 0 73324 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_780
timestamp 1607567185
transform 1 0 72864 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[34\]
timestamp 1607567185
transform 1 0 72036 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_766
timestamp 1607567185
transform 1 0 71576 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_763
timestamp 1607567185
transform 1 0 71300 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[21\]
timestamp 1607567185
transform 1 0 69644 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[31\]
timestamp 1607567185
transform 1 0 70472 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1607567185
transform 1 0 69552 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_738
timestamp 1607567185
transform 1 0 69000 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_754
timestamp 1607567185
transform 1 0 70472 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_742
timestamp 1607567185
transform 1 0 69368 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[19\]
timestamp 1607567185
transform 1 0 68540 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1607567185
transform 1 0 68448 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_726
timestamp 1607567185
transform 1 0 67896 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_727
timestamp 1607567185
transform 1 0 67988 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_731
timestamp 1607567185
transform 1 0 68356 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[18\]
timestamp 1607567185
transform 1 0 66056 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1607567185
transform 1 0 66700 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_707
timestamp 1607567185
transform 1 0 66148 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_714
timestamp 1607567185
transform 1 0 66792 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_698
timestamp 1607567185
transform 1 0 65320 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_715
timestamp 1607567185
transform 1 0 66884 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[27\]
timestamp 1607567185
transform 1 0 64492 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1607567185
transform 1 0 63848 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_681
timestamp 1607567185
transform 1 0 63756 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_683
timestamp 1607567185
transform 1 0 63940 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_695
timestamp 1607567185
transform 1 0 65044 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_681
timestamp 1607567185
transform 1 0 63756 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[23\]
timestamp 1607567185
transform 1 0 62928 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1607567185
transform 1 0 62836 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_661
timestamp 1607567185
transform 1 0 61916 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_673
timestamp 1607567185
transform 1 0 63020 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1607567185
transform 1 0 62284 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[16\]
timestamp 1607567185
transform 1 0 60352 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[9\]
timestamp 1607567185
transform 1 0 61088 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1607567185
transform 1 0 60996 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_653
timestamp 1607567185
transform 1 0 61180 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[14\]
timestamp 1607567185
transform 1 0 58788 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[15\]
timestamp 1607567185
transform 1 0 59064 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_629
timestamp 1607567185
transform 1 0 58972 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_639
timestamp 1607567185
transform 1 0 59892 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_626
timestamp 1607567185
transform 1 0 58696 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_636
timestamp 1607567185
transform 1 0 59616 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _596_
timestamp 1607567185
transform 1 0 57316 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1607567185
transform 1 0 58144 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1607567185
transform 1 0 57224 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_608
timestamp 1607567185
transform 1 0 57040 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_621
timestamp 1607567185
transform 1 0 58236 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_606
timestamp 1607567185
transform 1 0 56856 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_614
timestamp 1607567185
transform 1 0 57592 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[0\]
timestamp 1607567185
transform 1 0 56212 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[4\]
timestamp 1607567185
transform 1 0 54924 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1607567185
transform 1 0 55292 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_586
timestamp 1607567185
transform 1 0 55016 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_590
timestamp 1607567185
transform 1 0 55384 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_598
timestamp 1607567185
transform 1 0 56120 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_594
timestamp 1607567185
transform 1 0 55752 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1607567185
transform 1 0 54004 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[5\]
timestamp 1607567185
transform 1 0 53268 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_574
timestamp 1607567185
transform 1 0 53912 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1607567185
transform 1 0 54280 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_576
timestamp 1607567185
transform 1 0 54096 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_584
timestamp 1607567185
transform 1 0 54832 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _592_
timestamp 1607567185
transform 1 0 52532 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  user_to_mprj_in_buffers\[2\]
timestamp 1607567185
transform 1 0 51704 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1607567185
transform 1 0 52440 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1607567185
transform 1 0 51612 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_554
timestamp 1607567185
transform 1 0 52072 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_562
timestamp 1607567185
transform 1 0 52808 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_559
timestamp 1607567185
transform 1 0 52532 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _571_
timestamp 1607567185
transform 1 0 50692 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _587_
timestamp 1607567185
transform 1 0 50600 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_531
timestamp 1607567185
transform 1 0 49956 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_542
timestamp 1607567185
transform 1 0 50968 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_535
timestamp 1607567185
transform 1 0 50324 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_541
timestamp 1607567185
transform 1 0 50876 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _564_
timestamp 1607567185
transform 1 0 49680 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1607567185
transform 1 0 48208 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1607567185
transform 1 0 49588 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_521
timestamp 1607567185
transform 1 0 49036 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_515
timestamp 1607567185
transform 1 0 48484 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_527
timestamp 1607567185
transform 1 0 49588 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1607567185
transform 1 0 47196 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1607567185
transform 1 0 46736 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_497
timestamp 1607567185
transform 1 0 46828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_509
timestamp 1607567185
transform 1 0 47932 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_493
timestamp 1607567185
transform 1 0 46460 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_504
timestamp 1607567185
transform 1 0 47472 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _554_
timestamp 1607567185
transform 1 0 45356 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _566_
timestamp 1607567185
transform 1 0 46184 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1607567185
transform 1 0 46000 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_473
timestamp 1607567185
transform 1 0 44620 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_484
timestamp 1607567185
transform 1 0 45632 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_473
timestamp 1607567185
transform 1 0 44620 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_485
timestamp 1607567185
transform 1 0 45724 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_489
timestamp 1607567185
transform 1 0 46092 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_462
timestamp 1607567185
transform 1 0 43608 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_466
timestamp 1607567185
transform 1 0 43976 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1607567185
transform 1 0 43884 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _556_
timestamp 1607567185
transform 1 0 44344 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _552_
timestamp 1607567185
transform 1 0 44344 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_458
timestamp 1607567185
transform 1 0 43240 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_457
timestamp 1607567185
transform 1 0 43148 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_453
timestamp 1607567185
transform 1 0 42780 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _558_
timestamp 1607567185
transform 1 0 42872 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _550_
timestamp 1607567185
transform 1 0 43332 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp 1607567185
transform 1 0 42228 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_435
timestamp 1607567185
transform 1 0 41124 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_447
timestamp 1607567185
transform 1 0 42228 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_437
timestamp 1607567185
transform 1 0 41308 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_445
timestamp 1607567185
transform 1 0 42044 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_450
timestamp 1607567185
transform 1 0 42504 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[92\]
timestamp 1607567185
transform 1 0 40756 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[98\]
timestamp 1607567185
transform 1 0 40480 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607567185
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_425
timestamp 1607567185
transform 1 0 40204 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_423
timestamp 1607567185
transform 1 0 40020 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[154\]
timestamp 1607567185
transform 1 0 37720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607567185
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1607567185
transform 1 0 37996 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_413
timestamp 1607567185
transform 1 0 39100 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_399
timestamp 1607567185
transform 1 0 37812 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_411
timestamp 1607567185
transform 1 0 38916 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[84\]
timestamp 1607567185
transform 1 0 36156 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[158\]
timestamp 1607567185
transform 1 0 36064 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_383
timestamp 1607567185
transform 1 0 36340 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_395
timestamp 1607567185
transform 1 0 37444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_378
timestamp 1607567185
transform 1 0 35880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[145\]
timestamp 1607567185
transform 1 0 34868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[152\]
timestamp 1607567185
transform 1 0 35052 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607567185
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_361
timestamp 1607567185
transform 1 0 34316 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_372
timestamp 1607567185
transform 1 0 35328 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_363
timestamp 1607567185
transform 1 0 34500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_370
timestamp 1607567185
transform 1 0 35144 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[73\]
timestamp 1607567185
transform 1 0 32660 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_7_351
timestamp 1607567185
transform 1 0 33396 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[70\]
timestamp 1607567185
transform 1 0 31740 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[149\]
timestamp 1607567185
transform 1 0 30728 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607567185
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_321
timestamp 1607567185
transform 1 0 30636 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_325
timestamp 1607567185
transform 1 0 31004 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_333
timestamp 1607567185
transform 1 0 31740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_337
timestamp 1607567185
transform 1 0 32108 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_325
timestamp 1607567185
transform 1 0 31004 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[64\]
timestamp 1607567185
transform 1 0 29348 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607567185
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_313
timestamp 1607567185
transform 1 0 29900 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_306
timestamp 1607567185
transform 1 0 29256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  la_buf\[69\]
timestamp 1607567185
transform 1 0 28244 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_6_284
timestamp 1607567185
transform 1 0 27232 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_292
timestamp 1607567185
transform 1 0 27968 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_287
timestamp 1607567185
transform 1 0 27508 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_299
timestamp 1607567185
transform 1 0 28612 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[140\]
timestamp 1607567185
transform 1 0 26956 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607567185
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_269
timestamp 1607567185
transform 1 0 25852 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_276
timestamp 1607567185
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_280
timestamp 1607567185
transform 1 0 26864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_275
timestamp 1607567185
transform 1 0 26404 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[45\]
timestamp 1607567185
transform 1 0 23644 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_6_257
timestamp 1607567185
transform 1 0 24748 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_263
timestamp 1607567185
transform 1 0 25300 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[40\]
timestamp 1607567185
transform 1 0 23092 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607567185
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_229
timestamp 1607567185
transform 1 0 22172 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_237
timestamp 1607567185
transform 1 0 22908 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_238
timestamp 1607567185
transform 1 0 23000 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[113\]
timestamp 1607567185
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[117\]
timestamp 1607567185
transform 1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[118\]
timestamp 1607567185
transform 1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607567185
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1607567185
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_218
timestamp 1607567185
transform 1 0 21160 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1607567185
transform 1 0 20884 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_226
timestamp 1607567185
transform 1 0 21896 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[39\]
timestamp 1607567185
transform 1 0 19228 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[116\]
timestamp 1607567185
transform 1 0 19320 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 1607567185
transform 1 0 19228 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1607567185
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_196
timestamp 1607567185
transform 1 0 19136 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[112\]
timestamp 1607567185
transform 1 0 16744 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607567185
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_173
timestamp 1607567185
transform 1 0 17020 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_185
timestamp 1607567185
transform 1 0 18124 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1607567185
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1607567185
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[105\]
timestamp 1607567185
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607567185
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1607567185
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_157
timestamp 1607567185
transform 1 0 15548 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1607567185
transform 1 0 16652 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_167
timestamp 1607567185
transform 1 0 16468 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[31\]
timestamp 1607567185
transform 1 0 14812 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[101\]
timestamp 1607567185
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_136
timestamp 1607567185
transform 1 0 13616 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1607567185
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_141
timestamp 1607567185
transform 1 0 14076 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[27\]
timestamp 1607567185
transform 1 0 12420 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607567185
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_125
timestamp 1607567185
transform 1 0 12604 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1607567185
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  la_buf\[26\]
timestamp 1607567185
transform 1 0 10948 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[100\]
timestamp 1607567185
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_96
timestamp 1607567185
transform 1 0 9936 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_104
timestamp 1607567185
transform 1 0 10672 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_103
timestamp 1607567185
transform 1 0 10580 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_109
timestamp 1607567185
transform 1 0 11132 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[92\]
timestamp 1607567185
transform 1 0 9200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[99\]
timestamp 1607567185
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607567185
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_82
timestamp 1607567185
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1607567185
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_80
timestamp 1607567185
transform 1 0 8464 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_91
timestamp 1607567185
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[17\]
timestamp 1607567185
transform 1 0 6808 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  la_buf\[19\]
timestamp 1607567185
transform 1 0 6992 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607567185
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  la_buf\[10\]
timestamp 1607567185
transform 1 0 4600 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_6_56
timestamp 1607567185
transform 1 0 6256 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1607567185
transform 1 0 5980 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[14\]
timestamp 1607567185
transform 1 0 4324 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[84\]
timestamp 1607567185
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[88\]
timestamp 1607567185
transform 1 0 3312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607567185
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_19
timestamp 1607567185
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1607567185
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_32
timestamp 1607567185
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1607567185
transform 1 0 3588 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[93\]
timestamp 1607567185
transform 1 0 2300 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607567185
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607567185
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607567185
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1607567185
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1607567185
transform 1 0 1380 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1607567185
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_16
timestamp 1607567185
transform 1 0 2576 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[166\]
timestamp 1607567185
transform 1 0 40480 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1607567185
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_415
timestamp 1607567185
transform 1 0 39284 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_431
timestamp 1607567185
transform 1 0 40756 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_403
timestamp 1607567185
transform 1 0 38180 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1607567185
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_391
timestamp 1607567185
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1607567185
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_363
timestamp 1607567185
transform 1 0 34500 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1607567185
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[147\]
timestamp 1607567185
transform 1 0 33488 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_344
timestamp 1607567185
transform 1 0 32752 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_355
timestamp 1607567185
transform 1 0 33764 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[75\]
timestamp 1607567185
transform 1 0 31096 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_5_325
timestamp 1607567185
transform 1 0 31004 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[138\]
timestamp 1607567185
transform 1 0 29624 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1607567185
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_302
timestamp 1607567185
transform 1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_306
timestamp 1607567185
transform 1 0 29256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_313
timestamp 1607567185
transform 1 0 29900 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_294
timestamp 1607567185
transform 1 0 28152 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[66\]
timestamp 1607567185
transform 1 0 26496 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_5_275
timestamp 1607567185
transform 1 0 26404 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_8  la_buf\[48\]
timestamp 1607567185
transform 1 0 23644 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_5_263
timestamp 1607567185
transform 1 0 25300 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[119\]
timestamp 1607567185
transform 1 0 22540 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1607567185
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_230
timestamp 1607567185
transform 1 0 22264 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_236
timestamp 1607567185
transform 1 0 22816 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_218
timestamp 1607567185
transform 1 0 21160 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[59\]
timestamp 1607567185
transform 1 0 19504 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_5_196
timestamp 1607567185
transform 1 0 19136 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1607567185
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_173
timestamp 1607567185
transform 1 0 17020 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1607567185
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1607567185
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_161
timestamp 1607567185
transform 1 0 15916 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[103\]
timestamp 1607567185
transform 1 0 13432 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1607567185
transform 1 0 13708 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1607567185
transform 1 0 14812 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[102\]
timestamp 1607567185
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1607567185
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1607567185
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_126
timestamp 1607567185
transform 1 0 12696 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_111
timestamp 1607567185
transform 1 0 11316 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[25\]
timestamp 1607567185
transform 1 0 9660 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_5_85
timestamp 1607567185
transform 1 0 8924 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  la_buf\[23\]
timestamp 1607567185
transform 1 0 7268 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1607567185
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1607567185
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1607567185
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1607567185
transform 1 0 7176 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1607567185
transform 1 0 5244 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_48
timestamp 1607567185
transform 1 0 5520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _478_
timestamp 1607567185
transform 1 0 4232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _479_
timestamp 1607567185
transform 1 0 3220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_26
timestamp 1607567185
transform 1 0 3496 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_37
timestamp 1607567185
transform 1 0 4508 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607567185
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607567185
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1607567185
transform 1 0 2484 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_425
timestamp 1607567185
transform 1 0 40204 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _557_
timestamp 1607567185
transform 1 0 37720 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1607567185
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1607567185
transform 1 0 37996 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_413
timestamp 1607567185
transform 1 0 39100 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_383
timestamp 1607567185
transform 1 0 36340 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_395
timestamp 1607567185
transform 1 0 37444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_359
timestamp 1607567185
transform 1 0 34132 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_371
timestamp 1607567185
transform 1 0 35236 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[78\]
timestamp 1607567185
transform 1 0 32476 0 -1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1607567185
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_323
timestamp 1607567185
transform 1 0 30820 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1607567185
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_337
timestamp 1607567185
transform 1 0 32108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_311
timestamp 1607567185
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _533_
timestamp 1607567185
transform 1 0 27140 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[143\]
timestamp 1607567185
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_286
timestamp 1607567185
transform 1 0 27416 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_294
timestamp 1607567185
transform 1 0 28152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_299
timestamp 1607567185
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1607567185
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_273
timestamp 1607567185
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_276
timestamp 1607567185
transform 1 0 26496 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_282
timestamp 1607567185
transform 1 0 27048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _531_
timestamp 1607567185
transform 1 0 24840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[114\]
timestamp 1607567185
transform 1 0 23828 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_250
timestamp 1607567185
transform 1 0 24104 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_261
timestamp 1607567185
transform 1 0 25116 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[122\]
timestamp 1607567185
transform 1 0 22816 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_227
timestamp 1607567185
transform 1 0 21988 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_235
timestamp 1607567185
transform 1 0 22724 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_239
timestamp 1607567185
transform 1 0 23092 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1607567185
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1607567185
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _512_
timestamp 1607567185
transform 1 0 18768 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[133\]
timestamp 1607567185
transform 1 0 19780 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1607567185
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_195
timestamp 1607567185
transform 1 0 19044 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1607567185
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1607567185
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1607567185
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1607567185
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1607567185
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1607567185
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_140
timestamp 1607567185
transform 1 0 13984 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_128
timestamp 1607567185
transform 1 0 12880 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  la_buf\[29\]
timestamp 1607567185
transform 1 0 11224 0 -1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_4_96
timestamp 1607567185
transform 1 0 9936 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1607567185
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mprj_logic_high\[97\]
timestamp 1607567185
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1607567185
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_76
timestamp 1607567185
transform 1 0 8096 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1607567185
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _477_
timestamp 1607567185
transform 1 0 6532 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _490_
timestamp 1607567185
transform 1 0 7820 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_62
timestamp 1607567185
transform 1 0 6808 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_70
timestamp 1607567185
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1607567185
transform 1 0 5520 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_40
timestamp 1607567185
transform 1 0 4784 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1607567185
transform 1 0 5796 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1607567185
transform 1 0 4508 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1607567185
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607567185
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1607567185
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1607567185
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607567185
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607567185
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607567185
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_434
timestamp 1607567185
transform 1 0 41032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1607567185
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_415
timestamp 1607567185
transform 1 0 39284 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_428
timestamp 1607567185
transform 1 0 40480 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_403
timestamp 1607567185
transform 1 0 38180 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1607567185
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_391
timestamp 1607567185
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1607567185
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_364
timestamp 1607567185
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1607567185
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _542_
timestamp 1607567185
transform 1 0 33212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_341
timestamp 1607567185
transform 1 0 32476 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_352
timestamp 1607567185
transform 1 0 33488 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _547_
timestamp 1607567185
transform 1 0 32200 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_321
timestamp 1607567185
transform 1 0 30636 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_333
timestamp 1607567185
transform 1 0 31740 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_337
timestamp 1607567185
transform 1 0 32108 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _532_
timestamp 1607567185
transform 1 0 29256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1607567185
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_304
timestamp 1607567185
transform 1 0 29072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_309
timestamp 1607567185
transform 1 0 29532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_284
timestamp 1607567185
transform 1 0 27232 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_296
timestamp 1607567185
transform 1 0 28336 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _530_
timestamp 1607567185
transform 1 0 25392 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _538_
timestamp 1607567185
transform 1 0 26956 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_267
timestamp 1607567185
transform 1 0 25668 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_279
timestamp 1607567185
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _539_
timestamp 1607567185
transform 1 0 24380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1607567185
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_256
timestamp 1607567185
transform 1 0 24656 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1607567185
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_231
timestamp 1607567185
transform 1 0 22356 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1607567185
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _515_
timestamp 1607567185
transform 1 0 20976 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_215
timestamp 1607567185
transform 1 0 20884 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_219
timestamp 1607567185
transform 1 0 21252 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _513_
timestamp 1607567185
transform 1 0 19872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_196
timestamp 1607567185
transform 1 0 19136 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_207
timestamp 1607567185
transform 1 0 20148 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1607567185
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_176
timestamp 1607567185
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1607567185
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1607567185
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1607567185
transform 1 0 15088 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_164
timestamp 1607567185
transform 1 0 16192 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _499_
timestamp 1607567185
transform 1 0 13432 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _504_
timestamp 1607567185
transform 1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1607567185
transform 1 0 13708 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _497_
timestamp 1607567185
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1607567185
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_114
timestamp 1607567185
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_126
timestamp 1607567185
transform 1 0 12696 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _493_
timestamp 1607567185
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_99
timestamp 1607567185
transform 1 0 10212 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _491_
timestamp 1607567185
transform 1 0 8832 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_76
timestamp 1607567185
transform 1 0 8096 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_87
timestamp 1607567185
transform 1 0 9108 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1607567185
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _487_
timestamp 1607567185
transform 1 0 7820 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1607567185
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1607567185
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_65
timestamp 1607567185
transform 1 0 7084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 1607567185
transform 1 0 5520 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_40
timestamp 1607567185
transform 1 0 4784 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1607567185
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1607567185
transform 1 0 4508 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1607567185
transform 1 0 3588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1607567185
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607567185
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607567185
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1607567185
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_426
timestamp 1607567185
transform 1 0 40296 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _549_
timestamp 1607567185
transform 1 0 37812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1607567185
transform 1 0 37628 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_396
timestamp 1607567185
transform 1 0 37536 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_398
timestamp 1607567185
transform 1 0 37720 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_402
timestamp 1607567185
transform 1 0 38088 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_414
timestamp 1607567185
transform 1 0 39192 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _548_
timestamp 1607567185
transform 1 0 35788 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_380
timestamp 1607567185
transform 1 0 36064 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_392
timestamp 1607567185
transform 1 0 37168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_364
timestamp 1607567185
transform 1 0 34592 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_376
timestamp 1607567185
transform 1 0 35696 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _536_
timestamp 1607567185
transform 1 0 33212 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_352
timestamp 1607567185
transform 1 0 33488 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1607567185
transform 1 0 32016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_327
timestamp 1607567185
transform 1 0 31188 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_335
timestamp 1607567185
transform 1 0 31924 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_337
timestamp 1607567185
transform 1 0 32108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_303
timestamp 1607567185
transform 1 0 28980 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_315
timestamp 1607567185
transform 1 0 30084 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_291
timestamp 1607567185
transform 1 0 27876 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _528_
timestamp 1607567185
transform 1 0 26496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1607567185
transform 1 0 26404 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_279
timestamp 1607567185
transform 1 0 26772 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _524_
timestamp 1607567185
transform 1 0 23828 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _526_
timestamp 1607567185
transform 1 0 25024 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_250
timestamp 1607567185
transform 1 0 24104 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1607567185
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1607567185
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_229
timestamp 1607567185
transform 1 0 22172 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_241
timestamp 1607567185
transform 1 0 23276 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _510_
timestamp 1607567185
transform 1 0 20884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _517_
timestamp 1607567185
transform 1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1607567185
transform 1 0 20792 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1607567185
transform 1 0 20700 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_218
timestamp 1607567185
transform 1 0 21160 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_189
timestamp 1607567185
transform 1 0 18492 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1607567185
transform 1 0 19596 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 1607567185
transform 1 0 17112 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_173
timestamp 1607567185
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1607567185
transform 1 0 17388 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 1607567185
transform 1 0 15272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1607567185
transform 1 0 15180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_157
timestamp 1607567185
transform 1 0 15548 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_169
timestamp 1607567185
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _500_
timestamp 1607567185
transform 1 0 13800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_136
timestamp 1607567185
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1607567185
transform 1 0 14076 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_116
timestamp 1607567185
transform 1 0 11776 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_128
timestamp 1607567185
transform 1 0 12880 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _495_
timestamp 1607567185
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_105
timestamp 1607567185
transform 1 0 10764 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _489_
timestamp 1607567185
transform 1 0 8464 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1607567185
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_83
timestamp 1607567185
transform 1 0 8740 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1607567185
transform 1 0 9476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607567185
transform 1 0 9660 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _484_
timestamp 1607567185
transform 1 0 6440 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1607567185
transform 1 0 7452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_61
timestamp 1607567185
transform 1 0 6716 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_72
timestamp 1607567185
transform 1 0 7728 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _473_
timestamp 1607567185
transform 1 0 5428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp 1607567185
transform 1 0 5152 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_50
timestamp 1607567185
transform 1 0 5704 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1607567185
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607567185
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607567185
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607567185
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607567185
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607567185
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _555_
timestamp 1607567185
transform 1 0 41032 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1607567185
transform 1 0 41032 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _553_
timestamp 1607567185
transform 1 0 39284 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1607567185
transform 1 0 40388 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_415
timestamp 1607567185
transform 1 0 39284 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_427
timestamp 1607567185
transform 1 0 40388 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1607567185
transform 1 0 40940 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_418
timestamp 1607567185
transform 1 0 39560 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_426
timestamp 1607567185
transform 1 0 40296 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_428
timestamp 1607567185
transform 1 0 40480 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _543_
timestamp 1607567185
transform 1 0 37720 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _551_
timestamp 1607567185
transform 1 0 39008 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1607567185
transform 1 0 38180 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_400
timestamp 1607567185
transform 1 0 37904 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_404
timestamp 1607567185
transform 1 0 38272 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_397
timestamp 1607567185
transform 1 0 37628 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_401
timestamp 1607567185
transform 1 0 37996 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_413
timestamp 1607567185
transform 1 0 39100 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _546_
timestamp 1607567185
transform 1 0 36248 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_388
timestamp 1607567185
transform 1 0 36800 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_385
timestamp 1607567185
transform 1 0 36524 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _544_
timestamp 1607567185
transform 1 0 34868 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _545_
timestamp 1607567185
transform 1 0 35420 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1607567185
transform 1 0 35328 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1607567185
transform 1 0 34776 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_359
timestamp 1607567185
transform 1 0 34132 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_371
timestamp 1607567185
transform 1 0 35236 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_376
timestamp 1607567185
transform 1 0 35696 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_364
timestamp 1607567185
transform 1 0 34592 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_370
timestamp 1607567185
transform 1 0 35144 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _529_
timestamp 1607567185
transform 1 0 33856 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _534_
timestamp 1607567185
transform 1 0 33212 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _541_
timestamp 1607567185
transform 1 0 32844 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1607567185
transform 1 0 32476 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_342
timestamp 1607567185
transform 1 0 32568 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_348
timestamp 1607567185
transform 1 0 33120 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_341
timestamp 1607567185
transform 1 0 32476 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_352
timestamp 1607567185
transform 1 0 33488 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _537_
timestamp 1607567185
transform 1 0 31188 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _540_
timestamp 1607567185
transform 1 0 32200 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_323
timestamp 1607567185
transform 1 0 30820 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_335
timestamp 1607567185
transform 1 0 31924 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_330
timestamp 1607567185
transform 1 0 31464 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _535_
timestamp 1607567185
transform 1 0 30176 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1607567185
transform 1 0 29624 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1607567185
transform 1 0 29164 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_308
timestamp 1607567185
transform 1 0 29440 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_311
timestamp 1607567185
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_304
timestamp 1607567185
transform 1 0 29072 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_306
timestamp 1607567185
transform 1 0 29256 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_314
timestamp 1607567185
transform 1 0 29992 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_319
timestamp 1607567185
transform 1 0 30452 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _525_
timestamp 1607567185
transform 1 0 28428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_292
timestamp 1607567185
transform 1 0 27968 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_296
timestamp 1607567185
transform 1 0 28336 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1607567185
transform 1 0 28704 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_292
timestamp 1607567185
transform 1 0 27968 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _523_
timestamp 1607567185
transform 1 0 25576 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _527_
timestamp 1607567185
transform 1 0 26588 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1607567185
transform 1 0 26772 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_264
timestamp 1607567185
transform 1 0 25392 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_276
timestamp 1607567185
transform 1 0 26496 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1607567185
transform 1 0 26864 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1607567185
transform 1 0 25852 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_280
timestamp 1607567185
transform 1 0 26864 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _520_
timestamp 1607567185
transform 1 0 23644 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _521_
timestamp 1607567185
transform 1 0 24104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _522_
timestamp 1607567185
transform 1 0 25116 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1607567185
transform 1 0 23920 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_246
timestamp 1607567185
transform 1 0 23736 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_249
timestamp 1607567185
transform 1 0 24012 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1607567185
transform 1 0 24380 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_248
timestamp 1607567185
transform 1 0 23920 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_260
timestamp 1607567185
transform 1 0 25024 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _518_
timestamp 1607567185
transform 1 0 22356 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _519_
timestamp 1607567185
transform 1 0 22540 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1607567185
transform 1 0 23552 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_234
timestamp 1607567185
transform 1 0 22632 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_236
timestamp 1607567185
transform 1 0 22816 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1607567185
transform 1 0 21804 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_221
timestamp 1607567185
transform 1 0 21436 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_223
timestamp 1607567185
transform 1 0 21620 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1607567185
transform 1 0 21160 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1607567185
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _516_
timestamp 1607567185
transform 1 0 21344 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _511_
timestamp 1607567185
transform 1 0 21528 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_213
timestamp 1607567185
transform 1 0 20700 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 1607567185
transform 1 0 20332 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 1607567185
transform 1 0 20424 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _514_
timestamp 1607567185
transform 1 0 20056 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_199
timestamp 1607567185
transform 1 0 19412 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1607567185
transform 1 0 19964 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_199
timestamp 1607567185
transform 1 0 19412 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_207
timestamp 1607567185
transform 1 0 20148 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _503_
timestamp 1607567185
transform 1 0 16744 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _509_
timestamp 1607567185
transform 1 0 18032 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1607567185
transform 1 0 18216 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1607567185
transform 1 0 17940 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_173
timestamp 1607567185
transform 1 0 17020 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1607567185
transform 1 0 18124 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1607567185
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1607567185
transform 1 0 17572 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_187
timestamp 1607567185
transform 1 0 18308 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 1607567185
transform 1 0 16192 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _508_
timestamp 1607567185
transform 1 0 15732 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1607567185
transform 1 0 15364 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1607567185
transform 1 0 15456 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_162
timestamp 1607567185
transform 1 0 16008 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_152
timestamp 1607567185
transform 1 0 15088 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_167
timestamp 1607567185
transform 1 0 16468 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _498_
timestamp 1607567185
transform 1 0 13708 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1607567185
transform 1 0 13708 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1607567185
transform 1 0 14812 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_140
timestamp 1607567185
transform 1 0 13984 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _501_
timestamp 1607567185
transform 1 0 12696 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1607567185
transform 1 0 12512 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1607567185
transform 1 0 12328 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1607567185
transform 1 0 11960 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1607567185
transform 1 0 12604 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1607567185
transform 1 0 11592 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1607567185
transform 1 0 12420 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_129
timestamp 1607567185
transform 1 0 12972 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _494_
timestamp 1607567185
transform 1 0 9844 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _496_
timestamp 1607567185
transform 1 0 11316 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1607567185
transform 1 0 10856 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1607567185
transform 1 0 10120 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_110
timestamp 1607567185
transform 1 0 11224 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1607567185
transform 1 0 8832 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34
timestamp 1607567185
transform 1 0 9660 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_77
timestamp 1607567185
transform 1 0 8188 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1607567185
transform 1 0 9292 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1607567185
transform 1 0 9752 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_76
timestamp 1607567185
transform 1 0 8096 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_87
timestamp 1607567185
transform 1 0 9108 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66
timestamp 1607567185
transform 1 0 7176 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 1607567185
transform 1 0 7912 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _485_
timestamp 1607567185
transform 1 0 7820 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_65
timestamp 1607567185
transform 1 0 7084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1607567185
transform 1 0 6624 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1607567185
transform 1 0 6624 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1607567185
transform 1 0 6716 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_33
timestamp 1607567185
transform 1 0 6808 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _483_
timestamp 1607567185
transform 1 0 6808 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _482_
timestamp 1607567185
transform 1 0 6900 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1607567185
transform 1 0 5244 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _481_
timestamp 1607567185
transform 1 0 5244 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44
timestamp 1607567185
transform 1 0 5152 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_48
timestamp 1607567185
transform 1 0 5520 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_39
timestamp 1607567185
transform 1 0 4692 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_48
timestamp 1607567185
transform 1 0 5520 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_32
timestamp 1607567185
transform 1 0 3956 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1607567185
transform 1 0 3588 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607567185
transform 1 0 4048 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1607567185
transform 1 0 3588 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607567185
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1607567185
transform 1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1607567185
transform 1 0 1380 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607567185
transform 1 0 2484 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1607567185
transform 1 0 1380 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1607567185
transform 1 0 2484 0 1 1632
box -38 -48 1142 592
<< labels >>
rlabel metal3 s -400 1776 800 1896 4 caravel_clk
port 1 nsew
rlabel metal3 s -400 5448 800 5568 4 caravel_clk2
port 2 nsew
rlabel metal3 s -400 9120 800 9240 4 caravel_rstn
port 3 nsew
rlabel metal2 s 1858 10200 1914 11400 4 la_data_in_core[0]
port 4 nsew
rlabel metal2 s 45466 10200 45522 11400 4 la_data_in_core[100]
port 5 nsew
rlabel metal2 s 45926 10200 45982 11400 4 la_data_in_core[101]
port 6 nsew
rlabel metal2 s 46386 10200 46442 11400 4 la_data_in_core[102]
port 7 nsew
rlabel metal2 s 46754 10200 46810 11400 4 la_data_in_core[103]
port 8 nsew
rlabel metal2 s 47214 10200 47270 11400 4 la_data_in_core[104]
port 9 nsew
rlabel metal2 s 47674 10200 47730 11400 4 la_data_in_core[105]
port 10 nsew
rlabel metal2 s 48134 10200 48190 11400 4 la_data_in_core[106]
port 11 nsew
rlabel metal2 s 48502 10200 48558 11400 4 la_data_in_core[107]
port 12 nsew
rlabel metal2 s 48962 10200 49018 11400 4 la_data_in_core[108]
port 13 nsew
rlabel metal2 s 49422 10200 49478 11400 4 la_data_in_core[109]
port 14 nsew
rlabel metal2 s 6274 10200 6330 11400 4 la_data_in_core[10]
port 15 nsew
rlabel metal2 s 49790 10200 49846 11400 4 la_data_in_core[110]
port 16 nsew
rlabel metal2 s 50250 10200 50306 11400 4 la_data_in_core[111]
port 17 nsew
rlabel metal2 s 50710 10200 50766 11400 4 la_data_in_core[112]
port 18 nsew
rlabel metal2 s 51170 10200 51226 11400 4 la_data_in_core[113]
port 19 nsew
rlabel metal2 s 51538 10200 51594 11400 4 la_data_in_core[114]
port 20 nsew
rlabel metal2 s 51998 10200 52054 11400 4 la_data_in_core[115]
port 21 nsew
rlabel metal2 s 52458 10200 52514 11400 4 la_data_in_core[116]
port 22 nsew
rlabel metal2 s 52918 10200 52974 11400 4 la_data_in_core[117]
port 23 nsew
rlabel metal2 s 53286 10200 53342 11400 4 la_data_in_core[118]
port 24 nsew
rlabel metal2 s 53746 10200 53802 11400 4 la_data_in_core[119]
port 25 nsew
rlabel metal2 s 6734 10200 6790 11400 4 la_data_in_core[11]
port 26 nsew
rlabel metal2 s 54206 10200 54262 11400 4 la_data_in_core[120]
port 27 nsew
rlabel metal2 s 54666 10200 54722 11400 4 la_data_in_core[121]
port 28 nsew
rlabel metal2 s 55034 10200 55090 11400 4 la_data_in_core[122]
port 29 nsew
rlabel metal2 s 55494 10200 55550 11400 4 la_data_in_core[123]
port 30 nsew
rlabel metal2 s 55954 10200 56010 11400 4 la_data_in_core[124]
port 31 nsew
rlabel metal2 s 56322 10200 56378 11400 4 la_data_in_core[125]
port 32 nsew
rlabel metal2 s 56782 10200 56838 11400 4 la_data_in_core[126]
port 33 nsew
rlabel metal2 s 57242 10200 57298 11400 4 la_data_in_core[127]
port 34 nsew
rlabel metal2 s 7102 10200 7158 11400 4 la_data_in_core[12]
port 35 nsew
rlabel metal2 s 7562 10200 7618 11400 4 la_data_in_core[13]
port 36 nsew
rlabel metal2 s 8022 10200 8078 11400 4 la_data_in_core[14]
port 37 nsew
rlabel metal2 s 8390 10200 8446 11400 4 la_data_in_core[15]
port 38 nsew
rlabel metal2 s 8850 10200 8906 11400 4 la_data_in_core[16]
port 39 nsew
rlabel metal2 s 9310 10200 9366 11400 4 la_data_in_core[17]
port 40 nsew
rlabel metal2 s 9770 10200 9826 11400 4 la_data_in_core[18]
port 41 nsew
rlabel metal2 s 10138 10200 10194 11400 4 la_data_in_core[19]
port 42 nsew
rlabel metal2 s 2318 10200 2374 11400 4 la_data_in_core[1]
port 43 nsew
rlabel metal2 s 10598 10200 10654 11400 4 la_data_in_core[20]
port 44 nsew
rlabel metal2 s 11058 10200 11114 11400 4 la_data_in_core[21]
port 45 nsew
rlabel metal2 s 11518 10200 11574 11400 4 la_data_in_core[22]
port 46 nsew
rlabel metal2 s 11886 10200 11942 11400 4 la_data_in_core[23]
port 47 nsew
rlabel metal2 s 12346 10200 12402 11400 4 la_data_in_core[24]
port 48 nsew
rlabel metal2 s 12806 10200 12862 11400 4 la_data_in_core[25]
port 49 nsew
rlabel metal2 s 13266 10200 13322 11400 4 la_data_in_core[26]
port 50 nsew
rlabel metal2 s 13634 10200 13690 11400 4 la_data_in_core[27]
port 51 nsew
rlabel metal2 s 14094 10200 14150 11400 4 la_data_in_core[28]
port 52 nsew
rlabel metal2 s 14554 10200 14610 11400 4 la_data_in_core[29]
port 53 nsew
rlabel metal2 s 2778 10200 2834 11400 4 la_data_in_core[2]
port 54 nsew
rlabel metal2 s 15014 10200 15070 11400 4 la_data_in_core[30]
port 55 nsew
rlabel metal2 s 15382 10200 15438 11400 4 la_data_in_core[31]
port 56 nsew
rlabel metal2 s 15842 10200 15898 11400 4 la_data_in_core[32]
port 57 nsew
rlabel metal2 s 16302 10200 16358 11400 4 la_data_in_core[33]
port 58 nsew
rlabel metal2 s 16670 10200 16726 11400 4 la_data_in_core[34]
port 59 nsew
rlabel metal2 s 17130 10200 17186 11400 4 la_data_in_core[35]
port 60 nsew
rlabel metal2 s 17590 10200 17646 11400 4 la_data_in_core[36]
port 61 nsew
rlabel metal2 s 18050 10200 18106 11400 4 la_data_in_core[37]
port 62 nsew
rlabel metal2 s 18418 10200 18474 11400 4 la_data_in_core[38]
port 63 nsew
rlabel metal2 s 18878 10200 18934 11400 4 la_data_in_core[39]
port 64 nsew
rlabel metal2 s 3238 10200 3294 11400 4 la_data_in_core[3]
port 65 nsew
rlabel metal2 s 19338 10200 19394 11400 4 la_data_in_core[40]
port 66 nsew
rlabel metal2 s 19798 10200 19854 11400 4 la_data_in_core[41]
port 67 nsew
rlabel metal2 s 20166 10200 20222 11400 4 la_data_in_core[42]
port 68 nsew
rlabel metal2 s 20626 10200 20682 11400 4 la_data_in_core[43]
port 69 nsew
rlabel metal2 s 21086 10200 21142 11400 4 la_data_in_core[44]
port 70 nsew
rlabel metal2 s 21546 10200 21602 11400 4 la_data_in_core[45]
port 71 nsew
rlabel metal2 s 21914 10200 21970 11400 4 la_data_in_core[46]
port 72 nsew
rlabel metal2 s 22374 10200 22430 11400 4 la_data_in_core[47]
port 73 nsew
rlabel metal2 s 22834 10200 22890 11400 4 la_data_in_core[48]
port 74 nsew
rlabel metal2 s 23294 10200 23350 11400 4 la_data_in_core[49]
port 75 nsew
rlabel metal2 s 3606 10200 3662 11400 4 la_data_in_core[4]
port 76 nsew
rlabel metal2 s 23662 10200 23718 11400 4 la_data_in_core[50]
port 77 nsew
rlabel metal2 s 24122 10200 24178 11400 4 la_data_in_core[51]
port 78 nsew
rlabel metal2 s 24582 10200 24638 11400 4 la_data_in_core[52]
port 79 nsew
rlabel metal2 s 24950 10200 25006 11400 4 la_data_in_core[53]
port 80 nsew
rlabel metal2 s 25410 10200 25466 11400 4 la_data_in_core[54]
port 81 nsew
rlabel metal2 s 25870 10200 25926 11400 4 la_data_in_core[55]
port 82 nsew
rlabel metal2 s 26330 10200 26386 11400 4 la_data_in_core[56]
port 83 nsew
rlabel metal2 s 26698 10200 26754 11400 4 la_data_in_core[57]
port 84 nsew
rlabel metal2 s 27158 10200 27214 11400 4 la_data_in_core[58]
port 85 nsew
rlabel metal2 s 27618 10200 27674 11400 4 la_data_in_core[59]
port 86 nsew
rlabel metal2 s 4066 10200 4122 11400 4 la_data_in_core[5]
port 87 nsew
rlabel metal2 s 28078 10200 28134 11400 4 la_data_in_core[60]
port 88 nsew
rlabel metal2 s 28446 10200 28502 11400 4 la_data_in_core[61]
port 89 nsew
rlabel metal2 s 28906 10200 28962 11400 4 la_data_in_core[62]
port 90 nsew
rlabel metal2 s 29366 10200 29422 11400 4 la_data_in_core[63]
port 91 nsew
rlabel metal2 s 29826 10200 29882 11400 4 la_data_in_core[64]
port 92 nsew
rlabel metal2 s 30194 10200 30250 11400 4 la_data_in_core[65]
port 93 nsew
rlabel metal2 s 30654 10200 30710 11400 4 la_data_in_core[66]
port 94 nsew
rlabel metal2 s 31114 10200 31170 11400 4 la_data_in_core[67]
port 95 nsew
rlabel metal2 s 31574 10200 31630 11400 4 la_data_in_core[68]
port 96 nsew
rlabel metal2 s 31942 10200 31998 11400 4 la_data_in_core[69]
port 97 nsew
rlabel metal2 s 4526 10200 4582 11400 4 la_data_in_core[6]
port 98 nsew
rlabel metal2 s 32402 10200 32458 11400 4 la_data_in_core[70]
port 99 nsew
rlabel metal2 s 32862 10200 32918 11400 4 la_data_in_core[71]
port 100 nsew
rlabel metal2 s 33230 10200 33286 11400 4 la_data_in_core[72]
port 101 nsew
rlabel metal2 s 33690 10200 33746 11400 4 la_data_in_core[73]
port 102 nsew
rlabel metal2 s 34150 10200 34206 11400 4 la_data_in_core[74]
port 103 nsew
rlabel metal2 s 34610 10200 34666 11400 4 la_data_in_core[75]
port 104 nsew
rlabel metal2 s 34978 10200 35034 11400 4 la_data_in_core[76]
port 105 nsew
rlabel metal2 s 35438 10200 35494 11400 4 la_data_in_core[77]
port 106 nsew
rlabel metal2 s 35898 10200 35954 11400 4 la_data_in_core[78]
port 107 nsew
rlabel metal2 s 36358 10200 36414 11400 4 la_data_in_core[79]
port 108 nsew
rlabel metal2 s 4986 10200 5042 11400 4 la_data_in_core[7]
port 109 nsew
rlabel metal2 s 36726 10200 36782 11400 4 la_data_in_core[80]
port 110 nsew
rlabel metal2 s 37186 10200 37242 11400 4 la_data_in_core[81]
port 111 nsew
rlabel metal2 s 37646 10200 37702 11400 4 la_data_in_core[82]
port 112 nsew
rlabel metal2 s 38106 10200 38162 11400 4 la_data_in_core[83]
port 113 nsew
rlabel metal2 s 38474 10200 38530 11400 4 la_data_in_core[84]
port 114 nsew
rlabel metal2 s 38934 10200 38990 11400 4 la_data_in_core[85]
port 115 nsew
rlabel metal2 s 39394 10200 39450 11400 4 la_data_in_core[86]
port 116 nsew
rlabel metal2 s 39854 10200 39910 11400 4 la_data_in_core[87]
port 117 nsew
rlabel metal2 s 40222 10200 40278 11400 4 la_data_in_core[88]
port 118 nsew
rlabel metal2 s 40682 10200 40738 11400 4 la_data_in_core[89]
port 119 nsew
rlabel metal2 s 5354 10200 5410 11400 4 la_data_in_core[8]
port 120 nsew
rlabel metal2 s 41142 10200 41198 11400 4 la_data_in_core[90]
port 121 nsew
rlabel metal2 s 41510 10200 41566 11400 4 la_data_in_core[91]
port 122 nsew
rlabel metal2 s 41970 10200 42026 11400 4 la_data_in_core[92]
port 123 nsew
rlabel metal2 s 42430 10200 42486 11400 4 la_data_in_core[93]
port 124 nsew
rlabel metal2 s 42890 10200 42946 11400 4 la_data_in_core[94]
port 125 nsew
rlabel metal2 s 43258 10200 43314 11400 4 la_data_in_core[95]
port 126 nsew
rlabel metal2 s 43718 10200 43774 11400 4 la_data_in_core[96]
port 127 nsew
rlabel metal2 s 44178 10200 44234 11400 4 la_data_in_core[97]
port 128 nsew
rlabel metal2 s 44638 10200 44694 11400 4 la_data_in_core[98]
port 129 nsew
rlabel metal2 s 45006 10200 45062 11400 4 la_data_in_core[99]
port 130 nsew
rlabel metal2 s 5814 10200 5870 11400 4 la_data_in_core[9]
port 131 nsew
rlabel metal2 s 55954 -400 56010 800 4 la_data_in_mprj[0]
port 132 nsew
rlabel metal2 s 99470 -400 99526 800 4 la_data_in_mprj[100]
port 133 nsew
rlabel metal2 s 99930 -400 99986 800 4 la_data_in_mprj[101]
port 134 nsew
rlabel metal2 s 100390 -400 100446 800 4 la_data_in_mprj[102]
port 135 nsew
rlabel metal2 s 100850 -400 100906 800 4 la_data_in_mprj[103]
port 136 nsew
rlabel metal2 s 101218 -400 101274 800 4 la_data_in_mprj[104]
port 137 nsew
rlabel metal2 s 101678 -400 101734 800 4 la_data_in_mprj[105]
port 138 nsew
rlabel metal2 s 102138 -400 102194 800 4 la_data_in_mprj[106]
port 139 nsew
rlabel metal2 s 102598 -400 102654 800 4 la_data_in_mprj[107]
port 140 nsew
rlabel metal2 s 102966 -400 103022 800 4 la_data_in_mprj[108]
port 141 nsew
rlabel metal2 s 103426 -400 103482 800 4 la_data_in_mprj[109]
port 142 nsew
rlabel metal2 s 60278 -400 60334 800 4 la_data_in_mprj[10]
port 143 nsew
rlabel metal2 s 103886 -400 103942 800 4 la_data_in_mprj[110]
port 144 nsew
rlabel metal2 s 104254 -400 104310 800 4 la_data_in_mprj[111]
port 145 nsew
rlabel metal2 s 104714 -400 104770 800 4 la_data_in_mprj[112]
port 146 nsew
rlabel metal2 s 105174 -400 105230 800 4 la_data_in_mprj[113]
port 147 nsew
rlabel metal2 s 105634 -400 105690 800 4 la_data_in_mprj[114]
port 148 nsew
rlabel metal2 s 106002 -400 106058 800 4 la_data_in_mprj[115]
port 149 nsew
rlabel metal2 s 106462 -400 106518 800 4 la_data_in_mprj[116]
port 150 nsew
rlabel metal2 s 106922 -400 106978 800 4 la_data_in_mprj[117]
port 151 nsew
rlabel metal2 s 107382 -400 107438 800 4 la_data_in_mprj[118]
port 152 nsew
rlabel metal2 s 107750 -400 107806 800 4 la_data_in_mprj[119]
port 153 nsew
rlabel metal2 s 60738 -400 60794 800 4 la_data_in_mprj[11]
port 154 nsew
rlabel metal2 s 108210 -400 108266 800 4 la_data_in_mprj[120]
port 155 nsew
rlabel metal2 s 108670 -400 108726 800 4 la_data_in_mprj[121]
port 156 nsew
rlabel metal2 s 109130 -400 109186 800 4 la_data_in_mprj[122]
port 157 nsew
rlabel metal2 s 109498 -400 109554 800 4 la_data_in_mprj[123]
port 158 nsew
rlabel metal2 s 109958 -400 110014 800 4 la_data_in_mprj[124]
port 159 nsew
rlabel metal2 s 110418 -400 110474 800 4 la_data_in_mprj[125]
port 160 nsew
rlabel metal2 s 110878 -400 110934 800 4 la_data_in_mprj[126]
port 161 nsew
rlabel metal2 s 111246 -400 111302 800 4 la_data_in_mprj[127]
port 162 nsew
rlabel metal2 s 61198 -400 61254 800 4 la_data_in_mprj[12]
port 163 nsew
rlabel metal2 s 61566 -400 61622 800 4 la_data_in_mprj[13]
port 164 nsew
rlabel metal2 s 62026 -400 62082 800 4 la_data_in_mprj[14]
port 165 nsew
rlabel metal2 s 62486 -400 62542 800 4 la_data_in_mprj[15]
port 166 nsew
rlabel metal2 s 62946 -400 63002 800 4 la_data_in_mprj[16]
port 167 nsew
rlabel metal2 s 63314 -400 63370 800 4 la_data_in_mprj[17]
port 168 nsew
rlabel metal2 s 63774 -400 63830 800 4 la_data_in_mprj[18]
port 169 nsew
rlabel metal2 s 64234 -400 64290 800 4 la_data_in_mprj[19]
port 170 nsew
rlabel metal2 s 56322 -400 56378 800 4 la_data_in_mprj[1]
port 171 nsew
rlabel metal2 s 64602 -400 64658 800 4 la_data_in_mprj[20]
port 172 nsew
rlabel metal2 s 65062 -400 65118 800 4 la_data_in_mprj[21]
port 173 nsew
rlabel metal2 s 65522 -400 65578 800 4 la_data_in_mprj[22]
port 174 nsew
rlabel metal2 s 65982 -400 66038 800 4 la_data_in_mprj[23]
port 175 nsew
rlabel metal2 s 66350 -400 66406 800 4 la_data_in_mprj[24]
port 176 nsew
rlabel metal2 s 66810 -400 66866 800 4 la_data_in_mprj[25]
port 177 nsew
rlabel metal2 s 67270 -400 67326 800 4 la_data_in_mprj[26]
port 178 nsew
rlabel metal2 s 67730 -400 67786 800 4 la_data_in_mprj[27]
port 179 nsew
rlabel metal2 s 68098 -400 68154 800 4 la_data_in_mprj[28]
port 180 nsew
rlabel metal2 s 68558 -400 68614 800 4 la_data_in_mprj[29]
port 181 nsew
rlabel metal2 s 56782 -400 56838 800 4 la_data_in_mprj[2]
port 182 nsew
rlabel metal2 s 69018 -400 69074 800 4 la_data_in_mprj[30]
port 183 nsew
rlabel metal2 s 69478 -400 69534 800 4 la_data_in_mprj[31]
port 184 nsew
rlabel metal2 s 69846 -400 69902 800 4 la_data_in_mprj[32]
port 185 nsew
rlabel metal2 s 70306 -400 70362 800 4 la_data_in_mprj[33]
port 186 nsew
rlabel metal2 s 70766 -400 70822 800 4 la_data_in_mprj[34]
port 187 nsew
rlabel metal2 s 71226 -400 71282 800 4 la_data_in_mprj[35]
port 188 nsew
rlabel metal2 s 71594 -400 71650 800 4 la_data_in_mprj[36]
port 189 nsew
rlabel metal2 s 72054 -400 72110 800 4 la_data_in_mprj[37]
port 190 nsew
rlabel metal2 s 72514 -400 72570 800 4 la_data_in_mprj[38]
port 191 nsew
rlabel metal2 s 72882 -400 72938 800 4 la_data_in_mprj[39]
port 192 nsew
rlabel metal2 s 57242 -400 57298 800 4 la_data_in_mprj[3]
port 193 nsew
rlabel metal2 s 73342 -400 73398 800 4 la_data_in_mprj[40]
port 194 nsew
rlabel metal2 s 73802 -400 73858 800 4 la_data_in_mprj[41]
port 195 nsew
rlabel metal2 s 74262 -400 74318 800 4 la_data_in_mprj[42]
port 196 nsew
rlabel metal2 s 74630 -400 74686 800 4 la_data_in_mprj[43]
port 197 nsew
rlabel metal2 s 75090 -400 75146 800 4 la_data_in_mprj[44]
port 198 nsew
rlabel metal2 s 75550 -400 75606 800 4 la_data_in_mprj[45]
port 199 nsew
rlabel metal2 s 76010 -400 76066 800 4 la_data_in_mprj[46]
port 200 nsew
rlabel metal2 s 76378 -400 76434 800 4 la_data_in_mprj[47]
port 201 nsew
rlabel metal2 s 76838 -400 76894 800 4 la_data_in_mprj[48]
port 202 nsew
rlabel metal2 s 77298 -400 77354 800 4 la_data_in_mprj[49]
port 203 nsew
rlabel metal2 s 57702 -400 57758 800 4 la_data_in_mprj[4]
port 204 nsew
rlabel metal2 s 77758 -400 77814 800 4 la_data_in_mprj[50]
port 205 nsew
rlabel metal2 s 78126 -400 78182 800 4 la_data_in_mprj[51]
port 206 nsew
rlabel metal2 s 78586 -400 78642 800 4 la_data_in_mprj[52]
port 207 nsew
rlabel metal2 s 79046 -400 79102 800 4 la_data_in_mprj[53]
port 208 nsew
rlabel metal2 s 79506 -400 79562 800 4 la_data_in_mprj[54]
port 209 nsew
rlabel metal2 s 79874 -400 79930 800 4 la_data_in_mprj[55]
port 210 nsew
rlabel metal2 s 80334 -400 80390 800 4 la_data_in_mprj[56]
port 211 nsew
rlabel metal2 s 80794 -400 80850 800 4 la_data_in_mprj[57]
port 212 nsew
rlabel metal2 s 81162 -400 81218 800 4 la_data_in_mprj[58]
port 213 nsew
rlabel metal2 s 81622 -400 81678 800 4 la_data_in_mprj[59]
port 214 nsew
rlabel metal2 s 58070 -400 58126 800 4 la_data_in_mprj[5]
port 215 nsew
rlabel metal2 s 82082 -400 82138 800 4 la_data_in_mprj[60]
port 216 nsew
rlabel metal2 s 82542 -400 82598 800 4 la_data_in_mprj[61]
port 217 nsew
rlabel metal2 s 82910 -400 82966 800 4 la_data_in_mprj[62]
port 218 nsew
rlabel metal2 s 83370 -400 83426 800 4 la_data_in_mprj[63]
port 219 nsew
rlabel metal2 s 83830 -400 83886 800 4 la_data_in_mprj[64]
port 220 nsew
rlabel metal2 s 84290 -400 84346 800 4 la_data_in_mprj[65]
port 221 nsew
rlabel metal2 s 84658 -400 84714 800 4 la_data_in_mprj[66]
port 222 nsew
rlabel metal2 s 85118 -400 85174 800 4 la_data_in_mprj[67]
port 223 nsew
rlabel metal2 s 85578 -400 85634 800 4 la_data_in_mprj[68]
port 224 nsew
rlabel metal2 s 86038 -400 86094 800 4 la_data_in_mprj[69]
port 225 nsew
rlabel metal2 s 58530 -400 58586 800 4 la_data_in_mprj[6]
port 226 nsew
rlabel metal2 s 86406 -400 86462 800 4 la_data_in_mprj[70]
port 227 nsew
rlabel metal2 s 86866 -400 86922 800 4 la_data_in_mprj[71]
port 228 nsew
rlabel metal2 s 87326 -400 87382 800 4 la_data_in_mprj[72]
port 229 nsew
rlabel metal2 s 87786 -400 87842 800 4 la_data_in_mprj[73]
port 230 nsew
rlabel metal2 s 88154 -400 88210 800 4 la_data_in_mprj[74]
port 231 nsew
rlabel metal2 s 88614 -400 88670 800 4 la_data_in_mprj[75]
port 232 nsew
rlabel metal2 s 89074 -400 89130 800 4 la_data_in_mprj[76]
port 233 nsew
rlabel metal2 s 89442 -400 89498 800 4 la_data_in_mprj[77]
port 234 nsew
rlabel metal2 s 89902 -400 89958 800 4 la_data_in_mprj[78]
port 235 nsew
rlabel metal2 s 90362 -400 90418 800 4 la_data_in_mprj[79]
port 236 nsew
rlabel metal2 s 58990 -400 59046 800 4 la_data_in_mprj[7]
port 237 nsew
rlabel metal2 s 90822 -400 90878 800 4 la_data_in_mprj[80]
port 238 nsew
rlabel metal2 s 91190 -400 91246 800 4 la_data_in_mprj[81]
port 239 nsew
rlabel metal2 s 91650 -400 91706 800 4 la_data_in_mprj[82]
port 240 nsew
rlabel metal2 s 92110 -400 92166 800 4 la_data_in_mprj[83]
port 241 nsew
rlabel metal2 s 92570 -400 92626 800 4 la_data_in_mprj[84]
port 242 nsew
rlabel metal2 s 92938 -400 92994 800 4 la_data_in_mprj[85]
port 243 nsew
rlabel metal2 s 93398 -400 93454 800 4 la_data_in_mprj[86]
port 244 nsew
rlabel metal2 s 93858 -400 93914 800 4 la_data_in_mprj[87]
port 245 nsew
rlabel metal2 s 94318 -400 94374 800 4 la_data_in_mprj[88]
port 246 nsew
rlabel metal2 s 94686 -400 94742 800 4 la_data_in_mprj[89]
port 247 nsew
rlabel metal2 s 59450 -400 59506 800 4 la_data_in_mprj[8]
port 248 nsew
rlabel metal2 s 95146 -400 95202 800 4 la_data_in_mprj[90]
port 249 nsew
rlabel metal2 s 95606 -400 95662 800 4 la_data_in_mprj[91]
port 250 nsew
rlabel metal2 s 96066 -400 96122 800 4 la_data_in_mprj[92]
port 251 nsew
rlabel metal2 s 96434 -400 96490 800 4 la_data_in_mprj[93]
port 252 nsew
rlabel metal2 s 96894 -400 96950 800 4 la_data_in_mprj[94]
port 253 nsew
rlabel metal2 s 97354 -400 97410 800 4 la_data_in_mprj[95]
port 254 nsew
rlabel metal2 s 97722 -400 97778 800 4 la_data_in_mprj[96]
port 255 nsew
rlabel metal2 s 98182 -400 98238 800 4 la_data_in_mprj[97]
port 256 nsew
rlabel metal2 s 98642 -400 98698 800 4 la_data_in_mprj[98]
port 257 nsew
rlabel metal2 s 99102 -400 99158 800 4 la_data_in_mprj[99]
port 258 nsew
rlabel metal2 s 59818 -400 59874 800 4 la_data_in_mprj[9]
port 259 nsew
rlabel metal2 s 57702 10200 57758 11400 4 la_data_out_core[0]
port 260 nsew
rlabel metal2 s 101218 10200 101274 11400 4 la_data_out_core[100]
port 261 nsew
rlabel metal2 s 101678 10200 101734 11400 4 la_data_out_core[101]
port 262 nsew
rlabel metal2 s 102138 10200 102194 11400 4 la_data_out_core[102]
port 263 nsew
rlabel metal2 s 102598 10200 102654 11400 4 la_data_out_core[103]
port 264 nsew
rlabel metal2 s 102966 10200 103022 11400 4 la_data_out_core[104]
port 265 nsew
rlabel metal2 s 103426 10200 103482 11400 4 la_data_out_core[105]
port 266 nsew
rlabel metal2 s 103886 10200 103942 11400 4 la_data_out_core[106]
port 267 nsew
rlabel metal2 s 104254 10200 104310 11400 4 la_data_out_core[107]
port 268 nsew
rlabel metal2 s 104714 10200 104770 11400 4 la_data_out_core[108]
port 269 nsew
rlabel metal2 s 105174 10200 105230 11400 4 la_data_out_core[109]
port 270 nsew
rlabel metal2 s 62026 10200 62082 11400 4 la_data_out_core[10]
port 271 nsew
rlabel metal2 s 105634 10200 105690 11400 4 la_data_out_core[110]
port 272 nsew
rlabel metal2 s 106002 10200 106058 11400 4 la_data_out_core[111]
port 273 nsew
rlabel metal2 s 106462 10200 106518 11400 4 la_data_out_core[112]
port 274 nsew
rlabel metal2 s 106922 10200 106978 11400 4 la_data_out_core[113]
port 275 nsew
rlabel metal2 s 107382 10200 107438 11400 4 la_data_out_core[114]
port 276 nsew
rlabel metal2 s 107750 10200 107806 11400 4 la_data_out_core[115]
port 277 nsew
rlabel metal2 s 108210 10200 108266 11400 4 la_data_out_core[116]
port 278 nsew
rlabel metal2 s 108670 10200 108726 11400 4 la_data_out_core[117]
port 279 nsew
rlabel metal2 s 109130 10200 109186 11400 4 la_data_out_core[118]
port 280 nsew
rlabel metal2 s 109498 10200 109554 11400 4 la_data_out_core[119]
port 281 nsew
rlabel metal2 s 62486 10200 62542 11400 4 la_data_out_core[11]
port 282 nsew
rlabel metal2 s 109958 10200 110014 11400 4 la_data_out_core[120]
port 283 nsew
rlabel metal2 s 110418 10200 110474 11400 4 la_data_out_core[121]
port 284 nsew
rlabel metal2 s 110878 10200 110934 11400 4 la_data_out_core[122]
port 285 nsew
rlabel metal2 s 111246 10200 111302 11400 4 la_data_out_core[123]
port 286 nsew
rlabel metal2 s 111706 10200 111762 11400 4 la_data_out_core[124]
port 287 nsew
rlabel metal2 s 112166 10200 112222 11400 4 la_data_out_core[125]
port 288 nsew
rlabel metal2 s 112534 10200 112590 11400 4 la_data_out_core[126]
port 289 nsew
rlabel metal2 s 112994 10200 113050 11400 4 la_data_out_core[127]
port 290 nsew
rlabel metal2 s 62946 10200 63002 11400 4 la_data_out_core[12]
port 291 nsew
rlabel metal2 s 63314 10200 63370 11400 4 la_data_out_core[13]
port 292 nsew
rlabel metal2 s 63774 10200 63830 11400 4 la_data_out_core[14]
port 293 nsew
rlabel metal2 s 64234 10200 64290 11400 4 la_data_out_core[15]
port 294 nsew
rlabel metal2 s 64602 10200 64658 11400 4 la_data_out_core[16]
port 295 nsew
rlabel metal2 s 65062 10200 65118 11400 4 la_data_out_core[17]
port 296 nsew
rlabel metal2 s 65522 10200 65578 11400 4 la_data_out_core[18]
port 297 nsew
rlabel metal2 s 65982 10200 66038 11400 4 la_data_out_core[19]
port 298 nsew
rlabel metal2 s 58070 10200 58126 11400 4 la_data_out_core[1]
port 299 nsew
rlabel metal2 s 66350 10200 66406 11400 4 la_data_out_core[20]
port 300 nsew
rlabel metal2 s 66810 10200 66866 11400 4 la_data_out_core[21]
port 301 nsew
rlabel metal2 s 67270 10200 67326 11400 4 la_data_out_core[22]
port 302 nsew
rlabel metal2 s 67730 10200 67786 11400 4 la_data_out_core[23]
port 303 nsew
rlabel metal2 s 68098 10200 68154 11400 4 la_data_out_core[24]
port 304 nsew
rlabel metal2 s 68558 10200 68614 11400 4 la_data_out_core[25]
port 305 nsew
rlabel metal2 s 69018 10200 69074 11400 4 la_data_out_core[26]
port 306 nsew
rlabel metal2 s 69478 10200 69534 11400 4 la_data_out_core[27]
port 307 nsew
rlabel metal2 s 69846 10200 69902 11400 4 la_data_out_core[28]
port 308 nsew
rlabel metal2 s 70306 10200 70362 11400 4 la_data_out_core[29]
port 309 nsew
rlabel metal2 s 58530 10200 58586 11400 4 la_data_out_core[2]
port 310 nsew
rlabel metal2 s 70766 10200 70822 11400 4 la_data_out_core[30]
port 311 nsew
rlabel metal2 s 71226 10200 71282 11400 4 la_data_out_core[31]
port 312 nsew
rlabel metal2 s 71594 10200 71650 11400 4 la_data_out_core[32]
port 313 nsew
rlabel metal2 s 72054 10200 72110 11400 4 la_data_out_core[33]
port 314 nsew
rlabel metal2 s 72514 10200 72570 11400 4 la_data_out_core[34]
port 315 nsew
rlabel metal2 s 72882 10200 72938 11400 4 la_data_out_core[35]
port 316 nsew
rlabel metal2 s 73342 10200 73398 11400 4 la_data_out_core[36]
port 317 nsew
rlabel metal2 s 73802 10200 73858 11400 4 la_data_out_core[37]
port 318 nsew
rlabel metal2 s 74262 10200 74318 11400 4 la_data_out_core[38]
port 319 nsew
rlabel metal2 s 74630 10200 74686 11400 4 la_data_out_core[39]
port 320 nsew
rlabel metal2 s 58990 10200 59046 11400 4 la_data_out_core[3]
port 321 nsew
rlabel metal2 s 75090 10200 75146 11400 4 la_data_out_core[40]
port 322 nsew
rlabel metal2 s 75550 10200 75606 11400 4 la_data_out_core[41]
port 323 nsew
rlabel metal2 s 76010 10200 76066 11400 4 la_data_out_core[42]
port 324 nsew
rlabel metal2 s 76378 10200 76434 11400 4 la_data_out_core[43]
port 325 nsew
rlabel metal2 s 76838 10200 76894 11400 4 la_data_out_core[44]
port 326 nsew
rlabel metal2 s 77298 10200 77354 11400 4 la_data_out_core[45]
port 327 nsew
rlabel metal2 s 77758 10200 77814 11400 4 la_data_out_core[46]
port 328 nsew
rlabel metal2 s 78126 10200 78182 11400 4 la_data_out_core[47]
port 329 nsew
rlabel metal2 s 78586 10200 78642 11400 4 la_data_out_core[48]
port 330 nsew
rlabel metal2 s 79046 10200 79102 11400 4 la_data_out_core[49]
port 331 nsew
rlabel metal2 s 59450 10200 59506 11400 4 la_data_out_core[4]
port 332 nsew
rlabel metal2 s 79506 10200 79562 11400 4 la_data_out_core[50]
port 333 nsew
rlabel metal2 s 79874 10200 79930 11400 4 la_data_out_core[51]
port 334 nsew
rlabel metal2 s 80334 10200 80390 11400 4 la_data_out_core[52]
port 335 nsew
rlabel metal2 s 80794 10200 80850 11400 4 la_data_out_core[53]
port 336 nsew
rlabel metal2 s 81162 10200 81218 11400 4 la_data_out_core[54]
port 337 nsew
rlabel metal2 s 81622 10200 81678 11400 4 la_data_out_core[55]
port 338 nsew
rlabel metal2 s 82082 10200 82138 11400 4 la_data_out_core[56]
port 339 nsew
rlabel metal2 s 82542 10200 82598 11400 4 la_data_out_core[57]
port 340 nsew
rlabel metal2 s 82910 10200 82966 11400 4 la_data_out_core[58]
port 341 nsew
rlabel metal2 s 83370 10200 83426 11400 4 la_data_out_core[59]
port 342 nsew
rlabel metal2 s 59818 10200 59874 11400 4 la_data_out_core[5]
port 343 nsew
rlabel metal2 s 83830 10200 83886 11400 4 la_data_out_core[60]
port 344 nsew
rlabel metal2 s 84290 10200 84346 11400 4 la_data_out_core[61]
port 345 nsew
rlabel metal2 s 84658 10200 84714 11400 4 la_data_out_core[62]
port 346 nsew
rlabel metal2 s 85118 10200 85174 11400 4 la_data_out_core[63]
port 347 nsew
rlabel metal2 s 85578 10200 85634 11400 4 la_data_out_core[64]
port 348 nsew
rlabel metal2 s 86038 10200 86094 11400 4 la_data_out_core[65]
port 349 nsew
rlabel metal2 s 86406 10200 86462 11400 4 la_data_out_core[66]
port 350 nsew
rlabel metal2 s 86866 10200 86922 11400 4 la_data_out_core[67]
port 351 nsew
rlabel metal2 s 87326 10200 87382 11400 4 la_data_out_core[68]
port 352 nsew
rlabel metal2 s 87786 10200 87842 11400 4 la_data_out_core[69]
port 353 nsew
rlabel metal2 s 60278 10200 60334 11400 4 la_data_out_core[6]
port 354 nsew
rlabel metal2 s 88154 10200 88210 11400 4 la_data_out_core[70]
port 355 nsew
rlabel metal2 s 88614 10200 88670 11400 4 la_data_out_core[71]
port 356 nsew
rlabel metal2 s 89074 10200 89130 11400 4 la_data_out_core[72]
port 357 nsew
rlabel metal2 s 89442 10200 89498 11400 4 la_data_out_core[73]
port 358 nsew
rlabel metal2 s 89902 10200 89958 11400 4 la_data_out_core[74]
port 359 nsew
rlabel metal2 s 90362 10200 90418 11400 4 la_data_out_core[75]
port 360 nsew
rlabel metal2 s 90822 10200 90878 11400 4 la_data_out_core[76]
port 361 nsew
rlabel metal2 s 91190 10200 91246 11400 4 la_data_out_core[77]
port 362 nsew
rlabel metal2 s 91650 10200 91706 11400 4 la_data_out_core[78]
port 363 nsew
rlabel metal2 s 92110 10200 92166 11400 4 la_data_out_core[79]
port 364 nsew
rlabel metal2 s 60738 10200 60794 11400 4 la_data_out_core[7]
port 365 nsew
rlabel metal2 s 92570 10200 92626 11400 4 la_data_out_core[80]
port 366 nsew
rlabel metal2 s 92938 10200 92994 11400 4 la_data_out_core[81]
port 367 nsew
rlabel metal2 s 93398 10200 93454 11400 4 la_data_out_core[82]
port 368 nsew
rlabel metal2 s 93858 10200 93914 11400 4 la_data_out_core[83]
port 369 nsew
rlabel metal2 s 94318 10200 94374 11400 4 la_data_out_core[84]
port 370 nsew
rlabel metal2 s 94686 10200 94742 11400 4 la_data_out_core[85]
port 371 nsew
rlabel metal2 s 95146 10200 95202 11400 4 la_data_out_core[86]
port 372 nsew
rlabel metal2 s 95606 10200 95662 11400 4 la_data_out_core[87]
port 373 nsew
rlabel metal2 s 96066 10200 96122 11400 4 la_data_out_core[88]
port 374 nsew
rlabel metal2 s 96434 10200 96490 11400 4 la_data_out_core[89]
port 375 nsew
rlabel metal2 s 61198 10200 61254 11400 4 la_data_out_core[8]
port 376 nsew
rlabel metal2 s 96894 10200 96950 11400 4 la_data_out_core[90]
port 377 nsew
rlabel metal2 s 97354 10200 97410 11400 4 la_data_out_core[91]
port 378 nsew
rlabel metal2 s 97722 10200 97778 11400 4 la_data_out_core[92]
port 379 nsew
rlabel metal2 s 98182 10200 98238 11400 4 la_data_out_core[93]
port 380 nsew
rlabel metal2 s 98642 10200 98698 11400 4 la_data_out_core[94]
port 381 nsew
rlabel metal2 s 99102 10200 99158 11400 4 la_data_out_core[95]
port 382 nsew
rlabel metal2 s 99470 10200 99526 11400 4 la_data_out_core[96]
port 383 nsew
rlabel metal2 s 99930 10200 99986 11400 4 la_data_out_core[97]
port 384 nsew
rlabel metal2 s 100390 10200 100446 11400 4 la_data_out_core[98]
port 385 nsew
rlabel metal2 s 100850 10200 100906 11400 4 la_data_out_core[99]
port 386 nsew
rlabel metal2 s 61566 10200 61622 11400 4 la_data_out_core[9]
port 387 nsew
rlabel metal2 s 202 -400 258 800 4 la_data_out_mprj[0]
port 388 nsew
rlabel metal2 s 43718 -400 43774 800 4 la_data_out_mprj[100]
port 389 nsew
rlabel metal2 s 44178 -400 44234 800 4 la_data_out_mprj[101]
port 390 nsew
rlabel metal2 s 44638 -400 44694 800 4 la_data_out_mprj[102]
port 391 nsew
rlabel metal2 s 45006 -400 45062 800 4 la_data_out_mprj[103]
port 392 nsew
rlabel metal2 s 45466 -400 45522 800 4 la_data_out_mprj[104]
port 393 nsew
rlabel metal2 s 45926 -400 45982 800 4 la_data_out_mprj[105]
port 394 nsew
rlabel metal2 s 46386 -400 46442 800 4 la_data_out_mprj[106]
port 395 nsew
rlabel metal2 s 46754 -400 46810 800 4 la_data_out_mprj[107]
port 396 nsew
rlabel metal2 s 47214 -400 47270 800 4 la_data_out_mprj[108]
port 397 nsew
rlabel metal2 s 47674 -400 47730 800 4 la_data_out_mprj[109]
port 398 nsew
rlabel metal2 s 4526 -400 4582 800 4 la_data_out_mprj[10]
port 399 nsew
rlabel metal2 s 48134 -400 48190 800 4 la_data_out_mprj[110]
port 400 nsew
rlabel metal2 s 48502 -400 48558 800 4 la_data_out_mprj[111]
port 401 nsew
rlabel metal2 s 48962 -400 49018 800 4 la_data_out_mprj[112]
port 402 nsew
rlabel metal2 s 49422 -400 49478 800 4 la_data_out_mprj[113]
port 403 nsew
rlabel metal2 s 49790 -400 49846 800 4 la_data_out_mprj[114]
port 404 nsew
rlabel metal2 s 50250 -400 50306 800 4 la_data_out_mprj[115]
port 405 nsew
rlabel metal2 s 50710 -400 50766 800 4 la_data_out_mprj[116]
port 406 nsew
rlabel metal2 s 51170 -400 51226 800 4 la_data_out_mprj[117]
port 407 nsew
rlabel metal2 s 51538 -400 51594 800 4 la_data_out_mprj[118]
port 408 nsew
rlabel metal2 s 51998 -400 52054 800 4 la_data_out_mprj[119]
port 409 nsew
rlabel metal2 s 4986 -400 5042 800 4 la_data_out_mprj[11]
port 410 nsew
rlabel metal2 s 52458 -400 52514 800 4 la_data_out_mprj[120]
port 411 nsew
rlabel metal2 s 52918 -400 52974 800 4 la_data_out_mprj[121]
port 412 nsew
rlabel metal2 s 53286 -400 53342 800 4 la_data_out_mprj[122]
port 413 nsew
rlabel metal2 s 53746 -400 53802 800 4 la_data_out_mprj[123]
port 414 nsew
rlabel metal2 s 54206 -400 54262 800 4 la_data_out_mprj[124]
port 415 nsew
rlabel metal2 s 54666 -400 54722 800 4 la_data_out_mprj[125]
port 416 nsew
rlabel metal2 s 55034 -400 55090 800 4 la_data_out_mprj[126]
port 417 nsew
rlabel metal2 s 55494 -400 55550 800 4 la_data_out_mprj[127]
port 418 nsew
rlabel metal2 s 5354 -400 5410 800 4 la_data_out_mprj[12]
port 419 nsew
rlabel metal2 s 5814 -400 5870 800 4 la_data_out_mprj[13]
port 420 nsew
rlabel metal2 s 6274 -400 6330 800 4 la_data_out_mprj[14]
port 421 nsew
rlabel metal2 s 6734 -400 6790 800 4 la_data_out_mprj[15]
port 422 nsew
rlabel metal2 s 7102 -400 7158 800 4 la_data_out_mprj[16]
port 423 nsew
rlabel metal2 s 7562 -400 7618 800 4 la_data_out_mprj[17]
port 424 nsew
rlabel metal2 s 8022 -400 8078 800 4 la_data_out_mprj[18]
port 425 nsew
rlabel metal2 s 8390 -400 8446 800 4 la_data_out_mprj[19]
port 426 nsew
rlabel metal2 s 570 -400 626 800 4 la_data_out_mprj[1]
port 427 nsew
rlabel metal2 s 8850 -400 8906 800 4 la_data_out_mprj[20]
port 428 nsew
rlabel metal2 s 9310 -400 9366 800 4 la_data_out_mprj[21]
port 429 nsew
rlabel metal2 s 9770 -400 9826 800 4 la_data_out_mprj[22]
port 430 nsew
rlabel metal2 s 10138 -400 10194 800 4 la_data_out_mprj[23]
port 431 nsew
rlabel metal2 s 10598 -400 10654 800 4 la_data_out_mprj[24]
port 432 nsew
rlabel metal2 s 11058 -400 11114 800 4 la_data_out_mprj[25]
port 433 nsew
rlabel metal2 s 11518 -400 11574 800 4 la_data_out_mprj[26]
port 434 nsew
rlabel metal2 s 11886 -400 11942 800 4 la_data_out_mprj[27]
port 435 nsew
rlabel metal2 s 12346 -400 12402 800 4 la_data_out_mprj[28]
port 436 nsew
rlabel metal2 s 12806 -400 12862 800 4 la_data_out_mprj[29]
port 437 nsew
rlabel metal2 s 1030 -400 1086 800 4 la_data_out_mprj[2]
port 438 nsew
rlabel metal2 s 13266 -400 13322 800 4 la_data_out_mprj[30]
port 439 nsew
rlabel metal2 s 13634 -400 13690 800 4 la_data_out_mprj[31]
port 440 nsew
rlabel metal2 s 14094 -400 14150 800 4 la_data_out_mprj[32]
port 441 nsew
rlabel metal2 s 14554 -400 14610 800 4 la_data_out_mprj[33]
port 442 nsew
rlabel metal2 s 15014 -400 15070 800 4 la_data_out_mprj[34]
port 443 nsew
rlabel metal2 s 15382 -400 15438 800 4 la_data_out_mprj[35]
port 444 nsew
rlabel metal2 s 15842 -400 15898 800 4 la_data_out_mprj[36]
port 445 nsew
rlabel metal2 s 16302 -400 16358 800 4 la_data_out_mprj[37]
port 446 nsew
rlabel metal2 s 16670 -400 16726 800 4 la_data_out_mprj[38]
port 447 nsew
rlabel metal2 s 17130 -400 17186 800 4 la_data_out_mprj[39]
port 448 nsew
rlabel metal2 s 1490 -400 1546 800 4 la_data_out_mprj[3]
port 449 nsew
rlabel metal2 s 17590 -400 17646 800 4 la_data_out_mprj[40]
port 450 nsew
rlabel metal2 s 18050 -400 18106 800 4 la_data_out_mprj[41]
port 451 nsew
rlabel metal2 s 18418 -400 18474 800 4 la_data_out_mprj[42]
port 452 nsew
rlabel metal2 s 18878 -400 18934 800 4 la_data_out_mprj[43]
port 453 nsew
rlabel metal2 s 19338 -400 19394 800 4 la_data_out_mprj[44]
port 454 nsew
rlabel metal2 s 19798 -400 19854 800 4 la_data_out_mprj[45]
port 455 nsew
rlabel metal2 s 20166 -400 20222 800 4 la_data_out_mprj[46]
port 456 nsew
rlabel metal2 s 20626 -400 20682 800 4 la_data_out_mprj[47]
port 457 nsew
rlabel metal2 s 21086 -400 21142 800 4 la_data_out_mprj[48]
port 458 nsew
rlabel metal2 s 21546 -400 21602 800 4 la_data_out_mprj[49]
port 459 nsew
rlabel metal2 s 1858 -400 1914 800 4 la_data_out_mprj[4]
port 460 nsew
rlabel metal2 s 21914 -400 21970 800 4 la_data_out_mprj[50]
port 461 nsew
rlabel metal2 s 22374 -400 22430 800 4 la_data_out_mprj[51]
port 462 nsew
rlabel metal2 s 22834 -400 22890 800 4 la_data_out_mprj[52]
port 463 nsew
rlabel metal2 s 23294 -400 23350 800 4 la_data_out_mprj[53]
port 464 nsew
rlabel metal2 s 23662 -400 23718 800 4 la_data_out_mprj[54]
port 465 nsew
rlabel metal2 s 24122 -400 24178 800 4 la_data_out_mprj[55]
port 466 nsew
rlabel metal2 s 24582 -400 24638 800 4 la_data_out_mprj[56]
port 467 nsew
rlabel metal2 s 24950 -400 25006 800 4 la_data_out_mprj[57]
port 468 nsew
rlabel metal2 s 25410 -400 25466 800 4 la_data_out_mprj[58]
port 469 nsew
rlabel metal2 s 25870 -400 25926 800 4 la_data_out_mprj[59]
port 470 nsew
rlabel metal2 s 2318 -400 2374 800 4 la_data_out_mprj[5]
port 471 nsew
rlabel metal2 s 26330 -400 26386 800 4 la_data_out_mprj[60]
port 472 nsew
rlabel metal2 s 26698 -400 26754 800 4 la_data_out_mprj[61]
port 473 nsew
rlabel metal2 s 27158 -400 27214 800 4 la_data_out_mprj[62]
port 474 nsew
rlabel metal2 s 27618 -400 27674 800 4 la_data_out_mprj[63]
port 475 nsew
rlabel metal2 s 28078 -400 28134 800 4 la_data_out_mprj[64]
port 476 nsew
rlabel metal2 s 28446 -400 28502 800 4 la_data_out_mprj[65]
port 477 nsew
rlabel metal2 s 28906 -400 28962 800 4 la_data_out_mprj[66]
port 478 nsew
rlabel metal2 s 29366 -400 29422 800 4 la_data_out_mprj[67]
port 479 nsew
rlabel metal2 s 29826 -400 29882 800 4 la_data_out_mprj[68]
port 480 nsew
rlabel metal2 s 30194 -400 30250 800 4 la_data_out_mprj[69]
port 481 nsew
rlabel metal2 s 2778 -400 2834 800 4 la_data_out_mprj[6]
port 482 nsew
rlabel metal2 s 30654 -400 30710 800 4 la_data_out_mprj[70]
port 483 nsew
rlabel metal2 s 31114 -400 31170 800 4 la_data_out_mprj[71]
port 484 nsew
rlabel metal2 s 31574 -400 31630 800 4 la_data_out_mprj[72]
port 485 nsew
rlabel metal2 s 31942 -400 31998 800 4 la_data_out_mprj[73]
port 486 nsew
rlabel metal2 s 32402 -400 32458 800 4 la_data_out_mprj[74]
port 487 nsew
rlabel metal2 s 32862 -400 32918 800 4 la_data_out_mprj[75]
port 488 nsew
rlabel metal2 s 33230 -400 33286 800 4 la_data_out_mprj[76]
port 489 nsew
rlabel metal2 s 33690 -400 33746 800 4 la_data_out_mprj[77]
port 490 nsew
rlabel metal2 s 34150 -400 34206 800 4 la_data_out_mprj[78]
port 491 nsew
rlabel metal2 s 34610 -400 34666 800 4 la_data_out_mprj[79]
port 492 nsew
rlabel metal2 s 3238 -400 3294 800 4 la_data_out_mprj[7]
port 493 nsew
rlabel metal2 s 34978 -400 35034 800 4 la_data_out_mprj[80]
port 494 nsew
rlabel metal2 s 35438 -400 35494 800 4 la_data_out_mprj[81]
port 495 nsew
rlabel metal2 s 35898 -400 35954 800 4 la_data_out_mprj[82]
port 496 nsew
rlabel metal2 s 36358 -400 36414 800 4 la_data_out_mprj[83]
port 497 nsew
rlabel metal2 s 36726 -400 36782 800 4 la_data_out_mprj[84]
port 498 nsew
rlabel metal2 s 37186 -400 37242 800 4 la_data_out_mprj[85]
port 499 nsew
rlabel metal2 s 37646 -400 37702 800 4 la_data_out_mprj[86]
port 500 nsew
rlabel metal2 s 38106 -400 38162 800 4 la_data_out_mprj[87]
port 501 nsew
rlabel metal2 s 38474 -400 38530 800 4 la_data_out_mprj[88]
port 502 nsew
rlabel metal2 s 38934 -400 38990 800 4 la_data_out_mprj[89]
port 503 nsew
rlabel metal2 s 3606 -400 3662 800 4 la_data_out_mprj[8]
port 504 nsew
rlabel metal2 s 39394 -400 39450 800 4 la_data_out_mprj[90]
port 505 nsew
rlabel metal2 s 39854 -400 39910 800 4 la_data_out_mprj[91]
port 506 nsew
rlabel metal2 s 40222 -400 40278 800 4 la_data_out_mprj[92]
port 507 nsew
rlabel metal2 s 40682 -400 40738 800 4 la_data_out_mprj[93]
port 508 nsew
rlabel metal2 s 41142 -400 41198 800 4 la_data_out_mprj[94]
port 509 nsew
rlabel metal2 s 41510 -400 41566 800 4 la_data_out_mprj[95]
port 510 nsew
rlabel metal2 s 41970 -400 42026 800 4 la_data_out_mprj[96]
port 511 nsew
rlabel metal2 s 42430 -400 42486 800 4 la_data_out_mprj[97]
port 512 nsew
rlabel metal2 s 42890 -400 42946 800 4 la_data_out_mprj[98]
port 513 nsew
rlabel metal2 s 43258 -400 43314 800 4 la_data_out_mprj[99]
port 514 nsew
rlabel metal2 s 4066 -400 4122 800 4 la_data_out_mprj[9]
port 515 nsew
rlabel metal2 s 113454 10200 113510 11400 4 la_oen_core[0]
port 516 nsew
rlabel metal2 s 157062 10200 157118 11400 4 la_oen_core[100]
port 517 nsew
rlabel metal2 s 157430 10200 157486 11400 4 la_oen_core[101]
port 518 nsew
rlabel metal2 s 157890 10200 157946 11400 4 la_oen_core[102]
port 519 nsew
rlabel metal2 s 158350 10200 158406 11400 4 la_oen_core[103]
port 520 nsew
rlabel metal2 s 158810 10200 158866 11400 4 la_oen_core[104]
port 521 nsew
rlabel metal2 s 159178 10200 159234 11400 4 la_oen_core[105]
port 522 nsew
rlabel metal2 s 159638 10200 159694 11400 4 la_oen_core[106]
port 523 nsew
rlabel metal2 s 160098 10200 160154 11400 4 la_oen_core[107]
port 524 nsew
rlabel metal2 s 160466 10200 160522 11400 4 la_oen_core[108]
port 525 nsew
rlabel metal2 s 160926 10200 160982 11400 4 la_oen_core[109]
port 526 nsew
rlabel metal2 s 117778 10200 117834 11400 4 la_oen_core[10]
port 527 nsew
rlabel metal2 s 161386 10200 161442 11400 4 la_oen_core[110]
port 528 nsew
rlabel metal2 s 161846 10200 161902 11400 4 la_oen_core[111]
port 529 nsew
rlabel metal2 s 162214 10200 162270 11400 4 la_oen_core[112]
port 530 nsew
rlabel metal2 s 162674 10200 162730 11400 4 la_oen_core[113]
port 531 nsew
rlabel metal2 s 163134 10200 163190 11400 4 la_oen_core[114]
port 532 nsew
rlabel metal2 s 163594 10200 163650 11400 4 la_oen_core[115]
port 533 nsew
rlabel metal2 s 163962 10200 164018 11400 4 la_oen_core[116]
port 534 nsew
rlabel metal2 s 164422 10200 164478 11400 4 la_oen_core[117]
port 535 nsew
rlabel metal2 s 164882 10200 164938 11400 4 la_oen_core[118]
port 536 nsew
rlabel metal2 s 165342 10200 165398 11400 4 la_oen_core[119]
port 537 nsew
rlabel metal2 s 118238 10200 118294 11400 4 la_oen_core[11]
port 538 nsew
rlabel metal2 s 165710 10200 165766 11400 4 la_oen_core[120]
port 539 nsew
rlabel metal2 s 166170 10200 166226 11400 4 la_oen_core[121]
port 540 nsew
rlabel metal2 s 166630 10200 166686 11400 4 la_oen_core[122]
port 541 nsew
rlabel metal2 s 167090 10200 167146 11400 4 la_oen_core[123]
port 542 nsew
rlabel metal2 s 167458 10200 167514 11400 4 la_oen_core[124]
port 543 nsew
rlabel metal2 s 167918 10200 167974 11400 4 la_oen_core[125]
port 544 nsew
rlabel metal2 s 168378 10200 168434 11400 4 la_oen_core[126]
port 545 nsew
rlabel metal2 s 168746 10200 168802 11400 4 la_oen_core[127]
port 546 nsew
rlabel metal2 s 118698 10200 118754 11400 4 la_oen_core[12]
port 547 nsew
rlabel metal2 s 119158 10200 119214 11400 4 la_oen_core[13]
port 548 nsew
rlabel metal2 s 119526 10200 119582 11400 4 la_oen_core[14]
port 549 nsew
rlabel metal2 s 119986 10200 120042 11400 4 la_oen_core[15]
port 550 nsew
rlabel metal2 s 120446 10200 120502 11400 4 la_oen_core[16]
port 551 nsew
rlabel metal2 s 120814 10200 120870 11400 4 la_oen_core[17]
port 552 nsew
rlabel metal2 s 121274 10200 121330 11400 4 la_oen_core[18]
port 553 nsew
rlabel metal2 s 121734 10200 121790 11400 4 la_oen_core[19]
port 554 nsew
rlabel metal2 s 113914 10200 113970 11400 4 la_oen_core[1]
port 555 nsew
rlabel metal2 s 122194 10200 122250 11400 4 la_oen_core[20]
port 556 nsew
rlabel metal2 s 122562 10200 122618 11400 4 la_oen_core[21]
port 557 nsew
rlabel metal2 s 123022 10200 123078 11400 4 la_oen_core[22]
port 558 nsew
rlabel metal2 s 123482 10200 123538 11400 4 la_oen_core[23]
port 559 nsew
rlabel metal2 s 123942 10200 123998 11400 4 la_oen_core[24]
port 560 nsew
rlabel metal2 s 124310 10200 124366 11400 4 la_oen_core[25]
port 561 nsew
rlabel metal2 s 124770 10200 124826 11400 4 la_oen_core[26]
port 562 nsew
rlabel metal2 s 125230 10200 125286 11400 4 la_oen_core[27]
port 563 nsew
rlabel metal2 s 125690 10200 125746 11400 4 la_oen_core[28]
port 564 nsew
rlabel metal2 s 126058 10200 126114 11400 4 la_oen_core[29]
port 565 nsew
rlabel metal2 s 114282 10200 114338 11400 4 la_oen_core[2]
port 566 nsew
rlabel metal2 s 126518 10200 126574 11400 4 la_oen_core[30]
port 567 nsew
rlabel metal2 s 126978 10200 127034 11400 4 la_oen_core[31]
port 568 nsew
rlabel metal2 s 127438 10200 127494 11400 4 la_oen_core[32]
port 569 nsew
rlabel metal2 s 127806 10200 127862 11400 4 la_oen_core[33]
port 570 nsew
rlabel metal2 s 128266 10200 128322 11400 4 la_oen_core[34]
port 571 nsew
rlabel metal2 s 128726 10200 128782 11400 4 la_oen_core[35]
port 572 nsew
rlabel metal2 s 129094 10200 129150 11400 4 la_oen_core[36]
port 573 nsew
rlabel metal2 s 129554 10200 129610 11400 4 la_oen_core[37]
port 574 nsew
rlabel metal2 s 130014 10200 130070 11400 4 la_oen_core[38]
port 575 nsew
rlabel metal2 s 130474 10200 130530 11400 4 la_oen_core[39]
port 576 nsew
rlabel metal2 s 114742 10200 114798 11400 4 la_oen_core[3]
port 577 nsew
rlabel metal2 s 130842 10200 130898 11400 4 la_oen_core[40]
port 578 nsew
rlabel metal2 s 131302 10200 131358 11400 4 la_oen_core[41]
port 579 nsew
rlabel metal2 s 131762 10200 131818 11400 4 la_oen_core[42]
port 580 nsew
rlabel metal2 s 132222 10200 132278 11400 4 la_oen_core[43]
port 581 nsew
rlabel metal2 s 132590 10200 132646 11400 4 la_oen_core[44]
port 582 nsew
rlabel metal2 s 133050 10200 133106 11400 4 la_oen_core[45]
port 583 nsew
rlabel metal2 s 133510 10200 133566 11400 4 la_oen_core[46]
port 584 nsew
rlabel metal2 s 133970 10200 134026 11400 4 la_oen_core[47]
port 585 nsew
rlabel metal2 s 134338 10200 134394 11400 4 la_oen_core[48]
port 586 nsew
rlabel metal2 s 134798 10200 134854 11400 4 la_oen_core[49]
port 587 nsew
rlabel metal2 s 115202 10200 115258 11400 4 la_oen_core[4]
port 588 nsew
rlabel metal2 s 135258 10200 135314 11400 4 la_oen_core[50]
port 589 nsew
rlabel metal2 s 135718 10200 135774 11400 4 la_oen_core[51]
port 590 nsew
rlabel metal2 s 136086 10200 136142 11400 4 la_oen_core[52]
port 591 nsew
rlabel metal2 s 136546 10200 136602 11400 4 la_oen_core[53]
port 592 nsew
rlabel metal2 s 137006 10200 137062 11400 4 la_oen_core[54]
port 593 nsew
rlabel metal2 s 137374 10200 137430 11400 4 la_oen_core[55]
port 594 nsew
rlabel metal2 s 137834 10200 137890 11400 4 la_oen_core[56]
port 595 nsew
rlabel metal2 s 138294 10200 138350 11400 4 la_oen_core[57]
port 596 nsew
rlabel metal2 s 138754 10200 138810 11400 4 la_oen_core[58]
port 597 nsew
rlabel metal2 s 139122 10200 139178 11400 4 la_oen_core[59]
port 598 nsew
rlabel metal2 s 115662 10200 115718 11400 4 la_oen_core[5]
port 599 nsew
rlabel metal2 s 139582 10200 139638 11400 4 la_oen_core[60]
port 600 nsew
rlabel metal2 s 140042 10200 140098 11400 4 la_oen_core[61]
port 601 nsew
rlabel metal2 s 140502 10200 140558 11400 4 la_oen_core[62]
port 602 nsew
rlabel metal2 s 140870 10200 140926 11400 4 la_oen_core[63]
port 603 nsew
rlabel metal2 s 141330 10200 141386 11400 4 la_oen_core[64]
port 604 nsew
rlabel metal2 s 141790 10200 141846 11400 4 la_oen_core[65]
port 605 nsew
rlabel metal2 s 142250 10200 142306 11400 4 la_oen_core[66]
port 606 nsew
rlabel metal2 s 142618 10200 142674 11400 4 la_oen_core[67]
port 607 nsew
rlabel metal2 s 143078 10200 143134 11400 4 la_oen_core[68]
port 608 nsew
rlabel metal2 s 143538 10200 143594 11400 4 la_oen_core[69]
port 609 nsew
rlabel metal2 s 116030 10200 116086 11400 4 la_oen_core[6]
port 610 nsew
rlabel metal2 s 143998 10200 144054 11400 4 la_oen_core[70]
port 611 nsew
rlabel metal2 s 144366 10200 144422 11400 4 la_oen_core[71]
port 612 nsew
rlabel metal2 s 144826 10200 144882 11400 4 la_oen_core[72]
port 613 nsew
rlabel metal2 s 145286 10200 145342 11400 4 la_oen_core[73]
port 614 nsew
rlabel metal2 s 145654 10200 145710 11400 4 la_oen_core[74]
port 615 nsew
rlabel metal2 s 146114 10200 146170 11400 4 la_oen_core[75]
port 616 nsew
rlabel metal2 s 146574 10200 146630 11400 4 la_oen_core[76]
port 617 nsew
rlabel metal2 s 147034 10200 147090 11400 4 la_oen_core[77]
port 618 nsew
rlabel metal2 s 147402 10200 147458 11400 4 la_oen_core[78]
port 619 nsew
rlabel metal2 s 147862 10200 147918 11400 4 la_oen_core[79]
port 620 nsew
rlabel metal2 s 116490 10200 116546 11400 4 la_oen_core[7]
port 621 nsew
rlabel metal2 s 148322 10200 148378 11400 4 la_oen_core[80]
port 622 nsew
rlabel metal2 s 148782 10200 148838 11400 4 la_oen_core[81]
port 623 nsew
rlabel metal2 s 149150 10200 149206 11400 4 la_oen_core[82]
port 624 nsew
rlabel metal2 s 149610 10200 149666 11400 4 la_oen_core[83]
port 625 nsew
rlabel metal2 s 150070 10200 150126 11400 4 la_oen_core[84]
port 626 nsew
rlabel metal2 s 150530 10200 150586 11400 4 la_oen_core[85]
port 627 nsew
rlabel metal2 s 150898 10200 150954 11400 4 la_oen_core[86]
port 628 nsew
rlabel metal2 s 151358 10200 151414 11400 4 la_oen_core[87]
port 629 nsew
rlabel metal2 s 151818 10200 151874 11400 4 la_oen_core[88]
port 630 nsew
rlabel metal2 s 152186 10200 152242 11400 4 la_oen_core[89]
port 631 nsew
rlabel metal2 s 116950 10200 117006 11400 4 la_oen_core[8]
port 632 nsew
rlabel metal2 s 152646 10200 152702 11400 4 la_oen_core[90]
port 633 nsew
rlabel metal2 s 153106 10200 153162 11400 4 la_oen_core[91]
port 634 nsew
rlabel metal2 s 153566 10200 153622 11400 4 la_oen_core[92]
port 635 nsew
rlabel metal2 s 153934 10200 153990 11400 4 la_oen_core[93]
port 636 nsew
rlabel metal2 s 154394 10200 154450 11400 4 la_oen_core[94]
port 637 nsew
rlabel metal2 s 154854 10200 154910 11400 4 la_oen_core[95]
port 638 nsew
rlabel metal2 s 155314 10200 155370 11400 4 la_oen_core[96]
port 639 nsew
rlabel metal2 s 155682 10200 155738 11400 4 la_oen_core[97]
port 640 nsew
rlabel metal2 s 156142 10200 156198 11400 4 la_oen_core[98]
port 641 nsew
rlabel metal2 s 156602 10200 156658 11400 4 la_oen_core[99]
port 642 nsew
rlabel metal2 s 117410 10200 117466 11400 4 la_oen_core[9]
port 643 nsew
rlabel metal2 s 111706 -400 111762 800 4 la_oen_mprj[0]
port 644 nsew
rlabel metal2 s 155314 -400 155370 800 4 la_oen_mprj[100]
port 645 nsew
rlabel metal2 s 155682 -400 155738 800 4 la_oen_mprj[101]
port 646 nsew
rlabel metal2 s 156142 -400 156198 800 4 la_oen_mprj[102]
port 647 nsew
rlabel metal2 s 156602 -400 156658 800 4 la_oen_mprj[103]
port 648 nsew
rlabel metal2 s 157062 -400 157118 800 4 la_oen_mprj[104]
port 649 nsew
rlabel metal2 s 157430 -400 157486 800 4 la_oen_mprj[105]
port 650 nsew
rlabel metal2 s 157890 -400 157946 800 4 la_oen_mprj[106]
port 651 nsew
rlabel metal2 s 158350 -400 158406 800 4 la_oen_mprj[107]
port 652 nsew
rlabel metal2 s 158810 -400 158866 800 4 la_oen_mprj[108]
port 653 nsew
rlabel metal2 s 159178 -400 159234 800 4 la_oen_mprj[109]
port 654 nsew
rlabel metal2 s 116030 -400 116086 800 4 la_oen_mprj[10]
port 655 nsew
rlabel metal2 s 159638 -400 159694 800 4 la_oen_mprj[110]
port 656 nsew
rlabel metal2 s 160098 -400 160154 800 4 la_oen_mprj[111]
port 657 nsew
rlabel metal2 s 160466 -400 160522 800 4 la_oen_mprj[112]
port 658 nsew
rlabel metal2 s 160926 -400 160982 800 4 la_oen_mprj[113]
port 659 nsew
rlabel metal2 s 161386 -400 161442 800 4 la_oen_mprj[114]
port 660 nsew
rlabel metal2 s 161846 -400 161902 800 4 la_oen_mprj[115]
port 661 nsew
rlabel metal2 s 162214 -400 162270 800 4 la_oen_mprj[116]
port 662 nsew
rlabel metal2 s 162674 -400 162730 800 4 la_oen_mprj[117]
port 663 nsew
rlabel metal2 s 163134 -400 163190 800 4 la_oen_mprj[118]
port 664 nsew
rlabel metal2 s 163594 -400 163650 800 4 la_oen_mprj[119]
port 665 nsew
rlabel metal2 s 116490 -400 116546 800 4 la_oen_mprj[11]
port 666 nsew
rlabel metal2 s 163962 -400 164018 800 4 la_oen_mprj[120]
port 667 nsew
rlabel metal2 s 164422 -400 164478 800 4 la_oen_mprj[121]
port 668 nsew
rlabel metal2 s 164882 -400 164938 800 4 la_oen_mprj[122]
port 669 nsew
rlabel metal2 s 165342 -400 165398 800 4 la_oen_mprj[123]
port 670 nsew
rlabel metal2 s 165710 -400 165766 800 4 la_oen_mprj[124]
port 671 nsew
rlabel metal2 s 166170 -400 166226 800 4 la_oen_mprj[125]
port 672 nsew
rlabel metal2 s 166630 -400 166686 800 4 la_oen_mprj[126]
port 673 nsew
rlabel metal2 s 167090 -400 167146 800 4 la_oen_mprj[127]
port 674 nsew
rlabel metal2 s 116950 -400 117006 800 4 la_oen_mprj[12]
port 675 nsew
rlabel metal2 s 117410 -400 117466 800 4 la_oen_mprj[13]
port 676 nsew
rlabel metal2 s 117778 -400 117834 800 4 la_oen_mprj[14]
port 677 nsew
rlabel metal2 s 118238 -400 118294 800 4 la_oen_mprj[15]
port 678 nsew
rlabel metal2 s 118698 -400 118754 800 4 la_oen_mprj[16]
port 679 nsew
rlabel metal2 s 119158 -400 119214 800 4 la_oen_mprj[17]
port 680 nsew
rlabel metal2 s 119526 -400 119582 800 4 la_oen_mprj[18]
port 681 nsew
rlabel metal2 s 119986 -400 120042 800 4 la_oen_mprj[19]
port 682 nsew
rlabel metal2 s 112166 -400 112222 800 4 la_oen_mprj[1]
port 683 nsew
rlabel metal2 s 120446 -400 120502 800 4 la_oen_mprj[20]
port 684 nsew
rlabel metal2 s 120814 -400 120870 800 4 la_oen_mprj[21]
port 685 nsew
rlabel metal2 s 121274 -400 121330 800 4 la_oen_mprj[22]
port 686 nsew
rlabel metal2 s 121734 -400 121790 800 4 la_oen_mprj[23]
port 687 nsew
rlabel metal2 s 122194 -400 122250 800 4 la_oen_mprj[24]
port 688 nsew
rlabel metal2 s 122562 -400 122618 800 4 la_oen_mprj[25]
port 689 nsew
rlabel metal2 s 123022 -400 123078 800 4 la_oen_mprj[26]
port 690 nsew
rlabel metal2 s 123482 -400 123538 800 4 la_oen_mprj[27]
port 691 nsew
rlabel metal2 s 123942 -400 123998 800 4 la_oen_mprj[28]
port 692 nsew
rlabel metal2 s 124310 -400 124366 800 4 la_oen_mprj[29]
port 693 nsew
rlabel metal2 s 112534 -400 112590 800 4 la_oen_mprj[2]
port 694 nsew
rlabel metal2 s 124770 -400 124826 800 4 la_oen_mprj[30]
port 695 nsew
rlabel metal2 s 125230 -400 125286 800 4 la_oen_mprj[31]
port 696 nsew
rlabel metal2 s 125690 -400 125746 800 4 la_oen_mprj[32]
port 697 nsew
rlabel metal2 s 126058 -400 126114 800 4 la_oen_mprj[33]
port 698 nsew
rlabel metal2 s 126518 -400 126574 800 4 la_oen_mprj[34]
port 699 nsew
rlabel metal2 s 126978 -400 127034 800 4 la_oen_mprj[35]
port 700 nsew
rlabel metal2 s 127438 -400 127494 800 4 la_oen_mprj[36]
port 701 nsew
rlabel metal2 s 127806 -400 127862 800 4 la_oen_mprj[37]
port 702 nsew
rlabel metal2 s 128266 -400 128322 800 4 la_oen_mprj[38]
port 703 nsew
rlabel metal2 s 128726 -400 128782 800 4 la_oen_mprj[39]
port 704 nsew
rlabel metal2 s 112994 -400 113050 800 4 la_oen_mprj[3]
port 705 nsew
rlabel metal2 s 129094 -400 129150 800 4 la_oen_mprj[40]
port 706 nsew
rlabel metal2 s 129554 -400 129610 800 4 la_oen_mprj[41]
port 707 nsew
rlabel metal2 s 130014 -400 130070 800 4 la_oen_mprj[42]
port 708 nsew
rlabel metal2 s 130474 -400 130530 800 4 la_oen_mprj[43]
port 709 nsew
rlabel metal2 s 130842 -400 130898 800 4 la_oen_mprj[44]
port 710 nsew
rlabel metal2 s 131302 -400 131358 800 4 la_oen_mprj[45]
port 711 nsew
rlabel metal2 s 131762 -400 131818 800 4 la_oen_mprj[46]
port 712 nsew
rlabel metal2 s 132222 -400 132278 800 4 la_oen_mprj[47]
port 713 nsew
rlabel metal2 s 132590 -400 132646 800 4 la_oen_mprj[48]
port 714 nsew
rlabel metal2 s 133050 -400 133106 800 4 la_oen_mprj[49]
port 715 nsew
rlabel metal2 s 113454 -400 113510 800 4 la_oen_mprj[4]
port 716 nsew
rlabel metal2 s 133510 -400 133566 800 4 la_oen_mprj[50]
port 717 nsew
rlabel metal2 s 133970 -400 134026 800 4 la_oen_mprj[51]
port 718 nsew
rlabel metal2 s 134338 -400 134394 800 4 la_oen_mprj[52]
port 719 nsew
rlabel metal2 s 134798 -400 134854 800 4 la_oen_mprj[53]
port 720 nsew
rlabel metal2 s 135258 -400 135314 800 4 la_oen_mprj[54]
port 721 nsew
rlabel metal2 s 135718 -400 135774 800 4 la_oen_mprj[55]
port 722 nsew
rlabel metal2 s 136086 -400 136142 800 4 la_oen_mprj[56]
port 723 nsew
rlabel metal2 s 136546 -400 136602 800 4 la_oen_mprj[57]
port 724 nsew
rlabel metal2 s 137006 -400 137062 800 4 la_oen_mprj[58]
port 725 nsew
rlabel metal2 s 137374 -400 137430 800 4 la_oen_mprj[59]
port 726 nsew
rlabel metal2 s 113914 -400 113970 800 4 la_oen_mprj[5]
port 727 nsew
rlabel metal2 s 137834 -400 137890 800 4 la_oen_mprj[60]
port 728 nsew
rlabel metal2 s 138294 -400 138350 800 4 la_oen_mprj[61]
port 729 nsew
rlabel metal2 s 138754 -400 138810 800 4 la_oen_mprj[62]
port 730 nsew
rlabel metal2 s 139122 -400 139178 800 4 la_oen_mprj[63]
port 731 nsew
rlabel metal2 s 139582 -400 139638 800 4 la_oen_mprj[64]
port 732 nsew
rlabel metal2 s 140042 -400 140098 800 4 la_oen_mprj[65]
port 733 nsew
rlabel metal2 s 140502 -400 140558 800 4 la_oen_mprj[66]
port 734 nsew
rlabel metal2 s 140870 -400 140926 800 4 la_oen_mprj[67]
port 735 nsew
rlabel metal2 s 141330 -400 141386 800 4 la_oen_mprj[68]
port 736 nsew
rlabel metal2 s 141790 -400 141846 800 4 la_oen_mprj[69]
port 737 nsew
rlabel metal2 s 114282 -400 114338 800 4 la_oen_mprj[6]
port 738 nsew
rlabel metal2 s 142250 -400 142306 800 4 la_oen_mprj[70]
port 739 nsew
rlabel metal2 s 142618 -400 142674 800 4 la_oen_mprj[71]
port 740 nsew
rlabel metal2 s 143078 -400 143134 800 4 la_oen_mprj[72]
port 741 nsew
rlabel metal2 s 143538 -400 143594 800 4 la_oen_mprj[73]
port 742 nsew
rlabel metal2 s 143998 -400 144054 800 4 la_oen_mprj[74]
port 743 nsew
rlabel metal2 s 144366 -400 144422 800 4 la_oen_mprj[75]
port 744 nsew
rlabel metal2 s 144826 -400 144882 800 4 la_oen_mprj[76]
port 745 nsew
rlabel metal2 s 145286 -400 145342 800 4 la_oen_mprj[77]
port 746 nsew
rlabel metal2 s 145654 -400 145710 800 4 la_oen_mprj[78]
port 747 nsew
rlabel metal2 s 146114 -400 146170 800 4 la_oen_mprj[79]
port 748 nsew
rlabel metal2 s 114742 -400 114798 800 4 la_oen_mprj[7]
port 749 nsew
rlabel metal2 s 146574 -400 146630 800 4 la_oen_mprj[80]
port 750 nsew
rlabel metal2 s 147034 -400 147090 800 4 la_oen_mprj[81]
port 751 nsew
rlabel metal2 s 147402 -400 147458 800 4 la_oen_mprj[82]
port 752 nsew
rlabel metal2 s 147862 -400 147918 800 4 la_oen_mprj[83]
port 753 nsew
rlabel metal2 s 148322 -400 148378 800 4 la_oen_mprj[84]
port 754 nsew
rlabel metal2 s 148782 -400 148838 800 4 la_oen_mprj[85]
port 755 nsew
rlabel metal2 s 149150 -400 149206 800 4 la_oen_mprj[86]
port 756 nsew
rlabel metal2 s 149610 -400 149666 800 4 la_oen_mprj[87]
port 757 nsew
rlabel metal2 s 150070 -400 150126 800 4 la_oen_mprj[88]
port 758 nsew
rlabel metal2 s 150530 -400 150586 800 4 la_oen_mprj[89]
port 759 nsew
rlabel metal2 s 115202 -400 115258 800 4 la_oen_mprj[8]
port 760 nsew
rlabel metal2 s 150898 -400 150954 800 4 la_oen_mprj[90]
port 761 nsew
rlabel metal2 s 151358 -400 151414 800 4 la_oen_mprj[91]
port 762 nsew
rlabel metal2 s 151818 -400 151874 800 4 la_oen_mprj[92]
port 763 nsew
rlabel metal2 s 152186 -400 152242 800 4 la_oen_mprj[93]
port 764 nsew
rlabel metal2 s 152646 -400 152702 800 4 la_oen_mprj[94]
port 765 nsew
rlabel metal2 s 153106 -400 153162 800 4 la_oen_mprj[95]
port 766 nsew
rlabel metal2 s 153566 -400 153622 800 4 la_oen_mprj[96]
port 767 nsew
rlabel metal2 s 153934 -400 153990 800 4 la_oen_mprj[97]
port 768 nsew
rlabel metal2 s 154394 -400 154450 800 4 la_oen_mprj[98]
port 769 nsew
rlabel metal2 s 154854 -400 154910 800 4 la_oen_mprj[99]
port 770 nsew
rlabel metal2 s 115662 -400 115718 800 4 la_oen_mprj[9]
port 771 nsew
rlabel metal2 s 168746 -400 168802 800 4 mprj_adr_o_core[0]
port 772 nsew
rlabel metal2 s 179234 -400 179290 800 4 mprj_adr_o_core[10]
port 773 nsew
rlabel metal2 s 180154 -400 180210 800 4 mprj_adr_o_core[11]
port 774 nsew
rlabel metal2 s 180982 -400 181038 800 4 mprj_adr_o_core[12]
port 775 nsew
rlabel metal2 s 181902 -400 181958 800 4 mprj_adr_o_core[13]
port 776 nsew
rlabel metal2 s 182730 -400 182786 800 4 mprj_adr_o_core[14]
port 777 nsew
rlabel metal2 s 183650 -400 183706 800 4 mprj_adr_o_core[15]
port 778 nsew
rlabel metal2 s 184478 -400 184534 800 4 mprj_adr_o_core[16]
port 779 nsew
rlabel metal2 s 185306 -400 185362 800 4 mprj_adr_o_core[17]
port 780 nsew
rlabel metal2 s 186226 -400 186282 800 4 mprj_adr_o_core[18]
port 781 nsew
rlabel metal2 s 187054 -400 187110 800 4 mprj_adr_o_core[19]
port 782 nsew
rlabel metal2 s 170126 -400 170182 800 4 mprj_adr_o_core[1]
port 783 nsew
rlabel metal2 s 187974 -400 188030 800 4 mprj_adr_o_core[20]
port 784 nsew
rlabel metal2 s 188802 -400 188858 800 4 mprj_adr_o_core[21]
port 785 nsew
rlabel metal2 s 189722 -400 189778 800 4 mprj_adr_o_core[22]
port 786 nsew
rlabel metal2 s 190550 -400 190606 800 4 mprj_adr_o_core[23]
port 787 nsew
rlabel metal2 s 191470 -400 191526 800 4 mprj_adr_o_core[24]
port 788 nsew
rlabel metal2 s 192298 -400 192354 800 4 mprj_adr_o_core[25]
port 789 nsew
rlabel metal2 s 193218 -400 193274 800 4 mprj_adr_o_core[26]
port 790 nsew
rlabel metal2 s 194046 -400 194102 800 4 mprj_adr_o_core[27]
port 791 nsew
rlabel metal2 s 194966 -400 195022 800 4 mprj_adr_o_core[28]
port 792 nsew
rlabel metal2 s 195794 -400 195850 800 4 mprj_adr_o_core[29]
port 793 nsew
rlabel metal2 s 171414 -400 171470 800 4 mprj_adr_o_core[2]
port 794 nsew
rlabel metal2 s 196714 -400 196770 800 4 mprj_adr_o_core[30]
port 795 nsew
rlabel metal2 s 197542 -400 197598 800 4 mprj_adr_o_core[31]
port 796 nsew
rlabel metal2 s 172702 -400 172758 800 4 mprj_adr_o_core[3]
port 797 nsew
rlabel metal2 s 173990 -400 174046 800 4 mprj_adr_o_core[4]
port 798 nsew
rlabel metal2 s 174910 -400 174966 800 4 mprj_adr_o_core[5]
port 799 nsew
rlabel metal2 s 175738 -400 175794 800 4 mprj_adr_o_core[6]
port 800 nsew
rlabel metal2 s 176658 -400 176714 800 4 mprj_adr_o_core[7]
port 801 nsew
rlabel metal2 s 177486 -400 177542 800 4 mprj_adr_o_core[8]
port 802 nsew
rlabel metal2 s 178406 -400 178462 800 4 mprj_adr_o_core[9]
port 803 nsew
rlabel metal2 s 170494 10200 170550 11400 4 mprj_adr_o_user[0]
port 804 nsew
rlabel metal2 s 180982 10200 181038 11400 4 mprj_adr_o_user[10]
port 805 nsew
rlabel metal2 s 181902 10200 181958 11400 4 mprj_adr_o_user[11]
port 806 nsew
rlabel metal2 s 182730 10200 182786 11400 4 mprj_adr_o_user[12]
port 807 nsew
rlabel metal2 s 183650 10200 183706 11400 4 mprj_adr_o_user[13]
port 808 nsew
rlabel metal2 s 184478 10200 184534 11400 4 mprj_adr_o_user[14]
port 809 nsew
rlabel metal2 s 185306 10200 185362 11400 4 mprj_adr_o_user[15]
port 810 nsew
rlabel metal2 s 186226 10200 186282 11400 4 mprj_adr_o_user[16]
port 811 nsew
rlabel metal2 s 187054 10200 187110 11400 4 mprj_adr_o_user[17]
port 812 nsew
rlabel metal2 s 187974 10200 188030 11400 4 mprj_adr_o_user[18]
port 813 nsew
rlabel metal2 s 188802 10200 188858 11400 4 mprj_adr_o_user[19]
port 814 nsew
rlabel metal2 s 171874 10200 171930 11400 4 mprj_adr_o_user[1]
port 815 nsew
rlabel metal2 s 189722 10200 189778 11400 4 mprj_adr_o_user[20]
port 816 nsew
rlabel metal2 s 190550 10200 190606 11400 4 mprj_adr_o_user[21]
port 817 nsew
rlabel metal2 s 191470 10200 191526 11400 4 mprj_adr_o_user[22]
port 818 nsew
rlabel metal2 s 192298 10200 192354 11400 4 mprj_adr_o_user[23]
port 819 nsew
rlabel metal2 s 193218 10200 193274 11400 4 mprj_adr_o_user[24]
port 820 nsew
rlabel metal2 s 194046 10200 194102 11400 4 mprj_adr_o_user[25]
port 821 nsew
rlabel metal2 s 194966 10200 195022 11400 4 mprj_adr_o_user[26]
port 822 nsew
rlabel metal2 s 195794 10200 195850 11400 4 mprj_adr_o_user[27]
port 823 nsew
rlabel metal2 s 196714 10200 196770 11400 4 mprj_adr_o_user[28]
port 824 nsew
rlabel metal2 s 197542 10200 197598 11400 4 mprj_adr_o_user[29]
port 825 nsew
rlabel metal2 s 173162 10200 173218 11400 4 mprj_adr_o_user[2]
port 826 nsew
rlabel metal2 s 198462 10200 198518 11400 4 mprj_adr_o_user[30]
port 827 nsew
rlabel metal2 s 199290 10200 199346 11400 4 mprj_adr_o_user[31]
port 828 nsew
rlabel metal2 s 174450 10200 174506 11400 4 mprj_adr_o_user[3]
port 829 nsew
rlabel metal2 s 175738 10200 175794 11400 4 mprj_adr_o_user[4]
port 830 nsew
rlabel metal2 s 176658 10200 176714 11400 4 mprj_adr_o_user[5]
port 831 nsew
rlabel metal2 s 177486 10200 177542 11400 4 mprj_adr_o_user[6]
port 832 nsew
rlabel metal2 s 178406 10200 178462 11400 4 mprj_adr_o_user[7]
port 833 nsew
rlabel metal2 s 179234 10200 179290 11400 4 mprj_adr_o_user[8]
port 834 nsew
rlabel metal2 s 180154 10200 180210 11400 4 mprj_adr_o_user[9]
port 835 nsew
rlabel metal2 s 167458 -400 167514 800 4 mprj_cyc_o_core
port 836 nsew
rlabel metal2 s 169206 10200 169262 11400 4 mprj_cyc_o_user
port 837 nsew
rlabel metal2 s 169206 -400 169262 800 4 mprj_dat_o_core[0]
port 838 nsew
rlabel metal2 s 179694 -400 179750 800 4 mprj_dat_o_core[10]
port 839 nsew
rlabel metal2 s 180522 -400 180578 800 4 mprj_dat_o_core[11]
port 840 nsew
rlabel metal2 s 181442 -400 181498 800 4 mprj_dat_o_core[12]
port 841 nsew
rlabel metal2 s 182270 -400 182326 800 4 mprj_dat_o_core[13]
port 842 nsew
rlabel metal2 s 183190 -400 183246 800 4 mprj_dat_o_core[14]
port 843 nsew
rlabel metal2 s 184018 -400 184074 800 4 mprj_dat_o_core[15]
port 844 nsew
rlabel metal2 s 184938 -400 184994 800 4 mprj_dat_o_core[16]
port 845 nsew
rlabel metal2 s 185766 -400 185822 800 4 mprj_dat_o_core[17]
port 846 nsew
rlabel metal2 s 186686 -400 186742 800 4 mprj_dat_o_core[18]
port 847 nsew
rlabel metal2 s 187514 -400 187570 800 4 mprj_dat_o_core[19]
port 848 nsew
rlabel metal2 s 170494 -400 170550 800 4 mprj_dat_o_core[1]
port 849 nsew
rlabel metal2 s 188434 -400 188490 800 4 mprj_dat_o_core[20]
port 850 nsew
rlabel metal2 s 189262 -400 189318 800 4 mprj_dat_o_core[21]
port 851 nsew
rlabel metal2 s 190182 -400 190238 800 4 mprj_dat_o_core[22]
port 852 nsew
rlabel metal2 s 191010 -400 191066 800 4 mprj_dat_o_core[23]
port 853 nsew
rlabel metal2 s 191930 -400 191986 800 4 mprj_dat_o_core[24]
port 854 nsew
rlabel metal2 s 192758 -400 192814 800 4 mprj_dat_o_core[25]
port 855 nsew
rlabel metal2 s 193586 -400 193642 800 4 mprj_dat_o_core[26]
port 856 nsew
rlabel metal2 s 194506 -400 194562 800 4 mprj_dat_o_core[27]
port 857 nsew
rlabel metal2 s 195334 -400 195390 800 4 mprj_dat_o_core[28]
port 858 nsew
rlabel metal2 s 196254 -400 196310 800 4 mprj_dat_o_core[29]
port 859 nsew
rlabel metal2 s 171874 -400 171930 800 4 mprj_dat_o_core[2]
port 860 nsew
rlabel metal2 s 197082 -400 197138 800 4 mprj_dat_o_core[30]
port 861 nsew
rlabel metal2 s 198002 -400 198058 800 4 mprj_dat_o_core[31]
port 862 nsew
rlabel metal2 s 173162 -400 173218 800 4 mprj_dat_o_core[3]
port 863 nsew
rlabel metal2 s 174450 -400 174506 800 4 mprj_dat_o_core[4]
port 864 nsew
rlabel metal2 s 175370 -400 175426 800 4 mprj_dat_o_core[5]
port 865 nsew
rlabel metal2 s 176198 -400 176254 800 4 mprj_dat_o_core[6]
port 866 nsew
rlabel metal2 s 177026 -400 177082 800 4 mprj_dat_o_core[7]
port 867 nsew
rlabel metal2 s 177946 -400 178002 800 4 mprj_dat_o_core[8]
port 868 nsew
rlabel metal2 s 178774 -400 178830 800 4 mprj_dat_o_core[9]
port 869 nsew
rlabel metal2 s 170954 10200 171010 11400 4 mprj_dat_o_user[0]
port 870 nsew
rlabel metal2 s 181442 10200 181498 11400 4 mprj_dat_o_user[10]
port 871 nsew
rlabel metal2 s 182270 10200 182326 11400 4 mprj_dat_o_user[11]
port 872 nsew
rlabel metal2 s 183190 10200 183246 11400 4 mprj_dat_o_user[12]
port 873 nsew
rlabel metal2 s 184018 10200 184074 11400 4 mprj_dat_o_user[13]
port 874 nsew
rlabel metal2 s 184938 10200 184994 11400 4 mprj_dat_o_user[14]
port 875 nsew
rlabel metal2 s 185766 10200 185822 11400 4 mprj_dat_o_user[15]
port 876 nsew
rlabel metal2 s 186686 10200 186742 11400 4 mprj_dat_o_user[16]
port 877 nsew
rlabel metal2 s 187514 10200 187570 11400 4 mprj_dat_o_user[17]
port 878 nsew
rlabel metal2 s 188434 10200 188490 11400 4 mprj_dat_o_user[18]
port 879 nsew
rlabel metal2 s 189262 10200 189318 11400 4 mprj_dat_o_user[19]
port 880 nsew
rlabel metal2 s 172242 10200 172298 11400 4 mprj_dat_o_user[1]
port 881 nsew
rlabel metal2 s 190182 10200 190238 11400 4 mprj_dat_o_user[20]
port 882 nsew
rlabel metal2 s 191010 10200 191066 11400 4 mprj_dat_o_user[21]
port 883 nsew
rlabel metal2 s 191930 10200 191986 11400 4 mprj_dat_o_user[22]
port 884 nsew
rlabel metal2 s 192758 10200 192814 11400 4 mprj_dat_o_user[23]
port 885 nsew
rlabel metal2 s 193586 10200 193642 11400 4 mprj_dat_o_user[24]
port 886 nsew
rlabel metal2 s 194506 10200 194562 11400 4 mprj_dat_o_user[25]
port 887 nsew
rlabel metal2 s 195334 10200 195390 11400 4 mprj_dat_o_user[26]
port 888 nsew
rlabel metal2 s 196254 10200 196310 11400 4 mprj_dat_o_user[27]
port 889 nsew
rlabel metal2 s 197082 10200 197138 11400 4 mprj_dat_o_user[28]
port 890 nsew
rlabel metal2 s 198002 10200 198058 11400 4 mprj_dat_o_user[29]
port 891 nsew
rlabel metal2 s 173622 10200 173678 11400 4 mprj_dat_o_user[2]
port 892 nsew
rlabel metal2 s 198830 10200 198886 11400 4 mprj_dat_o_user[30]
port 893 nsew
rlabel metal2 s 199750 10200 199806 11400 4 mprj_dat_o_user[31]
port 894 nsew
rlabel metal2 s 174910 10200 174966 11400 4 mprj_dat_o_user[3]
port 895 nsew
rlabel metal2 s 176198 10200 176254 11400 4 mprj_dat_o_user[4]
port 896 nsew
rlabel metal2 s 177026 10200 177082 11400 4 mprj_dat_o_user[5]
port 897 nsew
rlabel metal2 s 177946 10200 178002 11400 4 mprj_dat_o_user[6]
port 898 nsew
rlabel metal2 s 178774 10200 178830 11400 4 mprj_dat_o_user[7]
port 899 nsew
rlabel metal2 s 179694 10200 179750 11400 4 mprj_dat_o_user[8]
port 900 nsew
rlabel metal2 s 180522 10200 180578 11400 4 mprj_dat_o_user[9]
port 901 nsew
rlabel metal2 s 169666 -400 169722 800 4 mprj_sel_o_core[0]
port 902 nsew
rlabel metal2 s 170954 -400 171010 800 4 mprj_sel_o_core[1]
port 903 nsew
rlabel metal2 s 172242 -400 172298 800 4 mprj_sel_o_core[2]
port 904 nsew
rlabel metal2 s 173622 -400 173678 800 4 mprj_sel_o_core[3]
port 905 nsew
rlabel metal2 s 171414 10200 171470 11400 4 mprj_sel_o_user[0]
port 906 nsew
rlabel metal2 s 172702 10200 172758 11400 4 mprj_sel_o_user[1]
port 907 nsew
rlabel metal2 s 173990 10200 174046 11400 4 mprj_sel_o_user[2]
port 908 nsew
rlabel metal2 s 175370 10200 175426 11400 4 mprj_sel_o_user[3]
port 909 nsew
rlabel metal2 s 167918 -400 167974 800 4 mprj_stb_o_core
port 910 nsew
rlabel metal2 s 169666 10200 169722 11400 4 mprj_stb_o_user
port 911 nsew
rlabel metal2 s 168378 -400 168434 800 4 mprj_we_o_core
port 912 nsew
rlabel metal2 s 170126 10200 170182 11400 4 mprj_we_o_user
port 913 nsew
rlabel metal2 s 198462 -400 198518 800 4 user1_vcc_powergood
port 914 nsew
rlabel metal2 s 198830 -400 198886 800 4 user1_vdd_powergood
port 915 nsew
rlabel metal2 s 199290 -400 199346 800 4 user2_vcc_powergood
port 916 nsew
rlabel metal2 s 199750 -400 199806 800 4 user2_vdd_powergood
port 917 nsew
rlabel metal2 s 202 10200 258 11400 4 user_clock
port 918 nsew
rlabel metal2 s 570 10200 626 11400 4 user_clock2
port 919 nsew
rlabel metal2 s 1030 10200 1086 11400 4 user_reset
port 920 nsew
rlabel metal2 s 1490 10200 1546 11400 4 user_resetn
port 921 nsew
rlabel metal3 s -326 11162 200242 11222 4 vccd1
port 922 nsew
rlabel metal3 s -326 -342 200242 -282 4 vccd1
port 922 nsew
rlabel metal4 s 164074 -482 164134 11362 4 vccd1
port 922 nsew
rlabel metal4 s 124074 -482 124134 11362 4 vccd1
port 922 nsew
rlabel metal4 s 84074 -482 84134 11362 4 vccd1
port 922 nsew
rlabel metal4 s 44074 -482 44134 11362 4 vccd1
port 922 nsew
rlabel metal4 s 4074 -482 4134 11362 4 vccd1
port 922 nsew
rlabel metal4 s 200182 -342 200242 11222 4 vccd1
port 922 nsew
rlabel metal4 s -326 -342 -266 11222 4 vccd1
port 922 nsew
rlabel metal3 s -466 11302 200382 11362 4 vssd1
port 923 nsew
rlabel metal3 s -466 -482 200382 -422 4 vssd1
port 923 nsew
rlabel metal4 s 200322 -482 200382 11362 4 vssd1
port 923 nsew
rlabel metal4 s 184074 -482 184134 11362 4 vssd1
port 923 nsew
rlabel metal4 s 144074 -482 144134 11362 4 vssd1
port 923 nsew
rlabel metal4 s 104074 -482 104134 11362 4 vssd1
port 923 nsew
rlabel metal4 s 64074 -482 64134 11362 4 vssd1
port 923 nsew
rlabel metal4 s 24074 -482 24134 11362 4 vssd1
port 923 nsew
rlabel metal4 s -466 -482 -406 11362 4 vssd1
port 923 nsew
rlabel metal3 s -606 11442 200522 11502 4 vccd
port 924 nsew
rlabel metal3 s -606 -622 200522 -562 4 vccd
port 924 nsew
rlabel metal4 s 164474 -762 164534 11642 4 vccd
port 924 nsew
rlabel metal4 s 124474 -762 124534 11642 4 vccd
port 924 nsew
rlabel metal4 s 84474 -762 84534 11642 4 vccd
port 924 nsew
rlabel metal4 s 44474 -762 44534 11642 4 vccd
port 924 nsew
rlabel metal4 s 4474 -762 4534 11642 4 vccd
port 924 nsew
rlabel metal4 s 200462 -622 200522 11502 4 vccd
port 924 nsew
rlabel metal4 s -606 -622 -546 11502 4 vccd
port 924 nsew
rlabel metal3 s -746 11582 200662 11642 4 vssd
port 925 nsew
rlabel metal3 s -746 -762 200662 -702 4 vssd
port 925 nsew
rlabel metal4 s 200602 -762 200662 11642 4 vssd
port 925 nsew
rlabel metal4 s 184474 -762 184534 11642 4 vssd
port 925 nsew
rlabel metal4 s 144474 -762 144534 11642 4 vssd
port 925 nsew
rlabel metal4 s 104474 -762 104534 11642 4 vssd
port 925 nsew
rlabel metal4 s 64474 -762 64534 11642 4 vssd
port 925 nsew
rlabel metal4 s 24474 -762 24534 11642 4 vssd
port 925 nsew
rlabel metal4 s -746 -762 -686 11642 4 vssd
port 925 nsew
rlabel metal3 s -886 11722 200802 11782 4 vccd2
port 926 nsew
rlabel metal3 s -886 -902 200802 -842 4 vccd2
port 926 nsew
rlabel metal4 s 164874 -1042 164934 11922 4 vccd2
port 926 nsew
rlabel metal4 s 124874 -1042 124934 11922 4 vccd2
port 926 nsew
rlabel metal4 s 84874 -1042 84934 11922 4 vccd2
port 926 nsew
rlabel metal4 s 44874 -1042 44934 11922 4 vccd2
port 926 nsew
rlabel metal4 s 4874 -1042 4934 11922 4 vccd2
port 926 nsew
rlabel metal4 s 200742 -902 200802 11782 4 vccd2
port 926 nsew
rlabel metal4 s -886 -902 -826 11782 4 vccd2
port 926 nsew
rlabel metal3 s -1026 11862 200942 11922 4 vssd2
port 927 nsew
rlabel metal3 s -1026 -1042 200942 -982 4 vssd2
port 927 nsew
rlabel metal4 s 200882 -1042 200942 11922 4 vssd2
port 927 nsew
rlabel metal4 s 184874 -1042 184934 11922 4 vssd2
port 927 nsew
rlabel metal4 s 144874 -1042 144934 11922 4 vssd2
port 927 nsew
rlabel metal4 s 104874 -1042 104934 11922 4 vssd2
port 927 nsew
rlabel metal4 s 64874 -1042 64934 11922 4 vssd2
port 927 nsew
rlabel metal4 s 24874 -1042 24934 11922 4 vssd2
port 927 nsew
rlabel metal4 s -1026 -1042 -966 11922 4 vssd2
port 927 nsew
rlabel metal3 s -1166 12002 201082 12062 4 vdda1
port 928 nsew
rlabel metal3 s -1166 -1182 201082 -1122 4 vdda1
port 928 nsew
rlabel metal4 s 165274 -1322 165334 12202 4 vdda1
port 928 nsew
rlabel metal4 s 125274 -1322 125334 12202 4 vdda1
port 928 nsew
rlabel metal4 s 85274 -1322 85334 12202 4 vdda1
port 928 nsew
rlabel metal4 s 45274 -1322 45334 12202 4 vdda1
port 928 nsew
rlabel metal4 s 5274 -1322 5334 12202 4 vdda1
port 928 nsew
rlabel metal4 s 201022 -1182 201082 12062 4 vdda1
port 928 nsew
rlabel metal4 s -1166 -1182 -1106 12062 4 vdda1
port 928 nsew
rlabel metal3 s -1306 12142 201222 12202 4 vssa1
port 929 nsew
rlabel metal3 s -1306 -1322 201222 -1262 4 vssa1
port 929 nsew
rlabel metal4 s 201162 -1322 201222 12202 4 vssa1
port 929 nsew
rlabel metal4 s 185274 -1322 185334 12202 4 vssa1
port 929 nsew
rlabel metal4 s 145274 -1322 145334 12202 4 vssa1
port 929 nsew
rlabel metal4 s 105274 -1322 105334 12202 4 vssa1
port 929 nsew
rlabel metal4 s 65274 -1322 65334 12202 4 vssa1
port 929 nsew
rlabel metal4 s 25274 -1322 25334 12202 4 vssa1
port 929 nsew
rlabel metal4 s -1306 -1322 -1246 12202 4 vssa1
port 929 nsew
rlabel metal3 s -1446 12282 201362 12342 4 vdda2
port 930 nsew
rlabel metal3 s -1446 -1462 201362 -1402 4 vdda2
port 930 nsew
rlabel metal4 s 165674 -1602 165734 12482 4 vdda2
port 930 nsew
rlabel metal4 s 125674 -1602 125734 12482 4 vdda2
port 930 nsew
rlabel metal4 s 85674 -1602 85734 12482 4 vdda2
port 930 nsew
rlabel metal4 s 45674 -1602 45734 12482 4 vdda2
port 930 nsew
rlabel metal4 s 5674 -1602 5734 12482 4 vdda2
port 930 nsew
rlabel metal4 s 201302 -1462 201362 12342 4 vdda2
port 930 nsew
rlabel metal4 s -1446 -1462 -1386 12342 4 vdda2
port 930 nsew
rlabel metal3 s -1586 12422 201502 12482 4 vssa2
port 931 nsew
rlabel metal3 s -1586 -1602 201502 -1542 4 vssa2
port 931 nsew
rlabel metal4 s 201442 -1602 201502 12482 4 vssa2
port 931 nsew
rlabel metal4 s 185674 -1602 185734 12482 4 vssa2
port 931 nsew
rlabel metal4 s 145674 -1602 145734 12482 4 vssa2
port 931 nsew
rlabel metal4 s 105674 -1602 105734 12482 4 vssa2
port 931 nsew
rlabel metal4 s 65674 -1602 65734 12482 4 vssa2
port 931 nsew
rlabel metal4 s 25674 -1602 25734 12482 4 vssa2
port 931 nsew
rlabel metal4 s -1586 -1602 -1526 12482 4 vssa2
port 931 nsew
<< properties >>
string FIXED_BBOX 0 0 200000 11000
<< end >>
