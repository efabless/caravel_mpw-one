magic
tech sky130A
magscale 1 2
timestamp 1619660031
<< metal2 >>
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< metal3 >>
rect 16836 710520 21836 712360
rect 68236 710520 73236 712360
rect 119636 710520 124636 712360
rect 166191 710521 170971 712360
rect 171271 710520 173471 712360
rect 173670 710520 175870 712360
rect 176170 710521 180950 712360
rect 217591 710521 222371 712360
rect 222671 710520 224871 712360
rect 225070 710520 227270 712360
rect 227570 710521 232350 712360
rect 319591 710521 324371 712360
rect 324671 710520 326871 712360
rect 327070 710520 329270 712360
rect 329570 710521 334350 712360
rect 413436 710520 418436 712360
rect 464836 710520 469836 712360
rect 510391 710434 515171 712360
rect 520370 710434 525150 712360
rect 566636 710520 571636 712360
rect -8960 689604 -7520 689844
rect 591520 688924 592960 689164
rect -9044 681426 -7546 686426
rect -8960 680220 -7520 680460
rect 591476 677938 593126 682938
rect 591530 676993 592970 677233
rect -8960 670836 -7520 671076
rect 591520 669068 592960 669308
rect -8960 661452 -7520 661692
rect 591520 659140 592960 659380
rect -8960 652068 -7520 652308
rect 591520 649212 592960 649452
rect -9044 643433 -7520 648222
rect -8960 642684 -7520 642924
rect 591492 638982 593126 643782
rect 591520 638284 592960 638524
rect -9044 633382 -7520 638182
rect -8960 632300 -7520 632540
rect 591492 628942 593126 633731
rect 591520 628356 592960 628596
rect -8960 623916 -7520 624156
rect 591520 619428 592960 619668
rect -8960 614532 -7520 614772
rect 591520 609500 592960 609740
rect -8960 605148 -7520 605388
rect 591520 599708 592960 599948
rect -8960 595764 -7520 596004
rect 591520 589780 592960 590020
rect -8960 586380 -7520 586620
rect 591520 579852 592960 580092
rect -8960 576996 -7520 577236
rect 591520 569924 592960 570164
rect -8960 567612 -7520 567852
rect -9044 558960 -7560 563740
rect 591520 559996 592960 560236
rect -8960 558228 -7520 558468
rect -9044 548981 -7560 553761
rect 591498 549803 593126 554583
rect 591520 549068 592960 549308
rect -8960 545844 -7520 546084
rect 591498 539824 593126 544604
rect -8960 539460 -7520 539700
rect 591520 539140 592960 539380
rect -8960 530076 -7520 530316
rect 591520 530212 592960 530452
rect -8960 520692 -7520 520932
rect 591520 520284 592960 520524
rect -8960 511308 -7520 511548
rect 591520 510356 592960 510596
rect -8960 501924 -7520 502164
rect 591520 500564 592960 500804
rect -8960 492540 -7520 492780
rect 591520 490636 592960 490876
rect -8960 483156 -7520 483396
rect 591520 480708 592960 480948
rect -8960 473772 -7520 474012
rect 591520 470780 592960 471020
rect -8960 464388 -7520 464628
rect 591520 460852 592960 461092
rect -8960 455004 -7520 455244
rect 591520 450924 592960 451164
rect -8960 445620 -7520 445860
rect 591520 440996 592960 441236
rect -8960 436236 -7520 436476
rect 591520 431068 592960 431308
rect -8960 426852 -7520 427092
rect 591520 421140 592960 421380
rect -8960 417468 -7520 417708
rect 591520 411212 592960 411452
rect -8960 408084 -7520 408324
rect 591520 401420 592960 401660
rect -8960 398700 -7520 398940
rect 591520 391492 592960 391732
rect -8960 389316 -7520 389556
rect 591520 381564 592960 381804
rect -8960 379932 -7520 380172
rect 591520 371636 592960 371876
rect -8960 370548 -7520 370788
rect 591520 361708 592960 361948
rect -8960 361164 -7520 361404
rect -8960 351780 -7520 352020
rect 591520 351780 592960 352020
rect -8960 342396 -7520 342636
rect 591520 341852 592960 342092
rect -8960 333012 -7520 333252
rect 591520 331924 592960 332164
rect -8960 323628 -7520 323868
rect 591520 321996 592960 322236
rect -8960 314244 -7520 314484
rect 591520 312068 592960 312308
rect -8960 304860 -7520 305100
rect 591520 302276 592960 302516
rect -8960 295476 -7520 295716
rect 591520 292348 592960 292588
rect -8960 286092 -7520 286332
rect 591520 282420 592960 282660
rect -8960 276708 -7520 276948
rect 591520 272492 592960 272732
rect -8960 267324 -7520 267564
rect 591520 262564 592960 262804
rect -8960 257940 -7520 258180
rect 591520 252636 592960 252876
rect -8960 248556 -7520 248796
rect 591520 242708 592960 242948
rect -8960 239172 -7520 239412
rect 591548 235203 593126 239983
rect 591520 232780 592960 233020
rect -8960 229788 -7520 230028
rect 591548 225224 593126 230004
rect 591520 222852 592960 223092
rect -8960 220404 -7520 220644
rect -9044 214360 -7514 219140
rect 591520 212924 592960 213164
rect -8960 211020 -7520 211260
rect -9044 204381 -7514 209161
rect 591520 203132 592960 203372
rect -8960 201636 -7520 201876
rect -8960 192252 -7520 192492
rect 591458 191182 593126 195982
rect 591520 190204 592960 190444
rect -8960 182868 -7520 183108
rect 591458 181142 593126 185931
rect 591520 180276 592960 180516
rect -9044 172233 -7644 177022
rect 591520 173348 592960 173588
rect -8960 170484 -7520 170724
rect -9044 162182 -7644 166982
rect 591520 163420 592960 163660
rect -8960 161100 -7520 161340
rect -8960 154716 -7520 154956
rect 591520 153492 592960 153732
rect 591488 147003 593126 151783
rect -8960 145332 -7520 145572
rect 591520 143564 592960 143804
rect 591488 137024 593126 141804
rect -8960 135948 -7520 136188
rect 591520 133636 592960 133876
rect -8960 126564 -7520 126804
rect 591520 123708 592960 123948
rect -8960 117180 -7520 117420
rect 591520 113780 592960 114020
rect -8960 107796 -7520 108036
rect 591520 103988 592960 104228
rect -8960 98412 -7520 98652
rect 591520 94060 592960 94300
rect -8960 89028 -7520 89268
rect 591520 84132 592960 84372
rect -8960 79644 -7520 79884
rect 591520 74204 592960 74444
rect -8960 70260 -7520 70500
rect 591520 64276 592960 64516
rect -8960 60876 -7520 61116
rect 591520 54348 592960 54588
rect -8960 51492 -7520 51732
rect 591520 44420 592960 44660
rect -8960 42108 -7520 42348
rect 591520 34492 592960 34732
rect -8960 32724 -7520 32964
rect 591520 24564 592960 24804
rect -8960 23340 -7520 23580
rect 591520 14636 592960 14876
rect -8960 13956 -7520 14196
rect 591520 4844 592960 5084
rect -8960 4572 -7520 4812
<< comment >>
rect -9044 712160 593126 712360
rect -9044 -708 -8844 712160
rect 592926 -708 593126 712160
rect -9044 -908 593126 -708
<< labels >>
flabel metal2 s 125846 -960 125958 480 0 FreeSans 1600 90 0 0 la_data_in[0]
port 161 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 1600 90 0 0 la_data_in[100]
port 162 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 1600 90 0 0 la_data_in[101]
port 163 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 1600 90 0 0 la_data_in[102]
port 164 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 1600 90 0 0 la_data_in[103]
port 165 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 1600 90 0 0 la_data_in[104]
port 166 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 1600 90 0 0 la_data_in[105]
port 167 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 1600 90 0 0 la_data_in[106]
port 168 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 1600 90 0 0 la_data_in[107]
port 169 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 1600 90 0 0 la_data_in[108]
port 170 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 1600 90 0 0 la_data_in[109]
port 171 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 1600 90 0 0 la_data_in[10]
port 172 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 1600 90 0 0 la_data_in[110]
port 173 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 1600 90 0 0 la_data_in[111]
port 174 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 1600 90 0 0 la_data_in[112]
port 175 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 1600 90 0 0 la_data_in[113]
port 176 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 1600 90 0 0 la_data_in[114]
port 177 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 1600 90 0 0 la_data_in[115]
port 178 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 1600 90 0 0 la_data_in[116]
port 179 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 1600 90 0 0 la_data_in[117]
port 180 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 1600 90 0 0 la_data_in[118]
port 181 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 1600 90 0 0 la_data_in[119]
port 182 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 1600 90 0 0 la_data_in[11]
port 183 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 1600 90 0 0 la_data_in[120]
port 184 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 1600 90 0 0 la_data_in[121]
port 185 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 1600 90 0 0 la_data_in[122]
port 186 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 1600 90 0 0 la_data_in[123]
port 187 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 1600 90 0 0 la_data_in[124]
port 188 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 1600 90 0 0 la_data_in[125]
port 189 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 1600 90 0 0 la_data_in[126]
port 190 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 1600 90 0 0 la_data_in[127]
port 191 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 1600 90 0 0 la_data_in[12]
port 192 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 1600 90 0 0 la_data_in[13]
port 193 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 1600 90 0 0 la_data_in[14]
port 194 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 1600 90 0 0 la_data_in[15]
port 195 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 1600 90 0 0 la_data_in[16]
port 196 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 1600 90 0 0 la_data_in[17]
port 197 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 1600 90 0 0 la_data_in[18]
port 198 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 1600 90 0 0 la_data_in[19]
port 199 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 1600 90 0 0 la_data_in[1]
port 200 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 1600 90 0 0 la_data_in[20]
port 201 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 1600 90 0 0 la_data_in[21]
port 202 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 1600 90 0 0 la_data_in[22]
port 203 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 1600 90 0 0 la_data_in[23]
port 204 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 1600 90 0 0 la_data_in[24]
port 205 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 1600 90 0 0 la_data_in[25]
port 206 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 1600 90 0 0 la_data_in[26]
port 207 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 1600 90 0 0 la_data_in[27]
port 208 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 1600 90 0 0 la_data_in[28]
port 209 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 1600 90 0 0 la_data_in[29]
port 210 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 1600 90 0 0 la_data_in[2]
port 211 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 1600 90 0 0 la_data_in[30]
port 212 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 1600 90 0 0 la_data_in[31]
port 213 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 1600 90 0 0 la_data_in[32]
port 214 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 1600 90 0 0 la_data_in[33]
port 215 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 1600 90 0 0 la_data_in[34]
port 216 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 1600 90 0 0 la_data_in[35]
port 217 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 1600 90 0 0 la_data_in[36]
port 218 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 1600 90 0 0 la_data_in[37]
port 219 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 1600 90 0 0 la_data_in[38]
port 220 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 1600 90 0 0 la_data_in[39]
port 221 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 1600 90 0 0 la_data_in[3]
port 222 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 1600 90 0 0 la_data_in[40]
port 223 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 1600 90 0 0 la_data_in[41]
port 224 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 1600 90 0 0 la_data_in[42]
port 225 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 1600 90 0 0 la_data_in[43]
port 226 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 1600 90 0 0 la_data_in[44]
port 227 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 1600 90 0 0 la_data_in[45]
port 228 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 1600 90 0 0 la_data_in[46]
port 229 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 1600 90 0 0 la_data_in[47]
port 230 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 1600 90 0 0 la_data_in[48]
port 231 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 1600 90 0 0 la_data_in[49]
port 232 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 1600 90 0 0 la_data_in[4]
port 233 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 1600 90 0 0 la_data_in[50]
port 234 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 1600 90 0 0 la_data_in[51]
port 235 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 1600 90 0 0 la_data_in[52]
port 236 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 1600 90 0 0 la_data_in[53]
port 237 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 1600 90 0 0 la_data_in[54]
port 238 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 1600 90 0 0 la_data_in[55]
port 239 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 1600 90 0 0 la_data_in[56]
port 240 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 1600 90 0 0 la_data_in[57]
port 241 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 1600 90 0 0 la_data_in[58]
port 242 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 1600 90 0 0 la_data_in[59]
port 243 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 1600 90 0 0 la_data_in[5]
port 244 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 1600 90 0 0 la_data_in[60]
port 245 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 1600 90 0 0 la_data_in[61]
port 246 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 1600 90 0 0 la_data_in[62]
port 247 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 1600 90 0 0 la_data_in[63]
port 248 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 1600 90 0 0 la_data_in[64]
port 249 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 1600 90 0 0 la_data_in[65]
port 250 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 1600 90 0 0 la_data_in[66]
port 251 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 1600 90 0 0 la_data_in[67]
port 252 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 1600 90 0 0 la_data_in[68]
port 253 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 1600 90 0 0 la_data_in[69]
port 254 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 1600 90 0 0 la_data_in[6]
port 255 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 1600 90 0 0 la_data_in[70]
port 256 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 1600 90 0 0 la_data_in[71]
port 257 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 1600 90 0 0 la_data_in[72]
port 258 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 1600 90 0 0 la_data_in[73]
port 259 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 1600 90 0 0 la_data_in[74]
port 260 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 1600 90 0 0 la_data_in[75]
port 261 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 1600 90 0 0 la_data_in[76]
port 262 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 1600 90 0 0 la_data_in[77]
port 263 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 1600 90 0 0 la_data_in[78]
port 264 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 1600 90 0 0 la_data_in[79]
port 265 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 1600 90 0 0 la_data_in[7]
port 266 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 1600 90 0 0 la_data_in[80]
port 267 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 1600 90 0 0 la_data_in[81]
port 268 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 1600 90 0 0 la_data_in[82]
port 269 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 1600 90 0 0 la_data_in[83]
port 270 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 1600 90 0 0 la_data_in[84]
port 271 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 1600 90 0 0 la_data_in[85]
port 272 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 1600 90 0 0 la_data_in[86]
port 273 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 1600 90 0 0 la_data_in[87]
port 274 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 1600 90 0 0 la_data_in[88]
port 275 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 1600 90 0 0 la_data_in[89]
port 276 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 1600 90 0 0 la_data_in[8]
port 277 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 1600 90 0 0 la_data_in[90]
port 278 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 1600 90 0 0 la_data_in[91]
port 279 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 1600 90 0 0 la_data_in[92]
port 280 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 1600 90 0 0 la_data_in[93]
port 281 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 1600 90 0 0 la_data_in[94]
port 282 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 1600 90 0 0 la_data_in[95]
port 283 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 1600 90 0 0 la_data_in[96]
port 284 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 1600 90 0 0 la_data_in[97]
port 285 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 1600 90 0 0 la_data_in[98]
port 286 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 1600 90 0 0 la_data_in[99]
port 287 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 1600 90 0 0 la_data_in[9]
port 288 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 1600 90 0 0 la_data_out[0]
port 289 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 1600 90 0 0 la_data_out[100]
port 290 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 1600 90 0 0 la_data_out[101]
port 291 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 1600 90 0 0 la_data_out[102]
port 292 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 1600 90 0 0 la_data_out[103]
port 293 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 1600 90 0 0 la_data_out[104]
port 294 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 1600 90 0 0 la_data_out[105]
port 295 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 1600 90 0 0 la_data_out[106]
port 296 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 1600 90 0 0 la_data_out[107]
port 297 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 1600 90 0 0 la_data_out[108]
port 298 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 1600 90 0 0 la_data_out[109]
port 299 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 1600 90 0 0 la_data_out[10]
port 300 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 1600 90 0 0 la_data_out[110]
port 301 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 1600 90 0 0 la_data_out[111]
port 302 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 1600 90 0 0 la_data_out[112]
port 303 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 1600 90 0 0 la_data_out[113]
port 304 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 1600 90 0 0 la_data_out[114]
port 305 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 1600 90 0 0 la_data_out[115]
port 306 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 1600 90 0 0 la_data_out[116]
port 307 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 1600 90 0 0 la_data_out[117]
port 308 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 1600 90 0 0 la_data_out[118]
port 309 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 1600 90 0 0 la_data_out[119]
port 310 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 1600 90 0 0 la_data_out[11]
port 311 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 1600 90 0 0 la_data_out[120]
port 312 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 1600 90 0 0 la_data_out[121]
port 313 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 1600 90 0 0 la_data_out[122]
port 314 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 1600 90 0 0 la_data_out[123]
port 315 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 1600 90 0 0 la_data_out[124]
port 316 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 1600 90 0 0 la_data_out[125]
port 317 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 1600 90 0 0 la_data_out[126]
port 318 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 1600 90 0 0 la_data_out[127]
port 319 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 1600 90 0 0 la_data_out[12]
port 320 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 1600 90 0 0 la_data_out[13]
port 321 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 1600 90 0 0 la_data_out[14]
port 322 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 1600 90 0 0 la_data_out[15]
port 323 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 1600 90 0 0 la_data_out[16]
port 324 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 1600 90 0 0 la_data_out[17]
port 325 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 1600 90 0 0 la_data_out[18]
port 326 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 1600 90 0 0 la_data_out[19]
port 327 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 1600 90 0 0 la_data_out[1]
port 328 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 1600 90 0 0 la_data_out[20]
port 329 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 1600 90 0 0 la_data_out[21]
port 330 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 1600 90 0 0 la_data_out[22]
port 331 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 1600 90 0 0 la_data_out[23]
port 332 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 1600 90 0 0 la_data_out[24]
port 333 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 1600 90 0 0 la_data_out[25]
port 334 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 1600 90 0 0 la_data_out[26]
port 335 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 1600 90 0 0 la_data_out[27]
port 336 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 1600 90 0 0 la_data_out[28]
port 337 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 1600 90 0 0 la_data_out[29]
port 338 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 1600 90 0 0 la_data_out[2]
port 339 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 1600 90 0 0 la_data_out[30]
port 340 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 1600 90 0 0 la_data_out[31]
port 341 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 1600 90 0 0 la_data_out[32]
port 342 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 1600 90 0 0 la_data_out[33]
port 343 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 1600 90 0 0 la_data_out[34]
port 344 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 1600 90 0 0 la_data_out[35]
port 345 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 1600 90 0 0 la_data_out[36]
port 346 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 1600 90 0 0 la_data_out[37]
port 347 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 1600 90 0 0 la_data_out[38]
port 348 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 1600 90 0 0 la_data_out[39]
port 349 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 1600 90 0 0 la_data_out[3]
port 350 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 1600 90 0 0 la_data_out[40]
port 351 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 1600 90 0 0 la_data_out[41]
port 352 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 1600 90 0 0 la_data_out[42]
port 353 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 1600 90 0 0 la_data_out[43]
port 354 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 1600 90 0 0 la_data_out[44]
port 355 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 1600 90 0 0 la_data_out[45]
port 356 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 1600 90 0 0 la_data_out[46]
port 357 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 1600 90 0 0 la_data_out[47]
port 358 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 1600 90 0 0 la_data_out[48]
port 359 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 1600 90 0 0 la_data_out[49]
port 360 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 1600 90 0 0 la_data_out[4]
port 361 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 1600 90 0 0 la_data_out[50]
port 362 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 1600 90 0 0 la_data_out[51]
port 363 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 1600 90 0 0 la_data_out[52]
port 364 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 1600 90 0 0 la_data_out[53]
port 365 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 1600 90 0 0 la_data_out[54]
port 366 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 1600 90 0 0 la_data_out[55]
port 367 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 1600 90 0 0 la_data_out[56]
port 368 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 1600 90 0 0 la_data_out[57]
port 369 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 1600 90 0 0 la_data_out[58]
port 370 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 1600 90 0 0 la_data_out[59]
port 371 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 1600 90 0 0 la_data_out[5]
port 372 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 1600 90 0 0 la_data_out[60]
port 373 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 1600 90 0 0 la_data_out[61]
port 374 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 1600 90 0 0 la_data_out[62]
port 375 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 1600 90 0 0 la_data_out[63]
port 376 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 1600 90 0 0 la_data_out[64]
port 377 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 1600 90 0 0 la_data_out[65]
port 378 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 1600 90 0 0 la_data_out[66]
port 379 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 1600 90 0 0 la_data_out[67]
port 380 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 1600 90 0 0 la_data_out[68]
port 381 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 1600 90 0 0 la_data_out[69]
port 382 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 1600 90 0 0 la_data_out[6]
port 383 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 1600 90 0 0 la_data_out[70]
port 384 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 1600 90 0 0 la_data_out[71]
port 385 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 1600 90 0 0 la_data_out[72]
port 386 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 1600 90 0 0 la_data_out[73]
port 387 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 1600 90 0 0 la_data_out[74]
port 388 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 1600 90 0 0 la_data_out[75]
port 389 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 1600 90 0 0 la_data_out[76]
port 390 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 1600 90 0 0 la_data_out[77]
port 391 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 1600 90 0 0 la_data_out[78]
port 392 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 1600 90 0 0 la_data_out[79]
port 393 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 1600 90 0 0 la_data_out[7]
port 394 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 1600 90 0 0 la_data_out[80]
port 395 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 1600 90 0 0 la_data_out[81]
port 396 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 1600 90 0 0 la_data_out[82]
port 397 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 1600 90 0 0 la_data_out[83]
port 398 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 1600 90 0 0 la_data_out[84]
port 399 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 1600 90 0 0 la_data_out[85]
port 400 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 1600 90 0 0 la_data_out[86]
port 401 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 1600 90 0 0 la_data_out[87]
port 402 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 1600 90 0 0 la_data_out[88]
port 403 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 1600 90 0 0 la_data_out[89]
port 404 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 1600 90 0 0 la_data_out[8]
port 405 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 1600 90 0 0 la_data_out[90]
port 406 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 1600 90 0 0 la_data_out[91]
port 407 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 1600 90 0 0 la_data_out[92]
port 408 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 1600 90 0 0 la_data_out[93]
port 409 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 1600 90 0 0 la_data_out[94]
port 410 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 1600 90 0 0 la_data_out[95]
port 411 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 1600 90 0 0 la_data_out[96]
port 412 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 1600 90 0 0 la_data_out[97]
port 413 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 1600 90 0 0 la_data_out[98]
port 414 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 1600 90 0 0 la_data_out[99]
port 415 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 1600 90 0 0 la_data_out[9]
port 416 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 1600 90 0 0 la_oenb[0]
port 417 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 1600 90 0 0 la_oenb[100]
port 418 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 1600 90 0 0 la_oenb[101]
port 419 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 1600 90 0 0 la_oenb[102]
port 420 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 1600 90 0 0 la_oenb[103]
port 421 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 1600 90 0 0 la_oenb[104]
port 422 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 1600 90 0 0 la_oenb[105]
port 423 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 1600 90 0 0 la_oenb[106]
port 424 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 1600 90 0 0 la_oenb[107]
port 425 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 1600 90 0 0 la_oenb[108]
port 426 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 1600 90 0 0 la_oenb[109]
port 427 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 1600 90 0 0 la_oenb[10]
port 428 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 1600 90 0 0 la_oenb[110]
port 429 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 1600 90 0 0 la_oenb[111]
port 430 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 1600 90 0 0 la_oenb[112]
port 431 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 1600 90 0 0 la_oenb[113]
port 432 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 1600 90 0 0 la_oenb[114]
port 433 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 1600 90 0 0 la_oenb[115]
port 434 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 1600 90 0 0 la_oenb[116]
port 435 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 1600 90 0 0 la_oenb[117]
port 436 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 1600 90 0 0 la_oenb[118]
port 437 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 1600 90 0 0 la_oenb[119]
port 438 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 1600 90 0 0 la_oenb[11]
port 439 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 1600 90 0 0 la_oenb[120]
port 440 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 1600 90 0 0 la_oenb[121]
port 441 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 1600 90 0 0 la_oenb[122]
port 442 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 1600 90 0 0 la_oenb[123]
port 443 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 1600 90 0 0 la_oenb[124]
port 444 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 1600 90 0 0 la_oenb[125]
port 445 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 1600 90 0 0 la_oenb[126]
port 446 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 1600 90 0 0 la_oenb[127]
port 447 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 1600 90 0 0 la_oenb[12]
port 448 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 1600 90 0 0 la_oenb[13]
port 449 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 1600 90 0 0 la_oenb[14]
port 450 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 1600 90 0 0 la_oenb[15]
port 451 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 1600 90 0 0 la_oenb[16]
port 452 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 1600 90 0 0 la_oenb[17]
port 453 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 1600 90 0 0 la_oenb[18]
port 454 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 1600 90 0 0 la_oenb[19]
port 455 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 1600 90 0 0 la_oenb[1]
port 456 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 1600 90 0 0 la_oenb[20]
port 457 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 1600 90 0 0 la_oenb[21]
port 458 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 1600 90 0 0 la_oenb[22]
port 459 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 1600 90 0 0 la_oenb[23]
port 460 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 1600 90 0 0 la_oenb[24]
port 461 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 1600 90 0 0 la_oenb[25]
port 462 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 1600 90 0 0 la_oenb[26]
port 463 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 1600 90 0 0 la_oenb[27]
port 464 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 1600 90 0 0 la_oenb[28]
port 465 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 1600 90 0 0 la_oenb[29]
port 466 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 1600 90 0 0 la_oenb[2]
port 467 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 1600 90 0 0 la_oenb[30]
port 468 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 1600 90 0 0 la_oenb[31]
port 469 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 1600 90 0 0 la_oenb[32]
port 470 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 1600 90 0 0 la_oenb[33]
port 471 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 1600 90 0 0 la_oenb[34]
port 472 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 1600 90 0 0 la_oenb[35]
port 473 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 1600 90 0 0 la_oenb[36]
port 474 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 1600 90 0 0 la_oenb[37]
port 475 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 1600 90 0 0 la_oenb[38]
port 476 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 1600 90 0 0 la_oenb[39]
port 477 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 1600 90 0 0 la_oenb[3]
port 478 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 1600 90 0 0 la_oenb[40]
port 479 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 1600 90 0 0 la_oenb[41]
port 480 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 1600 90 0 0 la_oenb[42]
port 481 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 1600 90 0 0 la_oenb[43]
port 482 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 1600 90 0 0 la_oenb[44]
port 483 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 1600 90 0 0 la_oenb[45]
port 484 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 1600 90 0 0 la_oenb[46]
port 485 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 1600 90 0 0 la_oenb[47]
port 486 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 1600 90 0 0 la_oenb[48]
port 487 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 1600 90 0 0 la_oenb[49]
port 488 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 1600 90 0 0 la_oenb[4]
port 489 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 1600 90 0 0 la_oenb[50]
port 490 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 1600 90 0 0 la_oenb[51]
port 491 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 1600 90 0 0 la_oenb[52]
port 492 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 1600 90 0 0 la_oenb[53]
port 493 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 1600 90 0 0 la_oenb[54]
port 494 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 1600 90 0 0 la_oenb[55]
port 495 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 1600 90 0 0 la_oenb[56]
port 496 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 1600 90 0 0 la_oenb[57]
port 497 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 1600 90 0 0 la_oenb[58]
port 498 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 1600 90 0 0 la_oenb[59]
port 499 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 1600 90 0 0 la_oenb[5]
port 500 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 1600 90 0 0 la_oenb[60]
port 501 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 1600 90 0 0 la_oenb[61]
port 502 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 1600 90 0 0 la_oenb[62]
port 503 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 1600 90 0 0 la_oenb[63]
port 504 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 1600 90 0 0 la_oenb[64]
port 505 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 1600 90 0 0 la_oenb[65]
port 506 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 1600 90 0 0 la_oenb[66]
port 507 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 1600 90 0 0 la_oenb[67]
port 508 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 1600 90 0 0 la_oenb[68]
port 509 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 1600 90 0 0 la_oenb[69]
port 510 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 1600 90 0 0 la_oenb[6]
port 511 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 1600 90 0 0 la_oenb[70]
port 512 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 1600 90 0 0 la_oenb[71]
port 513 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 1600 90 0 0 la_oenb[72]
port 514 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 1600 90 0 0 la_oenb[73]
port 515 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 1600 90 0 0 la_oenb[74]
port 516 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 1600 90 0 0 la_oenb[75]
port 517 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 1600 90 0 0 la_oenb[76]
port 518 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 1600 90 0 0 la_oenb[77]
port 519 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 1600 90 0 0 la_oenb[78]
port 520 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 1600 90 0 0 la_oenb[79]
port 521 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 1600 90 0 0 la_oenb[7]
port 522 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 1600 90 0 0 la_oenb[80]
port 523 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 1600 90 0 0 la_oenb[81]
port 524 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 1600 90 0 0 la_oenb[82]
port 525 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 1600 90 0 0 la_oenb[83]
port 526 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 1600 90 0 0 la_oenb[84]
port 527 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 1600 90 0 0 la_oenb[85]
port 528 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 1600 90 0 0 la_oenb[86]
port 529 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 1600 90 0 0 la_oenb[87]
port 530 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 1600 90 0 0 la_oenb[88]
port 531 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 1600 90 0 0 la_oenb[89]
port 532 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 1600 90 0 0 la_oenb[8]
port 533 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 1600 90 0 0 la_oenb[90]
port 534 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 1600 90 0 0 la_oenb[91]
port 535 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 1600 90 0 0 la_oenb[92]
port 536 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 1600 90 0 0 la_oenb[93]
port 537 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 1600 90 0 0 la_oenb[94]
port 538 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 1600 90 0 0 la_oenb[95]
port 539 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 1600 90 0 0 la_oenb[96]
port 540 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 1600 90 0 0 la_oenb[97]
port 541 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 1600 90 0 0 la_oenb[98]
port 542 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 1600 90 0 0 la_oenb[99]
port 543 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 1600 90 0 0 la_oenb[9]
port 544 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 1600 90 0 0 user_clock2
port 545 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 1600 90 0 0 user_irq[0]
port 546 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 1600 90 0 0 user_irq[1]
port 547 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 1600 90 0 0 user_irq[2]
port 548 nsew signal tristate
flabel metal2 s 542 -960 654 480 0 FreeSans 1600 90 0 0 wb_clk_i
port 549 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 1600 90 0 0 wbs_adr_i[10]
port 553 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 1600 90 0 0 wbs_adr_i[11]
port 554 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 1600 90 0 0 wbs_adr_i[12]
port 555 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 1600 90 0 0 wbs_adr_i[13]
port 556 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 1600 90 0 0 wbs_adr_i[14]
port 557 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 1600 90 0 0 wbs_adr_i[15]
port 558 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 1600 90 0 0 wbs_adr_i[16]
port 559 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 1600 90 0 0 wbs_adr_i[17]
port 560 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 1600 90 0 0 wbs_adr_i[18]
port 561 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 1600 90 0 0 wbs_adr_i[19]
port 562 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 1600 90 0 0 wbs_adr_i[1]
port 563 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 1600 90 0 0 wbs_adr_i[20]
port 564 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 1600 90 0 0 wbs_adr_i[21]
port 565 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 1600 90 0 0 wbs_adr_i[22]
port 566 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 1600 90 0 0 wbs_adr_i[23]
port 567 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 1600 90 0 0 wbs_adr_i[24]
port 568 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 1600 90 0 0 wbs_adr_i[25]
port 569 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 1600 90 0 0 wbs_adr_i[26]
port 570 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 1600 90 0 0 wbs_adr_i[27]
port 571 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 1600 90 0 0 wbs_adr_i[28]
port 572 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 1600 90 0 0 wbs_adr_i[29]
port 573 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 1600 90 0 0 wbs_adr_i[2]
port 574 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 1600 90 0 0 wbs_adr_i[30]
port 575 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 1600 90 0 0 wbs_adr_i[31]
port 576 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 1600 90 0 0 wbs_adr_i[3]
port 577 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 1600 90 0 0 wbs_adr_i[4]
port 578 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 1600 90 0 0 wbs_adr_i[5]
port 579 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 1600 90 0 0 wbs_adr_i[6]
port 580 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 1600 90 0 0 wbs_adr_i[7]
port 581 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 1600 90 0 0 wbs_adr_i[8]
port 582 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 1600 90 0 0 wbs_adr_i[9]
port 583 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 1600 90 0 0 wbs_dat_i[0]
port 585 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 1600 90 0 0 wbs_dat_i[10]
port 586 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 1600 90 0 0 wbs_dat_i[11]
port 587 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 1600 90 0 0 wbs_dat_i[12]
port 588 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 1600 90 0 0 wbs_dat_i[13]
port 589 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 1600 90 0 0 wbs_dat_i[14]
port 590 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 1600 90 0 0 wbs_dat_i[15]
port 591 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 1600 90 0 0 wbs_dat_i[16]
port 592 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 1600 90 0 0 wbs_dat_i[17]
port 593 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 1600 90 0 0 wbs_dat_i[18]
port 594 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 1600 90 0 0 wbs_dat_i[19]
port 595 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 1600 90 0 0 wbs_dat_i[1]
port 596 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 1600 90 0 0 wbs_dat_i[20]
port 597 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 1600 90 0 0 wbs_dat_i[21]
port 598 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 1600 90 0 0 wbs_dat_i[22]
port 599 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 1600 90 0 0 wbs_dat_i[23]
port 600 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 1600 90 0 0 wbs_dat_i[24]
port 601 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 1600 90 0 0 wbs_dat_i[25]
port 602 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 1600 90 0 0 wbs_dat_i[26]
port 603 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 1600 90 0 0 wbs_dat_i[27]
port 604 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 1600 90 0 0 wbs_dat_i[28]
port 605 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 1600 90 0 0 wbs_dat_i[29]
port 606 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 1600 90 0 0 wbs_dat_i[2]
port 607 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 1600 90 0 0 wbs_dat_i[30]
port 608 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 1600 90 0 0 wbs_dat_i[31]
port 609 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 1600 90 0 0 wbs_dat_i[3]
port 610 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 1600 90 0 0 wbs_dat_i[4]
port 611 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 1600 90 0 0 wbs_dat_i[5]
port 612 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 1600 90 0 0 wbs_dat_i[6]
port 613 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 1600 90 0 0 wbs_dat_i[7]
port 614 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 1600 90 0 0 wbs_dat_i[8]
port 615 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 1600 90 0 0 wbs_dat_i[9]
port 616 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 1600 90 0 0 wbs_dat_o[0]
port 617 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 1600 90 0 0 wbs_dat_o[10]
port 618 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 1600 90 0 0 wbs_dat_o[11]
port 619 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 1600 90 0 0 wbs_dat_o[12]
port 620 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 1600 90 0 0 wbs_dat_o[13]
port 621 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 1600 90 0 0 wbs_dat_o[14]
port 622 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 1600 90 0 0 wbs_dat_o[15]
port 623 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 1600 90 0 0 wbs_dat_o[16]
port 624 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 1600 90 0 0 wbs_dat_o[17]
port 625 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 1600 90 0 0 wbs_dat_o[18]
port 626 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 1600 90 0 0 wbs_dat_o[19]
port 627 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 1600 90 0 0 wbs_dat_o[1]
port 628 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 1600 90 0 0 wbs_dat_o[20]
port 629 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 1600 90 0 0 wbs_dat_o[21]
port 630 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 1600 90 0 0 wbs_dat_o[22]
port 631 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 1600 90 0 0 wbs_dat_o[23]
port 632 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 1600 90 0 0 wbs_dat_o[24]
port 633 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 1600 90 0 0 wbs_dat_o[25]
port 634 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 1600 90 0 0 wbs_dat_o[26]
port 635 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 1600 90 0 0 wbs_dat_o[27]
port 636 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 1600 90 0 0 wbs_dat_o[28]
port 637 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 1600 90 0 0 wbs_dat_o[29]
port 638 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 1600 90 0 0 wbs_dat_o[2]
port 639 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 1600 90 0 0 wbs_dat_o[30]
port 640 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 1600 90 0 0 wbs_dat_o[31]
port 641 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 1600 90 0 0 wbs_dat_o[3]
port 642 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 1600 90 0 0 wbs_dat_o[4]
port 643 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 1600 90 0 0 wbs_dat_o[5]
port 644 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 1600 90 0 0 wbs_dat_o[6]
port 645 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 1600 90 0 0 wbs_dat_o[7]
port 646 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 1600 90 0 0 wbs_dat_o[8]
port 647 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 1600 90 0 0 wbs_dat_o[9]
port 648 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 1600 90 0 0 wbs_sel_i[0]
port 649 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 1600 90 0 0 wbs_sel_i[1]
port 650 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 1600 90 0 0 wbs_sel_i[2]
port 651 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 1600 90 0 0 wbs_sel_i[3]
port 652 nsew signal input
flabel space 572491 272361 578029 279006 0 FreeSans 16000 0 0 0 IO7
flabel space 573045 317959 578583 324604 0 FreeSans 16000 0 0 0 IO8
flabel space 571119 364512 576657 371157 0 FreeSans 16000 0 0 0 IO9
flabel space 571304 409990 576842 416635 0 FreeSans 16000 0 0 0 IO10
flabel space 572321 453064 577859 459709 0 FreeSans 16000 0 0 0 IO11
flabel space 573615 497156 579153 503801 0 FreeSans 16000 0 0 0 IO12
flabel space 574447 587279 579985 593924 0 FreeSans 16000 0 0 0 IO13
flabel space 5619 37768 11157 44413 0 FreeSans 16000 0 0 0 IO34
flabel space 4855 80470 10393 87115 0 FreeSans 16000 0 0 0 IO33
flabel space 7945 121974 13483 128619 0 FreeSans 16000 0 0 0 IO32
flabel space 6264 249900 11802 256545 0 FreeSans 16000 0 0 0 IO31
flabel space 5718 294160 11256 300805 0 FreeSans 16000 0 0 0 IO30
flabel space 5429 337437 10967 344082 0 FreeSans 16000 0 0 0 IO29
flabel space 5806 379767 11344 386412 0 FreeSans 16000 0 0 0 IO28
flabel space 5602 423114 11140 429759 0 FreeSans 16000 0 0 0 IO27
flabel space 6992 466636 12530 473281 0 FreeSans 16000 0 0 0 IO26
flabel space 6648 510966 12186 517611 0 FreeSans 16000 0 0 0 IO25
flabel metal3 s -8960 558228 -7520 558468 0 FreeSans 1600 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -8960 501924 -7520 502164 0 FreeSans 1600 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -8960 445620 -7520 445860 0 FreeSans 1600 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -8960 389316 -7520 389556 0 FreeSans 1600 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -8960 333012 -7520 333252 0 FreeSans 1600 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -8960 276708 -7520 276948 0 FreeSans 1600 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -8960 220404 -7520 220644 0 FreeSans 1600 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -8960 689604 -7520 689844 0 FreeSans 1600 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -8960 670836 -7520 671076 0 FreeSans 1600 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -8960 614532 -7520 614772 0 FreeSans 1600 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s -8960 492540 -7520 492780 0 FreeSans 1600 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -8960 436236 -7520 436476 0 FreeSans 1600 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -8960 379932 -7520 380172 0 FreeSans 1600 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -8960 323628 -7520 323868 0 FreeSans 1600 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -8960 267324 -7520 267564 0 FreeSans 1600 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -8960 211020 -7520 211260 0 FreeSans 1600 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -8960 154716 -7520 154956 0 FreeSans 1600 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s -8960 680220 -7520 680460 0 FreeSans 1600 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -8960 661452 -7520 661692 0 FreeSans 1600 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -8960 642684 -7520 642924 0 FreeSans 1600 0 0 0 io_in[14]
port 63 nsew signal input
flabel metal3 s -8960 586380 -7520 586620 0 FreeSans 1600 0 0 0 io_in[15]
port 65 nsew signal input
flabel metal3 s -8960 576996 -7520 577236 0 FreeSans 1600 0 0 0 io_out[15]
port 66 nsew signal tristate
flabel metal3 s -8960 530076 -7520 530316 0 FreeSans 1600 0 0 0 io_in[16]
port 67 nsew signal input
flabel metal3 s -8960 520692 -7520 520932 0 FreeSans 1600 0 0 0 io_out[16]
port 68 nsew signal tristate
flabel metal3 s -8960 473772 -7520 474012 0 FreeSans 1600 0 0 0 io_in[17]
port 69 nsew signal input
flabel metal3 s -8960 464388 -7520 464628 0 FreeSans 1600 0 0 0 io_out[17]
port 70 nsew signal tristate
flabel metal3 s -8960 417468 -7520 417708 0 FreeSans 1600 0 0 0 io_in[18]
port 71 nsew signal input
flabel metal3 s -8960 408084 -7520 408324 0 FreeSans 1600 0 0 0 io_out[18]
port 72 nsew signal tristate
flabel metal3 s -8960 361164 -7520 361404 0 FreeSans 1600 0 0 0 io_in[19]
port 73 nsew signal input
flabel metal3 s -8960 351780 -7520 352020 0 FreeSans 1600 0 0 0 io_out[19]
port 74 nsew signal tristate
flabel metal3 s -8960 304860 -7520 305100 0 FreeSans 1600 0 0 0 io_in[20]
port 77 nsew signal input
flabel metal3 s -8960 295476 -7520 295716 0 FreeSans 1600 0 0 0 io_out[20]
port 78 nsew signal tristate
flabel metal3 s -8960 248556 -7520 248796 0 FreeSans 1600 0 0 0 io_in[21]
port 79 nsew signal input
flabel metal3 s -8960 239172 -7520 239412 0 FreeSans 1600 0 0 0 io_out[21]
port 80 nsew signal tristate
flabel metal3 s -8960 192252 -7520 192492 0 FreeSans 1600 0 0 0 io_in[22]
port 81 nsew signal input
flabel metal3 s -8960 182868 -7520 183108 0 FreeSans 1600 0 0 0 io_out[22]
port 82 nsew signal tristate
flabel metal3 s -8960 135948 -7520 136188 0 FreeSans 1600 0 0 0 io_in[23]
port 83 nsew signal input
flabel metal3 s -8960 126564 -7520 126804 0 FreeSans 1600 0 0 0 io_out[23]
port 84 nsew signal tristate
flabel metal3 s -8960 98412 -7520 98652 0 FreeSans 1600 0 0 0 io_in[24]
port 85 nsew signal input
flabel metal3 s -8960 89028 -7520 89268 0 FreeSans 1600 0 0 0 io_out[24]
port 86 nsew signal tristate
flabel metal3 s -8960 60876 -7520 61116 0 FreeSans 1600 0 0 0 io_in[25]
port 87 nsew signal input
flabel metal3 s -8960 51492 -7520 51732 0 FreeSans 1600 0 0 0 io_out[25]
port 88 nsew signal tristate
flabel metal3 s -8960 23340 -7520 23580 0 FreeSans 1600 0 0 0 io_in[26]
port 89 nsew signal input
flabel metal3 s -8960 13956 -7520 14196 0 FreeSans 1600 0 0 0 io_out[26]
port 90 nsew signal tristate
flabel metal3 s -8960 652068 -7520 652308 0 FreeSans 1600 0 0 0 io_in_3v3[14]
port 112 nsew signal input
flabel metal3 s -8960 539460 -7520 539700 0 FreeSans 1600 0 0 0 io_in_3v3[16]
port 114 nsew signal input
flabel metal3 s -8960 483156 -7520 483396 0 FreeSans 1600 0 0 0 io_in_3v3[17]
port 115 nsew signal input
flabel metal3 s -8960 426852 -7520 427092 0 FreeSans 1600 0 0 0 io_in_3v3[18]
port 116 nsew signal input
flabel metal3 s -8960 370548 -7520 370788 0 FreeSans 1600 0 0 0 io_in_3v3[19]
port 117 nsew signal input
flabel metal3 s -8960 314244 -7520 314484 0 FreeSans 1600 0 0 0 io_in_3v3[20]
port 119 nsew signal input
flabel metal3 s -8960 257940 -7520 258180 0 FreeSans 1600 0 0 0 io_in_3v3[21]
port 120 nsew signal input
flabel metal3 s -8960 201636 -7520 201876 0 FreeSans 1600 0 0 0 io_in_3v3[22]
port 121 nsew signal input
flabel metal3 s -8960 145332 -7520 145572 0 FreeSans 1600 0 0 0 io_in_3v3[23]
port 122 nsew signal input
flabel metal3 s -8960 107796 -7520 108036 0 FreeSans 1600 0 0 0 io_in_3v3[24]
port 123 nsew signal input
flabel metal3 s -8960 70260 -7520 70500 0 FreeSans 1600 0 0 0 io_in_3v3[25]
port 124 nsew signal input
flabel metal3 s -8960 32724 -7520 32964 0 FreeSans 1600 0 0 0 io_in_3v3[26]
port 125 nsew signal input
flabel metal3 s -8960 623916 -7520 624156 0 FreeSans 1600 0 0 0 io_oeb[14]
port 139 nsew signal tristate
flabel metal3 s -8960 567612 -7520 567852 0 FreeSans 1600 0 0 0 io_oeb[15]
port 140 nsew signal tristate
flabel metal3 s -8960 511308 -7520 511548 0 FreeSans 1600 0 0 0 io_oeb[16]
port 141 nsew signal tristate
flabel metal3 s -8960 455004 -7520 455244 0 FreeSans 1600 0 0 0 io_oeb[17]
port 142 nsew signal tristate
flabel metal3 s -8960 398700 -7520 398940 0 FreeSans 1600 0 0 0 io_oeb[18]
port 143 nsew signal tristate
flabel metal3 s -8960 342396 -7520 342636 0 FreeSans 1600 0 0 0 io_oeb[19]
port 144 nsew signal tristate
flabel metal3 s -8960 286092 -7520 286332 0 FreeSans 1600 0 0 0 io_oeb[20]
port 146 nsew signal tristate
flabel metal3 s -8960 229788 -7520 230028 0 FreeSans 1600 0 0 0 io_oeb[21]
port 147 nsew signal tristate
flabel metal3 s -8960 117180 -7520 117420 0 FreeSans 1600 0 0 0 io_oeb[23]
port 149 nsew signal tristate
flabel metal3 s -8960 79644 -7520 79884 0 FreeSans 1600 0 0 0 io_oeb[24]
port 150 nsew signal tristate
flabel metal3 s -8960 42108 -7520 42348 0 FreeSans 1600 0 0 0 io_oeb[25]
port 151 nsew signal tristate
flabel metal3 s -8960 4572 -7520 4812 0 FreeSans 1600 0 0 0 io_oeb[26]
port 152 nsew signal tristate
flabel metal3 s -8960 161100 -7520 161340 0 FreeSans 1600 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s -8960 170484 -7520 170724 0 FreeSans 1600 0 0 0 io_oeb[22]
port 148 nsew signal tristate
flabel metal3 s -8960 545844 -7520 546084 0 FreeSans 1600 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -8960 595764 -7520 596004 0 FreeSans 1600 0 0 0 io_in_3v3[15]
port 113 nsew signal input
flabel metal3 s -8960 605148 -7520 605388 0 FreeSans 1600 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s -8960 632300 -7520 632540 0 FreeSans 1600 0 0 0 io_out[14]
port 64 nsew signal tristate
flabel metal3 -7844 162182 -7644 166982 0 FreeSans 4000 0 0 0 VSSD2
port 689 nsew
flabel metal3 -7844 172233 -7644 177022 0 FreeSans 4000 0 0 0 VSSD2
port 690 nsew
flabel metal3 s 591520 282420 592960 282660 0 FreeSans 1600 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s 591520 341852 592960 342092 0 FreeSans 1600 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 591520 401420 592960 401660 0 FreeSans 1600 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 591520 460852 592960 461092 0 FreeSans 1600 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 591520 520284 592960 520524 0 FreeSans 1600 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 591520 579852 592960 580092 0 FreeSans 1600 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 591520 292348 592960 292588 0 FreeSans 1600 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s 591520 351780 592960 352020 0 FreeSans 1600 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 591520 411212 592960 411452 0 FreeSans 1600 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 591520 470780 592960 471020 0 FreeSans 1600 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 591520 530212 592960 530452 0 FreeSans 1600 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 591520 589780 592960 590020 0 FreeSans 1600 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 591520 649212 592960 649452 0 FreeSans 1600 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s 591520 14636 592960 14876 0 FreeSans 1600 0 0 0 io_in[0]
port 53 nsew signal input
flabel metal3 s 591520 24564 592960 24804 0 FreeSans 1600 0 0 0 io_out[0]
port 54 nsew signal tristate
flabel metal3 s 591520 490636 592960 490876 0 FreeSans 1600 0 0 0 io_in[10]
port 55 nsew signal input
flabel metal3 s 591520 500564 592960 500804 0 FreeSans 1600 0 0 0 io_out[10]
port 56 nsew signal tristate
flabel metal3 s 591520 559996 592960 560236 0 FreeSans 1600 0 0 0 io_out[11]
port 58 nsew signal tristate
flabel metal3 s 591520 609500 592960 609740 0 FreeSans 1600 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 591520 619428 592960 619668 0 FreeSans 1600 0 0 0 io_out[12]
port 60 nsew signal tristate
flabel metal3 s 591520 669068 592960 669308 0 FreeSans 1600 0 0 0 io_in[13]
port 61 nsew signal input
flabel metal3 s 591520 54348 592960 54588 0 FreeSans 1600 0 0 0 io_in[1]
port 75 nsew signal input
flabel metal3 s 591520 64276 592960 64516 0 FreeSans 1600 0 0 0 io_out[1]
port 76 nsew signal tristate
flabel metal3 s 591520 94060 592960 94300 0 FreeSans 1600 0 0 0 io_in[2]
port 91 nsew signal input
flabel metal3 s 591520 103988 592960 104228 0 FreeSans 1600 0 0 0 io_out[2]
port 92 nsew signal tristate
flabel metal3 s 591520 133636 592960 133876 0 FreeSans 1600 0 0 0 io_in[3]
port 93 nsew signal input
flabel metal3 s 591520 143564 592960 143804 0 FreeSans 1600 0 0 0 io_out[3]
port 94 nsew signal tristate
flabel metal3 s 591520 173348 592960 173588 0 FreeSans 1600 0 0 0 io_in[4]
port 95 nsew signal input
flabel metal3 s 591520 212924 592960 213164 0 FreeSans 1600 0 0 0 io_in[5]
port 97 nsew signal input
flabel metal3 s 591520 222852 592960 223092 0 FreeSans 1600 0 0 0 io_out[5]
port 98 nsew signal tristate
flabel metal3 s 591520 252636 592960 252876 0 FreeSans 1600 0 0 0 io_in[6]
port 99 nsew signal input
flabel metal3 s 591520 262564 592960 262804 0 FreeSans 1600 0 0 0 io_out[6]
port 100 nsew signal tristate
flabel metal3 s 591520 312068 592960 312308 0 FreeSans 1600 0 0 0 io_in[7]
port 101 nsew signal input
flabel metal3 s 591520 321996 592960 322236 0 FreeSans 1600 0 0 0 io_out[7]
port 102 nsew signal tristate
flabel metal3 s 591520 371636 592960 371876 0 FreeSans 1600 0 0 0 io_in[8]
port 103 nsew signal input
flabel metal3 s 591520 381564 592960 381804 0 FreeSans 1600 0 0 0 io_out[8]
port 104 nsew signal tristate
flabel metal3 s 591520 431068 592960 431308 0 FreeSans 1600 0 0 0 io_in[9]
port 105 nsew signal input
flabel metal3 s 591520 440996 592960 441236 0 FreeSans 1600 0 0 0 io_out[9]
port 106 nsew signal tristate
flabel metal3 s 591520 4844 592960 5084 0 FreeSans 1600 0 0 0 io_in_3v3[0]
port 107 nsew signal input
flabel metal3 s 591520 480708 592960 480948 0 FreeSans 1600 0 0 0 io_in_3v3[10]
port 108 nsew signal input
flabel metal3 s 591520 599708 592960 599948 0 FreeSans 1600 0 0 0 io_in_3v3[12]
port 110 nsew signal input
flabel metal3 s 591520 659140 592960 659380 0 FreeSans 1600 0 0 0 io_in_3v3[13]
port 111 nsew signal input
flabel metal3 s 591520 44420 592960 44660 0 FreeSans 1600 0 0 0 io_in_3v3[1]
port 118 nsew signal input
flabel metal3 s 591520 84132 592960 84372 0 FreeSans 1600 0 0 0 io_in_3v3[2]
port 126 nsew signal input
flabel metal3 s 591520 123708 592960 123948 0 FreeSans 1600 0 0 0 io_in_3v3[3]
port 127 nsew signal input
flabel metal3 s 591520 163420 592960 163660 0 FreeSans 1600 0 0 0 io_in_3v3[4]
port 128 nsew signal input
flabel metal3 s 591520 203132 592960 203372 0 FreeSans 1600 0 0 0 io_in_3v3[5]
port 129 nsew signal input
flabel metal3 s 591520 242708 592960 242948 0 FreeSans 1600 0 0 0 io_in_3v3[6]
port 130 nsew signal input
flabel metal3 s 591520 302276 592960 302516 0 FreeSans 1600 0 0 0 io_in_3v3[7]
port 131 nsew signal input
flabel metal3 s 591520 361708 592960 361948 0 FreeSans 1600 0 0 0 io_in_3v3[8]
port 132 nsew signal input
flabel metal3 s 591520 421140 592960 421380 0 FreeSans 1600 0 0 0 io_in_3v3[9]
port 133 nsew signal input
flabel metal3 s 591520 34492 592960 34732 0 FreeSans 1600 0 0 0 io_oeb[0]
port 134 nsew signal tristate
flabel metal3 s 591520 510356 592960 510596 0 FreeSans 1600 0 0 0 io_oeb[10]
port 135 nsew signal tristate
flabel metal3 s 591520 569924 592960 570164 0 FreeSans 1600 0 0 0 io_oeb[11]
port 136 nsew signal tristate
flabel metal3 s 591520 688924 592960 689164 0 FreeSans 1600 0 0 0 io_oeb[13]
port 138 nsew signal tristate
flabel metal3 s 591520 74204 592960 74444 0 FreeSans 1600 0 0 0 io_oeb[1]
port 145 nsew signal tristate
flabel metal3 s 591520 113780 592960 114020 0 FreeSans 1600 0 0 0 io_oeb[2]
port 153 nsew signal tristate
flabel metal3 s 591520 153492 592960 153732 0 FreeSans 1600 0 0 0 io_oeb[3]
port 154 nsew signal tristate
flabel metal3 s 591520 232780 592960 233020 0 FreeSans 1600 0 0 0 io_oeb[5]
port 156 nsew signal tristate
flabel metal3 s 591520 272492 592960 272732 0 FreeSans 1600 0 0 0 io_oeb[6]
port 157 nsew signal tristate
flabel metal3 s 591520 331924 592960 332164 0 FreeSans 1600 0 0 0 io_oeb[7]
port 158 nsew signal tristate
flabel metal3 s 591520 391492 592960 391732 0 FreeSans 1600 0 0 0 io_oeb[8]
port 159 nsew signal tristate
flabel metal3 s 591520 450924 592960 451164 0 FreeSans 1600 0 0 0 io_oeb[9]
port 160 nsew signal tristate
flabel metal3 s 591520 638284 592960 638524 0 FreeSans 1600 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s 591520 628356 592960 628596 0 FreeSans 1600 0 0 0 io_oeb[12]
port 137 nsew signal tristate
flabel metal3 s 591520 539140 592960 539380 0 FreeSans 1600 0 0 0 io_in_3v3[11]
port 109 nsew signal input
flabel metal3 s 591520 549068 592960 549308 0 FreeSans 1600 0 0 0 io_in[11]
port 57 nsew signal input
flabel metal3 s 591520 190204 592960 190444 0 FreeSans 1600 0 0 0 io_oeb[4]
port 155 nsew signal tristate
flabel metal3 s 591520 180276 592960 180516 0 FreeSans 1600 0 0 0 io_out[4]
port 96 nsew signal tristate
flabel metal3 s 591530 676993 592970 677233 0 FreeSans 1600 0 0 0 io_out[13]
port 62 nsew signal tristate
flabel metal3 591458 191182 591658 195982 0 FreeSans 4000 0 0 0 VSSD1
port 685 nsew
flabel metal3 591458 181142 591658 185931 0 FreeSans 4000 0 0 0 VSSD1
port 686 nsew
flabel metal3 566636 710520 571636 710720 0 FreeSans 4000 0 0 0 io_analog[1]
port 656 nsew
flabel metal3 464836 710520 469836 710720 0 FreeSans 4000 0 0 0 io_analog[2]
port 657 nsew
flabel metal3 413436 710520 418436 710720 0 FreeSans 4000 0 0 0 io_analog[3]
port 658 nsew
flabel metal3 119636 710520 124636 710720 0 FreeSans 4000 0 0 0 io_analog[7]
port 662 nsew
flabel metal3 68236 710520 73236 710720 0 FreeSans 4000 0 0 0 io_analog[8]
port 663 nsew
flabel metal3 16836 710520 21836 710720 0 FreeSans 4000 0 0 0 io_analog[9]
port 664 nsew
flabel metal3 171271 710520 173471 710720 0 FreeSans 1600 0 0 0 io_clamp_low[2]
port 673 nsew
flabel metal3 173670 710520 175870 710720 0 FreeSans 1600 0 0 0 io_clamp_high[2]
port 676 nsew
flabel metal3 176170 710521 180950 710721 0 FreeSans 4000 0 0 0 io_analog[6]
port 677 nsew
flabel metal3 166191 710521 170971 710721 0 FreeSans 4000 0 0 0 io_analog[6]
port 678 nsew
flabel metal3 217591 710521 222371 710721 0 FreeSans 4000 0 0 0 io_analog[6]
port 678 nsew
flabel metal3 227570 710521 232350 710721 0 FreeSans 4000 0 0 0 io_analog[5]
port 677 nsew
flabel metal3 222671 710520 224871 710720 0 FreeSans 1600 0 0 0 io_clamp_low[1]
port 673 nsew
flabel metal3 225070 710520 227270 710720 0 FreeSans 1600 0 0 0 io_clamp_high[1]
port 676 nsew
flabel metal3 510391 710434 515171 710634 0 FreeSans 8000 0 0 0 VSSA1
port 667 nsew
flabel metal3 520370 710434 525150 710634 0 FreeSans 8000 0 0 0 VSSA1
port 666 nsew
flabel metal3 591488 147003 591688 151783 0 FreeSans 4000 0 0 0 VSSA1
port 687 nsew
flabel metal3 591488 137024 591688 141804 0 FreeSans 4000 0 0 0 VSSA1
port 688 nsew
flabel metal3 591548 235203 591748 239983 0 FreeSans 4000 0 0 0 VDDA1
port 683 nsew
flabel metal3 591548 225224 591748 230004 0 FreeSans 4000 0 0 0 VDDA1
port 684 nsew
flabel metal3 591498 539824 591698 544604 0 FreeSans 4000 0 0 0 VDDA1
port 682 nsew
flabel metal3 591498 549803 591698 554583 0 FreeSans 4000 0 0 0 VDDA1
port 681 nsew
flabel metal3 591492 638982 591692 643782 0 FreeSans 4000 0 0 0 VCCD1
port 679 nsew
flabel metal3 591492 628942 591692 633731 0 FreeSans 4000 0 0 0 VCCD1
port 680 nsew
flabel metal3 -7720 633382 -7520 638182 0 FreeSans 4000 0 0 0 VCCD2
port 697 nsew
flabel metal3 -7720 643433 -7520 648222 0 FreeSans 4000 0 0 0 VCCD2
port 698 nsew
flabel metal3 -7760 558960 -7560 563740 0 FreeSans 4000 0 0 0 VSSA2
port 694 nsew
flabel metal3 -7760 548981 -7560 553761 0 FreeSans 4000 0 0 0 VSSA2
port 693 nsew
flabel metal3 -7714 204381 -7514 209161 0 FreeSans 4000 0 0 0 VDDA2
port 691 nsew
flabel metal3 -7714 214360 -7514 219140 0 FreeSans 4000 0 0 0 VDDA2
port 692 nsew
flabel metal2 s 6430 -960 6542 480 0 FreeSans 1600 90 0 0 wbs_we_i
port 654 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 1600 90 0 0 wbs_stb_i
port 653 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 1600 90 0 0 wbs_cyc_i
port 584 nsew signal input
flabel metal2 s 7626 -960 7738 480 0 FreeSans 1600 90 0 0 wbs_adr_i[0]
port 552 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 1600 90 0 0 wbs_ack_o
port 551 nsew signal tristate
flabel metal2 s 1646 -960 1758 480 0 FreeSans 1600 90 0 0 wb_rst_i
port 550 nsew signal input
flabel space 3823 979 9361 7624 0 FreeSans 16000 0 0 0 IO35
flabel metal3 319591 710521 324371 710721 0 FreeSans 4000 0 0 0 io_analog[4]
port 678 nsew
flabel metal3 329570 710521 334350 710721 0 FreeSans 4000 0 0 0 io_analog[4]
port 677 nsew
flabel metal3 324671 710520 326871 710720 0 FreeSans 1600 0 0 0 io_clamp_low[0]
port 673 nsew
flabel metal3 327070 710520 329270 710720 0 FreeSans 1600 0 0 0 io_clamp_high[0]
port 676 nsew
flabel metal3 591476 677938 591676 682938 0 FreeSans 4000 0 0 0 io_analog[0]
port 655 nsew
flabel metal3 -7746 681426 -7546 686426 0 FreeSans 4000 0 0 0 io_analog[10]
port 665 nsew
<< properties >>
string FIXED_BBOX -8844 -708 592926 712160
<< end >>
