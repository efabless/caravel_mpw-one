magic
tech sky130A
magscale 12 1
timestamp 1598776472
<< metal5 >>
rect 0 60 15 105
rect 30 60 45 75
rect 0 50 45 60
rect 0 45 40 50
rect 0 30 30 45
rect 0 25 40 30
rect 0 15 45 25
rect 0 0 15 15
rect 30 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
