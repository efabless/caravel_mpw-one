* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2
+ vssa2
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_oen_core[0] la_oen_core[100] la_oen_core[101] la_oen_core[102]
+ la_oen_core[103] la_oen_core[104] la_oen_core[105] la_oen_core[106] la_oen_core[107]
+ la_oen_core[108] la_oen_core[109] la_oen_core[10] la_oen_core[110] la_oen_core[111]
+ la_oen_core[112] la_oen_core[113] la_oen_core[114] la_oen_core[115] la_oen_core[116]
+ la_oen_core[117] la_oen_core[118] la_oen_core[119] la_oen_core[11] la_oen_core[120]
+ la_oen_core[121] la_oen_core[122] la_oen_core[123] la_oen_core[124] la_oen_core[125]
+ la_oen_core[126] la_oen_core[127] la_oen_core[12] la_oen_core[13] la_oen_core[14]
+ la_oen_core[15] la_oen_core[16] la_oen_core[17] la_oen_core[18] la_oen_core[19]
+ la_oen_core[1] la_oen_core[20] la_oen_core[21] la_oen_core[22] la_oen_core[23] la_oen_core[24]
+ la_oen_core[25] la_oen_core[26] la_oen_core[27] la_oen_core[28] la_oen_core[29]
+ la_oen_core[2] la_oen_core[30] la_oen_core[31] la_oen_core[32] la_oen_core[33] la_oen_core[34]
+ la_oen_core[35] la_oen_core[36] la_oen_core[37] la_oen_core[38] la_oen_core[39]
+ la_oen_core[3] la_oen_core[40] la_oen_core[41] la_oen_core[42] la_oen_core[43] la_oen_core[44]
+ la_oen_core[45] la_oen_core[46] la_oen_core[47] la_oen_core[48] la_oen_core[49]
+ la_oen_core[4] la_oen_core[50] la_oen_core[51] la_oen_core[52] la_oen_core[53] la_oen_core[54]
+ la_oen_core[55] la_oen_core[56] la_oen_core[57] la_oen_core[58] la_oen_core[59]
+ la_oen_core[5] la_oen_core[60] la_oen_core[61] la_oen_core[62] la_oen_core[63] la_oen_core[64]
+ la_oen_core[65] la_oen_core[66] la_oen_core[67] la_oen_core[68] la_oen_core[69]
+ la_oen_core[6] la_oen_core[70] la_oen_core[71] la_oen_core[72] la_oen_core[73] la_oen_core[74]
+ la_oen_core[75] la_oen_core[76] la_oen_core[77] la_oen_core[78] la_oen_core[79]
+ la_oen_core[7] la_oen_core[80] la_oen_core[81] la_oen_core[82] la_oen_core[83] la_oen_core[84]
+ la_oen_core[85] la_oen_core[86] la_oen_core[87] la_oen_core[88] la_oen_core[89]
+ la_oen_core[8] la_oen_core[90] la_oen_core[91] la_oen_core[92] la_oen_core[93] la_oen_core[94]
+ la_oen_core[95] la_oen_core[96] la_oen_core[97] la_oen_core[98] la_oen_core[99]
+ la_oen_core[9] la_oen_mprj[0] la_oen_mprj[100] la_oen_mprj[101] la_oen_mprj[102]
+ la_oen_mprj[103] la_oen_mprj[104] la_oen_mprj[105] la_oen_mprj[106] la_oen_mprj[107]
+ la_oen_mprj[108] la_oen_mprj[109] la_oen_mprj[10] la_oen_mprj[110] la_oen_mprj[111]
+ la_oen_mprj[112] la_oen_mprj[113] la_oen_mprj[114] la_oen_mprj[115] la_oen_mprj[116]
+ la_oen_mprj[117] la_oen_mprj[118] la_oen_mprj[119] la_oen_mprj[11] la_oen_mprj[120]
+ la_oen_mprj[121] la_oen_mprj[122] la_oen_mprj[123] la_oen_mprj[124] la_oen_mprj[125]
+ la_oen_mprj[126] la_oen_mprj[127] la_oen_mprj[12] la_oen_mprj[13] la_oen_mprj[14]
+ la_oen_mprj[15] la_oen_mprj[16] la_oen_mprj[17] la_oen_mprj[18] la_oen_mprj[19]
+ la_oen_mprj[1] la_oen_mprj[20] la_oen_mprj[21] la_oen_mprj[22] la_oen_mprj[23] la_oen_mprj[24]
+ la_oen_mprj[25] la_oen_mprj[26] la_oen_mprj[27] la_oen_mprj[28] la_oen_mprj[29]
+ la_oen_mprj[2] la_oen_mprj[30] la_oen_mprj[31] la_oen_mprj[32] la_oen_mprj[33] la_oen_mprj[34]
+ la_oen_mprj[35] la_oen_mprj[36] la_oen_mprj[37] la_oen_mprj[38] la_oen_mprj[39]
+ la_oen_mprj[3] la_oen_mprj[40] la_oen_mprj[41] la_oen_mprj[42] la_oen_mprj[43] la_oen_mprj[44]
+ la_oen_mprj[45] la_oen_mprj[46] la_oen_mprj[47] la_oen_mprj[48] la_oen_mprj[49]
+ la_oen_mprj[4] la_oen_mprj[50] la_oen_mprj[51] la_oen_mprj[52] la_oen_mprj[53] la_oen_mprj[54]
+ la_oen_mprj[55] la_oen_mprj[56] la_oen_mprj[57] la_oen_mprj[58] la_oen_mprj[59]
+ la_oen_mprj[5] la_oen_mprj[60] la_oen_mprj[61] la_oen_mprj[62] la_oen_mprj[63] la_oen_mprj[64]
+ la_oen_mprj[65] la_oen_mprj[66] la_oen_mprj[67] la_oen_mprj[68] la_oen_mprj[69]
+ la_oen_mprj[6] la_oen_mprj[70] la_oen_mprj[71] la_oen_mprj[72] la_oen_mprj[73] la_oen_mprj[74]
+ la_oen_mprj[75] la_oen_mprj[76] la_oen_mprj[77] la_oen_mprj[78] la_oen_mprj[79]
+ la_oen_mprj[7] la_oen_mprj[80] la_oen_mprj[81] la_oen_mprj[82] la_oen_mprj[83] la_oen_mprj[84]
+ la_oen_mprj[85] la_oen_mprj[86] la_oen_mprj[87] la_oen_mprj[88] la_oen_mprj[89]
+ la_oen_mprj[8] la_oen_mprj[90] la_oen_mprj[91] la_oen_mprj[92] la_oen_mprj[93] la_oen_mprj[94]
+ la_oen_mprj[95] la_oen_mprj[96] la_oen_mprj[97] la_oen_mprj[98] la_oen_mprj[99]
+ la_oen_mprj[9] mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12]
+ mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16]
+ mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20]
+ mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24]
+ mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28]
+ mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3]
+ mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8]
+ mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12]
+ mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16]
+ mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20]
+ mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24]
+ mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28]
+ mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3]
+ mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8]
+ mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_o_core[0] mprj_dat_o_core[10]
+ mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14]
+ mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18]
+ mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22]
+ mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26]
+ mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30]
+ mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6]
+ mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10]
+ mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14]
+ mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18]
+ mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22]
+ mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26]
+ mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30]
+ mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6]
+ mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_sel_o_core[0] mprj_sel_o_core[1]
+ mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2]
+ mprj_sel_o_user[3] mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user
+ user1_vcc_powergood user1_vdd_powergood user2_vcc_powergood user2_vdd_powergood
+ user_clock user_clock2 user_reset user_resetn vccd1 vssd1 vccd vssd vccd2 vssd2
+ vdda1 vssa1 vdda2 vssa2
XFILLER_11_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_432_ mprj_adr_o_core[25] vssd1 vssd1 vccd1 vccd1 _432_/Y sky130_fd_sc_hd__inv_2
X_501_ la_data_out_mprj[30] vssd1 vssd1 vccd1 vccd1 _501_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[299\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[299\]/HI mprj_logic_high\[299\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[36\] _507_/Y la_buf\[36\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[36]
+ sky130_fd_sc_hd__einvp_8
X_363_ la_oen_mprj[95] vssd1 vssd1 vccd1 vccd1 _363_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] mprj_logic_high\[355\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[25\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_2063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[76\] _344_/Y mprj_logic_high\[278\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[214\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[214\]/HI mprj_logic_high\[214\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[24\] _463_/Y mprj_dat_buf\[24\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_415_ mprj_adr_o_core[8] vssd1 vssd1 vccd1 vccd1 _415_/Y sky130_fd_sc_hd__inv_2
X_346_ la_oen_mprj[78] vssd1 vssd1 vccd1 vccd1 _346_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[75\] vssd1 vssd1 vccd1 vccd1 la_buf\[1\]/TE mprj_logic_high\[75\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[429\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[429\]/HI mprj_logic_high\[429\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[164\] vssd1 vssd1 vccd1 vccd1 la_buf\[90\]/TE mprj_logic_high\[164\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[331\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[331\]/HI mprj_logic_high\[331\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] mprj_logic_high\[422\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[92\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[39\] _638_/Y mprj_logic_high\[241\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[39] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[109\] _377_/Y mprj_logic_high\[311\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_1_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[281\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[281\]/HI mprj_logic_high\[281\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[379\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[379\]/HI mprj_logic_high\[379\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[62] sky130_fd_sc_hd__inv_8
XFILLER_15_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_2086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[38\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[28\]/TE mprj_logic_high\[38\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[127\] vssd1 vssd1 vccd1 vccd1 la_buf\[53\]/TE mprj_logic_high\[127\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xla_buf\[66\] _537_/Y la_buf\[66\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[66]
+ sky130_fd_sc_hd__einvp_8
X_594_ la_data_out_mprj[123] vssd1 vssd1 vccd1 vccd1 _594_/Y sky130_fd_sc_hd__inv_2
XPHY_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[122\] _593_/Y la_buf\[122\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[122]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_5 la_oen_mprj[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] mprj_logic_high\[385\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[55\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[244\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[244\]/HI mprj_logic_high\[244\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[411\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[411\]/HI mprj_logic_high\[411\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_577_ la_data_out_mprj[106] vssd1 vssd1 vccd1 vccd1 _577_/Y sky130_fd_sc_hd__inv_2
X_646_ la_oen_mprj[47] vssd1 vssd1 vccd1 vccd1 _646_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[25] sky130_fd_sc_hd__inv_8
XPHY_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_500_ la_data_out_mprj[29] vssd1 vssd1 vccd1 vccd1 _500_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[3\] _602_/Y mprj_logic_high\[205\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[3] sky130_fd_sc_hd__einvp_8
X_431_ mprj_adr_o_core[24] vssd1 vssd1 vccd1 vccd1 _431_/Y sky130_fd_sc_hd__inv_2
X_362_ la_oen_mprj[94] vssd1 vssd1 vccd1 vccd1 _362_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[21\] _620_/Y mprj_logic_high\[223\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[21] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[361\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[361\]/HI mprj_logic_high\[361\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[194\] vssd1 vssd1 vccd1 vccd1 la_buf\[120\]/TE mprj_logic_high\[194\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[29\] _500_/Y la_buf\[29\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_629_ la_oen_mprj[30] vssd1 vssd1 vccd1 vccd1 _629_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] mprj_logic_high\[348\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[18\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[20\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[10\]/TE mprj_logic_high\[20\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[69\] _337_/Y mprj_logic_high\[271\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[69] sky130_fd_sc_hd__einvp_8
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[17\] _456_/Y mprj_dat_buf\[17\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[207\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[207\]/HI mprj_logic_high\[207\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_414_ mprj_adr_o_core[7] vssd1 vssd1 vccd1 vccd1 _414_/Y sky130_fd_sc_hd__inv_2
X_345_ la_oen_mprj[77] vssd1 vssd1 vccd1 vccd1 _345_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[12\] _419_/Y mprj_adr_buf\[12\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[92] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[126] sky130_fd_sc_hd__inv_8
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[68\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[26\]/TE mprj_logic_high\[68\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[324\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[324\]/HI mprj_logic_high\[324\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[157\] vssd1 vssd1 vccd1 vccd1 la_buf\[83\]/TE mprj_logic_high\[157\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[96\] _567_/Y la_buf\[96\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[96]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] mprj_logic_high\[415\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[85\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[274\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[274\]/HI mprj_logic_high\[274\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[441\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[441\]/HI mprj_logic_high\[441\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[7\] _478_/Y la_buf\[7\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[7] sky130_fd_sc_hd__einvp_8
Xla_buf\[11\] _482_/Y la_buf\[11\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[11]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[4\] _411_/Y mprj_adr_buf\[4\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[55] sky130_fd_sc_hd__inv_8
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] mprj_logic_high\[441\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[111\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[121\] _389_/Y mprj_logic_high\[323\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[121] sky130_fd_sc_hd__einvp_8
XFILLER_4_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_sel_buf\[2\] _405_/Y mprj_sel_buf\[2\]/TE vssd1 vssd1 vccd1 vccd1 mprj_sel_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[51\] _650_/Y mprj_logic_high\[253\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[51] sky130_fd_sc_hd__einvp_8
XPHY_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[391\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[391\]/HI mprj_logic_high\[391\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[59\] _530_/Y la_buf\[59\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[59]
+ sky130_fd_sc_hd__einvp_8
X_593_ la_data_out_mprj[122] vssd1 vssd1 vccd1 vccd1 _593_/Y sky130_fd_sc_hd__inv_2
XPHY_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_6 la_oen_mprj[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[115\] _586_/Y la_buf\[115\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[115]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] mprj_logic_high\[378\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[48\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[50\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[8\]/TE mprj_logic_high\[50\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[99\] _367_/Y mprj_logic_high\[301\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[237\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[237\]/HI mprj_logic_high\[237\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[404\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[404\]/HI mprj_logic_high\[404\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj2_vdd_pwrgood mprj2_pwrgood/A vssd1 vssd1 vccd1 vccd1 user2_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_645_ la_oen_mprj[46] vssd1 vssd1 vccd1 vccd1 _645_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_576_ la_data_out_mprj[105] vssd1 vssd1 vccd1 vccd1 _576_/Y sky130_fd_sc_hd__inv_2
XPHY_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[18] sky130_fd_sc_hd__inv_8
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[98\] vssd1 vssd1 vccd1 vccd1 la_buf\[24\]/TE mprj_logic_high\[98\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[187\] vssd1 vssd1 vccd1 vccd1 la_buf\[113\]/TE mprj_logic_high\[187\]/LO
+ sky130_fd_sc_hd__conb_1
X_430_ mprj_adr_o_core[23] vssd1 vssd1 vccd1 vccd1 _430_/Y sky130_fd_sc_hd__inv_2
X_361_ la_oen_mprj[93] vssd1 vssd1 vccd1 vccd1 _361_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[14\] _613_/Y mprj_logic_high\[216\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[354\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[354\]/HI mprj_logic_high\[354\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_628_ la_oen_mprj[29] vssd1 vssd1 vccd1 vccd1 _628_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_559_ la_data_out_mprj[88] vssd1 vssd1 vccd1 vccd1 _559_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[13\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[3\]/TE mprj_logic_high\[13\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[102\] vssd1 vssd1 vccd1 vccd1 la_buf\[28\]/TE mprj_logic_high\[102\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_413_ mprj_adr_o_core[6] vssd1 vssd1 vccd1 vccd1 _413_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xla_buf\[41\] _512_/Y la_buf\[41\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[41]
+ sky130_fd_sc_hd__einvp_8
X_344_ la_oen_mprj[76] vssd1 vssd1 vccd1 vccd1 _344_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[85] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[119] sky130_fd_sc_hd__inv_8
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] mprj_logic_high\[360\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[30\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[317\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[317\]/HI mprj_logic_high\[317\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[81\] _349_/Y mprj_logic_high\[283\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[89\] _560_/Y la_buf\[89\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[89]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] mprj_logic_high\[408\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[78\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[80\] vssd1 vssd1 vccd1 vccd1 la_buf\[6\]/TE mprj_logic_high\[80\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[267\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[267\]/HI mprj_logic_high\[267\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[434\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[434\]/HI mprj_logic_high\[434\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[48] sky130_fd_sc_hd__inv_8
XFILLER_15_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] mprj_logic_high\[434\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[104\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[114\] _382_/Y mprj_logic_high\[316\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[44\] _643_/Y mprj_logic_high\[246\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_592_ la_data_out_mprj[121] vssd1 vssd1 vccd1 vccd1 _592_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[384\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[384\]/HI mprj_logic_high\[384\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 la_oen_mprj[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xla_buf\[108\] _579_/Y la_buf\[108\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[108]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[101] sky130_fd_sc_hd__inv_8
XFILLER_1_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[0\] _439_/Y mprj_dat_buf\[0\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[43\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[1\]/TE mprj_logic_high\[43\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[132\] vssd1 vssd1 vccd1 vccd1 la_buf\[58\]/TE mprj_logic_high\[132\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xla_buf\[71\] _542_/Y la_buf\[71\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[71]
+ sky130_fd_sc_hd__einvp_8
X_575_ la_data_out_mprj[104] vssd1 vssd1 vccd1 vccd1 _575_/Y sky130_fd_sc_hd__inv_2
X_644_ la_oen_mprj[45] vssd1 vssd1 vccd1 vccd1 _644_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] mprj_logic_high\[390\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[60\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_360_ la_oen_mprj[92] vssd1 vssd1 vccd1 vccd1 _360_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[347\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[347\]/HI mprj_logic_high\[347\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_558_ la_data_out_mprj[87] vssd1 vssd1 vccd1 vccd1 _558_/Y sky130_fd_sc_hd__inv_2
X_627_ la_oen_mprj[28] vssd1 vssd1 vccd1 vccd1 _627_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_489_ la_data_out_mprj[18] vssd1 vssd1 vccd1 vccd1 _489_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[30] sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[8\] vssd1 vssd1 vccd1 vccd1 mprj_sel_buf\[2\]/TE mprj_logic_high\[8\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[297\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[297\]/HI mprj_logic_high\[297\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_412_ mprj_adr_o_core[5] vssd1 vssd1 vccd1 vccd1 _412_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[34\] _505_/Y la_buf\[34\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[34]
+ sky130_fd_sc_hd__einvp_8
X_343_ la_oen_mprj[75] vssd1 vssd1 vccd1 vccd1 _343_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[78] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] mprj_logic_high\[353\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[23\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[74\] _342_/Y mprj_logic_high\[276\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[74] sky130_fd_sc_hd__einvp_8
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[212\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[212\]/HI mprj_logic_high\[212\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[22\] _461_/Y mprj_dat_buf\[22\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[73\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[31\]/TE mprj_logic_high\[73\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[427\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[427\]/HI mprj_logic_high\[427\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[162\] vssd1 vssd1 vccd1 vccd1 la_buf\[88\]/TE mprj_logic_high\[162\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] mprj_logic_high\[420\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[90\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[107\] _375_/Y mprj_logic_high\[309\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[107] sky130_fd_sc_hd__einvp_8
X_660_ la_oen_mprj[61] vssd1 vssd1 vccd1 vccd1 _660_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[37\] _636_/Y mprj_logic_high\[239\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[37] sky130_fd_sc_hd__einvp_8
X_591_ la_data_out_mprj[120] vssd1 vssd1 vccd1 vccd1 _591_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[377\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[377\]/HI mprj_logic_high\[377\]/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_8 la_oen_mprj[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[60] sky130_fd_sc_hd__inv_8
XFILLER_15_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[36\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[26\]/TE mprj_logic_high\[36\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[125\] vssd1 vssd1 vccd1 vccd1 la_buf\[51\]/TE mprj_logic_high\[125\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[64\] _535_/Y la_buf\[64\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[64]
+ sky130_fd_sc_hd__einvp_8
X_574_ la_data_out_mprj[103] vssd1 vssd1 vccd1 vccd1 _574_/Y sky130_fd_sc_hd__inv_2
X_643_ la_oen_mprj[44] vssd1 vssd1 vccd1 vccd1 _643_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_adr_buf\[28\] _435_/Y mprj_adr_buf\[28\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[28]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[120\] _591_/Y la_buf\[120\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[120]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] mprj_logic_high\[383\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[53\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[242\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[242\]/HI mprj_logic_high\[242\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_557_ la_data_out_mprj[86] vssd1 vssd1 vccd1 vccd1 _557_/Y sky130_fd_sc_hd__inv_2
X_488_ la_data_out_mprj[17] vssd1 vssd1 vccd1 vccd1 _488_/Y sky130_fd_sc_hd__inv_2
X_626_ la_oen_mprj[27] vssd1 vssd1 vccd1 vccd1 _626_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[23] sky130_fd_sc_hd__inv_8
XFILLER_1_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[192\] vssd1 vssd1 vccd1 vccd1 la_buf\[118\]/TE mprj_logic_high\[192\]/LO
+ sky130_fd_sc_hd__conb_1
X_411_ mprj_adr_o_core[4] vssd1 vssd1 vccd1 vccd1 _411_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[1\] _600_/Y mprj_logic_high\[203\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[1] sky130_fd_sc_hd__einvp_8
X_342_ la_oen_mprj[74] vssd1 vssd1 vccd1 vccd1 _342_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[457\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[457\]/HI mprj_logic_high\[457\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[27\] _498_/Y la_buf\[27\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[27]
+ sky130_fd_sc_hd__einvp_8
X_609_ la_oen_mprj[10] vssd1 vssd1 vccd1 vccd1 _609_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] mprj_logic_high\[346\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[16\]/Y sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] mprj_logic_high\[457\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[127\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[67\] _335_/Y mprj_logic_high\[269\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[67] sky130_fd_sc_hd__einvp_8
XFILLER_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[15\] _454_/Y mprj_dat_buf\[15\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[15]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[205\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[205\]/HI mprj_logic_high\[205\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[10\] _417_/Y mprj_adr_buf\[10\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[90] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[124] sky130_fd_sc_hd__inv_8
XFILLER_4_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[66\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[24\]/TE mprj_logic_high\[66\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[322\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[322\]/HI mprj_logic_high\[322\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[155\] vssd1 vssd1 vccd1 vccd1 la_buf\[81\]/TE mprj_logic_high\[155\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[94\] _565_/Y la_buf\[94\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[94]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] mprj_logic_high\[413\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[83\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_590_ la_data_out_mprj[119] vssd1 vssd1 vccd1 vccd1 _590_/Y sky130_fd_sc_hd__inv_2
XPHY_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[272\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[272\]/HI mprj_logic_high\[272\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[5\] _476_/Y la_buf\[5\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[5] sky130_fd_sc_hd__einvp_8
XFILLER_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 la_oen_mprj[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[2\] _409_/Y mprj_adr_buf\[2\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[53] sky130_fd_sc_hd__inv_8
XFILLER_15_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[29\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[19\]/TE mprj_logic_high\[29\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_sel_buf\[0\] _403_/Y mprj_sel_buf\[0\]/TE vssd1 vssd1 vccd1 vccd1 mprj_sel_o_user[0]
+ sky130_fd_sc_hd__einvp_8
X_642_ la_oen_mprj[43] vssd1 vssd1 vccd1 vccd1 _642_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[118\] vssd1 vssd1 vccd1 vccd1 la_buf\[44\]/TE mprj_logic_high\[118\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[57\] _528_/Y la_buf\[57\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[57]
+ sky130_fd_sc_hd__einvp_8
XPHY_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_573_ la_data_out_mprj[102] vssd1 vssd1 vccd1 vccd1 _573_/Y sky130_fd_sc_hd__inv_2
XPHY_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[113\] _584_/Y la_buf\[113\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[113]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] mprj_logic_high\[376\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[46\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_2130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] mprj_logic_high\[338\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[8\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[97\] _365_/Y mprj_logic_high\[299\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[97] sky130_fd_sc_hd__einvp_8
XFILLER_10_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[235\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[235\]/HI mprj_logic_high\[235\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[402\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[402\]/HI mprj_logic_high\[402\]/LO
+ sky130_fd_sc_hd__conb_1
X_625_ la_oen_mprj[26] vssd1 vssd1 vccd1 vccd1 _625_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_487_ la_data_out_mprj[16] vssd1 vssd1 vccd1 vccd1 _487_/Y sky130_fd_sc_hd__inv_2
X_556_ la_data_out_mprj[85] vssd1 vssd1 vccd1 vccd1 _556_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[16] sky130_fd_sc_hd__inv_8
XFILLER_5_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[96\] vssd1 vssd1 vccd1 vccd1 la_buf\[22\]/TE mprj_logic_high\[96\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[185\] vssd1 vssd1 vccd1 vccd1 la_buf\[111\]/TE mprj_logic_high\[185\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[12\] _611_/Y mprj_logic_high\[214\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[12] sky130_fd_sc_hd__einvp_8
X_410_ mprj_adr_o_core[3] vssd1 vssd1 vccd1 vccd1 _410_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[8] sky130_fd_sc_hd__inv_8
X_341_ la_oen_mprj[73] vssd1 vssd1 vccd1 vccd1 _341_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[352\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[352\]/HI mprj_logic_high\[352\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_stb_buf _401_/Y mprj_stb_buf/TE vssd1 vssd1 vccd1 vccd1 mprj_stb_o_user sky130_fd_sc_hd__einvp_8
XFILLER_2_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_608_ la_oen_mprj[9] vssd1 vssd1 vccd1 vccd1 _608_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_539_ la_data_out_mprj[68] vssd1 vssd1 vccd1 vccd1 _539_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[11\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[1\]/TE mprj_logic_high\[11\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[100\] vssd1 vssd1 vccd1 vccd1 la_buf\[26\]/TE mprj_logic_high\[100\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[83] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[117] sky130_fd_sc_hd__inv_8
XFILLER_0_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[59\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[17\]/TE mprj_logic_high\[59\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[148\] vssd1 vssd1 vccd1 vccd1 la_buf\[74\]/TE mprj_logic_high\[148\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[315\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[315\]/HI mprj_logic_high\[315\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[87\] _558_/Y la_buf\[87\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[87]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] mprj_logic_high\[406\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[76\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[265\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[265\]/HI mprj_logic_high\[265\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[432\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[432\]/HI mprj_logic_high\[432\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[46] sky130_fd_sc_hd__inv_8
XFILLER_15_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] mprj_logic_high\[432\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[102\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[112\] _380_/Y mprj_logic_high\[314\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[112] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[42\] _641_/Y mprj_logic_high\[244\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[42] sky130_fd_sc_hd__einvp_8
X_572_ la_data_out_mprj[101] vssd1 vssd1 vccd1 vccd1 _572_/Y sky130_fd_sc_hd__inv_2
X_641_ la_oen_mprj[42] vssd1 vssd1 vccd1 vccd1 _641_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[382\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[382\]/HI mprj_logic_high\[382\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[106\] _577_/Y la_buf\[106\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[106]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] mprj_logic_high\[369\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[39\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[41\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[31\]/TE mprj_logic_high\[41\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[130\] vssd1 vssd1 vccd1 vccd1 la_buf\[56\]/TE mprj_logic_high\[130\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[228\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[228\]/HI mprj_logic_high\[228\]/LO
+ sky130_fd_sc_hd__conb_1
X_555_ la_data_out_mprj[84] vssd1 vssd1 vccd1 vccd1 _555_/Y sky130_fd_sc_hd__inv_2
X_624_ la_oen_mprj[25] vssd1 vssd1 vccd1 vccd1 _624_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_we_buf _402_/Y mprj_we_buf/TE vssd1 vssd1 vccd1 vccd1 mprj_we_o_user sky130_fd_sc_hd__einvp_8
XFILLER_12_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_486_ la_data_out_mprj[15] vssd1 vssd1 vccd1 vccd1 _486_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_pwrgood mprj_pwrgood/A vssd1 vssd1 vccd1 vccd1 user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_4_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[178\] vssd1 vssd1 vccd1 vccd1 la_buf\[104\]/TE mprj_logic_high\[178\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[89\] vssd1 vssd1 vccd1 vccd1 la_buf\[15\]/TE mprj_logic_high\[89\]/LO
+ sky130_fd_sc_hd__conb_1
X_340_ la_oen_mprj[72] vssd1 vssd1 vccd1 vccd1 _340_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[345\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[345\]/HI mprj_logic_high\[345\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_538_ la_data_out_mprj[67] vssd1 vssd1 vccd1 vccd1 _538_/Y sky130_fd_sc_hd__inv_2
X_607_ la_oen_mprj[8] vssd1 vssd1 vccd1 vccd1 _607_/Y sky130_fd_sc_hd__inv_2
X_469_ mprj_dat_o_core[30] vssd1 vssd1 vccd1 vccd1 _469_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[6\] vssd1 vssd1 vccd1 vccd1 mprj_sel_buf\[0\]/TE mprj_logic_high\[6\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[295\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[295\]/HI mprj_logic_high\[295\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[32\] _503_/Y la_buf\[32\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[32]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[76] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] mprj_logic_high\[351\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[21\]/Y sky130_fd_sc_hd__nand2_4
Xmprj_dat_buf\[9\] _448_/Y mprj_dat_buf\[9\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[72\] _340_/Y mprj_logic_high\[274\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[72] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[210\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[210\]/HI mprj_logic_high\[210\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[20\] _459_/Y mprj_dat_buf\[20\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[20]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[308\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[308\]/HI mprj_logic_high\[308\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] mprj_logic_high\[399\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[69\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[71\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[29\]/TE mprj_logic_high\[71\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[258\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[258\]/HI mprj_logic_high\[258\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[160\] vssd1 vssd1 vccd1 vccd1 la_buf\[86\]/TE mprj_logic_high\[160\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[425\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[425\]/HI mprj_logic_high\[425\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_2078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[39] sky130_fd_sc_hd__inv_8
XFILLER_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[105\] _373_/Y mprj_logic_high\[307\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[105] sky130_fd_sc_hd__einvp_8
XFILLER_2_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[35\] _634_/Y mprj_logic_high\[237\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[35] sky130_fd_sc_hd__einvp_8
X_571_ la_data_out_mprj[100] vssd1 vssd1 vccd1 vccd1 _571_/Y sky130_fd_sc_hd__inv_2
X_640_ la_oen_mprj[41] vssd1 vssd1 vccd1 vccd1 _640_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[375\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[375\]/HI mprj_logic_high\[375\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[34\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[24\]/TE mprj_logic_high\[34\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[123\] vssd1 vssd1 vccd1 vccd1 la_buf\[49\]/TE mprj_logic_high\[123\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[62\] _533_/Y la_buf\[62\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[62]
+ sky130_fd_sc_hd__einvp_8
X_485_ la_data_out_mprj[14] vssd1 vssd1 vccd1 vccd1 _485_/Y sky130_fd_sc_hd__inv_2
X_554_ la_data_out_mprj[83] vssd1 vssd1 vccd1 vccd1 _554_/Y sky130_fd_sc_hd__inv_2
X_623_ la_oen_mprj[24] vssd1 vssd1 vccd1 vccd1 _623_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[26\] _433_/Y mprj_adr_buf\[26\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] mprj_logic_high\[381\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[51\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[240\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[240\]/HI mprj_logic_high\[240\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[338\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[338\]/HI mprj_logic_high\[338\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_468_ mprj_dat_o_core[29] vssd1 vssd1 vccd1 vccd1 _468_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_537_ la_data_out_mprj[66] vssd1 vssd1 vccd1 vccd1 _537_/Y sky130_fd_sc_hd__inv_2
X_606_ la_oen_mprj[7] vssd1 vssd1 vccd1 vccd1 _606_/Y sky130_fd_sc_hd__inv_2
X_399_ caravel_clk2 vssd1 vssd1 vccd1 vccd1 _399_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[21] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] mprj_logic_high\[429\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[99\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[288\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[288\]/HI mprj_logic_high\[288\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[190\] vssd1 vssd1 vccd1 vccd1 la_buf\[116\]/TE mprj_logic_high\[190\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_2110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[455\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[455\]/HI mprj_logic_high\[455\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xla_buf\[25\] _496_/Y la_buf\[25\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[69] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] mprj_logic_high\[344\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[14\]/Y sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] mprj_logic_high\[455\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[125\]/Y sky130_fd_sc_hd__nand2_4
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[65\] _333_/Y mprj_logic_high\[267\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[13\] _452_/Y mprj_dat_buf\[13\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[203\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[203\]/HI mprj_logic_high\[203\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[122] sky130_fd_sc_hd__inv_8
XFILLER_0_2016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[64\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[22\]/TE mprj_logic_high\[64\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[320\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[320\]/HI mprj_logic_high\[320\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[153\] vssd1 vssd1 vccd1 vccd1 la_buf\[79\]/TE mprj_logic_high\[153\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[418\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[418\]/HI mprj_logic_high\[418\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[92\] _563_/Y la_buf\[92\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[92]
+ sky130_fd_sc_hd__einvp_8
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A vssd1 vssd1 vccd1 vccd1 user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_1_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] mprj_logic_high\[411\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[81\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[28\] _627_/Y mprj_logic_high\[230\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[28] sky130_fd_sc_hd__einvp_8
XPHY_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_570_ la_data_out_mprj[99] vssd1 vssd1 vccd1 vccd1 _570_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[270\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[270\]/HI mprj_logic_high\[270\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[368\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[368\]/HI mprj_logic_high\[368\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[3\] _474_/Y la_buf\[3\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[3] sky130_fd_sc_hd__einvp_8
XFILLER_4_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_2144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[0\] _407_/Y mprj_adr_buf\[0\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[51] sky130_fd_sc_hd__inv_8
XFILLER_15_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[27\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[17\]/TE mprj_logic_high\[27\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[116\] vssd1 vssd1 vccd1 vccd1 la_buf\[42\]/TE mprj_logic_high\[116\]/LO
+ sky130_fd_sc_hd__conb_1
X_622_ la_oen_mprj[23] vssd1 vssd1 vccd1 vccd1 _622_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[55\] _526_/Y la_buf\[55\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[55]
+ sky130_fd_sc_hd__einvp_8
X_484_ la_data_out_mprj[13] vssd1 vssd1 vccd1 vccd1 _484_/Y sky130_fd_sc_hd__inv_2
X_553_ la_data_out_mprj[82] vssd1 vssd1 vccd1 vccd1 _553_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[19\] _426_/Y mprj_adr_buf\[19\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[19]
+ sky130_fd_sc_hd__einvp_8
XFILLER_10_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[111\] _582_/Y la_buf\[111\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[111]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[99] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] mprj_logic_high\[374\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[44\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] mprj_logic_high\[336\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[6\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[95\] _363_/Y mprj_logic_high\[297\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[233\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[233\]/HI mprj_logic_high\[233\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[400\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[400\]/HI mprj_logic_high\[400\]/LO
+ sky130_fd_sc_hd__conb_1
X_605_ la_oen_mprj[6] vssd1 vssd1 vccd1 vccd1 _605_/Y sky130_fd_sc_hd__inv_2
X_467_ mprj_dat_o_core[28] vssd1 vssd1 vccd1 vccd1 _467_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_398_ caravel_clk vssd1 vssd1 vccd1 vccd1 _398_/Y sky130_fd_sc_hd__inv_2
X_536_ la_data_out_mprj[65] vssd1 vssd1 vccd1 vccd1 _536_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[14] sky130_fd_sc_hd__inv_8
XFILLER_4_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[94\] vssd1 vssd1 vccd1 vccd1 la_buf\[20\]/TE mprj_logic_high\[94\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[6] sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[183\] vssd1 vssd1 vccd1 vccd1 la_buf\[109\]/TE mprj_logic_high\[183\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[10\] _609_/Y mprj_logic_high\[212\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_13_2133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[448\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[448\]/HI mprj_logic_high\[448\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[350\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[350\]/HI mprj_logic_high\[350\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[18\] _489_/Y la_buf\[18\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[18]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_519_ la_data_out_mprj[48] vssd1 vssd1 vccd1 vccd1 _519_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] mprj_logic_high\[448\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[118\]/Y sky130_fd_sc_hd__nand2_4
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[58\] _657_/Y mprj_logic_high\[260\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[58] sky130_fd_sc_hd__einvp_8
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[398\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[398\]/HI mprj_logic_high\[398\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[81] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[115] sky130_fd_sc_hd__inv_8
XFILLER_14_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[57\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[15\]/TE mprj_logic_high\[57\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[146\] vssd1 vssd1 vccd1 vccd1 la_buf\[72\]/TE mprj_logic_high\[146\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[313\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[313\]/HI mprj_logic_high\[313\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[85\] _556_/Y la_buf\[85\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[85]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] mprj_logic_high\[404\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[74\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[263\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[263\]/HI mprj_logic_high\[263\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[430\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[430\]/HI mprj_logic_high\[430\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_2134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[44] sky130_fd_sc_hd__inv_8
XFILLER_15_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] mprj_logic_high\[430\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[100\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[110\] _378_/Y mprj_logic_high\[312\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[110] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[40\] _639_/Y mprj_logic_high\[242\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[40] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[109\] vssd1 vssd1 vccd1 vccd1 la_buf\[35\]/TE mprj_logic_high\[109\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_621_ la_oen_mprj[22] vssd1 vssd1 vccd1 vccd1 _621_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[380\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[380\]/HI mprj_logic_high\[380\]/LO
+ sky130_fd_sc_hd__conb_1
X_483_ la_data_out_mprj[12] vssd1 vssd1 vccd1 vccd1 _483_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[48\] _519_/Y la_buf\[48\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[48]
+ sky130_fd_sc_hd__einvp_8
X_552_ la_data_out_mprj[81] vssd1 vssd1 vccd1 vccd1 _552_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[104\] _575_/Y la_buf\[104\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[104]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] mprj_logic_high\[367\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[37\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[88\] _356_/Y mprj_logic_high\[290\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[88] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[226\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[226\]/HI mprj_logic_high\[226\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_535_ la_data_out_mprj[64] vssd1 vssd1 vccd1 vccd1 _535_/Y sky130_fd_sc_hd__inv_2
X_604_ la_oen_mprj[5] vssd1 vssd1 vccd1 vccd1 _604_/Y sky130_fd_sc_hd__inv_2
X_466_ mprj_dat_o_core[27] vssd1 vssd1 vccd1 vccd1 _466_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_397_ user_resetn vssd1 vssd1 vccd1 vccd1 user_reset sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[31\] _438_/Y mprj_adr_buf\[31\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[176\] vssd1 vssd1 vccd1 vccd1 la_buf\[102\]/TE mprj_logic_high\[176\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[87\] vssd1 vssd1 vccd1 vccd1 la_buf\[13\]/TE mprj_logic_high\[87\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[343\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[343\]/HI mprj_logic_high\[343\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_2092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_518_ la_data_out_mprj[47] vssd1 vssd1 vccd1 vccd1 _518_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_449_ mprj_dat_o_core[10] vssd1 vssd1 vccd1 vccd1 _449_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[4\] vssd1 vssd1 vccd1 vccd1 mprj_stb_buf/TE mprj_logic_high\[4\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[293\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[293\]/HI mprj_logic_high\[293\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[30\] _501_/Y la_buf\[30\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_13_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[108] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[74] sky130_fd_sc_hd__inv_8
Xmprj_dat_buf\[7\] _446_/Y mprj_dat_buf\[7\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XPHY_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[70\] _338_/Y mprj_logic_high\[272\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[70] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[139\] vssd1 vssd1 vccd1 vccd1 la_buf\[65\]/TE mprj_logic_high\[139\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[306\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[306\]/HI mprj_logic_high\[306\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[78\] _549_/Y la_buf\[78\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[78]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] mprj_logic_high\[397\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[67\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_2092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[256\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[256\]/HI mprj_logic_high\[256\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[423\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[423\]/HI mprj_logic_high\[423\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[37] sky130_fd_sc_hd__inv_8
XFILLER_8_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[103\] _371_/Y mprj_logic_high\[305\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[103] sky130_fd_sc_hd__einvp_8
XFILLER_2_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[33\] _632_/Y mprj_logic_high\[235\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[33] sky130_fd_sc_hd__einvp_8
X_551_ la_data_out_mprj[80] vssd1 vssd1 vccd1 vccd1 _551_/Y sky130_fd_sc_hd__inv_2
X_620_ la_oen_mprj[21] vssd1 vssd1 vccd1 vccd1 _620_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[373\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[373\]/HI mprj_logic_high\[373\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_482_ la_data_out_mprj[11] vssd1 vssd1 vccd1 vccd1 _482_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[32\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[22\]/TE mprj_logic_high\[32\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[29\] _468_/Y mprj_dat_buf\[29\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[29]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[219\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[219\]/HI mprj_logic_high\[219\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[121\] vssd1 vssd1 vccd1 vccd1 la_buf\[47\]/TE mprj_logic_high\[121\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[60\] _531_/Y la_buf\[60\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[60]
+ sky130_fd_sc_hd__einvp_8
X_465_ mprj_dat_o_core[26] vssd1 vssd1 vccd1 vccd1 _465_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_534_ la_data_out_mprj[63] vssd1 vssd1 vccd1 vccd1 _534_/Y sky130_fd_sc_hd__inv_2
X_603_ la_oen_mprj[4] vssd1 vssd1 vccd1 vccd1 _603_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_396_ caravel_rstn vssd1 vssd1 vccd1 vccd1 _396_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[24\] _431_/Y mprj_adr_buf\[24\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[169\] vssd1 vssd1 vccd1 vccd1 la_buf\[95\]/TE mprj_logic_high\[169\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[336\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[336\]/HI mprj_logic_high\[336\]/LO
+ sky130_fd_sc_hd__conb_1
X_448_ mprj_dat_o_core[9] vssd1 vssd1 vccd1 vccd1 _448_/Y sky130_fd_sc_hd__inv_2
X_517_ la_data_out_mprj[46] vssd1 vssd1 vccd1 vccd1 _517_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_379_ la_oen_mprj[111] vssd1 vssd1 vccd1 vccd1 _379_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] mprj_logic_high\[427\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[97\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[286\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[286\]/HI mprj_logic_high\[286\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[453\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[453\]/HI mprj_logic_high\[453\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[23\] _494_/Y la_buf\[23\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[23]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[67] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] mprj_logic_high\[342\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[12\]/Y sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] mprj_logic_high\[453\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[123\]/Y sky130_fd_sc_hd__nand2_4
XPHY_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[63\] _331_/Y mprj_logic_high\[265\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[63] sky130_fd_sc_hd__einvp_8
XFILLER_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[11\] _450_/Y mprj_dat_buf\[11\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[11]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[201\] vssd1 vssd1 vccd1 vccd1 la_buf\[127\]/TE mprj_logic_high\[201\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_2016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[127\] _598_/Y la_buf\[127\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[127]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[120] sky130_fd_sc_hd__inv_8
XFILLER_0_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[62\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[20\]/TE mprj_logic_high\[62\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[249\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[249\]/HI mprj_logic_high\[249\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[151\] vssd1 vssd1 vccd1 vccd1 la_buf\[77\]/TE mprj_logic_high\[151\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[416\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[416\]/HI mprj_logic_high\[416\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[90\] _561_/Y la_buf\[90\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[90]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_2136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[8\] _607_/Y mprj_logic_high\[210\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[8] sky130_fd_sc_hd__einvp_8
X_481_ la_data_out_mprj[10] vssd1 vssd1 vccd1 vccd1 _481_/Y sky130_fd_sc_hd__inv_2
X_550_ la_data_out_mprj[79] vssd1 vssd1 vccd1 vccd1 _550_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[199\] vssd1 vssd1 vccd1 vccd1 la_buf\[125\]/TE mprj_logic_high\[199\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[26\] _625_/Y mprj_logic_high\[228\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[366\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[366\]/HI mprj_logic_high\[366\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[1\] _472_/Y la_buf\[1\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_5_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[25\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[15\]/TE mprj_logic_high\[25\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[114\] vssd1 vssd1 vccd1 vccd1 la_buf\[40\]/TE mprj_logic_high\[114\]/LO
+ sky130_fd_sc_hd__conb_1
X_602_ la_oen_mprj[3] vssd1 vssd1 vccd1 vccd1 _602_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[53\] _524_/Y la_buf\[53\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[53]
+ sky130_fd_sc_hd__einvp_8
X_464_ mprj_dat_o_core[25] vssd1 vssd1 vccd1 vccd1 _464_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_533_ la_data_out_mprj[62] vssd1 vssd1 vccd1 vccd1 _533_/Y sky130_fd_sc_hd__inv_2
X_395_ la_oen_mprj[127] vssd1 vssd1 vccd1 vccd1 _395_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[17\] _424_/Y mprj_adr_buf\[17\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[97] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] mprj_logic_high\[372\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[42\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] mprj_logic_high\[334\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[4\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_13_2136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[329\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[329\]/HI mprj_logic_high\[329\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[93\] _361_/Y mprj_logic_high\[295\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[231\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[231\]/HI mprj_logic_high\[231\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_378_ la_oen_mprj[110] vssd1 vssd1 vccd1 vccd1 _378_/Y sky130_fd_sc_hd__inv_2
X_447_ mprj_dat_o_core[8] vssd1 vssd1 vccd1 vccd1 _447_/Y sky130_fd_sc_hd__inv_2
X_516_ la_data_out_mprj[45] vssd1 vssd1 vccd1 vccd1 _516_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[12] sky130_fd_sc_hd__inv_8
XFILLER_7_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[279\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[279\]/HI mprj_logic_high\[279\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[181\] vssd1 vssd1 vccd1 vccd1 la_buf\[107\]/TE mprj_logic_high\[181\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[92\] vssd1 vssd1 vccd1 vccd1 la_buf\[18\]/TE mprj_logic_high\[92\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[4] sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[446\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[446\]/HI mprj_logic_high\[446\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xla_buf\[16\] _487_/Y la_buf\[16\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[16]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[9\] _416_/Y mprj_adr_buf\[9\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] mprj_logic_high\[446\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[116\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[126\] _394_/Y mprj_logic_high\[328\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[126] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[56\] _655_/Y mprj_logic_high\[258\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[56] sky130_fd_sc_hd__einvp_8
XFILLER_10_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[396\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[396\]/HI mprj_logic_high\[396\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[113] sky130_fd_sc_hd__inv_8
XFILLER_4_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[55\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[13\]/TE mprj_logic_high\[55\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[144\] vssd1 vssd1 vccd1 vccd1 la_buf\[70\]/TE mprj_logic_high\[144\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[311\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[311\]/HI mprj_logic_high\[311\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[409\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[409\]/HI mprj_logic_high\[409\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[83\] _554_/Y la_buf\[83\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[83]
+ sky130_fd_sc_hd__einvp_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] mprj_logic_high\[402\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[72\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[19\] _618_/Y mprj_logic_high\[221\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[19] sky130_fd_sc_hd__einvp_8
X_480_ la_data_out_mprj[9] vssd1 vssd1 vccd1 vccd1 _480_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[261\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[261\]/HI mprj_logic_high\[261\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[359\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[359\]/HI mprj_logic_high\[359\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[42] sky130_fd_sc_hd__inv_8
XFILLER_1_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[18\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[8\]/TE mprj_logic_high\[18\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[107\] vssd1 vssd1 vccd1 vccd1 la_buf\[33\]/TE mprj_logic_high\[107\]/LO
+ sky130_fd_sc_hd__conb_1
X_601_ la_oen_mprj[2] vssd1 vssd1 vccd1 vccd1 _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xla_buf\[46\] _517_/Y la_buf\[46\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[46]
+ sky130_fd_sc_hd__einvp_8
X_463_ mprj_dat_o_core[24] vssd1 vssd1 vccd1 vccd1 _463_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_394_ la_oen_mprj[126] vssd1 vssd1 vccd1 vccd1 _394_/Y sky130_fd_sc_hd__inv_2
X_532_ la_data_out_mprj[61] vssd1 vssd1 vccd1 vccd1 _532_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xla_buf\[102\] _573_/Y la_buf\[102\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[102]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] mprj_logic_high\[365\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[35\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[86\] _354_/Y mprj_logic_high\[288\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[224\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[224\]/HI mprj_logic_high\[224\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_2084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_515_ la_data_out_mprj[44] vssd1 vssd1 vccd1 vccd1 _515_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_446_ mprj_dat_o_core[7] vssd1 vssd1 vccd1 vccd1 _446_/Y sky130_fd_sc_hd__inv_2
X_377_ la_oen_mprj[109] vssd1 vssd1 vccd1 vccd1 _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[174\] vssd1 vssd1 vccd1 vccd1 la_buf\[100\]/TE mprj_logic_high\[174\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[85\] vssd1 vssd1 vccd1 vccd1 la_buf\[11\]/TE mprj_logic_high\[85\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[341\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[341\]/HI mprj_logic_high\[341\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[439\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[439\]/HI mprj_logic_high\[439\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_429_ mprj_adr_o_core[22] vssd1 vssd1 vccd1 vccd1 _429_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[2\] vssd1 vssd1 vccd1 vccd1 mprj_clk2_buf/TE mprj_logic_high\[2\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] mprj_logic_high\[439\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[109\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[119\] _387_/Y mprj_logic_high\[321\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_15_2007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[291\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[291\]/HI mprj_logic_high\[291\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[389\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[389\]/HI mprj_logic_high\[389\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[49\] _648_/Y mprj_logic_high\[251\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[72] sky130_fd_sc_hd__inv_8
XFILLER_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[106] sky130_fd_sc_hd__inv_8
XFILLER_0_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[5\] _444_/Y mprj_dat_buf\[5\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[137\] vssd1 vssd1 vccd1 vccd1 la_buf\[63\]/TE mprj_logic_high\[137\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[48\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[6\]/TE mprj_logic_high\[48\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[304\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[304\]/HI mprj_logic_high\[304\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[76\] _547_/Y la_buf\[76\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[76]
+ sky130_fd_sc_hd__einvp_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] mprj_logic_high\[395\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[65\]/Y sky130_fd_sc_hd__nand2_4
Xmprj_logic_high\[254\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[254\]/HI mprj_logic_high\[254\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[421\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[421\]/HI mprj_logic_high\[421\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[35] sky130_fd_sc_hd__inv_8
XFILLER_1_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[101\] _369_/Y mprj_logic_high\[303\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_2_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[31\] _630_/Y mprj_logic_high\[233\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[31] sky130_fd_sc_hd__einvp_8
X_531_ la_data_out_mprj[60] vssd1 vssd1 vccd1 vccd1 _531_/Y sky130_fd_sc_hd__inv_2
X_600_ la_oen_mprj[1] vssd1 vssd1 vccd1 vccd1 _600_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[371\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[371\]/HI mprj_logic_high\[371\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_462_ mprj_dat_o_core[23] vssd1 vssd1 vccd1 vccd1 _462_/Y sky130_fd_sc_hd__inv_2
X_393_ la_oen_mprj[125] vssd1 vssd1 vccd1 vccd1 _393_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[39\] _510_/Y la_buf\[39\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[39]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] mprj_logic_high\[358\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[28\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[30\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[20\]/TE mprj_logic_high\[30\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[27\] _466_/Y mprj_dat_buf\[27\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[27]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[79\] _347_/Y mprj_logic_high\[281\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[217\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[217\]/HI mprj_logic_high\[217\]/LO
+ sky130_fd_sc_hd__conb_1
X_514_ la_data_out_mprj[43] vssd1 vssd1 vccd1 vccd1 _514_/Y sky130_fd_sc_hd__inv_2
X_445_ mprj_dat_o_core[6] vssd1 vssd1 vccd1 vccd1 _445_/Y sky130_fd_sc_hd__inv_2
X_376_ la_oen_mprj[108] vssd1 vssd1 vccd1 vccd1 _376_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[22\] _429_/Y mprj_adr_buf\[22\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[167\] vssd1 vssd1 vccd1 vccd1 la_buf\[93\]/TE mprj_logic_high\[167\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[78\] vssd1 vssd1 vccd1 vccd1 la_buf\[4\]/TE mprj_logic_high\[78\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[334\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[334\]/HI mprj_logic_high\[334\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_428_ mprj_adr_o_core[21] vssd1 vssd1 vccd1 vccd1 _428_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_359_ la_oen_mprj[91] vssd1 vssd1 vccd1 vccd1 _359_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] mprj_logic_high\[425\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[95\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[284\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[284\]/HI mprj_logic_high\[284\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xla_buf\[21\] _492_/Y la_buf\[21\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[21]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[451\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[451\]/HI mprj_logic_high\[451\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[65] sky130_fd_sc_hd__inv_8
XFILLER_4_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] mprj_logic_high\[340\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[10\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] mprj_logic_high\[451\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[121\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_13_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[61\] _660_/Y mprj_logic_high\[263\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[61] sky130_fd_sc_hd__einvp_8
XFILLER_5_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xla_buf\[69\] _540_/Y la_buf\[69\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[69]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[125\] _596_/Y la_buf\[125\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[125]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] mprj_logic_high\[388\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[58\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[60\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[18\]/TE mprj_logic_high\[60\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[247\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[247\]/HI mprj_logic_high\[247\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[414\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[414\]/HI mprj_logic_high\[414\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[28] sky130_fd_sc_hd__inv_8
XFILLER_12_1888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[24\] _623_/Y mprj_logic_high\[226\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[24] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[6\] _605_/Y mprj_logic_high\[208\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[6] sky130_fd_sc_hd__einvp_8
X_461_ mprj_dat_o_core[22] vssd1 vssd1 vccd1 vccd1 _461_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_530_ la_data_out_mprj[59] vssd1 vssd1 vccd1 vccd1 _530_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[197\] vssd1 vssd1 vccd1 vccd1 la_buf\[123\]/TE mprj_logic_high\[197\]/LO
+ sky130_fd_sc_hd__conb_1
X_392_ la_oen_mprj[124] vssd1 vssd1 vccd1 vccd1 _392_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[364\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[364\]/HI mprj_logic_high\[364\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_659_ la_oen_mprj[60] vssd1 vssd1 vccd1 vccd1 _659_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[23\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[13\]/TE mprj_logic_high\[23\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[112\] vssd1 vssd1 vccd1 vccd1 la_buf\[38\]/TE mprj_logic_high\[112\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[51\] _522_/Y la_buf\[51\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[51]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_444_ mprj_dat_o_core[5] vssd1 vssd1 vccd1 vccd1 _444_/Y sky130_fd_sc_hd__inv_2
X_513_ la_data_out_mprj[42] vssd1 vssd1 vccd1 vccd1 _513_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_375_ la_oen_mprj[107] vssd1 vssd1 vccd1 vccd1 _375_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[15\] _422_/Y mprj_adr_buf\[15\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[95] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] mprj_logic_high\[370\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[40\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] mprj_logic_high\[332\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[2\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_13_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[327\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[327\]/HI mprj_logic_high\[327\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[91\] _359_/Y mprj_logic_high\[293\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_13_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[99\] _570_/Y la_buf\[99\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[99]
+ sky130_fd_sc_hd__einvp_8
X_427_ mprj_adr_o_core[20] vssd1 vssd1 vccd1 vccd1 _427_/Y sky130_fd_sc_hd__inv_2
X_358_ la_oen_mprj[90] vssd1 vssd1 vccd1 vccd1 _358_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[10] sky130_fd_sc_hd__inv_8
XFILLER_6_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] mprj_logic_high\[418\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[88\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[277\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[277\]/HI mprj_logic_high\[277\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[90\] vssd1 vssd1 vccd1 vccd1 la_buf\[16\]/TE mprj_logic_high\[90\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[2] sky130_fd_sc_hd__inv_8
Xmprj_logic_high\[444\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[444\]/HI mprj_logic_high\[444\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[14\] _485_/Y la_buf\[14\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[14]
+ sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[7\] _414_/Y mprj_adr_buf\[7\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[58] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] mprj_logic_high\[444\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[114\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[124\] _392_/Y mprj_logic_high\[326\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[124] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[54\] _653_/Y mprj_logic_high\[256\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_1_2118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[394\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[394\]/HI mprj_logic_high\[394\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[118\] _589_/Y la_buf\[118\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[118]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[111] sky130_fd_sc_hd__inv_8
XFILLER_0_2140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[53\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[11\]/TE mprj_logic_high\[53\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[142\] vssd1 vssd1 vccd1 vccd1 la_buf\[68\]/TE mprj_logic_high\[142\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[407\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[407\]/HI mprj_logic_high\[407\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[81\] _552_/Y la_buf\[81\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[81]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] mprj_logic_high\[400\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[70\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_clk_buf _398_/Y mprj_clk_buf/TE vssd1 vssd1 vccd1 vccd1 user_clock sky130_fd_sc_hd__einvp_8
XFILLER_1_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[17\] _616_/Y mprj_logic_high\[219\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[17] sky130_fd_sc_hd__einvp_8
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_460_ mprj_dat_o_core[21] vssd1 vssd1 vccd1 vccd1 _460_/Y sky130_fd_sc_hd__inv_2
X_391_ la_oen_mprj[123] vssd1 vssd1 vccd1 vccd1 _391_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[357\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[357\]/HI mprj_logic_high\[357\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_658_ la_oen_mprj[59] vssd1 vssd1 vccd1 vccd1 _658_/Y sky130_fd_sc_hd__inv_2
X_589_ la_data_out_mprj[118] vssd1 vssd1 vccd1 vccd1 _589_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[40] sky130_fd_sc_hd__inv_8
XFILLER_1_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[16\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[6\]/TE mprj_logic_high\[16\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[105\] vssd1 vssd1 vccd1 vccd1 la_buf\[31\]/TE mprj_logic_high\[105\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[44\] _515_/Y la_buf\[44\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[44]
+ sky130_fd_sc_hd__einvp_8
X_443_ mprj_dat_o_core[4] vssd1 vssd1 vccd1 vccd1 _443_/Y sky130_fd_sc_hd__inv_2
X_374_ la_oen_mprj[106] vssd1 vssd1 vccd1 vccd1 _374_/Y sky130_fd_sc_hd__inv_2
X_512_ la_data_out_mprj[41] vssd1 vssd1 vccd1 vccd1 _512_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[100\] _571_/Y la_buf\[100\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[100]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] mprj_logic_high\[363\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[33\]/Y sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[88] sky130_fd_sc_hd__inv_8
XFILLER_3_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[84\] _352_/Y mprj_logic_high\[286\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[84] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[222\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[222\]/HI mprj_logic_high\[222\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_426_ mprj_adr_o_core[19] vssd1 vssd1 vccd1 vccd1 _426_/Y sky130_fd_sc_hd__inv_2
X_357_ la_oen_mprj[89] vssd1 vssd1 vccd1 vccd1 _357_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[83\] vssd1 vssd1 vccd1 vccd1 la_buf\[9\]/TE mprj_logic_high\[83\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[172\] vssd1 vssd1 vccd1 vccd1 la_buf\[98\]/TE mprj_logic_high\[172\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[437\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[437\]/HI mprj_logic_high\[437\]/LO
+ sky130_fd_sc_hd__conb_1
X_409_ mprj_adr_o_core[2] vssd1 vssd1 vccd1 vccd1 _409_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[0\] vssd1 vssd1 vccd1 vccd1 mprj_rstn_buf/TE mprj_logic_high\[0\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] mprj_logic_high\[437\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[107\]/Y sky130_fd_sc_hd__nand2_4
XPHY_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[117\] _385_/Y mprj_logic_high\[319\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[117] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[47\] _646_/Y mprj_logic_high\[249\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[47] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[387\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[387\]/HI mprj_logic_high\[387\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[70] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[104] sky130_fd_sc_hd__inv_8
XFILLER_15_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[3\] _442_/Y mprj_dat_buf\[3\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_14_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[46\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[4\]/TE mprj_logic_high\[46\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[135\] vssd1 vssd1 vccd1 vccd1 la_buf\[61\]/TE mprj_logic_high\[135\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[302\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[302\]/HI mprj_logic_high\[302\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[74\] _545_/Y la_buf\[74\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[74]
+ sky130_fd_sc_hd__einvp_8
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] mprj_logic_high\[393\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[63\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_390_ la_oen_mprj[122] vssd1 vssd1 vccd1 vccd1 _390_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[252\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[252\]/HI mprj_logic_high\[252\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_657_ la_oen_mprj[58] vssd1 vssd1 vccd1 vccd1 _657_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_588_ la_data_out_mprj[117] vssd1 vssd1 vccd1 vccd1 _588_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[33] sky130_fd_sc_hd__inv_8
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_511_ la_data_out_mprj[40] vssd1 vssd1 vccd1 vccd1 _511_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[37\] _508_/Y la_buf\[37\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[37]
+ sky130_fd_sc_hd__einvp_8
X_442_ mprj_dat_o_core[3] vssd1 vssd1 vccd1 vccd1 _442_/Y sky130_fd_sc_hd__inv_2
X_373_ la_oen_mprj[105] vssd1 vssd1 vccd1 vccd1 _373_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] mprj_logic_high\[356\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[26\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[25\] _464_/Y mprj_dat_buf\[25\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[25]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[77\] _345_/Y mprj_logic_high\[279\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[77] sky130_fd_sc_hd__einvp_8
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[215\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[215\]/HI mprj_logic_high\[215\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_425_ mprj_adr_o_core[18] vssd1 vssd1 vccd1 vccd1 _425_/Y sky130_fd_sc_hd__inv_2
X_356_ la_oen_mprj[88] vssd1 vssd1 vccd1 vccd1 _356_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[20\] _427_/Y mprj_adr_buf\[20\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[165\] vssd1 vssd1 vccd1 vccd1 la_buf\[91\]/TE mprj_logic_high\[165\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[76\] vssd1 vssd1 vccd1 vccd1 la_buf\[2\]/TE mprj_logic_high\[76\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[332\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[332\]/HI mprj_logic_high\[332\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_408_ mprj_adr_o_core[1] vssd1 vssd1 vccd1 vccd1 _408_/Y sky130_fd_sc_hd__inv_2
X_339_ la_oen_mprj[71] vssd1 vssd1 vccd1 vccd1 _339_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] mprj_logic_high\[423\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[93\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_2066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_10 la_oen_mprj[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[282\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[282\]/HI mprj_logic_high\[282\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[63] sky130_fd_sc_hd__inv_8
XFILLER_4_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[39\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[29\]/TE mprj_logic_high\[39\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[128\] vssd1 vssd1 vccd1 vccd1 la_buf\[54\]/TE mprj_logic_high\[128\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[67\] _538_/Y la_buf\[67\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[67]
+ sky130_fd_sc_hd__einvp_8
XFILLER_10_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[123\] _594_/Y la_buf\[123\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[123]
+ sky130_fd_sc_hd__einvp_8
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] mprj_logic_high\[386\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[56\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[245\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[245\]/HI mprj_logic_high\[245\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[412\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[412\]/HI mprj_logic_high\[412\]/LO
+ sky130_fd_sc_hd__conb_1
X_656_ la_oen_mprj[57] vssd1 vssd1 vccd1 vccd1 _656_/Y sky130_fd_sc_hd__inv_2
X_587_ la_data_out_mprj[116] vssd1 vssd1 vccd1 vccd1 _587_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[26] sky130_fd_sc_hd__inv_8
XFILLER_12_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[4\] _603_/Y mprj_logic_high\[206\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[4] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[195\] vssd1 vssd1 vccd1 vccd1 la_buf\[121\]/TE mprj_logic_high\[195\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_2056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_441_ mprj_dat_o_core[2] vssd1 vssd1 vccd1 vccd1 _441_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[22\] _621_/Y mprj_logic_high\[224\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[22] sky130_fd_sc_hd__einvp_8
X_510_ la_data_out_mprj[39] vssd1 vssd1 vccd1 vccd1 _510_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[362\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[362\]/HI mprj_logic_high\[362\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_372_ la_oen_mprj[104] vssd1 vssd1 vccd1 vccd1 _372_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_639_ la_oen_mprj[40] vssd1 vssd1 vccd1 vccd1 _639_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] mprj_logic_high\[349\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[19\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[21\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[11\]/TE mprj_logic_high\[21\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[18\] _457_/Y mprj_dat_buf\[18\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[18]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[110\] vssd1 vssd1 vccd1 vccd1 la_buf\[36\]/TE mprj_logic_high\[110\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[208\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[208\]/HI mprj_logic_high\[208\]/LO
+ sky130_fd_sc_hd__conb_1
X_424_ mprj_adr_o_core[17] vssd1 vssd1 vccd1 vccd1 _424_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_355_ la_oen_mprj[87] vssd1 vssd1 vccd1 vccd1 _355_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[13\] _420_/Y mprj_adr_buf\[13\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[93] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[127] sky130_fd_sc_hd__inv_8
XFILLER_14_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] mprj_logic_high\[330\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[0\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[69\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[27\]/TE mprj_logic_high\[69\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[158\] vssd1 vssd1 vccd1 vccd1 la_buf\[84\]/TE mprj_logic_high\[158\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[325\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[325\]/HI mprj_logic_high\[325\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[97\] _568_/Y la_buf\[97\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[97]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ mprj_adr_o_core[0] vssd1 vssd1 vccd1 vccd1 _407_/Y sky130_fd_sc_hd__inv_2
X_338_ la_oen_mprj[70] vssd1 vssd1 vccd1 vccd1 _338_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] mprj_logic_high\[416\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[86\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_11 la_oen_mprj[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[275\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[275\]/HI mprj_logic_high\[275\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[0] sky130_fd_sc_hd__inv_8
Xla_buf\[8\] _479_/Y la_buf\[8\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[8] sky130_fd_sc_hd__einvp_8
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[12\] _483_/Y la_buf\[12\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[12]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[442\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[442\]/HI mprj_logic_high\[442\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_adr_buf\[5\] _412_/Y mprj_adr_buf\[5\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[56] sky130_fd_sc_hd__inv_8
XFILLER_11_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] mprj_logic_high\[442\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[112\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_sel_buf\[3\] _406_/Y mprj_sel_buf\[3\]/TE vssd1 vssd1 vccd1 vccd1 mprj_sel_o_user[3]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[122\] _390_/Y mprj_logic_high\[324\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[122] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[52\] _651_/Y mprj_logic_high\[254\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[52] sky130_fd_sc_hd__einvp_8
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[392\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[392\]/HI mprj_logic_high\[392\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[116\] _587_/Y la_buf\[116\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[116]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] mprj_logic_high\[379\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[49\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_2140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[51\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[9\]/TE mprj_logic_high\[51\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[238\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[238\]/HI mprj_logic_high\[238\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[140\] vssd1 vssd1 vccd1 vccd1 la_buf\[66\]/TE mprj_logic_high\[140\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[405\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[405\]/HI mprj_logic_high\[405\]/LO
+ sky130_fd_sc_hd__conb_1
X_655_ la_oen_mprj[56] vssd1 vssd1 vccd1 vccd1 _655_/Y sky130_fd_sc_hd__inv_2
X_586_ la_data_out_mprj[115] vssd1 vssd1 vccd1 vccd1 _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[19] sky130_fd_sc_hd__inv_8
XPHY_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_2002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[188\] vssd1 vssd1 vccd1 vccd1 la_buf\[114\]/TE mprj_logic_high\[188\]/LO
+ sky130_fd_sc_hd__conb_1
X_440_ mprj_dat_o_core[1] vssd1 vssd1 vccd1 vccd1 _440_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_371_ la_oen_mprj[103] vssd1 vssd1 vccd1 vccd1 _371_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[99\] vssd1 vssd1 vccd1 vccd1 la_buf\[25\]/TE mprj_logic_high\[99\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[15\] _614_/Y mprj_logic_high\[217\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_0_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[355\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[355\]/HI mprj_logic_high\[355\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_638_ la_oen_mprj[39] vssd1 vssd1 vccd1 vccd1 _638_/Y sky130_fd_sc_hd__inv_2
X_569_ la_data_out_mprj[98] vssd1 vssd1 vccd1 vccd1 _569_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[14\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[4\]/TE mprj_logic_high\[14\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[103\] vssd1 vssd1 vccd1 vccd1 la_buf\[29\]/TE mprj_logic_high\[103\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[42\] _513_/Y la_buf\[42\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[42]
+ sky130_fd_sc_hd__einvp_8
X_423_ mprj_adr_o_core[16] vssd1 vssd1 vccd1 vccd1 _423_/Y sky130_fd_sc_hd__inv_2
X_354_ la_oen_mprj[86] vssd1 vssd1 vccd1 vccd1 _354_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[86] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] mprj_logic_high\[361\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[31\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[30\] _469_/Y mprj_dat_buf\[30\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[30]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[318\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[318\]/HI mprj_logic_high\[318\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[82\] _350_/Y mprj_logic_high\[284\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[82] sky130_fd_sc_hd__einvp_8
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[220\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[220\]/HI mprj_logic_high\[220\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_337_ la_oen_mprj[69] vssd1 vssd1 vccd1 vccd1 _337_/Y sky130_fd_sc_hd__inv_2
X_406_ mprj_sel_o_core[3] vssd1 vssd1 vccd1 vccd1 _406_/Y sky130_fd_sc_hd__inv_2
XPHY_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] mprj_logic_high\[409\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[79\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_12 la_oen_mprj[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[268\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[268\]/HI mprj_logic_high\[268\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[170\] vssd1 vssd1 vccd1 vccd1 la_buf\[96\]/TE mprj_logic_high\[170\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[81\] vssd1 vssd1 vccd1 vccd1 la_buf\[7\]/TE mprj_logic_high\[81\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[435\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[435\]/HI mprj_logic_high\[435\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[49] sky130_fd_sc_hd__inv_8
XFILLER_4_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] mprj_logic_high\[435\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[105\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[115\] _383_/Y mprj_logic_high\[317\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[115] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[45\] _644_/Y mprj_logic_high\[247\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[45] sky130_fd_sc_hd__einvp_8
XFILLER_5_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[385\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[385\]/HI mprj_logic_high\[385\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[109\] _580_/Y la_buf\[109\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[109]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[102] sky130_fd_sc_hd__inv_8
XFILLER_15_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[1\] _440_/Y mprj_dat_buf\[1\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[44\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[2\]/TE mprj_logic_high\[44\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[133\] vssd1 vssd1 vccd1 vccd1 la_buf\[59\]/TE mprj_logic_high\[133\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[300\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[300\]/HI mprj_logic_high\[300\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_654_ la_oen_mprj[55] vssd1 vssd1 vccd1 vccd1 _654_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[72\] _543_/Y la_buf\[72\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[72]
+ sky130_fd_sc_hd__einvp_8
XPHY_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_585_ la_data_out_mprj[114] vssd1 vssd1 vccd1 vccd1 _585_/Y sky130_fd_sc_hd__inv_2
XPHY_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] mprj_logic_high\[391\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[61\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_370_ la_oen_mprj[102] vssd1 vssd1 vccd1 vccd1 _370_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[250\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[250\]/HI mprj_logic_high\[250\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[348\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[348\]/HI mprj_logic_high\[348\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_637_ la_oen_mprj[38] vssd1 vssd1 vccd1 vccd1 _637_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_499_ la_data_out_mprj[28] vssd1 vssd1 vccd1 vccd1 _499_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[31] sky130_fd_sc_hd__inv_8
X_568_ la_data_out_mprj[97] vssd1 vssd1 vccd1 vccd1 _568_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[9\] vssd1 vssd1 vccd1 vccd1 mprj_sel_buf\[3\]/TE mprj_logic_high\[9\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[298\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[298\]/HI mprj_logic_high\[298\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[35\] _506_/Y la_buf\[35\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[35]
+ sky130_fd_sc_hd__einvp_8
X_422_ mprj_adr_o_core[15] vssd1 vssd1 vccd1 vccd1 _422_/Y sky130_fd_sc_hd__inv_2
X_353_ la_oen_mprj[85] vssd1 vssd1 vccd1 vccd1 _353_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[79] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] mprj_logic_high\[354\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[24\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[23\] _462_/Y mprj_dat_buf\[23\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[23]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[75\] _343_/Y mprj_logic_high\[277\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[75] sky130_fd_sc_hd__einvp_8
XFILLER_8_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[213\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[213\]/HI mprj_logic_high\[213\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ mprj_sel_o_core[2] vssd1 vssd1 vccd1 vccd1 _405_/Y sky130_fd_sc_hd__inv_2
XPHY_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ la_oen_mprj[68] vssd1 vssd1 vccd1 vccd1 _336_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_13 la_oen_mprj[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[163\] vssd1 vssd1 vccd1 vccd1 la_buf\[89\]/TE mprj_logic_high\[163\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[74\] vssd1 vssd1 vccd1 vccd1 la_buf\[0\]/TE mprj_logic_high\[74\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[330\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[330\]/HI mprj_logic_high\[330\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[428\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[428\]/HI mprj_logic_high\[428\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xpowergood_check mprj2_pwrgood/A mprj_vdd_pwrgood/A vccd vssd vdda1 vssa1 vdda2 vssa2
+ mgmt_protect_hv
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] mprj_logic_high\[421\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[91\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[108\] _376_/Y mprj_logic_high\[310\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[108] sky130_fd_sc_hd__einvp_8
XFILLER_5_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[280\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[280\]/HI mprj_logic_high\[280\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[378\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[378\]/HI mprj_logic_high\[378\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[38\] _637_/Y mprj_logic_high\[240\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_1_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[61] sky130_fd_sc_hd__inv_8
XFILLER_15_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[37\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[27\]/TE mprj_logic_high\[37\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[126\] vssd1 vssd1 vccd1 vccd1 la_buf\[52\]/TE mprj_logic_high\[126\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_653_ la_oen_mprj[54] vssd1 vssd1 vccd1 vccd1 _653_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[65\] _536_/Y la_buf\[65\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[65]
+ sky130_fd_sc_hd__einvp_8
XPHY_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_584_ la_data_out_mprj[113] vssd1 vssd1 vccd1 vccd1 _584_/Y sky130_fd_sc_hd__inv_2
XPHY_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_adr_buf\[29\] _436_/Y mprj_adr_buf\[29\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[121\] _592_/Y la_buf\[121\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[121]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] mprj_logic_high\[384\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[54\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[243\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[243\]/HI mprj_logic_high\[243\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[410\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[410\]/HI mprj_logic_high\[410\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_636_ la_oen_mprj[37] vssd1 vssd1 vccd1 vccd1 _636_/Y sky130_fd_sc_hd__inv_2
X_567_ la_data_out_mprj[96] vssd1 vssd1 vccd1 vccd1 _567_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_498_ la_data_out_mprj[27] vssd1 vssd1 vccd1 vccd1 _498_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[24] sky130_fd_sc_hd__inv_8
XFILLER_5_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[20\] _619_/Y mprj_logic_high\[222\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[20] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[2\] _601_/Y mprj_logic_high\[204\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[2] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[193\] vssd1 vssd1 vccd1 vccd1 la_buf\[119\]/TE mprj_logic_high\[193\]/LO
+ sky130_fd_sc_hd__conb_1
X_421_ mprj_adr_o_core[14] vssd1 vssd1 vccd1 vccd1 _421_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[360\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[360\]/HI mprj_logic_high\[360\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[458\] vssd1 vssd1 vccd1 vccd1 mprj_pwrgood/A mprj_logic_high\[458\]/LO
+ sky130_fd_sc_hd__conb_1
X_352_ la_oen_mprj[84] vssd1 vssd1 vccd1 vccd1 _352_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[28\] _499_/Y la_buf\[28\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[28]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_619_ la_oen_mprj[20] vssd1 vssd1 vccd1 vccd1 _619_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] mprj_logic_high\[347\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[17\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[16\] _455_/Y mprj_dat_buf\[16\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[16]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[206\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[206\]/HI mprj_logic_high\[206\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[68\] _336_/Y mprj_logic_high\[270\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[68] sky130_fd_sc_hd__einvp_8
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_404_ mprj_sel_o_core[1] vssd1 vssd1 vccd1 vccd1 _404_/Y sky130_fd_sc_hd__inv_2
XPHY_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ la_oen_mprj[67] vssd1 vssd1 vccd1 vccd1 _335_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[11\] _418_/Y mprj_adr_buf\[11\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[11]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[125] sky130_fd_sc_hd__inv_8
XFILLER_1_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[91] sky130_fd_sc_hd__inv_8
XFILLER_14_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_14 la_oen_mprj[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[156\] vssd1 vssd1 vccd1 vccd1 la_buf\[82\]/TE mprj_logic_high\[156\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[67\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[25\]/TE mprj_logic_high\[67\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[323\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[323\]/HI mprj_logic_high\[323\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xla_buf\[95\] _566_/Y la_buf\[95\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[95]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] mprj_logic_high\[414\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[84\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[273\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[273\]/HI mprj_logic_high\[273\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[6\] _477_/Y la_buf\[6\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[6] sky130_fd_sc_hd__einvp_8
Xla_buf\[10\] _481_/Y la_buf\[10\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[440\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[440\]/HI mprj_logic_high\[440\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_adr_buf\[3\] _410_/Y mprj_adr_buf\[3\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[54] sky130_fd_sc_hd__inv_8
XFILLER_15_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] mprj_logic_high\[440\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[110\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[120\] _388_/Y mprj_logic_high\[322\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[120] sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[1\] _404_/Y mprj_sel_buf\[1\]/TE vssd1 vssd1 vccd1 vccd1 mprj_sel_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[119\] vssd1 vssd1 vccd1 vccd1 la_buf\[45\]/TE mprj_logic_high\[119\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[390\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[390\]/HI mprj_logic_high\[390\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[50\] _649_/Y mprj_logic_high\[252\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[50] sky130_fd_sc_hd__einvp_8
X_652_ la_oen_mprj[53] vssd1 vssd1 vccd1 vccd1 _652_/Y sky130_fd_sc_hd__inv_2
X_583_ la_data_out_mprj[112] vssd1 vssd1 vccd1 vccd1 _583_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[58\] _529_/Y la_buf\[58\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[58]
+ sky130_fd_sc_hd__einvp_8
XPHY_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[114\] _585_/Y la_buf\[114\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[114]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] mprj_logic_high\[377\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[47\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] mprj_logic_high\[339\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[9\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[98\] _366_/Y mprj_logic_high\[300\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_6_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[236\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[236\]/HI mprj_logic_high\[236\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[403\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[403\]/HI mprj_logic_high\[403\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_566_ la_data_out_mprj[95] vssd1 vssd1 vccd1 vccd1 _566_/Y sky130_fd_sc_hd__inv_2
X_635_ la_oen_mprj[36] vssd1 vssd1 vccd1 vccd1 _635_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_2124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_497_ la_data_out_mprj[26] vssd1 vssd1 vccd1 vccd1 _497_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[17] sky130_fd_sc_hd__inv_8
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[13\] _612_/Y mprj_logic_high\[215\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[13] sky130_fd_sc_hd__einvp_8
X_420_ mprj_adr_o_core[13] vssd1 vssd1 vccd1 vccd1 _420_/Y sky130_fd_sc_hd__inv_2
X_351_ la_oen_mprj[83] vssd1 vssd1 vccd1 vccd1 _351_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[97\] vssd1 vssd1 vccd1 vccd1 la_buf\[23\]/TE mprj_logic_high\[97\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[186\] vssd1 vssd1 vccd1 vccd1 la_buf\[112\]/TE mprj_logic_high\[186\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[353\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[353\]/HI mprj_logic_high\[353\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[9] sky130_fd_sc_hd__inv_8
XFILLER_13_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_549_ la_data_out_mprj[78] vssd1 vssd1 vccd1 vccd1 _549_/Y sky130_fd_sc_hd__inv_2
X_618_ la_oen_mprj[19] vssd1 vssd1 vccd1 vccd1 _618_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[12\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[2\]/TE mprj_logic_high\[12\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[101\] vssd1 vssd1 vccd1 vccd1 la_buf\[27\]/TE mprj_logic_high\[101\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ mprj_sel_o_core[0] vssd1 vssd1 vccd1 vccd1 _403_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[40\] _511_/Y la_buf\[40\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[40]
+ sky130_fd_sc_hd__einvp_8
XPHY_50 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ la_oen_mprj[66] vssd1 vssd1 vccd1 vccd1 _334_/Y sky130_fd_sc_hd__inv_2
XPHY_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[118] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[84] sky130_fd_sc_hd__inv_8
XFILLER_14_2027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_15 mprj_sel_o_core[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[149\] vssd1 vssd1 vccd1 vccd1 la_buf\[75\]/TE mprj_logic_high\[149\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[316\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[316\]/HI mprj_logic_high\[316\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[80\] _348_/Y mprj_logic_high\[282\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[80] sky130_fd_sc_hd__einvp_8
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[88\] _559_/Y la_buf\[88\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[88]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] mprj_logic_high\[407\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[77\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[266\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[266\]/HI mprj_logic_high\[266\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[433\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[433\]/HI mprj_logic_high\[433\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_2100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[47] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] mprj_logic_high\[433\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[103\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[113\] _381_/Y mprj_logic_high\[315\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[113] sky130_fd_sc_hd__einvp_8
Xmprj_clk2_buf _399_/Y mprj_clk2_buf/TE vssd1 vssd1 vccd1 vccd1 user_clock2 sky130_fd_sc_hd__einvp_8
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_651_ la_oen_mprj[52] vssd1 vssd1 vccd1 vccd1 _651_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[43\] _642_/Y mprj_logic_high\[245\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[43] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[383\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[383\]/HI mprj_logic_high\[383\]/LO
+ sky130_fd_sc_hd__conb_1
X_582_ la_data_out_mprj[111] vssd1 vssd1 vccd1 vccd1 _582_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xla_buf\[107\] _578_/Y la_buf\[107\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[107]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[100] sky130_fd_sc_hd__inv_8
XFILLER_15_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[42\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[0\]/TE mprj_logic_high\[42\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[131\] vssd1 vssd1 vccd1 vccd1 la_buf\[57\]/TE mprj_logic_high\[131\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[229\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[229\]/HI mprj_logic_high\[229\]/LO
+ sky130_fd_sc_hd__conb_1
X_634_ la_oen_mprj[35] vssd1 vssd1 vccd1 vccd1 _634_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_496_ la_data_out_mprj[25] vssd1 vssd1 vccd1 vccd1 _496_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[70\] _541_/Y la_buf\[70\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[70]
+ sky130_fd_sc_hd__einvp_8
X_565_ la_data_out_mprj[94] vssd1 vssd1 vccd1 vccd1 _565_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_350_ la_oen_mprj[82] vssd1 vssd1 vccd1 vccd1 _350_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[179\] vssd1 vssd1 vccd1 vccd1 la_buf\[105\]/TE mprj_logic_high\[179\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[346\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[346\]/HI mprj_logic_high\[346\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_617_ la_oen_mprj[18] vssd1 vssd1 vccd1 vccd1 _617_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_479_ la_data_out_mprj[8] vssd1 vssd1 vccd1 vccd1 _479_/Y sky130_fd_sc_hd__inv_2
X_548_ la_data_out_mprj[77] vssd1 vssd1 vccd1 vccd1 _548_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[7\] vssd1 vssd1 vccd1 vccd1 mprj_sel_buf\[1\]/TE mprj_logic_high\[7\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[296\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[296\]/HI mprj_logic_high\[296\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ mprj_we_o_core vssd1 vssd1 vccd1 vccd1 _402_/Y sky130_fd_sc_hd__inv_2
XPHY_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_333_ la_oen_mprj[65] vssd1 vssd1 vccd1 vccd1 _333_/Y sky130_fd_sc_hd__inv_2
XPHY_40 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[33\] _504_/Y la_buf\[33\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[33]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[77] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] mprj_logic_high\[352\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[22\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_16 mprj_we_o_core vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[21\] _460_/Y mprj_dat_buf\[21\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[21]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[309\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[309\]/HI mprj_logic_high\[309\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[73\] _341_/Y mprj_logic_high\[275\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[73] sky130_fd_sc_hd__einvp_8
XFILLER_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[211\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[211\]/HI mprj_logic_high\[211\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[72\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[30\]/TE mprj_logic_high\[72\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[161\] vssd1 vssd1 vccd1 vccd1 la_buf\[87\]/TE mprj_logic_high\[161\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[259\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[259\]/HI mprj_logic_high\[259\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[426\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[426\]/HI mprj_logic_high\[426\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[106\] _374_/Y mprj_logic_high\[308\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[106] sky130_fd_sc_hd__einvp_8
X_650_ la_oen_mprj[51] vssd1 vssd1 vccd1 vccd1 _650_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[36\] _635_/Y mprj_logic_high\[238\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[36] sky130_fd_sc_hd__einvp_8
XPHY_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_581_ la_data_out_mprj[110] vssd1 vssd1 vccd1 vccd1 _581_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[376\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[376\]/HI mprj_logic_high\[376\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[35\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[25\]/TE mprj_logic_high\[35\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[124\] vssd1 vssd1 vccd1 vccd1 la_buf\[50\]/TE mprj_logic_high\[124\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_633_ la_oen_mprj[34] vssd1 vssd1 vccd1 vccd1 _633_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[63\] _534_/Y la_buf\[63\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[63]
+ sky130_fd_sc_hd__einvp_8
X_495_ la_data_out_mprj[24] vssd1 vssd1 vccd1 vccd1 _495_/Y sky130_fd_sc_hd__inv_2
X_564_ la_data_out_mprj[93] vssd1 vssd1 vccd1 vccd1 _564_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[27\] _434_/Y mprj_adr_buf\[27\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] mprj_logic_high\[382\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[52\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_2062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_2051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[241\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[241\]/HI mprj_logic_high\[241\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[339\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[339\]/HI mprj_logic_high\[339\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_547_ la_data_out_mprj[76] vssd1 vssd1 vccd1 vccd1 _547_/Y sky130_fd_sc_hd__inv_2
X_616_ la_oen_mprj[17] vssd1 vssd1 vccd1 vccd1 _616_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_478_ la_data_out_mprj[7] vssd1 vssd1 vccd1 vccd1 _478_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[22] sky130_fd_sc_hd__inv_8
XFILLER_12_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[191\] vssd1 vssd1 vccd1 vccd1 la_buf\[117\]/TE mprj_logic_high\[191\]/LO
+ sky130_fd_sc_hd__conb_1
X_401_ mprj_stb_o_core vssd1 vssd1 vccd1 vccd1 _401_/Y sky130_fd_sc_hd__inv_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[0\] _599_/Y mprj_logic_high\[202\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[0] sky130_fd_sc_hd__einvp_8
XPHY_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[456\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[456\]/HI mprj_logic_high\[456\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[289\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[289\]/HI mprj_logic_high\[289\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_332_ la_oen_mprj[64] vssd1 vssd1 vccd1 vccd1 _332_/Y sky130_fd_sc_hd__inv_2
XPHY_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xla_buf\[26\] _497_/Y la_buf\[26\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_14_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] mprj_logic_high\[345\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[15\]/Y sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] mprj_logic_high\[456\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[126\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[14\] _453_/Y mprj_dat_buf\[14\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[14]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[66\] _334_/Y mprj_logic_high\[268\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[66] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[204\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[204\]/HI mprj_logic_high\[204\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[123] sky130_fd_sc_hd__inv_8
XFILLER_4_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[65\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[23\]/TE mprj_logic_high\[65\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[154\] vssd1 vssd1 vccd1 vccd1 la_buf\[80\]/TE mprj_logic_high\[154\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[419\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[419\]/HI mprj_logic_high\[419\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[321\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[321\]/HI mprj_logic_high\[321\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[93\] _564_/Y la_buf\[93\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[93]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] mprj_logic_high\[412\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[82\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_580_ la_data_out_mprj[109] vssd1 vssd1 vccd1 vccd1 _580_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[271\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[271\]/HI mprj_logic_high\[271\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[369\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[369\]/HI mprj_logic_high\[369\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[29\] _628_/Y mprj_logic_high\[231\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[29] sky130_fd_sc_hd__einvp_8
XPHY_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xla_buf\[4\] _475_/Y la_buf\[4\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[4] sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[1\] _408_/Y mprj_adr_buf\[1\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[52] sky130_fd_sc_hd__inv_8
XFILLER_6_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[28\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[18\]/TE mprj_logic_high\[28\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[117\] vssd1 vssd1 vccd1 vccd1 la_buf\[43\]/TE mprj_logic_high\[117\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_632_ la_oen_mprj[33] vssd1 vssd1 vccd1 vccd1 _632_/Y sky130_fd_sc_hd__inv_2
X_563_ la_data_out_mprj[92] vssd1 vssd1 vccd1 vccd1 _563_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xla_buf\[56\] _527_/Y la_buf\[56\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[56]
+ sky130_fd_sc_hd__einvp_8
X_494_ la_data_out_mprj[23] vssd1 vssd1 vccd1 vccd1 _494_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[112\] _583_/Y la_buf\[112\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[112]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] mprj_logic_high\[375\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[45\]/Y sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] mprj_logic_high\[337\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[7\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[96\] _364_/Y mprj_logic_high\[298\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[96] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[234\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[234\]/HI mprj_logic_high\[234\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[401\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[401\]/HI mprj_logic_high\[401\]/LO
+ sky130_fd_sc_hd__conb_1
X_546_ la_data_out_mprj[75] vssd1 vssd1 vccd1 vccd1 _546_/Y sky130_fd_sc_hd__inv_2
X_615_ la_oen_mprj[16] vssd1 vssd1 vccd1 vccd1 _615_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_477_ la_data_out_mprj[6] vssd1 vssd1 vccd1 vccd1 _477_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[15] sky130_fd_sc_hd__inv_8
XFILLER_3_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj2_pwrgood mprj2_pwrgood/A vssd1 vssd1 vccd1 vccd1 user2_vcc_powergood sky130_fd_sc_hd__buf_8
Xuser_to_mprj_oen_buffers\[11\] _610_/Y mprj_logic_high\[213\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[11] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[95\] vssd1 vssd1 vccd1 vccd1 la_buf\[21\]/TE mprj_logic_high\[95\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_400_ mprj_cyc_o_core vssd1 vssd1 vccd1 vccd1 _400_/Y sky130_fd_sc_hd__inv_2
X_331_ la_oen_mprj[63] vssd1 vssd1 vccd1 vccd1 _331_/Y sky130_fd_sc_hd__inv_2
XPHY_42 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[351\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[351\]/HI mprj_logic_high\[351\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[449\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[449\]/HI mprj_logic_high\[449\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[184\] vssd1 vssd1 vccd1 vccd1 la_buf\[110\]/TE mprj_logic_high\[184\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[7] sky130_fd_sc_hd__inv_8
XFILLER_13_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[19\] _490_/Y la_buf\[19\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[19]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_529_ la_data_out_mprj[58] vssd1 vssd1 vccd1 vccd1 _529_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] mprj_logic_high\[449\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[119\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[10\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[0\]/TE mprj_logic_high\[10\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[59\] _658_/Y mprj_logic_high\[261\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[59] sky130_fd_sc_hd__einvp_8
XFILLER_8_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[399\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[399\]/HI mprj_logic_high\[399\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[116] sky130_fd_sc_hd__inv_8
XFILLER_4_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[82] sky130_fd_sc_hd__inv_8
XFILLER_9_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[58\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[16\]/TE mprj_logic_high\[58\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[147\] vssd1 vssd1 vccd1 vccd1 la_buf\[73\]/TE mprj_logic_high\[147\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[314\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[314\]/HI mprj_logic_high\[314\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[86\] _557_/Y la_buf\[86\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[86]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] mprj_logic_high\[405\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[75\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[264\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[264\]/HI mprj_logic_high\[264\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[431\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[431\]/HI mprj_logic_high\[431\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[45] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] mprj_logic_high\[431\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[101\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[111\] _379_/Y mprj_logic_high\[313\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[111] sky130_fd_sc_hd__einvp_8
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[41\] _640_/Y mprj_logic_high\[243\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[41] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[381\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[381\]/HI mprj_logic_high\[381\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_631_ la_oen_mprj[32] vssd1 vssd1 vccd1 vccd1 _631_/Y sky130_fd_sc_hd__inv_2
X_493_ la_data_out_mprj[22] vssd1 vssd1 vccd1 vccd1 _493_/Y sky130_fd_sc_hd__inv_2
X_562_ la_data_out_mprj[91] vssd1 vssd1 vccd1 vccd1 _562_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[49\] _520_/Y la_buf\[49\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[49]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[105\] _576_/Y la_buf\[105\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[105]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] mprj_logic_high\[368\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[38\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_2075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[40\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[30\]/TE mprj_logic_high\[40\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[89\] _357_/Y mprj_logic_high\[291\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_2_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[227\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[227\]/HI mprj_logic_high\[227\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_476_ la_data_out_mprj[5] vssd1 vssd1 vccd1 vccd1 _476_/Y sky130_fd_sc_hd__inv_2
X_545_ la_data_out_mprj[74] vssd1 vssd1 vccd1 vccd1 _545_/Y sky130_fd_sc_hd__inv_2
X_614_ la_oen_mprj[15] vssd1 vssd1 vccd1 vccd1 _614_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_330_ la_oen_mprj[62] vssd1 vssd1 vccd1 vccd1 _330_/Y sky130_fd_sc_hd__inv_2
XPHY_43 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[88\] vssd1 vssd1 vccd1 vccd1 la_buf\[14\]/TE mprj_logic_high\[88\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_54 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[344\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[344\]/HI mprj_logic_high\[344\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[177\] vssd1 vssd1 vccd1 vccd1 la_buf\[103\]/TE mprj_logic_high\[177\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_459_ mprj_dat_o_core[20] vssd1 vssd1 vccd1 vccd1 _459_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_528_ la_data_out_mprj[57] vssd1 vssd1 vccd1 vccd1 _528_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[5\] vssd1 vssd1 vccd1 vccd1 mprj_we_buf/TE mprj_logic_high\[5\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[294\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[294\]/HI mprj_logic_high\[294\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xla_buf\[31\] _502_/Y la_buf\[31\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[109] sky130_fd_sc_hd__inv_8
XFILLER_4_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[75] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] mprj_logic_high\[350\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[20\]/Y sky130_fd_sc_hd__nand2_4
Xmprj_dat_buf\[8\] _447_/Y mprj_dat_buf\[8\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[307\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[307\]/HI mprj_logic_high\[307\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[71\] _339_/Y mprj_logic_high\[273\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[71] sky130_fd_sc_hd__einvp_8
Xla_buf\[79\] _550_/Y la_buf\[79\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[79]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] mprj_logic_high\[398\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[68\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[257\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[257\]/HI mprj_logic_high\[257\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[70\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[28\]/TE mprj_logic_high\[70\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[424\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[424\]/HI mprj_logic_high\[424\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[38] sky130_fd_sc_hd__inv_8
XFILLER_6_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[104\] _372_/Y mprj_logic_high\[306\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_630_ la_oen_mprj[31] vssd1 vssd1 vccd1 vccd1 _630_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[34\] _633_/Y mprj_logic_high\[236\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[34] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[374\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[374\]/HI mprj_logic_high\[374\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_492_ la_data_out_mprj[21] vssd1 vssd1 vccd1 vccd1 _492_/Y sky130_fd_sc_hd__inv_2
X_561_ la_data_out_mprj[90] vssd1 vssd1 vccd1 vccd1 _561_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[33\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[23\]/TE mprj_logic_high\[33\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[122\] vssd1 vssd1 vccd1 vccd1 la_buf\[48\]/TE mprj_logic_high\[122\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_613_ la_oen_mprj[14] vssd1 vssd1 vccd1 vccd1 _613_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[61\] _532_/Y la_buf\[61\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[61]
+ sky130_fd_sc_hd__einvp_8
X_475_ la_data_out_mprj[4] vssd1 vssd1 vccd1 vccd1 _475_/Y sky130_fd_sc_hd__inv_2
X_544_ la_data_out_mprj[73] vssd1 vssd1 vccd1 vccd1 _544_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[25\] _432_/Y mprj_adr_buf\[25\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] mprj_logic_high\[380\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[50\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[337\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[337\]/HI mprj_logic_high\[337\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_527_ la_data_out_mprj[56] vssd1 vssd1 vccd1 vccd1 _527_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_458_ mprj_dat_o_core[19] vssd1 vssd1 vccd1 vccd1 _458_/Y sky130_fd_sc_hd__inv_2
X_389_ la_oen_mprj[121] vssd1 vssd1 vccd1 vccd1 _389_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[20] sky130_fd_sc_hd__inv_8
XFILLER_9_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] mprj_logic_high\[428\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[98\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[454\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[454\]/HI mprj_logic_high\[454\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[287\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[287\]/HI mprj_logic_high\[287\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[24\] _495_/Y la_buf\[24\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[68] sky130_fd_sc_hd__inv_8
XFILLER_14_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] mprj_logic_high\[343\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[13\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] mprj_logic_high\[454\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[124\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[12\] _451_/Y mprj_dat_buf\[12\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[12]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[64\] _332_/Y mprj_logic_high\[266\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[64] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[202\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[202\]/HI mprj_logic_high\[202\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[121] sky130_fd_sc_hd__inv_8
XPHY_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[63\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[21\]/TE mprj_logic_high\[63\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[152\] vssd1 vssd1 vccd1 vccd1 la_buf\[78\]/TE mprj_logic_high\[152\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[417\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[417\]/HI mprj_logic_high\[417\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xla_buf\[91\] _562_/Y la_buf\[91\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[91]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] mprj_logic_high\[410\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[80\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_560_ la_data_out_mprj[89] vssd1 vssd1 vccd1 vccd1 _560_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[27\] _626_/Y mprj_logic_high\[229\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[27] sky130_fd_sc_hd__einvp_8
X_491_ la_data_out_mprj[20] vssd1 vssd1 vccd1 vccd1 _491_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[367\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[367\]/HI mprj_logic_high\[367\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[9\] _608_/Y mprj_logic_high\[211\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[9] sky130_fd_sc_hd__einvp_8
Xla_buf\[2\] _473_/Y la_buf\[2\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[2] sky130_fd_sc_hd__einvp_8
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_2033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[50] sky130_fd_sc_hd__inv_8
XFILLER_12_1941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[26\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[16\]/TE mprj_logic_high\[26\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[115\] vssd1 vssd1 vccd1 vccd1 la_buf\[41\]/TE mprj_logic_high\[115\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_543_ la_data_out_mprj[72] vssd1 vssd1 vccd1 vccd1 _543_/Y sky130_fd_sc_hd__inv_2
X_612_ la_oen_mprj[13] vssd1 vssd1 vccd1 vccd1 _612_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[54\] _525_/Y la_buf\[54\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[54]
+ sky130_fd_sc_hd__einvp_8
X_474_ la_data_out_mprj[3] vssd1 vssd1 vccd1 vccd1 _474_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[18\] _425_/Y mprj_adr_buf\[18\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xla_buf\[110\] _581_/Y la_buf\[110\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[110]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[98] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] mprj_logic_high\[373\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[43\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] mprj_logic_high\[335\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[5\]/Y sky130_fd_sc_hd__nand2_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[94\] _362_/Y mprj_logic_high\[296\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_13_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[232\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[232\]/HI mprj_logic_high\[232\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_526_ la_data_out_mprj[55] vssd1 vssd1 vccd1 vccd1 _526_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_457_ mprj_dat_o_core[18] vssd1 vssd1 vccd1 vccd1 _457_/Y sky130_fd_sc_hd__inv_2
X_388_ la_oen_mprj[120] vssd1 vssd1 vccd1 vccd1 _388_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[13] sky130_fd_sc_hd__inv_8
XFILLER_9_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[93\] vssd1 vssd1 vccd1 vccd1 la_buf\[19\]/TE mprj_logic_high\[93\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[447\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[447\]/HI mprj_logic_high\[447\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[182\] vssd1 vssd1 vccd1 vccd1 la_buf\[108\]/TE mprj_logic_high\[182\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[5] sky130_fd_sc_hd__inv_8
XFILLER_7_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[17\] _488_/Y la_buf\[17\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_509_ la_data_out_mprj[38] vssd1 vssd1 vccd1 vccd1 _509_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] mprj_logic_high\[447\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[117\]/Y sky130_fd_sc_hd__nand2_4
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[127\] _395_/Y mprj_logic_high\[329\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[127] sky130_fd_sc_hd__einvp_8
XFILLER_4_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[57\] _656_/Y mprj_logic_high\[259\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[57] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[397\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[397\]/HI mprj_logic_high\[397\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[114] sky130_fd_sc_hd__inv_8
XFILLER_4_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[80] sky130_fd_sc_hd__inv_8
XFILLER_0_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[56\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[14\]/TE mprj_logic_high\[56\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[145\] vssd1 vssd1 vccd1 vccd1 la_buf\[71\]/TE mprj_logic_high\[145\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[312\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[312\]/HI mprj_logic_high\[312\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[84\] _555_/Y la_buf\[84\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[84]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] mprj_logic_high\[403\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[73\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[262\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[262\]/HI mprj_logic_high\[262\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_490_ la_data_out_mprj[19] vssd1 vssd1 vccd1 vccd1 _490_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[43] sky130_fd_sc_hd__inv_8
XFILLER_12_1975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[19\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[9\]/TE mprj_logic_high\[19\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[108\] vssd1 vssd1 vccd1 vccd1 la_buf\[34\]/TE mprj_logic_high\[108\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_542_ la_data_out_mprj[71] vssd1 vssd1 vccd1 vccd1 _542_/Y sky130_fd_sc_hd__inv_2
X_473_ la_data_out_mprj[2] vssd1 vssd1 vccd1 vccd1 _473_/Y sky130_fd_sc_hd__inv_2
X_611_ la_oen_mprj[12] vssd1 vssd1 vccd1 vccd1 _611_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[47\] _518_/Y la_buf\[47\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[47]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[103\] _574_/Y la_buf\[103\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[103]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] mprj_logic_high\[366\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[36\]/Y sky130_fd_sc_hd__nand2_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[87\] _355_/Y mprj_logic_high\[289\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_11_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[225\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[225\]/HI mprj_logic_high\[225\]/LO
+ sky130_fd_sc_hd__conb_1
X_456_ mprj_dat_o_core[17] vssd1 vssd1 vccd1 vccd1 _456_/Y sky130_fd_sc_hd__inv_2
X_525_ la_data_out_mprj[54] vssd1 vssd1 vccd1 vccd1 _525_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[30\] _437_/Y mprj_adr_buf\[30\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[30]
+ sky130_fd_sc_hd__einvp_8
X_387_ la_oen_mprj[119] vssd1 vssd1 vccd1 vccd1 _387_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[86\] vssd1 vssd1 vccd1 vccd1 la_buf\[12\]/TE mprj_logic_high\[86\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_2078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[342\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[342\]/HI mprj_logic_high\[342\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[175\] vssd1 vssd1 vccd1 vccd1 la_buf\[101\]/TE mprj_logic_high\[175\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_439_ mprj_dat_o_core[0] vssd1 vssd1 vccd1 vccd1 _439_/Y sky130_fd_sc_hd__inv_2
X_508_ la_data_out_mprj[37] vssd1 vssd1 vccd1 vccd1 _508_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[3\] vssd1 vssd1 vccd1 vccd1 mprj_cyc_buf/TE mprj_logic_high\[3\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[292\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[292\]/HI mprj_logic_high\[292\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[107] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[73] sky130_fd_sc_hd__inv_8
XFILLER_15_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[6\] _445_/Y mprj_dat_buf\[6\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[49\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[7\]/TE mprj_logic_high\[49\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[305\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[305\]/HI mprj_logic_high\[305\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[138\] vssd1 vssd1 vccd1 vccd1 la_buf\[64\]/TE mprj_logic_high\[138\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[77\] _548_/Y la_buf\[77\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[77]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] mprj_logic_high\[396\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[66\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[255\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[255\]/HI mprj_logic_high\[255\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[422\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[422\]/HI mprj_logic_high\[422\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[36] sky130_fd_sc_hd__inv_8
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[102\] _370_/Y mprj_logic_high\[304\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_610_ la_oen_mprj[11] vssd1 vssd1 vccd1 vccd1 _610_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[372\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[372\]/HI mprj_logic_high\[372\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[32\] _631_/Y mprj_logic_high\[234\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[32] sky130_fd_sc_hd__einvp_8
X_472_ la_data_out_mprj[1] vssd1 vssd1 vccd1 vccd1 _472_/Y sky130_fd_sc_hd__inv_2
X_541_ la_data_out_mprj[70] vssd1 vssd1 vccd1 vccd1 _541_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] mprj_logic_high\[359\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[29\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[31\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[21\]/TE mprj_logic_high\[31\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[28\] _467_/Y mprj_dat_buf\[28\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[28]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[218\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[218\]/HI mprj_logic_high\[218\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[120\] vssd1 vssd1 vccd1 vccd1 la_buf\[46\]/TE mprj_logic_high\[120\]/LO
+ sky130_fd_sc_hd__conb_1
X_455_ mprj_dat_o_core[16] vssd1 vssd1 vccd1 vccd1 _455_/Y sky130_fd_sc_hd__inv_2
X_386_ la_oen_mprj[118] vssd1 vssd1 vccd1 vccd1 _386_/Y sky130_fd_sc_hd__inv_2
X_524_ la_data_out_mprj[53] vssd1 vssd1 vccd1 vccd1 _524_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[23\] _430_/Y mprj_adr_buf\[23\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[79\] vssd1 vssd1 vccd1 vccd1 la_buf\[5\]/TE mprj_logic_high\[79\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[168\] vssd1 vssd1 vccd1 vccd1 la_buf\[94\]/TE mprj_logic_high\[168\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[335\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[335\]/HI mprj_logic_high\[335\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_438_ mprj_adr_o_core[31] vssd1 vssd1 vccd1 vccd1 _438_/Y sky130_fd_sc_hd__inv_2
X_369_ la_oen_mprj[101] vssd1 vssd1 vccd1 vccd1 _369_/Y sky130_fd_sc_hd__inv_2
X_507_ la_data_out_mprj[36] vssd1 vssd1 vccd1 vccd1 _507_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] mprj_logic_high\[426\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[96\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[285\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[285\]/HI mprj_logic_high\[285\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[452\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[452\]/HI mprj_logic_high\[452\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[22\] _493_/Y la_buf\[22\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[66] sky130_fd_sc_hd__inv_8
XFILLER_15_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] mprj_logic_high\[341\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[11\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] mprj_logic_high\[452\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[122\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[10\] _449_/Y mprj_dat_buf\[10\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[10]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[62\] _330_/Y mprj_logic_high\[264\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[62] sky130_fd_sc_hd__einvp_8
XFILLER_0_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[200\] vssd1 vssd1 vccd1 vccd1 la_buf\[126\]/TE mprj_logic_high\[200\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[126\] _597_/Y la_buf\[126\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[126]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] mprj_logic_high\[389\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[59\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[150\] vssd1 vssd1 vccd1 vccd1 la_buf\[76\]/TE mprj_logic_high\[150\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[61\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[19\]/TE mprj_logic_high\[61\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[248\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[248\]/HI mprj_logic_high\[248\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[415\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[415\]/HI mprj_logic_high\[415\]/LO
+ sky130_fd_sc_hd__conb_1
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[29] sky130_fd_sc_hd__inv_8
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_540_ la_data_out_mprj[69] vssd1 vssd1 vccd1 vccd1 _540_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[365\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[365\]/HI mprj_logic_high\[365\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[7\] _606_/Y mprj_logic_high\[209\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[7] sky130_fd_sc_hd__einvp_8
XFILLER_2_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[25\] _624_/Y mprj_logic_high\[227\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[25] sky130_fd_sc_hd__einvp_8
X_471_ la_data_out_mprj[0] vssd1 vssd1 vccd1 vccd1 _471_/Y sky130_fd_sc_hd__inv_2
Xmprj_logic_high\[198\] vssd1 vssd1 vccd1 vccd1 la_buf\[124\]/TE mprj_logic_high\[198\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[0\] _471_/Y la_buf\[0\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[0] sky130_fd_sc_hd__einvp_8
XFILLER_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[24\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[14\]/TE mprj_logic_high\[24\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[113\] vssd1 vssd1 vccd1 vccd1 la_buf\[39\]/TE mprj_logic_high\[113\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_523_ la_data_out_mprj[52] vssd1 vssd1 vccd1 vccd1 _523_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[52\] _523_/Y la_buf\[52\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[52]
+ sky130_fd_sc_hd__einvp_8
X_454_ mprj_dat_o_core[15] vssd1 vssd1 vccd1 vccd1 _454_/Y sky130_fd_sc_hd__inv_2
X_385_ la_oen_mprj[117] vssd1 vssd1 vccd1 vccd1 _385_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[16\] _423_/Y mprj_adr_buf\[16\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_rstn_buf _396_/Y mprj_rstn_buf/TE vssd1 vssd1 vccd1 vccd1 user_resetn sky130_fd_sc_hd__einvp_8
XFILLER_1_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[96] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] mprj_logic_high\[371\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[41\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] mprj_logic_high\[333\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[3\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_2058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[328\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[328\]/HI mprj_logic_high\[328\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[92\] _360_/Y mprj_logic_high\[294\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[92] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[230\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[230\]/HI mprj_logic_high\[230\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_506_ la_data_out_mprj[35] vssd1 vssd1 vccd1 vccd1 _506_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_437_ mprj_adr_o_core[30] vssd1 vssd1 vccd1 vccd1 _437_/Y sky130_fd_sc_hd__inv_2
X_368_ la_oen_mprj[100] vssd1 vssd1 vccd1 vccd1 _368_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[11] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] mprj_logic_high\[419\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[89\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_cyc_buf _400_/Y mprj_cyc_buf/TE vssd1 vssd1 vccd1 vccd1 mprj_cyc_o_user sky130_fd_sc_hd__einvp_8
XFILLER_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[91\] vssd1 vssd1 vccd1 vccd1 la_buf\[17\]/TE mprj_logic_high\[91\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[445\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[445\]/HI mprj_logic_high\[445\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[278\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[278\]/HI mprj_logic_high\[278\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[180\] vssd1 vssd1 vccd1 vccd1 la_buf\[106\]/TE mprj_logic_high\[180\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[3] sky130_fd_sc_hd__inv_8
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[15\] _486_/Y la_buf\[15\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[8\] _415_/Y mprj_adr_buf\[8\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[59] sky130_fd_sc_hd__inv_8
XFILLER_9_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] mprj_logic_high\[445\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[115\]/Y sky130_fd_sc_hd__nand2_4
XPHY_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[125\] _393_/Y mprj_logic_high\[327\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_4_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[55\] _654_/Y mprj_logic_high\[257\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[55] sky130_fd_sc_hd__einvp_8
XFILLER_5_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[395\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[395\]/HI mprj_logic_high\[395\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[119\] _590_/Y la_buf\[119\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[119]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[112] sky130_fd_sc_hd__inv_8
XFILLER_4_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[54\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[12\]/TE mprj_logic_high\[54\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[310\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[310\]/HI mprj_logic_high\[310\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[143\] vssd1 vssd1 vccd1 vccd1 la_buf\[69\]/TE mprj_logic_high\[143\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[408\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[408\]/HI mprj_logic_high\[408\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[82\] _553_/Y la_buf\[82\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[82]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] mprj_logic_high\[401\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[71\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_470_ mprj_dat_o_core[31] vssd1 vssd1 vccd1 vccd1 _470_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[18\] _617_/Y mprj_logic_high\[220\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[260\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[260\]/HI mprj_logic_high\[260\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[358\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[358\]/HI mprj_logic_high\[358\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_599_ la_oen_mprj[0] vssd1 vssd1 vccd1 vccd1 _599_/Y sky130_fd_sc_hd__inv_2
XPHY_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[41] sky130_fd_sc_hd__inv_8
XANTENNA_0 la_oen_mprj[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_49 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[17\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[7\]/TE mprj_logic_high\[17\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[106\] vssd1 vssd1 vccd1 vccd1 la_buf\[32\]/TE mprj_logic_high\[106\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_453_ mprj_dat_o_core[14] vssd1 vssd1 vccd1 vccd1 _453_/Y sky130_fd_sc_hd__inv_2
X_522_ la_data_out_mprj[51] vssd1 vssd1 vccd1 vccd1 _522_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_384_ la_oen_mprj[116] vssd1 vssd1 vccd1 vccd1 _384_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[45\] _516_/Y la_buf\[45\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[45]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[101\] _572_/Y la_buf\[101\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[101]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[89] sky130_fd_sc_hd__inv_8
XFILLER_0_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] mprj_logic_high\[364\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[34\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[85\] _353_/Y mprj_logic_high\[287\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_11_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[223\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[223\]/HI mprj_logic_high\[223\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_436_ mprj_adr_o_core[29] vssd1 vssd1 vccd1 vccd1 _436_/Y sky130_fd_sc_hd__inv_2
X_505_ la_data_out_mprj[34] vssd1 vssd1 vccd1 vccd1 _505_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_367_ la_oen_mprj[99] vssd1 vssd1 vccd1 vccd1 _367_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[84\] vssd1 vssd1 vccd1 vccd1 la_buf\[10\]/TE mprj_logic_high\[84\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[340\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[340\]/HI mprj_logic_high\[340\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[173\] vssd1 vssd1 vccd1 vccd1 la_buf\[99\]/TE mprj_logic_high\[173\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[438\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[438\]/HI mprj_logic_high\[438\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_419_ mprj_adr_o_core[12] vssd1 vssd1 vccd1 vccd1 _419_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[1\] vssd1 vssd1 vccd1 vccd1 mprj_clk_buf/TE mprj_logic_high\[1\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] mprj_logic_high\[438\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[108\]/Y sky130_fd_sc_hd__nand2_4
XPHY_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_2143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[118\] _386_/Y mprj_logic_high\[320\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_0_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[48\] _647_/Y mprj_logic_high\[250\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[48] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[290\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[290\]/HI mprj_logic_high\[290\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[388\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[388\]/HI mprj_logic_high\[388\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[105] sky130_fd_sc_hd__inv_8
XFILLER_4_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[71] sky130_fd_sc_hd__inv_8
XFILLER_11_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[4\] _443_/Y mprj_dat_buf\[4\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[47\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[5\]/TE mprj_logic_high\[47\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[303\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[303\]/HI mprj_logic_high\[303\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[136\] vssd1 vssd1 vccd1 vccd1 la_buf\[62\]/TE mprj_logic_high\[136\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_2005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xla_buf\[75\] _546_/Y la_buf\[75\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[75]
+ sky130_fd_sc_hd__einvp_8
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] mprj_logic_high\[394\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[64\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[253\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[253\]/HI mprj_logic_high\[253\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[420\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[420\]/HI mprj_logic_high\[420\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_598_ la_data_out_mprj[127] vssd1 vssd1 vccd1 vccd1 _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1 la_oen_mprj[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[34] sky130_fd_sc_hd__inv_8
XFILLER_6_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[100\] _368_/Y mprj_logic_high\[302\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[370\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[370\]/HI mprj_logic_high\[370\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_452_ mprj_dat_o_core[13] vssd1 vssd1 vccd1 vccd1 _452_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_383_ la_oen_mprj[115] vssd1 vssd1 vccd1 vccd1 _383_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[30\] _629_/Y mprj_logic_high\[232\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[30] sky130_fd_sc_hd__einvp_8
X_521_ la_data_out_mprj[50] vssd1 vssd1 vccd1 vccd1 _521_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[38\] _509_/Y la_buf\[38\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[38]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] mprj_logic_high\[357\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[27\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_13_2005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[26\] _465_/Y mprj_dat_buf\[26\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[26]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[78\] _346_/Y mprj_logic_high\[280\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[78] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[216\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[216\]/HI mprj_logic_high\[216\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_435_ mprj_adr_o_core[28] vssd1 vssd1 vccd1 vccd1 _435_/Y sky130_fd_sc_hd__inv_2
X_366_ la_oen_mprj[98] vssd1 vssd1 vccd1 vccd1 _366_/Y sky130_fd_sc_hd__inv_2
X_504_ la_data_out_mprj[33] vssd1 vssd1 vccd1 vccd1 _504_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[21\] _428_/Y mprj_adr_buf\[21\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[77\] vssd1 vssd1 vccd1 vccd1 la_buf\[3\]/TE mprj_logic_high\[77\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[333\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[333\]/HI mprj_logic_high\[333\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[166\] vssd1 vssd1 vccd1 vccd1 la_buf\[92\]/TE mprj_logic_high\[166\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_418_ mprj_adr_o_core[11] vssd1 vssd1 vccd1 vccd1 _418_/Y sky130_fd_sc_hd__inv_2
X_349_ la_oen_mprj[81] vssd1 vssd1 vccd1 vccd1 _349_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] mprj_logic_high\[424\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[94\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[283\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[283\]/HI mprj_logic_high\[283\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[450\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[450\]/HI mprj_logic_high\[450\]/LO
+ sky130_fd_sc_hd__conb_1
Xla_buf\[20\] _491_/Y la_buf\[20\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[20]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[64] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] mprj_logic_high\[450\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[120\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[129\] vssd1 vssd1 vccd1 vccd1 la_buf\[55\]/TE mprj_logic_high\[129\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[60\] _659_/Y mprj_logic_high\[262\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[60] sky130_fd_sc_hd__einvp_8
Xla_buf\[68\] _539_/Y la_buf\[68\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[68]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xla_buf\[124\] _595_/Y la_buf\[124\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[124]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] mprj_logic_high\[387\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[57\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[246\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[246\]/HI mprj_logic_high\[246\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[413\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[413\]/HI mprj_logic_high\[413\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_597_ la_data_out_mprj[126] vssd1 vssd1 vccd1 vccd1 _597_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2 la_oen_mprj[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[27] sky130_fd_sc_hd__inv_8
XFILLER_4_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_520_ la_data_out_mprj[49] vssd1 vssd1 vccd1 vccd1 _520_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[196\] vssd1 vssd1 vccd1 vccd1 la_buf\[122\]/TE mprj_logic_high\[196\]/LO
+ sky130_fd_sc_hd__conb_1
Xuser_to_mprj_oen_buffers\[5\] _604_/Y mprj_logic_high\[207\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[5] sky130_fd_sc_hd__einvp_8
X_451_ mprj_dat_o_core[12] vssd1 vssd1 vccd1 vccd1 _451_/Y sky130_fd_sc_hd__inv_2
X_382_ la_oen_mprj[114] vssd1 vssd1 vccd1 vccd1 _382_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[23\] _622_/Y mprj_logic_high\[225\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[23] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[363\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[363\]/HI mprj_logic_high\[363\]/LO
+ sky130_fd_sc_hd__conb_1
X_649_ la_oen_mprj[50] vssd1 vssd1 vccd1 vccd1 _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[22\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[12\]/TE mprj_logic_high\[22\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[111\] vssd1 vssd1 vccd1 vccd1 la_buf\[37\]/TE mprj_logic_high\[111\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[209\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[209\]/HI mprj_logic_high\[209\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_dat_buf\[19\] _458_/Y mprj_dat_buf\[19\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[19]
+ sky130_fd_sc_hd__einvp_8
X_503_ la_data_out_mprj[32] vssd1 vssd1 vccd1 vccd1 _503_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[50\] _521_/Y la_buf\[50\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[50]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_434_ mprj_adr_o_core[27] vssd1 vssd1 vccd1 vccd1 _434_/Y sky130_fd_sc_hd__inv_2
X_365_ la_oen_mprj[97] vssd1 vssd1 vccd1 vccd1 _365_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[14\] _421_/Y mprj_adr_buf\[14\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[94] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] mprj_logic_high\[331\]/HI vssd1 vssd1
+ vccd1 vccd1 user_to_mprj_in_gates\[1\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[326\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[326\]/HI mprj_logic_high\[326\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[159\] vssd1 vssd1 vccd1 vccd1 la_buf\[85\]/TE mprj_logic_high\[159\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[90\] _358_/Y mprj_logic_high\[292\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[90] sky130_fd_sc_hd__einvp_8
Xla_buf\[98\] _569_/Y la_buf\[98\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[98]
+ sky130_fd_sc_hd__einvp_8
XFILLER_15_1945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_417_ mprj_adr_o_core[10] vssd1 vssd1 vccd1 vccd1 _417_/Y sky130_fd_sc_hd__inv_2
X_348_ la_oen_mprj[80] vssd1 vssd1 vccd1 vccd1 _348_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] mprj_logic_high\[417\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[87\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_logic_high\[443\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[443\]/HI mprj_logic_high\[443\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[276\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[276\]/HI mprj_logic_high\[276\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[1] sky130_fd_sc_hd__inv_8
XFILLER_7_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xla_buf\[9\] _480_/Y la_buf\[9\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[9] sky130_fd_sc_hd__einvp_8
Xla_buf\[13\] _484_/Y la_buf\[13\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[6\] _413_/Y mprj_adr_buf\[6\]/TE vssd1 vssd1 vccd1 vccd1 mprj_adr_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[57] sky130_fd_sc_hd__inv_8
XFILLER_15_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] mprj_logic_high\[443\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[113\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[123\] _391_/Y mprj_logic_high\[325\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[123] sky130_fd_sc_hd__einvp_8
XFILLER_14_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[53\] _652_/Y mprj_logic_high\[255\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_1_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[393\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[393\]/HI mprj_logic_high\[393\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[117\] _588_/Y la_buf\[117\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[117]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[110] sky130_fd_sc_hd__inv_8
XFILLER_6_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_2062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmprj_logic_high\[52\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[10\]/TE mprj_logic_high\[52\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[406\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[406\]/HI mprj_logic_high\[406\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[141\] vssd1 vssd1 vccd1 vccd1 la_buf\[67\]/TE mprj_logic_high\[141\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[239\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[239\]/HI mprj_logic_high\[239\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xla_buf\[80\] _551_/Y la_buf\[80\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[80]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_596_ la_data_out_mprj[125] vssd1 vssd1 vccd1 vccd1 _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_3 la_oen_mprj[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_450_ mprj_dat_o_core[11] vssd1 vssd1 vccd1 vccd1 _450_/Y sky130_fd_sc_hd__inv_2
X_381_ la_oen_mprj[113] vssd1 vssd1 vccd1 vccd1 _381_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[16\] _615_/Y mprj_logic_high\[218\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[16] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[189\] vssd1 vssd1 vccd1 vccd1 la_buf\[115\]/TE mprj_logic_high\[189\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[356\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[356\]/HI mprj_logic_high\[356\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_648_ la_oen_mprj[49] vssd1 vssd1 vccd1 vccd1 _648_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_579_ la_data_out_mprj[108] vssd1 vssd1 vccd1 vccd1 _579_/Y sky130_fd_sc_hd__inv_2
XPHY_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmprj_logic_high\[15\] vssd1 vssd1 vccd1 vccd1 mprj_adr_buf\[5\]/TE mprj_logic_high\[15\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmprj_logic_high\[104\] vssd1 vssd1 vccd1 vccd1 la_buf\[30\]/TE mprj_logic_high\[104\]/LO
+ sky130_fd_sc_hd__conb_1
X_433_ mprj_adr_o_core[26] vssd1 vssd1 vccd1 vccd1 _433_/Y sky130_fd_sc_hd__inv_2
X_502_ la_data_out_mprj[31] vssd1 vssd1 vccd1 vccd1 _502_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xla_buf\[43\] _514_/Y la_buf\[43\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[43]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_364_ la_oen_mprj[96] vssd1 vssd1 vccd1 vccd1 _364_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[87] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] mprj_logic_high\[362\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[32\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[31\] _470_/Y mprj_dat_buf\[31\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[31]
+ sky130_fd_sc_hd__einvp_8
Xmprj_logic_high\[319\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[319\]/HI mprj_logic_high\[319\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[83\] _351_/Y mprj_logic_high\[285\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[83] sky130_fd_sc_hd__einvp_8
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[221\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[221\]/HI mprj_logic_high\[221\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_416_ mprj_adr_o_core[9] vssd1 vssd1 vccd1 vccd1 _416_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_347_ la_oen_mprj[79] vssd1 vssd1 vccd1 vccd1 _347_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_2135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[82\] vssd1 vssd1 vccd1 vccd1 la_buf\[8\]/TE mprj_logic_high\[82\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[269\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[269\]/HI mprj_logic_high\[269\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[171\] vssd1 vssd1 vccd1 vccd1 la_buf\[97\]/TE mprj_logic_high\[171\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[436\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[436\]/HI mprj_logic_high\[436\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] mprj_logic_high\[436\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[106\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[116\] _384_/Y mprj_logic_high\[318\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_9_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[46\] _645_/Y mprj_logic_high\[248\]/HI vssd1 vssd1 vccd1
+ vccd1 la_oen_core[46] sky130_fd_sc_hd__einvp_8
XFILLER_5_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high\[386\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[386\]/HI mprj_logic_high\[386\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[103] sky130_fd_sc_hd__inv_8
Xmprj_dat_buf\[2\] _441_/Y mprj_dat_buf\[2\]/TE vssd1 vssd1 vccd1 vccd1 mprj_dat_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmprj_logic_high\[45\] vssd1 vssd1 vccd1 vccd1 mprj_dat_buf\[3\]/TE mprj_logic_high\[45\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xmprj_logic_high\[301\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[301\]/HI mprj_logic_high\[301\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[134\] vssd1 vssd1 vccd1 vccd1 la_buf\[60\]/TE mprj_logic_high\[134\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xla_buf\[73\] _544_/Y la_buf\[73\]/TE vssd1 vssd1 vccd1 vccd1 la_data_in_core[73]
+ sky130_fd_sc_hd__einvp_8
X_595_ la_data_out_mprj[124] vssd1 vssd1 vccd1 vccd1 _595_/Y sky130_fd_sc_hd__inv_2
XPHY_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 la_oen_mprj[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] mprj_logic_high\[392\]/HI vssd1
+ vssd1 vccd1 vccd1 user_to_mprj_in_gates\[62\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_380_ la_oen_mprj[112] vssd1 vssd1 vccd1 vccd1 _380_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmprj_logic_high\[251\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[251\]/HI mprj_logic_high\[251\]/LO
+ sky130_fd_sc_hd__conb_1
Xmprj_logic_high\[349\] vssd1 vssd1 vccd1 vccd1 mprj_logic_high\[349\]/HI mprj_logic_high\[349\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_647_ la_oen_mprj[48] vssd1 vssd1 vccd1 vccd1 _647_/Y sky130_fd_sc_hd__inv_2
X_578_ la_data_out_mprj[107] vssd1 vssd1 vccd1 vccd1 _578_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y vssd1 vssd1 vccd1 vccd1
+ la_data_in_mprj[32] sky130_fd_sc_hd__inv_8
XPHY_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

