magic
tech sky130A
magscale 1 2
timestamp 1606424343
<< metal3 >>
rect -5178 1572 -1806 1600
rect -5178 -1572 -1890 1572
rect -1826 -1572 -1806 1572
rect -5178 -1600 -1806 -1572
rect -1686 1572 1686 1600
rect -1686 -1572 1602 1572
rect 1666 -1572 1686 1572
rect -1686 -1600 1686 -1572
rect 1806 1572 5178 1600
rect 1806 -1572 5094 1572
rect 5158 -1572 5178 1572
rect 1806 -1600 5178 -1572
<< via3 >>
rect -1890 -1572 -1826 1572
rect 1602 -1572 1666 1572
rect 5094 -1572 5158 1572
<< mimcap >>
rect -5078 1460 -2078 1500
rect -5078 -1460 -5038 1460
rect -2118 -1460 -2078 1460
rect -5078 -1500 -2078 -1460
rect -1586 1460 1414 1500
rect -1586 -1460 -1546 1460
rect 1374 -1460 1414 1460
rect -1586 -1500 1414 -1460
rect 1906 1460 4906 1500
rect 1906 -1460 1946 1460
rect 4866 -1460 4906 1460
rect 1906 -1500 4906 -1460
<< mimcapcontact >>
rect -5038 -1460 -2118 1460
rect -1546 -1460 1374 1460
rect 1946 -1460 4866 1460
<< metal4 >>
rect -1906 1572 -1810 1588
rect -5039 1460 -2117 1461
rect -5039 -1460 -5038 1460
rect -2118 -1460 -2117 1460
rect -5039 -1461 -2117 -1460
rect -1906 -1572 -1890 1572
rect -1826 -1572 -1810 1572
rect 1586 1572 1682 1588
rect -1547 1460 1375 1461
rect -1547 -1460 -1546 1460
rect 1374 -1460 1375 1460
rect -1547 -1461 1375 -1460
rect -1906 -1588 -1810 -1572
rect 1586 -1572 1602 1572
rect 1666 -1572 1682 1572
rect 5078 1572 5174 1588
rect 1945 1460 4867 1461
rect 1945 -1460 1946 1460
rect 4866 -1460 4867 1460
rect 1945 -1461 4867 -1460
rect 1586 -1588 1682 -1572
rect 5078 -1572 5094 1572
rect 5158 -1572 5174 1572
rect 5078 -1588 5174 -1572
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 1806 -1600 5006 1600
string parameters w 15.0 l 15.0 val 235.2 carea 1.00 cperi 0.17 nx 3 ny 1 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string library sky130
<< end >>
